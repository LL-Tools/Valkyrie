

module b17_C_gen_AntiSAT_k_256_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510;

  AOI22_X1 U11261 ( .A1(n15235), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14249), .B2(n14248), .ZN(n14252) );
  INV_X1 U11262 ( .A(n20313), .ZN(n20288) );
  AND2_X1 U11263 ( .A1(n10401), .A2(n14330), .ZN(n10396) );
  CLKBUF_X2 U11264 ( .A(n15010), .Z(n9843) );
  CLKBUF_X2 U11265 ( .A(n16764), .Z(n9840) );
  OR2_X1 U11266 ( .A1(n13480), .A2(n13476), .ZN(n19899) );
  NAND2_X1 U11267 ( .A1(n11557), .A2(n11586), .ZN(n12986) );
  INV_X1 U11268 ( .A(n17344), .ZN(n13275) );
  INV_X2 U11269 ( .A(n9838), .ZN(n9833) );
  CLKBUF_X2 U11270 ( .A(n17416), .Z(n17398) );
  NOR4_X1 U11271 ( .A1(n15811), .A2(n10412), .A3(n15810), .A4(n15809), .ZN(
        n15812) );
  AND2_X1 U11272 ( .A1(n11061), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12478) );
  AND2_X1 U11273 ( .A1(n9834), .A2(n16502), .ZN(n12479) );
  AND2_X1 U11274 ( .A1(n11020), .A2(n16502), .ZN(n10732) );
  AND2_X1 U11275 ( .A1(n10724), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11087) );
  AND2_X1 U11276 ( .A1(n9827), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12480) );
  INV_X2 U11277 ( .A(n15793), .ZN(n9829) );
  OR4_X1 U11278 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n13107), .ZN(n9846) );
  INV_X1 U11279 ( .A(n11503), .ZN(n11962) );
  INV_X1 U11280 ( .A(n9876), .ZN(n17359) );
  INV_X1 U11281 ( .A(n11449), .ZN(n11456) );
  NAND2_X1 U11282 ( .A1(n10588), .A2(n10587), .ZN(n10620) );
  MUX2_X1 U11283 ( .A(n10574), .B(n10564), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19541) );
  AND2_X2 U11284 ( .A1(n10519), .A2(n10518), .ZN(n12569) );
  INV_X2 U11286 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16502) );
  CLKBUF_X2 U11287 ( .A(n11319), .Z(n13298) );
  AND2_X1 U11288 ( .A1(n11221), .A2(n13291), .ZN(n11402) );
  AND2_X1 U11289 ( .A1(n11227), .A2(n11221), .ZN(n11401) );
  NAND2_X2 U11290 ( .A1(n15675), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11036) );
  AND2_X1 U11291 ( .A1(n13291), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13299) );
  INV_X1 U11293 ( .A(n21510), .ZN(n9818) );
  INV_X1 U11294 ( .A(n11418), .ZN(n12136) );
  INV_X2 U11295 ( .A(n11037), .ZN(n10723) );
  NAND2_X1 U11296 ( .A1(n15664), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9895) );
  AND2_X1 U11297 ( .A1(n10613), .A2(n12575), .ZN(n11113) );
  AND2_X1 U11298 ( .A1(n10723), .A2(n16502), .ZN(n12487) );
  AND2_X1 U11299 ( .A1(n10723), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10747) );
  OR2_X1 U11300 ( .A1(n19156), .A2(n14110), .ZN(n14174) );
  AND2_X1 U11301 ( .A1(n16445), .A2(n16443), .ZN(n13911) );
  AND3_X1 U11302 ( .A1(n10177), .A2(n9945), .A3(n10178), .ZN(n13783) );
  AND2_X1 U11303 ( .A1(n10889), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12488) );
  NOR2_X2 U11304 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U11305 ( .A1(n13502), .A2(n13482), .ZN(n13787) );
  BUF_X1 U11306 ( .A(n13454), .Z(n13500) );
  NAND2_X2 U11307 ( .A1(n11355), .A2(n20423), .ZN(n12318) );
  AND2_X1 U11308 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13012) );
  BUF_X1 U11309 ( .A(n12254), .Z(n13619) );
  AND2_X1 U11310 ( .A1(n12218), .A2(n20478), .ZN(n13632) );
  AND2_X1 U11311 ( .A1(n15070), .A2(n15059), .ZN(n15061) );
  OAI21_X1 U11312 ( .B1(n14185), .B2(n14184), .A(n14187), .ZN(n16346) );
  OAI21_X1 U11313 ( .B1(n15044), .B2(n10259), .A(n10258), .ZN(n15026) );
  INV_X1 U11314 ( .A(n10604), .ZN(n12467) );
  AND2_X1 U11315 ( .A1(n13982), .A2(n15111), .ZN(n15112) );
  AND2_X1 U11316 ( .A1(n15254), .A2(n9875), .ZN(n14225) );
  NAND2_X1 U11317 ( .A1(n10142), .A2(n10141), .ZN(n15292) );
  INV_X2 U11318 ( .A(n9965), .ZN(n9828) );
  INV_X2 U11319 ( .A(n17396), .ZN(n17363) );
  OR3_X1 U11320 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n17118), .ZN(n17238) );
  CLKBUF_X3 U11321 ( .A(n17418), .Z(n9822) );
  INV_X1 U11322 ( .A(n20318), .ZN(n20270) );
  OR2_X1 U11323 ( .A1(n13603), .A2(n13602), .ZN(n13605) );
  AND2_X1 U11324 ( .A1(n15061), .A2(n15050), .ZN(n15052) );
  AND2_X1 U11325 ( .A1(n13992), .A2(n9944), .ZN(n15070) );
  AND2_X1 U11326 ( .A1(n15052), .A2(n15039), .ZN(n15041) );
  NOR2_X1 U11327 ( .A1(n16385), .A2(n15937), .ZN(n15940) );
  OAI21_X1 U11328 ( .B1(n15347), .B2(n15348), .A(n15298), .ZN(n15339) );
  INV_X2 U11329 ( .A(n13155), .ZN(n17376) );
  OAI22_X1 U11330 ( .A1(n18273), .A2(n18088), .B1(n17992), .B2(n17902), .ZN(
        n17974) );
  INV_X1 U11331 ( .A(n13971), .ZN(n15125) );
  OAI21_X1 U11332 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n16288) );
  AOI211_X1 U11333 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n15800), .B(n15799), .ZN(n17584) );
  AND2_X1 U11334 ( .A1(n19541), .A2(n12569), .ZN(n9819) );
  INV_X1 U11335 ( .A(n10419), .ZN(n17418) );
  INV_X1 U11336 ( .A(n9839), .ZN(n20223) );
  OR2_X4 U11337 ( .A1(n12376), .A2(n10407), .ZN(n10646) );
  NAND2_X1 U11338 ( .A1(n12868), .A2(n20423), .ZN(n21104) );
  NOR2_X1 U11339 ( .A1(n14093), .A2(n10280), .ZN(n13434) );
  NOR2_X2 U11341 ( .A1(n14465), .A2(n10318), .ZN(n14429) );
  NAND2_X2 U11342 ( .A1(n17460), .A2(n18449), .ZN(n17596) );
  AOI21_X2 U11343 ( .B1(n16002), .B2(n16001), .A(n19078), .ZN(n17460) );
  NOR2_X2 U11344 ( .A1(n10427), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10429) );
  NOR2_X2 U11345 ( .A1(n16346), .A2(n14110), .ZN(n14186) );
  NAND2_X2 U11346 ( .A1(n11416), .A2(n11383), .ZN(n10308) );
  INV_X2 U11347 ( .A(n12569), .ZN(n19565) );
  BUF_X2 U11348 ( .A(n18894), .Z(n9820) );
  INV_X2 U11349 ( .A(n12070), .ZN(n9821) );
  INV_X4 U11350 ( .A(n12153), .ZN(n9823) );
  INV_X1 U11351 ( .A(n9823), .ZN(n9824) );
  NAND2_X1 U11352 ( .A1(n14971), .A2(n10058), .ZN(n12153) );
  AND2_X4 U11353 ( .A1(n15948), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11227) );
  CLKBUF_X3 U11354 ( .A(n11319), .Z(n12163) );
  INV_X1 U11355 ( .A(n18068), .ZN(n9825) );
  INV_X1 U11356 ( .A(n9825), .ZN(n9826) );
  INV_X1 U11357 ( .A(n11027), .ZN(n9827) );
  NAND2_X2 U11358 ( .A1(n13012), .A2(n10428), .ZN(n11027) );
  CLKBUF_X1 U11359 ( .A(n11036), .Z(n9837) );
  AOI21_X2 U11361 ( .B1(n15339), .B2(n15300), .A(n15299), .ZN(n15316) );
  NOR3_X4 U11362 ( .A1(n13721), .A2(n10255), .A3(n10252), .ZN(n13982) );
  OAI21_X1 U11363 ( .B1(n13583), .B2(n14183), .A(n15000), .ZN(n13549) );
  AOI211_X2 U11364 ( .C1(n16314), .C2(n19510), .A(n15259), .B(n15258), .ZN(
        n15260) );
  NAND2_X2 U11365 ( .A1(n9998), .A2(n9996), .ZN(n15022) );
  NAND2_X2 U11366 ( .A1(n15032), .A2(n11026), .ZN(n9998) );
  OR2_X1 U11367 ( .A1(n15044), .A2(n15043), .ZN(n10262) );
  OAI21_X1 U11368 ( .B1(n14784), .B2(n14337), .A(n14334), .ZN(n14759) );
  AOI21_X2 U11369 ( .B1(n15292), .B2(n14179), .A(n14178), .ZN(n15451) );
  NOR2_X1 U11370 ( .A1(n15128), .A2(n15120), .ZN(n14401) );
  XNOR2_X1 U11371 ( .A(n15128), .B(n10249), .ZN(n16268) );
  AND2_X1 U11372 ( .A1(n15130), .A2(n14292), .ZN(n16290) );
  NAND2_X1 U11373 ( .A1(n13725), .A2(n10886), .ZN(n10921) );
  AND2_X1 U11374 ( .A1(n14023), .A2(n14024), .ZN(n15199) );
  XNOR2_X1 U11375 ( .A(n13783), .B(n13782), .ZN(n13872) );
  INV_X1 U11376 ( .A(n14336), .ZN(n14833) );
  AND2_X1 U11377 ( .A1(n12546), .A2(n13609), .ZN(n13655) );
  OAI22_X1 U11378 ( .A1(n13515), .A2(n19899), .B1(n19938), .B2(n13514), .ZN(
        n13518) );
  OR2_X1 U11380 ( .A1(n13480), .A2(n13471), .ZN(n20011) );
  INV_X1 U11381 ( .A(n13787), .ZN(n19672) );
  NOR2_X2 U11382 ( .A1(n19547), .A2(n19564), .ZN(n19548) );
  OR2_X1 U11383 ( .A1(n13497), .A2(n13496), .ZN(n19572) );
  OR2_X1 U11384 ( .A1(n13497), .A2(n13476), .ZN(n19516) );
  OR2_X1 U11385 ( .A1(n13497), .A2(n13471), .ZN(n19636) );
  AND4_X1 U11386 ( .A1(n10070), .A2(n10071), .A3(n10069), .A4(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17993) );
  NAND2_X1 U11387 ( .A1(n9879), .A2(n14194), .ZN(n14112) );
  NAND2_X1 U11388 ( .A1(n10703), .A2(n10702), .ZN(n19350) );
  OAI21_X1 U11389 ( .B1(n18878), .B2(n18437), .A(n15736), .ZN(n18883) );
  NAND2_X1 U11390 ( .A1(n13926), .A2(n13924), .ZN(n14096) );
  BUF_X2 U11391 ( .A(n11113), .Z(n14227) );
  XOR2_X1 U11392 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16567), .Z(
        n16764) );
  INV_X2 U11393 ( .A(n11196), .ZN(n14228) );
  NAND2_X2 U11394 ( .A1(n12367), .A2(n15745), .ZN(n12376) );
  NOR2_X1 U11395 ( .A1(n11359), .A2(n11369), .ZN(n11302) );
  CLKBUF_X2 U11396 ( .A(n12467), .Z(n9838) );
  INV_X2 U11397 ( .A(n20463), .ZN(n12218) );
  INV_X2 U11398 ( .A(n20446), .ZN(n12965) );
  INV_X2 U11399 ( .A(n11576), .ZN(n20471) );
  OAI211_X1 U11400 ( .C1(n13155), .C2(n17406), .A(n13210), .B(n13209), .ZN(
        n18416) );
  NAND2_X2 U11401 ( .A1(n20217), .A2(n10604), .ZN(n12581) );
  CLKBUF_X2 U11402 ( .A(n12402), .Z(n14208) );
  NAND2_X1 U11403 ( .A1(n19554), .A2(n12402), .ZN(n12507) );
  NAND2_X1 U11404 ( .A1(n18765), .A2(n18713), .ZN(n18797) );
  CLKBUF_X2 U11405 ( .A(n10718), .Z(n11057) );
  CLKBUF_X2 U11406 ( .A(n11422), .Z(n12076) );
  INV_X4 U11407 ( .A(n12070), .ZN(n12137) );
  INV_X1 U11408 ( .A(n11308), .ZN(n12155) );
  INV_X4 U11409 ( .A(n12018), .ZN(n11900) );
  INV_X4 U11410 ( .A(n10541), .ZN(n10718) );
  INV_X4 U11411 ( .A(n17238), .ZN(n17417) );
  INV_X4 U11412 ( .A(n9846), .ZN(n17318) );
  INV_X4 U11413 ( .A(n17328), .ZN(n9830) );
  INV_X4 U11414 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19037) );
  XNOR2_X1 U11415 ( .A(n10138), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14851) );
  AND2_X1 U11416 ( .A1(n15543), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15515) );
  NOR2_X1 U11417 ( .A1(n15555), .A2(n15549), .ZN(n15543) );
  AND2_X1 U11418 ( .A1(n10261), .A2(n11011), .ZN(n9855) );
  NAND2_X1 U11419 ( .A1(n10346), .A2(n10351), .ZN(n15274) );
  OR2_X1 U11420 ( .A1(n15578), .A2(n15563), .ZN(n15555) );
  AOI21_X1 U11421 ( .B1(n16268), .B2(n16485), .A(n10247), .ZN(n15374) );
  NAND2_X1 U11422 ( .A1(n15047), .A2(n10405), .ZN(n10986) );
  NAND2_X1 U11423 ( .A1(n15049), .A2(n15048), .ZN(n15047) );
  AND2_X1 U11424 ( .A1(n15121), .A2(n10272), .ZN(n10271) );
  OR2_X1 U11425 ( .A1(n15019), .A2(n14257), .ZN(n15031) );
  AND2_X1 U11426 ( .A1(n14327), .A2(n10402), .ZN(n10401) );
  NAND2_X1 U11427 ( .A1(n13881), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13916) );
  AND2_X1 U11428 ( .A1(n15076), .A2(n10940), .ZN(n10922) );
  INV_X1 U11429 ( .A(n10393), .ZN(n10394) );
  NOR2_X1 U11430 ( .A1(n10393), .A2(n10135), .ZN(n10133) );
  OR2_X1 U11431 ( .A1(n10066), .A2(n14321), .ZN(n10393) );
  NOR2_X1 U11432 ( .A1(n16071), .A2(n14802), .ZN(n14335) );
  INV_X1 U11433 ( .A(n17757), .ZN(n10044) );
  NOR2_X1 U11434 ( .A1(n14246), .A2(n14203), .ZN(n14206) );
  NAND2_X1 U11435 ( .A1(n10388), .A2(n10389), .ZN(n16107) );
  OR2_X1 U11436 ( .A1(n17770), .A2(n15863), .ZN(n17756) );
  AND2_X1 U11437 ( .A1(n13919), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14218) );
  XNOR2_X1 U11438 ( .A(n10921), .B(n10940), .ZN(n15065) );
  AND2_X1 U11439 ( .A1(n15142), .A2(n15143), .ZN(n15145) );
  OR2_X1 U11440 ( .A1(n10400), .A2(n10399), .ZN(n10398) );
  OR2_X1 U11441 ( .A1(n14790), .A2(n16080), .ZN(n16071) );
  AND3_X1 U11442 ( .A1(n10081), .A2(n9873), .A3(n17854), .ZN(n17757) );
  OR3_X1 U11443 ( .A1(n14821), .A2(n14820), .A3(n14814), .ZN(n14804) );
  NAND2_X1 U11444 ( .A1(n17854), .A2(n10080), .ZN(n17781) );
  NAND2_X1 U11445 ( .A1(n14196), .A2(n10202), .ZN(n14201) );
  NAND2_X1 U11446 ( .A1(n17780), .A2(n17816), .ZN(n17854) );
  AND2_X1 U11447 ( .A1(n10123), .A2(n10387), .ZN(n13680) );
  AND2_X1 U11448 ( .A1(n14783), .A2(n9972), .ZN(n10129) );
  OR2_X1 U11449 ( .A1(n13869), .A2(n16497), .ZN(n16444) );
  INV_X2 U11450 ( .A(n14833), .ZN(n14805) );
  NAND2_X1 U11451 ( .A1(n15199), .A2(n15198), .ZN(n15200) );
  NOR2_X1 U11452 ( .A1(n16784), .A2(n16785), .ZN(n16783) );
  NAND2_X1 U11453 ( .A1(n13783), .A2(n13782), .ZN(n13821) );
  NAND2_X1 U11454 ( .A1(n13655), .A2(n13654), .ZN(n13721) );
  NOR2_X1 U11455 ( .A1(n13101), .A2(n13383), .ZN(n11610) );
  NOR2_X1 U11456 ( .A1(n14189), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14193) );
  NOR3_X1 U11457 ( .A1(n18919), .A2(n19078), .A3(n10019), .ZN(n19028) );
  AND2_X1 U11458 ( .A1(n13861), .A2(n13860), .ZN(n13862) );
  OR2_X1 U11459 ( .A1(n10213), .A2(n14146), .ZN(n10212) );
  AND2_X1 U11460 ( .A1(n12547), .A2(n13435), .ZN(n12546) );
  OAI21_X1 U11461 ( .B1(n18077), .B2(n17823), .A(n18797), .ZN(n17926) );
  NOR2_X1 U11462 ( .A1(n14132), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10213) );
  AND2_X1 U11463 ( .A1(n13368), .A2(n9863), .ZN(n13435) );
  NAND2_X1 U11464 ( .A1(n10275), .A2(n9857), .ZN(n10004) );
  NAND2_X2 U11465 ( .A1(n14674), .A2(n13633), .ZN(n14672) );
  NAND2_X1 U11466 ( .A1(n10137), .A2(n9940), .ZN(n11635) );
  INV_X1 U11467 ( .A(n11597), .ZN(n10137) );
  NOR2_X1 U11468 ( .A1(n14158), .A2(n14128), .ZN(n14141) );
  NAND2_X1 U11469 ( .A1(n12627), .A2(n20204), .ZN(n16477) );
  NAND2_X1 U11470 ( .A1(n13932), .A2(n16468), .ZN(n16467) );
  NOR2_X1 U11471 ( .A1(n17539), .A2(n17713), .ZN(n17535) );
  NAND2_X1 U11472 ( .A1(n13500), .A2(n13490), .ZN(n13531) );
  NOR2_X1 U11473 ( .A1(n13588), .A2(n13587), .ZN(n14082) );
  NAND2_X1 U11474 ( .A1(n13500), .A2(n13501), .ZN(n13784) );
  NAND2_X1 U11475 ( .A1(n13500), .A2(n13489), .ZN(n19868) );
  AND2_X1 U11476 ( .A1(n14157), .A2(n14148), .ZN(n19185) );
  NAND2_X1 U11477 ( .A1(n9992), .A2(n9955), .ZN(n14158) );
  NAND2_X1 U11478 ( .A1(n10057), .A2(n13347), .ZN(n11597) );
  NAND2_X1 U11479 ( .A1(n18083), .A2(n18044), .ZN(n18078) );
  NAND2_X1 U11480 ( .A1(n13500), .A2(n13482), .ZN(n19786) );
  NOR2_X2 U11481 ( .A1(n19535), .A2(n20019), .ZN(n19536) );
  NOR2_X2 U11482 ( .A1(n19435), .A2(n20019), .ZN(n13458) );
  NOR2_X2 U11483 ( .A1(n19531), .A2(n20019), .ZN(n19532) );
  OR2_X1 U11484 ( .A1(n13497), .A2(n13495), .ZN(n13805) );
  NOR2_X2 U11485 ( .A1(n19526), .A2(n20019), .ZN(n19527) );
  NOR2_X1 U11486 ( .A1(n13971), .A2(n13462), .ZN(n19559) );
  NOR2_X1 U11487 ( .A1(n15125), .A2(n13462), .ZN(n19558) );
  NOR2_X2 U11488 ( .A1(n19542), .A2(n20019), .ZN(n19543) );
  INV_X1 U11489 ( .A(n14153), .ZN(n9992) );
  INV_X2 U11490 ( .A(n14824), .ZN(n20365) );
  NOR2_X2 U11491 ( .A1(n19549), .A2(n20019), .ZN(n19550) );
  NAND2_X1 U11492 ( .A1(n10001), .A2(n10695), .ZN(n10712) );
  INV_X2 U11493 ( .A(n15104), .ZN(n9831) );
  AND2_X1 U11494 ( .A1(n14060), .A2(n14059), .ZN(n14607) );
  AND2_X1 U11495 ( .A1(n13893), .A2(n13892), .ZN(n13895) );
  NAND2_X1 U11496 ( .A1(n18870), .A2(n16557), .ZN(n18086) );
  NAND2_X1 U11497 ( .A1(n18870), .A2(n18920), .ZN(n16733) );
  NAND2_X1 U11498 ( .A1(n12791), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12981) );
  AND2_X1 U11499 ( .A1(n11435), .A2(n11434), .ZN(n12962) );
  OR2_X1 U11500 ( .A1(n11129), .A2(n10674), .ZN(n10679) );
  AND2_X1 U11501 ( .A1(n11485), .A2(n11484), .ZN(n11563) );
  NOR2_X1 U11502 ( .A1(n18016), .A2(n15835), .ZN(n15849) );
  OR2_X1 U11503 ( .A1(n13479), .A2(n15653), .ZN(n13476) );
  NOR3_X1 U11504 ( .A1(n18416), .A2(n10172), .A3(n18874), .ZN(n10171) );
  AND2_X1 U11505 ( .A1(n12837), .A2(n10232), .ZN(n16481) );
  OR2_X1 U11506 ( .A1(n11483), .A2(n11482), .ZN(n11485) );
  NAND2_X1 U11507 ( .A1(n20551), .A2(n11415), .ZN(n20890) );
  CLKBUF_X1 U11508 ( .A(n11416), .Z(n11417) );
  NAND2_X1 U11509 ( .A1(n11575), .A2(n11574), .ZN(n20513) );
  NAND2_X1 U11510 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  NAND2_X1 U11511 ( .A1(n10175), .A2(n15889), .ZN(n18892) );
  OR2_X1 U11512 ( .A1(n18883), .A2(n15890), .ZN(n10175) );
  NAND2_X1 U11513 ( .A1(n9991), .A2(n9952), .ZN(n14105) );
  NAND2_X1 U11514 ( .A1(n10701), .A2(n10700), .ZN(n10703) );
  NOR2_X1 U11515 ( .A1(n15821), .A2(n15820), .ZN(n15822) );
  NOR2_X2 U11516 ( .A1(n18883), .A2(n10201), .ZN(n18881) );
  XNOR2_X1 U11517 ( .A(n11136), .B(n11137), .ZN(n11134) );
  OR2_X1 U11518 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  AND2_X1 U11519 ( .A1(n11438), .A2(n11436), .ZN(n11414) );
  XNOR2_X1 U11520 ( .A(n11367), .B(n11380), .ZN(n11413) );
  INV_X1 U11521 ( .A(n14096), .ZN(n9991) );
  OAI211_X1 U11522 ( .C1(n15976), .C2(n20764), .A(n11390), .B(n11389), .ZN(
        n11391) );
  OAI21_X1 U11523 ( .B1(n11112), .B2(n13547), .A(n10617), .ZN(n11136) );
  OAI211_X1 U11524 ( .C1(n11112), .C2(n15654), .A(n10413), .B(n10658), .ZN(
        n10701) );
  OR2_X1 U11525 ( .A1(n10042), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U11526 ( .A1(n11491), .A2(n11490), .ZN(n20588) );
  NAND2_X1 U11527 ( .A1(n9890), .A2(n10642), .ZN(n10691) );
  OAI21_X1 U11528 ( .B1(n15735), .B2(n15890), .A(n15889), .ZN(n18878) );
  OR2_X1 U11529 ( .A1(n12780), .A2(n12779), .ZN(n12782) );
  OR2_X1 U11530 ( .A1(n11384), .A2(n11208), .ZN(n11390) );
  NOR2_X1 U11531 ( .A1(n10657), .A2(n10414), .ZN(n10658) );
  AND2_X1 U11532 ( .A1(n10648), .A2(n10647), .ZN(n10669) );
  AOI21_X1 U11533 ( .B1(n10661), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10643), .ZN(n11131) );
  NAND2_X2 U11534 ( .A1(n18915), .A2(n17648), .ZN(n17712) );
  NAND2_X1 U11535 ( .A1(n9914), .A2(n10002), .ZN(n10661) );
  NOR2_X1 U11536 ( .A1(n10160), .A2(n10157), .ZN(n15732) );
  NAND2_X1 U11537 ( .A1(n10165), .A2(n10164), .ZN(n15736) );
  OR2_X1 U11538 ( .A1(n15726), .A2(n9877), .ZN(n10165) );
  OR2_X1 U11539 ( .A1(n15723), .A2(n10161), .ZN(n10160) );
  NOR2_X1 U11540 ( .A1(n12827), .A2(n12829), .ZN(n13546) );
  NAND2_X1 U11541 ( .A1(n20223), .A2(n13364), .ZN(n10688) );
  NAND2_X2 U11542 ( .A1(n10611), .A2(n9889), .ZN(n11196) );
  OAI21_X1 U11543 ( .B1(n10622), .B2(n10623), .A(n10621), .ZN(n10339) );
  INV_X4 U11544 ( .A(n12473), .ZN(n14399) );
  OR2_X1 U11545 ( .A1(n15721), .A2(n18426), .ZN(n10158) );
  AND2_X1 U11546 ( .A1(n11358), .A2(n11373), .ZN(n12879) );
  AND3_X1 U11547 ( .A1(n11302), .A2(n11303), .A3(n10103), .ZN(n12642) );
  AND2_X1 U11548 ( .A1(n18449), .A2(n17068), .ZN(n15721) );
  AND3_X1 U11549 ( .A1(n9819), .A2(n10605), .A3(n10628), .ZN(n12575) );
  OAI211_X1 U11550 ( .C1(n9847), .C2(n12581), .A(n9986), .B(n9984), .ZN(n12587) );
  INV_X1 U11551 ( .A(n12563), .ZN(n12607) );
  INV_X1 U11552 ( .A(n17068), .ZN(n18412) );
  INV_X1 U11553 ( .A(n15715), .ZN(n18437) );
  INV_X1 U11554 ( .A(n15872), .ZN(n18432) );
  AND2_X1 U11555 ( .A1(n11360), .A2(n20452), .ZN(n11369) );
  NAND2_X1 U11556 ( .A1(n17068), .A2(n18416), .ZN(n15887) );
  INV_X1 U11557 ( .A(n15734), .ZN(n18426) );
  OR2_X1 U11558 ( .A1(n12401), .A2(n12400), .ZN(n12847) );
  OR2_X1 U11559 ( .A1(n10573), .A2(n10572), .ZN(n10588) );
  AND2_X1 U11560 ( .A1(n19554), .A2(n10552), .ZN(n10605) );
  INV_X1 U11561 ( .A(n18443), .ZN(n17463) );
  OR2_X1 U11562 ( .A1(n12413), .A2(n12412), .ZN(n13511) );
  NAND2_X1 U11563 ( .A1(n13394), .A2(n20440), .ZN(n13403) );
  INV_X2 U11564 ( .A(n18416), .ZN(n19084) );
  AND2_X1 U11565 ( .A1(n10618), .A2(n12614), .ZN(n10628) );
  OR2_X1 U11566 ( .A1(n11455), .A2(n11454), .ZN(n13771) );
  OR2_X1 U11567 ( .A1(n12497), .A2(n12496), .ZN(n12722) );
  OAI211_X1 U11568 ( .C1(n17238), .C2(n18446), .A(n13183), .B(n13182), .ZN(
        n18443) );
  OAI211_X1 U11569 ( .C1(n10419), .C2(n17262), .A(n13163), .B(n13162), .ZN(
        n18421) );
  AND2_X1 U11570 ( .A1(n10470), .A2(n10469), .ZN(n12614) );
  INV_X1 U11571 ( .A(n19554), .ZN(n10714) );
  INV_X1 U11572 ( .A(n20440), .ZN(n12868) );
  INV_X2 U11573 ( .A(n20217), .ZN(n16528) );
  INV_X1 U11574 ( .A(n20423), .ZN(n13394) );
  AND3_X2 U11575 ( .A1(n9858), .A2(n11235), .A3(n11233), .ZN(n11354) );
  OR2_X2 U11576 ( .A1(n11288), .A2(n11287), .ZN(n20452) );
  NAND2_X2 U11577 ( .A1(n10013), .A2(n10012), .ZN(n20217) );
  NAND2_X1 U11578 ( .A1(n10551), .A2(n10550), .ZN(n12402) );
  OR2_X1 U11579 ( .A1(n11274), .A2(n11273), .ZN(n20446) );
  OR2_X2 U11580 ( .A1(n16682), .A2(n16633), .ZN(n16685) );
  AND2_X1 U11581 ( .A1(n17927), .A2(n9926), .ZN(n17824) );
  NAND2_X1 U11582 ( .A1(n10580), .A2(n16502), .ZN(n10518) );
  NOR2_X1 U11583 ( .A1(n10517), .A2(n10516), .ZN(n10580) );
  NOR2_X1 U11584 ( .A1(n10528), .A2(n10527), .ZN(n10579) );
  NOR2_X1 U11585 ( .A1(n10538), .A2(n10537), .ZN(n10565) );
  AND4_X1 U11586 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11259) );
  OR2_X1 U11587 ( .A1(n12155), .A2(n11327), .ZN(n11331) );
  BUF_X2 U11588 ( .A(n15837), .Z(n17411) );
  NOR2_X1 U11590 ( .A1(n19273), .A2(n12362), .ZN(n12364) );
  INV_X2 U11591 ( .A(n11036), .ZN(n10724) );
  INV_X2 U11592 ( .A(n12128), .ZN(n12164) );
  AND2_X2 U11593 ( .A1(n9834), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12481) );
  NAND2_X2 U11594 ( .A1(n19092), .A2(n18953), .ZN(n19011) );
  CLKBUF_X2 U11595 ( .A(n17637), .Z(n19079) );
  NAND2_X1 U11596 ( .A1(n13292), .A2(n13291), .ZN(n12128) );
  INV_X2 U11597 ( .A(n16721), .ZN(n16723) );
  NOR2_X1 U11598 ( .A1(n19042), .A2(n18936), .ZN(n17637) );
  NAND2_X2 U11599 ( .A1(n15663), .A2(n11072), .ZN(n10541) );
  NAND2_X1 U11600 ( .A1(n11226), .A2(n13292), .ZN(n12018) );
  CLKBUF_X1 U11601 ( .A(n11037), .Z(n9836) );
  OR2_X1 U11602 ( .A1(n13110), .A2(n13111), .ZN(n17377) );
  NAND2_X1 U11603 ( .A1(n13107), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13111) );
  NAND2_X1 U11604 ( .A1(n19037), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13110) );
  NAND3_X1 U11605 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n19055), .ZN(n13108) );
  NAND2_X1 U11606 ( .A1(n13184), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13112) );
  AND2_X1 U11607 ( .A1(n10431), .A2(n15665), .ZN(n15663) );
  INV_X2 U11608 ( .A(n18388), .ZN(n9832) );
  NOR2_X2 U11609 ( .A1(n11208), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13295) );
  AND2_X1 U11610 ( .A1(n11221), .A2(n14971), .ZN(n11949) );
  AND2_X1 U11611 ( .A1(n12893), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11226) );
  INV_X1 U11612 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12893) );
  INV_X1 U11613 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11072) );
  INV_X1 U11614 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10428) );
  INV_X1 U11615 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15665) );
  INV_X1 U11616 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13469) );
  OR2_X2 U11617 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17118) );
  NAND2_X1 U11618 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18879) );
  INV_X1 U11619 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19055) );
  AND2_X1 U11620 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10058) );
  OR2_X2 U11621 ( .A1(n15266), .A2(n10146), .ZN(n15246) );
  NOR2_X1 U11622 ( .A1(n17858), .A2(n17929), .ZN(n18068) );
  INV_X2 U11623 ( .A(n11028), .ZN(n9834) );
  OAI21_X1 U11624 ( .B1(n13583), .B2(n13582), .A(n13585), .ZN(n13871) );
  AND2_X1 U11625 ( .A1(n15653), .A2(n10696), .ZN(n13489) );
  NOR2_X1 U11626 ( .A1(n17118), .A2(n13110), .ZN(n9835) );
  NOR2_X1 U11627 ( .A1(n17118), .A2(n13110), .ZN(n17360) );
  NAND3_X2 U11628 ( .A1(n10431), .A2(n10427), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11037) );
  BUF_X4 U11629 ( .A(n12467), .Z(n9839) );
  AND2_X1 U11630 ( .A1(n9833), .A2(n12466), .ZN(n9841) );
  AND2_X1 U11631 ( .A1(n9833), .A2(n12466), .ZN(n9842) );
  AND2_X2 U11632 ( .A1(n11057), .A2(n16502), .ZN(n12416) );
  NAND2_X1 U11633 ( .A1(n12969), .A2(n12968), .ZN(n12983) );
  INV_X1 U11634 ( .A(n12457), .ZN(n14110) );
  NAND2_X1 U11635 ( .A1(n18449), .A2(n18426), .ZN(n15729) );
  INV_X1 U11636 ( .A(n15887), .ZN(n10164) );
  AND2_X1 U11637 ( .A1(n12892), .A2(n12218), .ZN(n12239) );
  INV_X1 U11638 ( .A(n13905), .ZN(n10066) );
  INV_X1 U11639 ( .A(n11586), .ZN(n10057) );
  AND2_X1 U11640 ( .A1(n13295), .A2(n11226), .ZN(n11422) );
  NAND2_X1 U11641 ( .A1(n20588), .A2(n10062), .ZN(n10114) );
  NAND2_X1 U11642 ( .A1(n13819), .A2(n9907), .ZN(n13917) );
  INV_X1 U11643 ( .A(n13821), .ZN(n13819) );
  AND2_X1 U11644 ( .A1(n9839), .A2(n12466), .ZN(n12468) );
  NAND2_X1 U11645 ( .A1(n12507), .A2(n12614), .ZN(n10619) );
  NAND2_X1 U11646 ( .A1(n15819), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10075) );
  AOI21_X1 U11647 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18405), .A(
        n13194), .ZN(n15712) );
  NAND2_X1 U11648 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  OR2_X1 U11649 ( .A1(n18432), .A2(n16003), .ZN(n10162) );
  NAND2_X1 U11650 ( .A1(n15724), .A2(n15725), .ZN(n10163) );
  NAND2_X1 U11651 ( .A1(n15722), .A2(n18432), .ZN(n10159) );
  OAI21_X1 U11652 ( .B1(n15734), .B2(n15733), .A(n15732), .ZN(n15738) );
  NAND2_X1 U11653 ( .A1(n14441), .A2(n10322), .ZN(n10321) );
  INV_X1 U11654 ( .A(n14455), .ZN(n10322) );
  NAND2_X1 U11655 ( .A1(n16107), .A2(n16105), .ZN(n10136) );
  NAND2_X1 U11656 ( .A1(n11361), .A2(n12736), .ZN(n14368) );
  NOR2_X1 U11657 ( .A1(n11334), .A2(n11333), .ZN(n11350) );
  INV_X1 U11658 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11332) );
  INV_X1 U11659 ( .A(n10688), .ZN(n11008) );
  NAND2_X1 U11660 ( .A1(n10239), .A2(n14000), .ZN(n10238) );
  INV_X1 U11661 ( .A(n15545), .ZN(n10239) );
  AOI21_X1 U11662 ( .B1(n10661), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10637), .ZN(n11137) );
  AND2_X1 U11663 ( .A1(n14194), .A2(n14243), .ZN(n14213) );
  NAND2_X1 U11664 ( .A1(n10203), .A2(n14201), .ZN(n10371) );
  NAND2_X1 U11665 ( .A1(n9887), .A2(n10143), .ZN(n10141) );
  NOR2_X1 U11666 ( .A1(n10184), .A2(n16421), .ZN(n10183) );
  OR2_X1 U11667 ( .A1(n13112), .A2(n13111), .ZN(n9876) );
  NOR2_X2 U11668 ( .A1(n18879), .A2(n13110), .ZN(n17416) );
  AOI21_X1 U11669 ( .B1(n15736), .B2(n10030), .A(n15738), .ZN(n15889) );
  AND2_X1 U11670 ( .A1(n15729), .A2(n18416), .ZN(n10030) );
  OR2_X1 U11671 ( .A1(n13620), .A2(n12740), .ZN(n12914) );
  INV_X2 U11672 ( .A(n11633), .ZN(n12180) );
  AND2_X1 U11673 ( .A1(n15976), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13627) );
  NOR2_X1 U11674 ( .A1(n11216), .A2(n11215), .ZN(n11235) );
  INV_X1 U11675 ( .A(n14956), .ZN(n13690) );
  INV_X1 U11676 ( .A(n12217), .ZN(n10310) );
  BUF_X1 U11677 ( .A(n11112), .Z(n14232) );
  AND4_X1 U11678 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12455) );
  AND4_X1 U11679 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12453) );
  AND4_X1 U11680 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12454) );
  OR2_X1 U11681 ( .A1(n15243), .A2(n15263), .ZN(n10146) );
  XNOR2_X1 U11682 ( .A(n10703), .B(n10696), .ZN(n13479) );
  AND2_X1 U11683 ( .A1(n12603), .A2(n16551), .ZN(n12627) );
  XNOR2_X1 U11684 ( .A(n15655), .B(n10707), .ZN(n13357) );
  OR2_X1 U11685 ( .A1(n13112), .A2(n17118), .ZN(n17328) );
  NAND2_X1 U11686 ( .A1(n10035), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10032) );
  AND2_X1 U11687 ( .A1(n10029), .A2(n10027), .ZN(n17068) );
  INV_X1 U11688 ( .A(n13129), .ZN(n10029) );
  NOR2_X1 U11689 ( .A1(n13130), .A2(n10028), .ZN(n10027) );
  OAI21_X1 U11690 ( .B1(n18881), .B2(n10200), .A(n10199), .ZN(n16002) );
  NOR2_X1 U11691 ( .A1(n16731), .A2(n18938), .ZN(n10199) );
  OAI22_X2 U11692 ( .A1(n18869), .A2(n10170), .B1(n18863), .B2(n16556), .ZN(
        n18870) );
  NAND2_X1 U11693 ( .A1(n10044), .A2(n15863), .ZN(n10422) );
  NAND2_X1 U11694 ( .A1(n10084), .A2(n18190), .ZN(n17799) );
  INV_X1 U11695 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20199) );
  NOR2_X2 U11696 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20169) );
  INV_X1 U11697 ( .A(n11375), .ZN(n10109) );
  NAND2_X1 U11698 ( .A1(n12252), .A2(n12737), .ZN(n10378) );
  NOR2_X2 U11699 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11221) );
  NAND2_X1 U11700 ( .A1(n11226), .A2(n11221), .ZN(n12070) );
  NOR2_X1 U11701 ( .A1(n12893), .A2(n10062), .ZN(n10107) );
  NAND2_X1 U11702 ( .A1(n11366), .A2(n10107), .ZN(n10105) );
  INV_X1 U11703 ( .A(n13820), .ZN(n13818) );
  AND2_X1 U11704 ( .A1(n11543), .A2(n11542), .ZN(n11545) );
  NAND2_X1 U11705 ( .A1(n11626), .A2(n11625), .ZN(n11636) );
  INV_X1 U11706 ( .A(n11544), .ZN(n11596) );
  NOR2_X1 U11707 ( .A1(n15948), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U11708 ( .A1(n11366), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11380) );
  NOR2_X1 U11709 ( .A1(n10211), .A2(n14182), .ZN(n10210) );
  INV_X1 U11710 ( .A(n14184), .ZN(n10211) );
  INV_X1 U11711 ( .A(n15055), .ZN(n10279) );
  AND2_X1 U11712 ( .A1(n10279), .A2(n15064), .ZN(n10277) );
  AND2_X1 U11713 ( .A1(n15617), .A2(n10357), .ZN(n10356) );
  INV_X1 U11714 ( .A(n15632), .ZN(n10357) );
  NAND2_X1 U11715 ( .A1(n10014), .A2(n10618), .ZN(n12563) );
  INV_X1 U11716 ( .A(n19541), .ZN(n12568) );
  INV_X1 U11717 ( .A(n10056), .ZN(n15801) );
  OR2_X1 U11718 ( .A1(n17591), .A2(n15903), .ZN(n10056) );
  INV_X1 U11719 ( .A(n13141), .ZN(n10026) );
  INV_X1 U11720 ( .A(n12148), .ZN(n12175) );
  AND2_X1 U11721 ( .A1(n10324), .A2(n14494), .ZN(n10323) );
  NOR2_X1 U11722 ( .A1(n14509), .A2(n10325), .ZN(n10324) );
  INV_X1 U11723 ( .A(n10326), .ZN(n10325) );
  NOR2_X1 U11724 ( .A1(n14521), .A2(n10327), .ZN(n10326) );
  INV_X1 U11725 ( .A(n14575), .ZN(n10327) );
  OR2_X1 U11726 ( .A1(n13978), .A2(n14035), .ZN(n10317) );
  AND2_X1 U11727 ( .A1(n14039), .A2(n14049), .ZN(n11763) );
  INV_X1 U11728 ( .A(n11762), .ZN(n11796) );
  INV_X1 U11729 ( .A(n10129), .ZN(n10128) );
  NAND2_X1 U11730 ( .A1(n12293), .A2(n10337), .ZN(n10336) );
  OR2_X1 U11731 ( .A1(n13734), .A2(n14070), .ZN(n10333) );
  OR2_X1 U11732 ( .A1(n13754), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13752) );
  NAND2_X1 U11733 ( .A1(n13671), .A2(n13766), .ZN(n13678) );
  INV_X1 U11734 ( .A(n16117), .ZN(n13679) );
  NAND2_X1 U11735 ( .A1(n11414), .A2(n11413), .ZN(n11416) );
  OAI21_X1 U11736 ( .B1(n21105), .B2(n13321), .A(n14986), .ZN(n20422) );
  AOI21_X1 U11737 ( .B1(n10780), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(n9888), .ZN(n9985) );
  OR3_X1 U11738 ( .A1(n11100), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n16517), .ZN(n12368) );
  NOR2_X1 U11739 ( .A1(n9994), .A2(n14123), .ZN(n9993) );
  INV_X1 U11740 ( .A(n14111), .ZN(n9994) );
  NAND2_X1 U11741 ( .A1(n13440), .A2(n10207), .ZN(n10206) );
  NAND2_X1 U11742 ( .A1(n13865), .A2(n13823), .ZN(n9989) );
  NOR2_X1 U11743 ( .A1(n9990), .A2(n9988), .ZN(n13866) );
  INV_X1 U11744 ( .A(n13823), .ZN(n9988) );
  NAND2_X1 U11745 ( .A1(n13546), .A2(n13545), .ZN(n13579) );
  NAND2_X1 U11746 ( .A1(n11129), .A2(n11131), .ZN(n11132) );
  OAI21_X1 U11747 ( .B1(n11129), .B2(n11131), .A(n11130), .ZN(n11133) );
  INV_X1 U11748 ( .A(n12514), .ZN(n13542) );
  NAND2_X1 U11749 ( .A1(n9911), .A2(n10003), .ZN(n10002) );
  INV_X1 U11750 ( .A(n10659), .ZN(n10003) );
  INV_X1 U11751 ( .A(n15225), .ZN(n10365) );
  AND2_X1 U11752 ( .A1(n15448), .A2(n15449), .ZN(n10352) );
  INV_X1 U11753 ( .A(n15286), .ZN(n9995) );
  INV_X1 U11754 ( .A(n9956), .ZN(n10254) );
  INV_X1 U11755 ( .A(n13722), .ZN(n10253) );
  AND2_X1 U11756 ( .A1(n19219), .A2(n14183), .ZN(n14172) );
  OR2_X1 U11757 ( .A1(n10244), .A2(n12544), .ZN(n10243) );
  INV_X1 U11758 ( .A(n13826), .ZN(n10342) );
  NAND2_X1 U11759 ( .A1(n14994), .A2(n19509), .ZN(n13480) );
  NAND2_X1 U11760 ( .A1(n10583), .A2(n16502), .ZN(n10469) );
  NAND2_X1 U11761 ( .A1(n10563), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10470) );
  INV_X1 U11762 ( .A(n17716), .ZN(n10095) );
  INV_X1 U11763 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15792) );
  INV_X1 U11764 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15752) );
  NOR2_X1 U11765 ( .A1(n18432), .A2(n18426), .ZN(n15716) );
  NOR2_X1 U11766 ( .A1(n17727), .A2(n10091), .ZN(n10090) );
  NOR2_X1 U11767 ( .A1(n17584), .A2(n15823), .ZN(n15836) );
  NAND2_X1 U11768 ( .A1(n9912), .A2(n17780), .ZN(n10081) );
  NAND2_X1 U11769 ( .A1(n18040), .A2(n10075), .ZN(n10074) );
  NAND2_X1 U11770 ( .A1(n9920), .A2(n10043), .ZN(n10042) );
  INV_X1 U11771 ( .A(n18052), .ZN(n10043) );
  INV_X1 U11772 ( .A(n15818), .ZN(n10076) );
  XNOR2_X1 U11773 ( .A(n10056), .B(n15898), .ZN(n15819) );
  XNOR2_X1 U11774 ( .A(n15802), .B(n17597), .ZN(n15814) );
  NAND2_X1 U11775 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  NOR2_X1 U11776 ( .A1(n15728), .A2(n15737), .ZN(n15726) );
  NOR2_X1 U11777 ( .A1(n15724), .A2(n15719), .ZN(n15869) );
  INV_X1 U11778 ( .A(n18880), .ZN(n10035) );
  NAND2_X1 U11779 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15704) );
  INV_X1 U11780 ( .A(n18865), .ZN(n16731) );
  OR3_X1 U11781 ( .A1(n15729), .A2(n15879), .A3(n15735), .ZN(n15888) );
  INV_X1 U11782 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17262) );
  AOI21_X1 U11783 ( .B1(n19053), .B2(n10016), .A(n9896), .ZN(n18900) );
  NAND2_X1 U11784 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  OR3_X1 U11785 ( .A1(n21108), .A2(n20380), .A3(n13393), .ZN(n20277) );
  NAND2_X1 U11786 ( .A1(n20277), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13404) );
  AND2_X1 U11787 ( .A1(n12239), .A2(n13400), .ZN(n13622) );
  AND2_X1 U11788 ( .A1(n21028), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14378) );
  NAND2_X1 U11789 ( .A1(n14377), .A2(n10320), .ZN(n10319) );
  INV_X1 U11790 ( .A(n10320), .ZN(n10318) );
  NAND2_X1 U11791 ( .A1(n11983), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12034) );
  AND2_X1 U11792 ( .A1(n11706), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11707) );
  AND2_X2 U11793 ( .A1(n13731), .A2(n13730), .ZN(n13979) );
  NAND2_X1 U11794 ( .A1(n13903), .A2(n13902), .ZN(n10395) );
  AND2_X1 U11795 ( .A1(n11562), .A2(n11585), .ZN(n10403) );
  NAND2_X1 U11796 ( .A1(n10063), .A2(n9938), .ZN(n14690) );
  NAND2_X1 U11797 ( .A1(n14714), .A2(n9931), .ZN(n10063) );
  AOI21_X1 U11798 ( .B1(n14699), .B2(n14722), .A(n14888), .ZN(n14711) );
  AOI21_X1 U11799 ( .B1(n10394), .B2(n10392), .A(n9910), .ZN(n10391) );
  NAND2_X1 U11800 ( .A1(n10136), .A2(n16104), .ZN(n13903) );
  NAND2_X1 U11801 ( .A1(n10384), .A2(n13665), .ZN(n10123) );
  NAND2_X1 U11802 ( .A1(n13680), .A2(n13679), .ZN(n16114) );
  AND2_X1 U11803 ( .A1(n12939), .A2(n13627), .ZN(n12954) );
  INV_X1 U11804 ( .A(n11485), .ZN(n11486) );
  NAND2_X1 U11805 ( .A1(n10308), .A2(n10120), .ZN(n10119) );
  AND2_X1 U11806 ( .A1(n10122), .A2(n11391), .ZN(n10120) );
  INV_X1 U11807 ( .A(n10308), .ZN(n10118) );
  OR2_X1 U11808 ( .A1(n11384), .A2(n11214), .ZN(n11491) );
  NAND2_X1 U11809 ( .A1(n11303), .A2(n11302), .ZN(n12872) );
  OR2_X1 U11810 ( .A1(n13316), .A2(n20513), .ZN(n20742) );
  AND4_X1 U11811 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11326) );
  NOR2_X1 U11812 ( .A1(n11314), .A2(n11313), .ZN(n11325) );
  AND4_X1 U11813 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11348) );
  AND4_X1 U11814 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11349) );
  INV_X1 U11815 ( .A(n11414), .ZN(n11415) );
  NOR2_X1 U11816 ( .A1(n20594), .A2(n20593), .ZN(n20940) );
  INV_X1 U11817 ( .A(n20742), .ZN(n20887) );
  NAND2_X1 U11818 ( .A1(n13316), .A2(n20513), .ZN(n20933) );
  NOR2_X1 U11819 ( .A1(n14105), .A2(n10206), .ZN(n14109) );
  NAND2_X1 U11820 ( .A1(n10263), .A2(n10260), .ZN(n10259) );
  NAND2_X1 U11821 ( .A1(n10406), .A2(n10263), .ZN(n10258) );
  INV_X1 U11822 ( .A(n15043), .ZN(n10260) );
  NAND2_X1 U11823 ( .A1(n10283), .A2(n10282), .ZN(n10281) );
  INV_X1 U11824 ( .A(n10284), .ZN(n10282) );
  NAND2_X1 U11825 ( .A1(n13040), .A2(n10713), .ZN(n13009) );
  INV_X1 U11826 ( .A(n15160), .ZN(n10240) );
  OR2_X1 U11827 ( .A1(n10238), .A2(n14018), .ZN(n10237) );
  AND2_X1 U11828 ( .A1(n13968), .A2(n13967), .ZN(n15545) );
  AND2_X1 U11829 ( .A1(n12523), .A2(n10233), .ZN(n10232) );
  NOR2_X1 U11830 ( .A1(n10234), .A2(n12529), .ZN(n10233) );
  INV_X1 U11831 ( .A(n13591), .ZN(n10234) );
  AOI21_X1 U11832 ( .B1(n10372), .B2(n10373), .A(n10371), .ZN(n10368) );
  NAND2_X1 U11833 ( .A1(n14392), .A2(n15381), .ZN(n10373) );
  NAND2_X1 U11834 ( .A1(n14250), .A2(n9974), .ZN(n10369) );
  NAND2_X1 U11835 ( .A1(n15254), .A2(n10374), .ZN(n15223) );
  INV_X1 U11836 ( .A(n10371), .ZN(n14241) );
  NAND2_X1 U11837 ( .A1(n10147), .A2(n10148), .ZN(n15266) );
  NAND2_X1 U11838 ( .A1(n10349), .A2(n10347), .ZN(n10147) );
  NAND2_X1 U11839 ( .A1(n15274), .A2(n15278), .ZN(n10148) );
  AOI21_X1 U11840 ( .B1(n10351), .B2(n10348), .A(n15272), .ZN(n10347) );
  AND2_X1 U11841 ( .A1(n15320), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15452) );
  AND2_X1 U11842 ( .A1(n15637), .A2(n10377), .ZN(n15320) );
  AND2_X1 U11843 ( .A1(n9872), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U11844 ( .A1(n15637), .A2(n9872), .ZN(n15324) );
  NAND2_X1 U11845 ( .A1(n15637), .A2(n14275), .ZN(n15343) );
  NOR2_X1 U11846 ( .A1(n9927), .A2(n10145), .ZN(n10144) );
  INV_X1 U11847 ( .A(n14102), .ZN(n10145) );
  OR2_X2 U11848 ( .A1(n16467), .A2(n10242), .ZN(n15607) );
  OR2_X1 U11849 ( .A1(n10243), .A2(n10246), .ZN(n10242) );
  INV_X1 U11850 ( .A(n15606), .ZN(n10246) );
  OR2_X1 U11851 ( .A1(n16394), .A2(n16397), .ZN(n15597) );
  OR2_X1 U11852 ( .A1(n13917), .A2(n14110), .ZN(n14220) );
  NAND2_X1 U11853 ( .A1(n13916), .A2(n9906), .ZN(n10185) );
  INV_X1 U11854 ( .A(n14218), .ZN(n10182) );
  NAND2_X1 U11855 ( .A1(n13875), .A2(n13874), .ZN(n16445) );
  NAND2_X1 U11856 ( .A1(n13548), .A2(n13547), .ZN(n13577) );
  INV_X1 U11857 ( .A(n13549), .ZN(n13548) );
  AOI21_X1 U11858 ( .B1(n13479), .B2(n10699), .A(n10698), .ZN(n13356) );
  NAND2_X1 U11859 ( .A1(n13356), .A2(n13357), .ZN(n13359) );
  AOI21_X2 U11860 ( .B1(n15656), .B2(n13453), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19975) );
  AND2_X1 U11861 ( .A1(n20174), .A2(n20184), .ZN(n20023) );
  NAND2_X1 U11862 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19975), .ZN(n19564) );
  INV_X1 U11863 ( .A(n19975), .ZN(n20019) );
  OR2_X1 U11864 ( .A1(n17118), .A2(n15704), .ZN(n9885) );
  NAND2_X1 U11865 ( .A1(n17602), .A2(n10194), .ZN(n17571) );
  AND2_X1 U11866 ( .A1(n17461), .A2(n9970), .ZN(n10194) );
  NAND2_X1 U11867 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10049) );
  NOR2_X1 U11868 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  OR2_X2 U11869 ( .A1(n13111), .A2(n15704), .ZN(n17396) );
  INV_X1 U11870 ( .A(n15775), .ZN(n10292) );
  INV_X1 U11871 ( .A(n15773), .ZN(n10293) );
  NAND2_X1 U11872 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10298) );
  NAND2_X1 U11873 ( .A1(n9965), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10296) );
  NAND3_X1 U11874 ( .A1(n15774), .A2(n15771), .A3(n10299), .ZN(n10288) );
  AOI21_X1 U11875 ( .B1(n15736), .B2(n17647), .A(n19082), .ZN(n17610) );
  NAND2_X1 U11876 ( .A1(n10168), .A2(n10167), .ZN(n10166) );
  NOR2_X1 U11877 ( .A1(n17068), .A2(n18437), .ZN(n10168) );
  INV_X1 U11878 ( .A(n15731), .ZN(n10167) );
  INV_X1 U11879 ( .A(n17836), .ZN(n10099) );
  INV_X1 U11880 ( .A(n17926), .ZN(n17875) );
  NOR2_X1 U11881 ( .A1(n15985), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10031) );
  INV_X1 U11882 ( .A(n10081), .ZN(n17770) );
  NAND3_X1 U11883 ( .A1(n15857), .A2(n15856), .A3(n9937), .ZN(n17859) );
  NOR2_X1 U11884 ( .A1(n10045), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17906) );
  NOR2_X1 U11885 ( .A1(n17966), .A2(n9969), .ZN(n10047) );
  OAI211_X1 U11886 ( .C1(n15787), .C2(n17144), .A(n15847), .B(n15846), .ZN(
        n16619) );
  NAND2_X1 U11887 ( .A1(n10302), .A2(n9901), .ZN(n15854) );
  NAND2_X1 U11888 ( .A1(n15854), .A2(n17951), .ZN(n10083) );
  NAND2_X1 U11889 ( .A1(n15853), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17902) );
  INV_X1 U11890 ( .A(n13199), .ZN(n18869) );
  NAND2_X1 U11891 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U11892 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13210) );
  AOI211_X1 U11893 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n13208), .B(n13207), .ZN(n13209) );
  INV_X1 U11894 ( .A(n18920), .ZN(n19078) );
  INV_X1 U11895 ( .A(n12217), .ZN(n13400) );
  NAND2_X1 U11896 ( .A1(n12867), .A2(n12701), .ZN(n21108) );
  INV_X1 U11897 ( .A(n20297), .ZN(n20315) );
  NAND2_X1 U11898 ( .A1(n12241), .A2(n13627), .ZN(n14600) );
  NAND2_X1 U11899 ( .A1(n12914), .A2(n12240), .ZN(n12241) );
  INV_X1 U11900 ( .A(n14600), .ZN(n14612) );
  INV_X1 U11901 ( .A(n14647), .ZN(n14383) );
  INV_X1 U11902 ( .A(n16219), .ZN(n16134) );
  AND2_X1 U11903 ( .A1(n14887), .A2(n14363), .ZN(n14873) );
  INV_X1 U11904 ( .A(n16211), .ZN(n20404) );
  NAND2_X1 U11905 ( .A1(n11417), .A2(n20890), .ZN(n20932) );
  CLKBUF_X1 U11906 ( .A(n12871), .Z(n20845) );
  OR2_X1 U11907 ( .A1(n20555), .A2(n20813), .ZN(n20596) );
  NOR2_X1 U11908 ( .A1(n12367), .A2(n12373), .ZN(n12638) );
  AND2_X1 U11909 ( .A1(n19481), .A2(n12714), .ZN(n19290) );
  XNOR2_X1 U11910 ( .A(n14234), .B(n14233), .ZN(n16263) );
  NAND2_X1 U11911 ( .A1(n10775), .A2(n10774), .ZN(n13653) );
  INV_X1 U11912 ( .A(n20184), .ZN(n19667) );
  NOR2_X1 U11913 ( .A1(n10274), .A2(n10273), .ZN(n10272) );
  INV_X1 U11914 ( .A(n15123), .ZN(n10273) );
  INV_X1 U11915 ( .A(n15122), .ZN(n10274) );
  NAND2_X1 U11916 ( .A1(n10268), .A2(n10270), .ZN(n10266) );
  NOR2_X1 U11917 ( .A1(n9997), .A2(n11046), .ZN(n9996) );
  INV_X1 U11918 ( .A(n15020), .ZN(n9997) );
  AND2_X1 U11919 ( .A1(n13948), .A2(n16551), .ZN(n19391) );
  AND2_X1 U11920 ( .A1(n19391), .A2(n13949), .ZN(n19429) );
  AND2_X1 U11921 ( .A1(n19514), .A2(n12721), .ZN(n16442) );
  AOI21_X1 U11922 ( .B1(n19361), .B2(n16485), .A(n14402), .ZN(n14403) );
  NAND2_X1 U11923 ( .A1(n16263), .A2(n16492), .ZN(n10251) );
  NAND2_X1 U11924 ( .A1(n10358), .A2(n15216), .ZN(n14216) );
  AOI211_X1 U11925 ( .C1(n15371), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15366), .B(n9892), .ZN(n10248) );
  INV_X1 U11926 ( .A(n15120), .ZN(n10249) );
  NAND2_X1 U11927 ( .A1(n10361), .A2(n10359), .ZN(n15218) );
  INV_X1 U11928 ( .A(n15517), .ZN(n15620) );
  OR2_X1 U11929 ( .A1(n15527), .A2(n16477), .ZN(n10011) );
  NOR2_X1 U11930 ( .A1(n9899), .A2(n10008), .ZN(n10007) );
  OAI211_X1 U11931 ( .C1(n19184), .C2(n16469), .A(n10010), .B(n10009), .ZN(
        n10008) );
  INV_X1 U11932 ( .A(n15522), .ZN(n10009) );
  AND2_X1 U11933 ( .A1(n12627), .A2(n12620), .ZN(n16485) );
  AND2_X1 U11934 ( .A1(n12627), .A2(n20203), .ZN(n16493) );
  NAND2_X1 U11935 ( .A1(n10706), .A2(n10705), .ZN(n15655) );
  OR2_X1 U11936 ( .A1(n19350), .A2(n12716), .ZN(n10706) );
  NOR2_X1 U11937 ( .A1(n16783), .A2(n9840), .ZN(n16775) );
  INV_X1 U11938 ( .A(n16776), .ZN(n10098) );
  NAND2_X1 U11939 ( .A1(n17460), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17603) );
  OR2_X1 U11940 ( .A1(n16625), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10306) );
  INV_X1 U11941 ( .A(n16601), .ZN(n10307) );
  NAND2_X1 U11942 ( .A1(n17730), .A2(n17729), .ZN(n10086) );
  NAND2_X1 U11943 ( .A1(n17794), .A2(n17725), .ZN(n10085) );
  OR2_X1 U11944 ( .A1(n17723), .A2(n17722), .ZN(n10089) );
  NOR2_X1 U11945 ( .A1(n18140), .A2(n17882), .ZN(n17794) );
  NAND2_X1 U11946 ( .A1(n10156), .A2(n10151), .ZN(n10150) );
  AOI21_X1 U11947 ( .B1(n17813), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n10152), .ZN(n10151) );
  NAND2_X1 U11948 ( .A1(n17819), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10156) );
  NAND2_X1 U11949 ( .A1(n10155), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U11950 ( .A1(n18190), .A2(n17974), .ZN(n17882) );
  INV_X1 U11951 ( .A(n17911), .ZN(n17992) );
  XNOR2_X1 U11952 ( .A(n15868), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16593) );
  NAND2_X1 U11953 ( .A1(n17902), .A2(n15854), .ZN(n18312) );
  OAI21_X1 U11954 ( .B1(n10023), .B2(n10022), .A(n10020), .ZN(n18919) );
  INV_X1 U11955 ( .A(n18910), .ZN(n10022) );
  AOI21_X1 U11956 ( .B1(n18907), .B2(n18908), .A(n10021), .ZN(n10020) );
  INV_X1 U11957 ( .A(n18909), .ZN(n10023) );
  NOR2_X1 U11958 ( .A1(n19028), .A2(n18924), .ZN(n18927) );
  INV_X1 U11959 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13851) );
  INV_X1 U11960 ( .A(n12733), .ZN(n10311) );
  AND2_X1 U11961 ( .A1(n12195), .A2(n12194), .ZN(n12202) );
  AOI22_X1 U11962 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10542) );
  INV_X1 U11963 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13498) );
  OR2_X1 U11964 ( .A1(n11036), .A2(n13487), .ZN(n10455) );
  OR2_X1 U11965 ( .A1(n11037), .A2(n13504), .ZN(n10457) );
  INV_X1 U11966 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13840) );
  INV_X1 U11967 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13838) );
  INV_X1 U11968 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13831) );
  INV_X1 U11969 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13844) );
  INV_X1 U11970 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13849) );
  INV_X1 U11971 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13837) );
  OAI21_X1 U11972 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13184), .A(
        n13186), .ZN(n13187) );
  OR2_X1 U11973 ( .A1(n16081), .A2(n14329), .ZN(n10400) );
  INV_X1 U11974 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12066) );
  INV_X1 U11975 ( .A(n11360), .ZN(n12736) );
  INV_X1 U11976 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U11977 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11255) );
  BUF_X1 U11978 ( .A(n11319), .Z(n11729) );
  NAND2_X1 U11979 ( .A1(n13299), .A2(n11214), .ZN(n11938) );
  NAND2_X1 U11980 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  OR3_X1 U11981 ( .A1(n12229), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20414), .ZN(n12196) );
  AOI21_X1 U11982 ( .B1(n12583), .B2(n11071), .A(n11070), .ZN(n11093) );
  INV_X1 U11983 ( .A(n13824), .ZN(n9990) );
  OR2_X1 U11984 ( .A1(n10541), .A2(n10506), .ZN(n10510) );
  AOI22_X1 U11985 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U11986 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10889), .ZN(n11055) );
  CLKBUF_X1 U11987 ( .A(n10498), .Z(n10900) );
  AOI22_X1 U11988 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11033) );
  INV_X1 U11989 ( .A(n15583), .ZN(n10143) );
  NOR2_X1 U11990 ( .A1(n12569), .A2(n12402), .ZN(n10005) );
  NOR2_X1 U11991 ( .A1(n10620), .A2(n20217), .ZN(n10621) );
  OR2_X1 U11992 ( .A1(n11036), .A2(n13498), .ZN(n10463) );
  OR2_X1 U11993 ( .A1(n11037), .A2(n13499), .ZN(n10465) );
  NAND2_X1 U11994 ( .A1(n13481), .A2(n13468), .ZN(n13497) );
  INV_X1 U11995 ( .A(n13476), .ZN(n13482) );
  OR2_X1 U11996 ( .A1(n10498), .A2(n10443), .ZN(n10448) );
  OR2_X1 U11997 ( .A1(n10498), .A2(n10430), .ZN(n10436) );
  OR2_X1 U11998 ( .A1(n10541), .A2(n10988), .ZN(n10474) );
  OR2_X1 U11999 ( .A1(n10541), .A2(n10997), .ZN(n10485) );
  OR2_X1 U12000 ( .A1(n10541), .A2(n13840), .ZN(n10532) );
  OR2_X1 U12001 ( .A1(n11037), .A2(n13838), .ZN(n10535) );
  OR2_X1 U12002 ( .A1(n11036), .A2(n13831), .ZN(n10533) );
  OR2_X1 U12003 ( .A1(n10541), .A2(n13844), .ZN(n10523) );
  OR2_X1 U12004 ( .A1(n11036), .A2(n13849), .ZN(n10524) );
  OR2_X1 U12005 ( .A1(n11037), .A2(n13837), .ZN(n10526) );
  INV_X1 U12006 ( .A(n19057), .ZN(n10018) );
  NOR2_X1 U12007 ( .A1(n18898), .A2(n18897), .ZN(n10017) );
  INV_X1 U12008 ( .A(n12196), .ZN(n12646) );
  NOR2_X1 U12009 ( .A1(n14430), .A2(n10321), .ZN(n10320) );
  OR2_X1 U12010 ( .A1(n14583), .A2(n14586), .ZN(n11882) );
  AND2_X1 U12011 ( .A1(n11804), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11824) );
  NOR2_X1 U12012 ( .A1(n11803), .A2(n10316), .ZN(n10314) );
  AND2_X1 U12013 ( .A1(n11627), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11639) );
  AND2_X1 U12014 ( .A1(n11549), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11627) );
  AND2_X1 U12015 ( .A1(n11547), .A2(n11635), .ZN(n13671) );
  AND2_X1 U12016 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11548), .ZN(
        n11587) );
  NAND2_X1 U12017 ( .A1(n10331), .A2(n14442), .ZN(n10330) );
  INV_X1 U12018 ( .A(n14473), .ZN(n10331) );
  NOR2_X1 U12019 ( .A1(n14596), .A2(n10338), .ZN(n10337) );
  NAND2_X1 U12020 ( .A1(n10065), .A2(n11636), .ZN(n13769) );
  INV_X1 U12021 ( .A(n11635), .ZN(n10065) );
  INV_X1 U12022 ( .A(n16104), .ZN(n10135) );
  INV_X1 U12023 ( .A(n13902), .ZN(n10392) );
  OR2_X1 U12024 ( .A1(n11524), .A2(n11523), .ZN(n13672) );
  NAND2_X1 U12025 ( .A1(n12327), .A2(n13619), .ZN(n12315) );
  NAND2_X1 U12026 ( .A1(n12985), .A2(n12984), .ZN(n13326) );
  AND4_X1 U12027 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(
        n11234) );
  AND2_X1 U12028 ( .A1(n20423), .A2(n20440), .ZN(n12254) );
  OR2_X1 U12029 ( .A1(n11471), .A2(n11470), .ZN(n12964) );
  OR2_X1 U12030 ( .A1(n11433), .A2(n11432), .ZN(n12963) );
  INV_X1 U12031 ( .A(n11492), .ZN(n13767) );
  NAND2_X1 U12032 ( .A1(n20423), .A2(n10379), .ZN(n12226) );
  NOR2_X1 U12033 ( .A1(n11354), .A2(n10062), .ZN(n10379) );
  OR2_X1 U12034 ( .A1(n20423), .A2(n21026), .ZN(n11493) );
  NAND2_X1 U12035 ( .A1(n11354), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11492) );
  NAND3_X1 U12036 ( .A1(n10060), .A2(n10059), .A3(n11368), .ZN(n11438) );
  NAND2_X1 U12037 ( .A1(n13299), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11319) );
  NOR2_X1 U12038 ( .A1(n10313), .A2(n12737), .ZN(n12904) );
  NAND2_X1 U12039 ( .A1(n13632), .A2(n11352), .ZN(n10313) );
  AND2_X1 U12040 ( .A1(n12238), .A2(n12877), .ZN(n12882) );
  INV_X1 U12041 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11209) );
  INV_X1 U12042 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11208) );
  AND2_X1 U12043 ( .A1(n10113), .A2(n10111), .ZN(n10117) );
  NOR2_X1 U12044 ( .A1(n12226), .A2(n13756), .ZN(n12235) );
  NAND2_X1 U12045 ( .A1(n11493), .A2(n11492), .ZN(n12232) );
  OR2_X1 U12046 ( .A1(n12229), .A2(n12228), .ZN(n12231) );
  OR2_X1 U12047 ( .A1(n12388), .A2(n12387), .ZN(n12514) );
  NAND2_X1 U12048 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20199), .ZN(
        n11075) );
  NAND2_X1 U12049 ( .A1(n10212), .A2(n9953), .ZN(n14189) );
  NAND2_X1 U12050 ( .A1(n10212), .A2(n10210), .ZN(n14187) );
  INV_X1 U12051 ( .A(n14182), .ZN(n10209) );
  NAND2_X1 U12052 ( .A1(n14141), .A2(n14129), .ZN(n14132) );
  NAND2_X1 U12053 ( .A1(n10215), .A2(n10214), .ZN(n12829) );
  NAND2_X1 U12054 ( .A1(n19547), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12055 ( .A1(n12584), .A2(n14208), .ZN(n10215) );
  NOR2_X1 U12056 ( .A1(n10505), .A2(n10504), .ZN(n10566) );
  OR2_X1 U12057 ( .A1(n10541), .A2(n10492), .ZN(n10496) );
  NAND2_X1 U12058 ( .A1(n10922), .A2(n10279), .ZN(n10278) );
  INV_X1 U12059 ( .A(n15167), .ZN(n10241) );
  AND2_X1 U12060 ( .A1(n10863), .A2(n15082), .ZN(n15075) );
  OR2_X1 U12061 ( .A1(n10634), .A2(n12614), .ZN(n10635) );
  OR2_X1 U12062 ( .A1(n12426), .A2(n12425), .ZN(n13814) );
  NOR2_X1 U12063 ( .A1(n16345), .A2(n10228), .ZN(n10227) );
  AND2_X1 U12064 ( .A1(n9934), .A2(n15078), .ZN(n10257) );
  NOR2_X1 U12065 ( .A1(n16374), .A2(n10225), .ZN(n10224) );
  INV_X1 U12066 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U12067 ( .A1(n19252), .A2(n10222), .ZN(n10221) );
  INV_X1 U12068 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12069 ( .A1(n15381), .A2(n14392), .ZN(n10376) );
  NOR2_X1 U12070 ( .A1(n10188), .A2(n15401), .ZN(n10187) );
  INV_X1 U12071 ( .A(n10189), .ZN(n10188) );
  AND2_X1 U12072 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10202) );
  NOR2_X1 U12073 ( .A1(n15278), .A2(n15437), .ZN(n10189) );
  INV_X1 U12074 ( .A(n15631), .ZN(n10355) );
  INV_X1 U12075 ( .A(n10356), .ZN(n10354) );
  OR2_X1 U12076 ( .A1(n15639), .A2(n10245), .ZN(n10244) );
  INV_X1 U12077 ( .A(n15623), .ZN(n10245) );
  NAND2_X1 U12078 ( .A1(n10355), .A2(n10356), .ZN(n16396) );
  AND2_X1 U12079 ( .A1(n9852), .A2(n13375), .ZN(n10256) );
  OAI21_X1 U12080 ( .B1(n13868), .B2(n14183), .A(n19286), .ZN(n13923) );
  NAND2_X1 U12081 ( .A1(n10341), .A2(n19296), .ZN(n13828) );
  INV_X1 U12082 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U12083 ( .A1(n10014), .A2(n10606), .ZN(n10607) );
  NAND2_X1 U12084 ( .A1(n10633), .A2(n12564), .ZN(n12609) );
  NAND2_X1 U12085 ( .A1(n19509), .A2(n10699), .ZN(n10001) );
  NAND3_X1 U12086 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20169), .A3(n19975), 
        .ZN(n13462) );
  NOR4_X1 U12087 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13107), .A4(n19037), .ZN(
        n13132) );
  NAND2_X1 U12088 ( .A1(n9965), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10055) );
  NAND2_X1 U12089 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10053) );
  NAND2_X1 U12090 ( .A1(n15837), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10054) );
  NOR2_X1 U12091 ( .A1(n10408), .A2(n17362), .ZN(n10051) );
  NAND2_X1 U12092 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10299) );
  INV_X1 U12093 ( .A(n15760), .ZN(n15764) );
  AND2_X1 U12094 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10028) );
  NAND2_X1 U12095 ( .A1(n17747), .A2(n9866), .ZN(n16596) );
  AND2_X1 U12096 ( .A1(n10102), .A2(n10101), .ZN(n10100) );
  INV_X1 U12097 ( .A(n17876), .ZN(n10101) );
  INV_X1 U12098 ( .A(n17799), .ZN(n15861) );
  AND2_X1 U12099 ( .A1(n15862), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10080) );
  NAND2_X1 U12100 ( .A1(n17902), .A2(n10083), .ZN(n10084) );
  INV_X1 U12101 ( .A(n18017), .ZN(n10301) );
  NAND2_X1 U12102 ( .A1(n10042), .A2(n9904), .ZN(n10038) );
  NAND2_X1 U12103 ( .A1(n10037), .A2(n15820), .ZN(n10036) );
  INV_X1 U12104 ( .A(n10074), .ZN(n10037) );
  OAI21_X1 U12105 ( .B1(n13196), .B2(n13195), .A(n15712), .ZN(n15874) );
  NOR2_X1 U12106 ( .A1(n15738), .A2(n15737), .ZN(n15885) );
  NOR2_X1 U12107 ( .A1(n13140), .A2(n10024), .ZN(n15734) );
  NAND2_X1 U12108 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U12109 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10025) );
  AOI211_X1 U12110 ( .C1(n13275), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n13152), .B(n13151), .ZN(n15715) );
  NOR2_X2 U12111 ( .A1(n14488), .A2(n10328), .ZN(n14431) );
  NAND2_X1 U12112 ( .A1(n14451), .A2(n10329), .ZN(n10328) );
  NOR2_X1 U12113 ( .A1(n10330), .A2(n14432), .ZN(n10329) );
  NAND2_X1 U12114 ( .A1(n14607), .A2(n14606), .ZN(n14609) );
  AND2_X1 U12115 ( .A1(n11927), .A2(n11926), .ZN(n14575) );
  NOR2_X1 U12116 ( .A1(n14383), .A2(n13629), .ZN(n14382) );
  AND2_X1 U12117 ( .A1(n14681), .A2(n13391), .ZN(n12181) );
  AND2_X1 U12118 ( .A1(n14698), .A2(n13391), .ZN(n12116) );
  AND2_X1 U12119 ( .A1(n12088), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12089) );
  NAND2_X1 U12120 ( .A1(n12089), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12119) );
  NOR2_X1 U12121 ( .A1(n14465), .A2(n14455), .ZN(n14454) );
  AND2_X1 U12122 ( .A1(n12035), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12036) );
  AND2_X1 U12123 ( .A1(n12041), .A2(n12040), .ZN(n14480) );
  OR2_X1 U12124 ( .A1(n14738), .A2(n12178), .ZN(n12040) );
  AND2_X1 U12125 ( .A1(n14747), .A2(n13391), .ZN(n12008) );
  OR2_X1 U12126 ( .A1(n14755), .A2(n12178), .ZN(n11986) );
  AND2_X1 U12127 ( .A1(n14576), .A2(n10324), .ZN(n14508) );
  NAND2_X1 U12128 ( .A1(n14576), .A2(n10326), .ZN(n14519) );
  NAND2_X1 U12129 ( .A1(n14576), .A2(n14575), .ZN(n14574) );
  AND2_X1 U12130 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11922), .ZN(
        n11923) );
  NAND2_X1 U12131 ( .A1(n11923), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11982) );
  AND2_X1 U12132 ( .A1(n11878), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11879) );
  NAND2_X1 U12133 ( .A1(n11879), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11921) );
  CLKBUF_X1 U12134 ( .A(n14532), .Z(n14584) );
  NAND2_X1 U12135 ( .A1(n10067), .A2(n10397), .ZN(n14784) );
  NAND2_X1 U12136 ( .A1(n10396), .A2(n9893), .ZN(n10067) );
  CLKBUF_X1 U12137 ( .A(n14542), .Z(n14593) );
  NAND2_X1 U12138 ( .A1(n11824), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11841) );
  AND2_X1 U12139 ( .A1(n11783), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11804) );
  INV_X1 U12140 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11725) );
  AND2_X1 U12141 ( .A1(n11796), .A2(n11724), .ZN(n14035) );
  INV_X1 U12142 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11701) );
  AOI21_X1 U12143 ( .B1(n13908), .B2(n12145), .A(n11687), .ZN(n13711) );
  NOR2_X2 U12144 ( .A1(n13712), .A2(n13711), .ZN(n13731) );
  AND2_X1 U12145 ( .A1(n11639), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11669) );
  AOI21_X1 U12146 ( .B1(n13683), .B2(n11796), .A(n11634), .ZN(n13606) );
  AOI21_X1 U12147 ( .B1(n13669), .B2(n11796), .A(n11609), .ZN(n13383) );
  NAND2_X1 U12148 ( .A1(n12974), .A2(n11585), .ZN(n13103) );
  CLKBUF_X1 U12149 ( .A(n13101), .Z(n13384) );
  INV_X1 U12150 ( .A(n12973), .ZN(n11584) );
  NAND2_X1 U12151 ( .A1(n12970), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12985) );
  NOR3_X1 U12152 ( .A1(n14488), .A2(n12317), .A3(n14473), .ZN(n14453) );
  NAND2_X1 U12153 ( .A1(n14711), .A2(n14733), .ZN(n10140) );
  NOR2_X1 U12154 ( .A1(n14488), .A2(n14473), .ZN(n14475) );
  INV_X1 U12155 ( .A(n10124), .ZN(n10127) );
  NAND2_X1 U12156 ( .A1(n10132), .A2(n10397), .ZN(n10131) );
  NOR2_X1 U12157 ( .A1(n14597), .A2(n10335), .ZN(n14587) );
  INV_X1 U12158 ( .A(n10337), .ZN(n10335) );
  NOR2_X1 U12159 ( .A1(n14597), .A2(n14596), .ZN(n14599) );
  NAND2_X1 U12160 ( .A1(n9893), .A2(n14327), .ZN(n14793) );
  OR2_X1 U12161 ( .A1(n14336), .A2(n16173), .ZN(n14803) );
  AND2_X1 U12162 ( .A1(n14336), .A2(n14818), .ZN(n14820) );
  OR2_X1 U12163 ( .A1(n10333), .A2(n14040), .ZN(n10332) );
  NOR2_X1 U12164 ( .A1(n13735), .A2(n13734), .ZN(n14014) );
  NAND2_X1 U12165 ( .A1(n10395), .A2(n10394), .ZN(n14832) );
  AOI21_X1 U12166 ( .B1(n13752), .B2(n10390), .A(n9909), .ZN(n10389) );
  INV_X1 U12167 ( .A(n13682), .ZN(n10390) );
  OR2_X1 U12168 ( .A1(n13387), .A2(n13386), .ZN(n13603) );
  NAND2_X1 U12169 ( .A1(n16242), .A2(n21026), .ZN(n12795) );
  OR2_X1 U12170 ( .A1(n20411), .A2(n20412), .ZN(n13696) );
  NAND2_X1 U12171 ( .A1(n13379), .A2(n13378), .ZN(n13387) );
  CLKBUF_X1 U12172 ( .A(n12252), .Z(n14341) );
  NAND2_X1 U12173 ( .A1(n14370), .A2(n21026), .ZN(n11575) );
  XNOR2_X1 U12174 ( .A(n10308), .B(n11391), .ZN(n12871) );
  XNOR2_X1 U12175 ( .A(n11586), .B(n13347), .ZN(n20419) );
  AND2_X2 U12176 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13291) );
  CLKBUF_X1 U12177 ( .A(n12887), .Z(n12888) );
  NAND2_X1 U12178 ( .A1(n10308), .A2(n11391), .ZN(n13309) );
  AND3_X1 U12179 ( .A1(n12923), .A2(n12922), .A3(n12921), .ZN(n15949) );
  INV_X1 U12180 ( .A(n11354), .ZN(n10380) );
  AOI21_X1 U12181 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20889), .A(n20593), 
        .ZN(n20974) );
  INV_X1 U12182 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20804) );
  AND2_X1 U12183 ( .A1(n13620), .A2(n12787), .ZN(n15965) );
  NOR2_X1 U12184 ( .A1(n12605), .A2(n12604), .ZN(n16533) );
  NAND2_X1 U12185 ( .A1(n12581), .A2(n12368), .ZN(n9986) );
  NAND2_X1 U12186 ( .A1(n11091), .A2(n12624), .ZN(n9984) );
  OAI21_X1 U12187 ( .B1(n12514), .B2(n12581), .A(n10216), .ZN(n12584) );
  NAND2_X1 U12188 ( .A1(n12581), .A2(n12389), .ZN(n10216) );
  NAND2_X1 U12189 ( .A1(n14198), .A2(n14242), .ZN(n14246) );
  NAND2_X1 U12190 ( .A1(n10205), .A2(n11122), .ZN(n10204) );
  INV_X1 U12191 ( .A(n10206), .ZN(n10205) );
  NAND2_X1 U12192 ( .A1(n14112), .A2(n14111), .ZN(n14124) );
  AND2_X1 U12193 ( .A1(n16529), .A2(n16551), .ZN(n12632) );
  NAND2_X1 U12194 ( .A1(n10285), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10284) );
  INV_X1 U12195 ( .A(n10717), .ZN(n10285) );
  NOR2_X1 U12196 ( .A1(n11069), .A2(n11050), .ZN(n10267) );
  INV_X1 U12197 ( .A(n11069), .ZN(n10270) );
  NAND2_X1 U12198 ( .A1(n15145), .A2(n14291), .ZN(n15130) );
  INV_X1 U12199 ( .A(n10406), .ZN(n10261) );
  NAND2_X1 U12200 ( .A1(n15176), .A2(n9950), .ZN(n15169) );
  NAND2_X1 U12201 ( .A1(n15176), .A2(n9949), .ZN(n15441) );
  AND2_X1 U12202 ( .A1(n15176), .A2(n15177), .ZN(n15439) );
  AND2_X1 U12203 ( .A1(n14279), .A2(n14278), .ZN(n15186) );
  NAND2_X1 U12204 ( .A1(n10236), .A2(n15208), .ZN(n10235) );
  INV_X1 U12205 ( .A(n10237), .ZN(n10236) );
  NAND2_X1 U12206 ( .A1(n15083), .A2(n15082), .ZN(n13997) );
  INV_X1 U12207 ( .A(n10635), .ZN(n13945) );
  AND2_X1 U12208 ( .A1(n19554), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13364) );
  AND2_X1 U12209 ( .A1(n19391), .A2(n13970), .ZN(n19368) );
  INV_X1 U12210 ( .A(n12357), .ZN(n13971) );
  AND2_X1 U12211 ( .A1(n15228), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15229) );
  NOR2_X1 U12212 ( .A1(n15236), .A2(n14253), .ZN(n15228) );
  NAND2_X1 U12213 ( .A1(n15248), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15236) );
  AND2_X1 U12214 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n15267), .ZN(
        n15248) );
  AND2_X1 U12215 ( .A1(n15935), .A2(n10226), .ZN(n15267) );
  AND2_X1 U12216 ( .A1(n9868), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U12217 ( .A1(n15935), .A2(n9868), .ZN(n15276) );
  NAND2_X1 U12218 ( .A1(n15935), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15934) );
  NOR2_X1 U12219 ( .A1(n19127), .A2(n15317), .ZN(n15935) );
  AND2_X1 U12220 ( .A1(n13992), .A2(n9934), .ZN(n15088) );
  NOR2_X1 U12221 ( .A1(n15332), .A2(n15340), .ZN(n15330) );
  NAND2_X1 U12222 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n15330), .ZN(
        n15317) );
  AND2_X1 U12223 ( .A1(n13992), .A2(n15099), .ZN(n15100) );
  AND2_X1 U12224 ( .A1(n15940), .A2(n10223), .ZN(n15349) );
  AND2_X1 U12225 ( .A1(n9867), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10223) );
  NAND2_X1 U12226 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n15349), .ZN(
        n15340) );
  NAND2_X1 U12227 ( .A1(n15940), .A2(n9867), .ZN(n15360) );
  NAND2_X1 U12228 ( .A1(n15940), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15939) );
  AND2_X1 U12229 ( .A1(n11168), .A2(n11167), .ZN(n13722) );
  NAND2_X1 U12230 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n15938), .ZN(
        n15937) );
  AND2_X1 U12231 ( .A1(n12364), .A2(n10220), .ZN(n15938) );
  AND2_X1 U12232 ( .A1(n9851), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10220) );
  NAND2_X1 U12233 ( .A1(n12364), .A2(n9851), .ZN(n12365) );
  NAND2_X1 U12234 ( .A1(n12364), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12363) );
  NAND3_X1 U12235 ( .A1(n10231), .A2(n10229), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12362) );
  NOR2_X1 U12236 ( .A1(n19295), .A2(n10230), .ZN(n10229) );
  NAND2_X1 U12237 ( .A1(n11140), .A2(n11139), .ZN(n13588) );
  AND2_X1 U12238 ( .A1(n11145), .A2(n11144), .ZN(n13587) );
  NOR2_X1 U12239 ( .A1(n12359), .A2(n14995), .ZN(n12361) );
  NAND2_X1 U12240 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U12241 ( .A1(n10667), .A2(n10666), .ZN(n10700) );
  AOI21_X1 U12242 ( .B1(n10665), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10664), 
        .ZN(n10666) );
  OAI22_X1 U12243 ( .A1(n10661), .A2(n10660), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14228), .ZN(n10667) );
  NOR2_X1 U12244 ( .A1(n10375), .A2(n15382), .ZN(n10374) );
  INV_X1 U12245 ( .A(n10376), .ZN(n10375) );
  NAND2_X1 U12246 ( .A1(n15246), .A2(n10362), .ZN(n10361) );
  NOR2_X1 U12247 ( .A1(n10367), .A2(n15224), .ZN(n10362) );
  INV_X1 U12248 ( .A(n10368), .ZN(n10367) );
  INV_X1 U12249 ( .A(n10364), .ZN(n10360) );
  AOI21_X1 U12250 ( .B1(n10366), .B2(n10368), .A(n10365), .ZN(n10364) );
  INV_X1 U12251 ( .A(n10369), .ZN(n10366) );
  NAND2_X1 U12252 ( .A1(n15454), .A2(n9971), .ZN(n15238) );
  INV_X1 U12253 ( .A(n14248), .ZN(n14247) );
  AND2_X1 U12254 ( .A1(n14200), .A2(n14199), .ZN(n15263) );
  NAND2_X1 U12255 ( .A1(n15454), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15284) );
  NAND2_X1 U12256 ( .A1(n15451), .A2(n9849), .ZN(n10346) );
  OR3_X1 U12257 ( .A1(n14176), .A2(n14110), .A3(n15479), .ZN(n15303) );
  NAND2_X1 U12258 ( .A1(n19177), .A2(n16492), .ZN(n10010) );
  NOR3_X1 U12259 ( .A1(n13721), .A2(n9956), .A3(n13722), .ZN(n14009) );
  AND2_X1 U12260 ( .A1(n12472), .A2(n12471), .ZN(n12544) );
  OR2_X1 U12261 ( .A1(n16467), .A2(n10244), .ZN(n15624) );
  AND2_X1 U12262 ( .A1(n14116), .A2(n15643), .ZN(n15632) );
  NAND2_X1 U12263 ( .A1(n14103), .A2(n14102), .ZN(n15631) );
  OR2_X1 U12264 ( .A1(n13917), .A2(n14222), .ZN(n14223) );
  NAND2_X1 U12265 ( .A1(n10185), .A2(n10183), .ZN(n10186) );
  NOR2_X1 U12266 ( .A1(n16467), .A2(n15639), .ZN(n15638) );
  NAND2_X1 U12267 ( .A1(n13368), .A2(n10256), .ZN(n13436) );
  AND2_X1 U12268 ( .A1(n13368), .A2(n9852), .ZN(n13374) );
  NAND2_X1 U12269 ( .A1(n13368), .A2(n13369), .ZN(n13367) );
  NAND2_X1 U12270 ( .A1(n16484), .A2(n12533), .ZN(n13893) );
  NAND2_X1 U12271 ( .A1(n10345), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10344) );
  INV_X1 U12272 ( .A(n19308), .ZN(n10345) );
  XNOR2_X1 U12273 ( .A(n13828), .B(n16497), .ZN(n16447) );
  NAND2_X1 U12274 ( .A1(n10177), .A2(n13513), .ZN(n13581) );
  NAND2_X1 U12275 ( .A1(n10178), .A2(n13544), .ZN(n13580) );
  OAI21_X1 U12276 ( .B1(n12473), .B2(n19341), .A(n12502), .ZN(n12621) );
  INV_X1 U12277 ( .A(n10699), .ZN(n12716) );
  INV_X1 U12278 ( .A(n9843), .ZN(n19315) );
  NAND2_X1 U12279 ( .A1(n12597), .A2(n11107), .ZN(n13028) );
  OR2_X1 U12280 ( .A1(n20222), .A2(n12589), .ZN(n11107) );
  AND3_X1 U12281 ( .A1(n14204), .A2(n10014), .A3(n12569), .ZN(n10603) );
  AOI21_X1 U12282 ( .B1(n14237), .B2(n20218), .A(n10217), .ZN(n15010) );
  AND2_X1 U12283 ( .A1(n14231), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10217) );
  XNOR2_X1 U12284 ( .A(n10712), .B(n10710), .ZN(n13038) );
  AND2_X1 U12285 ( .A1(n13359), .A2(n10709), .ZN(n13037) );
  NAND2_X1 U12286 ( .A1(n13038), .A2(n13037), .ZN(n13040) );
  INV_X1 U12287 ( .A(n19969), .ZN(n19835) );
  INV_X1 U12288 ( .A(n19936), .ZN(n19864) );
  INV_X1 U12289 ( .A(n19559), .ZN(n19560) );
  INV_X1 U12290 ( .A(n19558), .ZN(n19562) );
  OR2_X1 U12291 ( .A1(n19583), .A2(n19582), .ZN(n19969) );
  INV_X1 U12292 ( .A(n20023), .ZN(n19968) );
  OR2_X1 U12293 ( .A1(n20078), .A2(n20013), .ZN(n19106) );
  NOR3_X1 U12294 ( .A1(n9877), .A2(n16748), .A3(n18881), .ZN(n18866) );
  INV_X1 U12295 ( .A(n15736), .ZN(n16748) );
  NAND2_X1 U12296 ( .A1(n9840), .A2(n10095), .ZN(n10092) );
  AND2_X1 U12297 ( .A1(n10095), .A2(n17735), .ZN(n10094) );
  OR2_X1 U12298 ( .A1(n16816), .A2(n9840), .ZN(n10096) );
  NOR2_X1 U12299 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16985), .ZN(n16970) );
  INV_X1 U12300 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16981) );
  NOR2_X1 U12301 ( .A1(n18866), .A2(n17609), .ZN(n17067) );
  NOR2_X1 U12302 ( .A1(n17667), .A2(n10197), .ZN(n10196) );
  INV_X1 U12303 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17406) );
  NAND2_X1 U12304 ( .A1(n10287), .A2(n10286), .ZN(n17415) );
  NOR2_X1 U12305 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10286) );
  INV_X1 U12306 ( .A(n18879), .ZN(n10287) );
  OAI211_X1 U12307 ( .C1(n15787), .C2(n17343), .A(n15786), .B(n15785), .ZN(
        n15898) );
  NAND2_X1 U12308 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n15806) );
  INV_X1 U12309 ( .A(n17609), .ZN(n17648) );
  AND2_X1 U12310 ( .A1(n17747), .A2(n9870), .ZN(n16595) );
  NAND2_X1 U12311 ( .A1(n17747), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17726) );
  NOR2_X1 U12312 ( .A1(n17760), .A2(n17761), .ZN(n17747) );
  NOR2_X1 U12313 ( .A1(n17805), .A2(n17806), .ZN(n16760) );
  INV_X1 U12314 ( .A(n10154), .ZN(n10153) );
  NAND2_X1 U12315 ( .A1(n17929), .A2(n17804), .ZN(n10155) );
  NAND2_X1 U12316 ( .A1(n17927), .A2(n9853), .ZN(n17835) );
  NAND2_X1 U12317 ( .A1(n17927), .A2(n10102), .ZN(n17874) );
  NOR3_X2 U12318 ( .A1(n17981), .A2(n17940), .A3(n16981), .ZN(n17927) );
  NAND2_X1 U12319 ( .A1(n18015), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17981) );
  NOR2_X1 U12320 ( .A1(n18024), .A2(n17055), .ZN(n18015) );
  AND2_X1 U12321 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18045) );
  NOR2_X1 U12322 ( .A1(n19078), .A2(n19084), .ZN(n16557) );
  NOR2_X1 U12323 ( .A1(n15882), .A2(n15870), .ZN(n16620) );
  OAI21_X1 U12324 ( .B1(n10079), .B2(n17781), .A(n10078), .ZN(n10077) );
  NAND2_X1 U12325 ( .A1(n15864), .A2(n18119), .ZN(n10078) );
  NAND2_X1 U12326 ( .A1(n10081), .A2(n9869), .ZN(n10079) );
  NOR2_X1 U12327 ( .A1(n17745), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17744) );
  NOR2_X1 U12328 ( .A1(n18218), .A2(n15922), .ZN(n18131) );
  AND2_X1 U12329 ( .A1(n15889), .A2(n10174), .ZN(n10173) );
  INV_X1 U12330 ( .A(n10173), .ZN(n10172) );
  INV_X1 U12331 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10046) );
  INV_X1 U12332 ( .A(n10084), .ZN(n17952) );
  NOR2_X1 U12333 ( .A1(n15919), .A2(n17979), .ZN(n18273) );
  NAND2_X1 U12334 ( .A1(n18016), .A2(n15848), .ZN(n10069) );
  NAND2_X1 U12335 ( .A1(n10068), .A2(n9856), .ZN(n10070) );
  NAND2_X1 U12336 ( .A1(n15848), .A2(n15835), .ZN(n10071) );
  NAND2_X1 U12337 ( .A1(n10042), .A2(n10074), .ZN(n15821) );
  NOR2_X1 U12338 ( .A1(n18027), .A2(n18028), .ZN(n18026) );
  AOI211_X1 U12339 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n13173), .B(n13172), .ZN(n15872) );
  INV_X1 U12340 ( .A(n16620), .ZN(n18863) );
  NOR2_X1 U12341 ( .A1(n18892), .A2(n18893), .ZN(n18896) );
  NAND2_X1 U12342 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10035), .ZN(
        n17101) );
  AOI21_X1 U12343 ( .B1(n15740), .B2(n17610), .A(n15739), .ZN(n18901) );
  NOR3_X1 U12344 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19083), .ZN(n18713) );
  AOI211_X1 U12345 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n13161), .B(n13160), .ZN(n13162) );
  AOI211_X1 U12346 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n13181), .B(n13180), .ZN(n13182) );
  INV_X1 U12347 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18897) );
  INV_X1 U12348 ( .A(n18797), .ZN(n18741) );
  NAND2_X1 U12349 ( .A1(n13413), .A2(n13396), .ZN(n20318) );
  AND2_X1 U12350 ( .A1(n20277), .A2(n13405), .ZN(n20264) );
  AND2_X1 U12351 ( .A1(n20318), .A2(n20277), .ZN(n20279) );
  NAND2_X1 U12352 ( .A1(n13413), .A2(n13409), .ZN(n20297) );
  INV_X1 U12353 ( .A(n14386), .ZN(n14668) );
  AND2_X1 U12354 ( .A1(n14382), .A2(n20416), .ZN(n14669) );
  INV_X1 U12355 ( .A(n14800), .ZN(n14673) );
  INV_X1 U12356 ( .A(n14383), .ZN(n14674) );
  OR2_X1 U12357 ( .A1(n13626), .A2(n13625), .ZN(n13628) );
  NOR2_X2 U12358 ( .A1(n13630), .A2(n14382), .ZN(n14676) );
  INV_X1 U12359 ( .A(n14666), .ZN(n13630) );
  OAI22_X1 U12360 ( .A1(n12867), .A2(n15970), .B1(n12920), .B2(n20235), .ZN(
        n20328) );
  INV_X1 U12361 ( .A(n14320), .ZN(n20362) );
  OR2_X1 U12362 ( .A1(n20361), .A2(n12868), .ZN(n13043) );
  NAND2_X1 U12363 ( .A1(n10395), .A2(n13905), .ZN(n14322) );
  AND2_X1 U12364 ( .A1(n12801), .A2(n20842), .ZN(n14411) );
  INV_X1 U12365 ( .A(n14411), .ZN(n20417) );
  INV_X1 U12366 ( .A(n20370), .ZN(n20242) );
  AND2_X1 U12367 ( .A1(n14904), .A2(n14361), .ZN(n14887) );
  XNOR2_X1 U12368 ( .A(n10381), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14413) );
  NAND2_X1 U12369 ( .A1(n10383), .A2(n10382), .ZN(n10381) );
  NAND2_X1 U12370 ( .A1(n14690), .A2(n14339), .ZN(n10383) );
  NAND2_X1 U12371 ( .A1(n14679), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U12372 ( .A1(n16114), .A2(n13682), .ZN(n13753) );
  OR2_X1 U12373 ( .A1(n12795), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16210) );
  INV_X1 U12374 ( .A(n13680), .ZN(n16116) );
  NAND2_X1 U12375 ( .A1(n13665), .A2(n13664), .ZN(n20368) );
  OR2_X1 U12376 ( .A1(n14958), .A2(n14956), .ZN(n20396) );
  AND2_X1 U12377 ( .A1(n12954), .A2(n12943), .ZN(n20405) );
  INV_X1 U12378 ( .A(n13005), .ZN(n13006) );
  NAND2_X1 U12379 ( .A1(n12954), .A2(n12945), .ZN(n16211) );
  INV_X1 U12380 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20889) );
  INV_X1 U12381 ( .A(n11563), .ZN(n11565) );
  INV_X1 U12382 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20764) );
  OR2_X1 U12383 ( .A1(n11556), .A2(n11555), .ZN(n11557) );
  NAND2_X1 U12384 ( .A1(n10119), .A2(n9942), .ZN(n20710) );
  NAND2_X1 U12385 ( .A1(n10118), .A2(n20588), .ZN(n10116) );
  OAI21_X1 U12386 ( .B1(n13315), .B2(n16252), .A(n20593), .ZN(n20413) );
  NOR2_X1 U12387 ( .A1(n12872), .A2(n12808), .ZN(n14373) );
  INV_X2 U12388 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15948) );
  NAND2_X1 U12389 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13620), .ZN(n14986) );
  NOR2_X1 U12390 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16242) );
  OAI21_X1 U12391 ( .B1(n20612), .B2(n20595), .A(n20940), .ZN(n20614) );
  OR2_X1 U12392 ( .A1(n20686), .A2(n20933), .ZN(n20708) );
  INV_X1 U12393 ( .A(n20700), .ZN(n20732) );
  INV_X1 U12394 ( .A(n20798), .ZN(n20766) );
  NAND2_X1 U12395 ( .A1(n20815), .A2(n20887), .ZN(n20798) );
  INV_X1 U12396 ( .A(n20829), .ZN(n20834) );
  NAND2_X1 U12397 ( .A1(n20479), .A2(n10380), .ZN(n20867) );
  OR2_X1 U12398 ( .A1(n20934), .A2(n20838), .ZN(n20894) );
  OAI211_X1 U12399 ( .C1(n20957), .C2(n20941), .A(n20940), .B(n20939), .ZN(
        n20959) );
  INV_X1 U12400 ( .A(n20840), .ZN(n20969) );
  INV_X1 U12401 ( .A(n20855), .ZN(n20982) );
  INV_X1 U12402 ( .A(n20859), .ZN(n20987) );
  INV_X1 U12403 ( .A(n20863), .ZN(n20993) );
  INV_X1 U12404 ( .A(n20867), .ZN(n20999) );
  INV_X1 U12405 ( .A(n20871), .ZN(n21004) );
  INV_X1 U12406 ( .A(n20875), .ZN(n21010) );
  OR2_X1 U12407 ( .A1(n20934), .A2(n20933), .ZN(n21023) );
  INV_X1 U12408 ( .A(n20976), .ZN(n21019) );
  INV_X1 U12409 ( .A(n20880), .ZN(n21018) );
  AND2_X1 U12410 ( .A1(n21025), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15976) );
  INV_X2 U12411 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21028) );
  INV_X1 U12412 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21025) );
  INV_X1 U12413 ( .A(n19325), .ZN(n19343) );
  NOR2_X1 U12414 ( .A1(n14105), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14107) );
  OR2_X1 U12415 ( .A1(n20214), .A2(n12378), .ZN(n19342) );
  INV_X1 U12416 ( .A(n19342), .ZN(n19323) );
  INV_X1 U12417 ( .A(n19339), .ZN(n19303) );
  OR4_X1 U12418 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n20079), .ZN(n19339) );
  NOR2_X1 U12419 ( .A1(n9843), .A2(n19339), .ZN(n19335) );
  INV_X1 U12420 ( .A(n19324), .ZN(n19353) );
  AND2_X1 U12421 ( .A1(n9998), .A2(n15027), .ZN(n15021) );
  OR2_X1 U12422 ( .A1(n10884), .A2(n10883), .ZN(n13962) );
  AND2_X1 U12423 ( .A1(n13725), .A2(n13962), .ZN(n15083) );
  OR2_X1 U12424 ( .A1(n10753), .A2(n10752), .ZN(n13433) );
  OR2_X1 U12425 ( .A1(n10281), .A2(n13372), .ZN(n10280) );
  CLKBUF_X1 U12426 ( .A(n13432), .Z(n13613) );
  OR2_X1 U12427 ( .A1(n14093), .A2(n10281), .ZN(n13373) );
  XNOR2_X1 U12428 ( .A(n13009), .B(n13010), .ZN(n19583) );
  AND2_X1 U12429 ( .A1(n15104), .A2(n12569), .ZN(n15110) );
  INV_X1 U12430 ( .A(n10262), .ZN(n15042) );
  NOR2_X1 U12431 ( .A1(n9891), .A2(n10922), .ZN(n15056) );
  AND2_X1 U12432 ( .A1(n19368), .A2(n15125), .ZN(n19360) );
  NOR2_X1 U12433 ( .A1(n15565), .A2(n15545), .ZN(n13999) );
  INV_X1 U12434 ( .A(n19428), .ZN(n19365) );
  AND2_X1 U12435 ( .A1(n19391), .A2(n9898), .ZN(n19367) );
  NAND2_X1 U12436 ( .A1(n10275), .A2(n10715), .ZN(n14091) );
  AND2_X1 U12437 ( .A1(n19391), .A2(n19565), .ZN(n19428) );
  INV_X1 U12438 ( .A(n19391), .ZN(n19427) );
  NAND2_X1 U12439 ( .A1(n19476), .A2(n20211), .ZN(n19443) );
  INV_X2 U12440 ( .A(n19443), .ZN(n19473) );
  AND2_X1 U12441 ( .A1(n12638), .A2(n12551), .ZN(n19481) );
  XNOR2_X1 U12442 ( .A(n10219), .B(n10218), .ZN(n14237) );
  INV_X1 U12443 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12444 ( .A1(n15229), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10219) );
  INV_X1 U12445 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16374) );
  INV_X1 U12446 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19252) );
  INV_X1 U12447 ( .A(n16442), .ZN(n19503) );
  NAND2_X1 U12448 ( .A1(n19108), .A2(n12707), .ZN(n19514) );
  INV_X1 U12449 ( .A(n19514), .ZN(n19490) );
  INV_X1 U12450 ( .A(n19493), .ZN(n19504) );
  INV_X1 U12451 ( .A(n19510), .ZN(n16438) );
  NAND2_X1 U12452 ( .A1(n10363), .A2(n10368), .ZN(n15227) );
  OAI21_X1 U12453 ( .B1(n15451), .B2(n15448), .A(n15449), .ZN(n15285) );
  AOI21_X1 U12454 ( .B1(n14103), .B2(n10144), .A(n9887), .ZN(n15585) );
  NAND2_X1 U12455 ( .A1(n10185), .A2(n14217), .ZN(n16420) );
  NAND2_X1 U12456 ( .A1(n10343), .A2(n13577), .ZN(n13827) );
  INV_X1 U12457 ( .A(n16485), .ZN(n16469) );
  INV_X1 U12458 ( .A(n19582), .ZN(n20194) );
  INV_X1 U12459 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20190) );
  INV_X1 U12460 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20181) );
  NAND2_X1 U12461 ( .A1(n12837), .A2(n12523), .ZN(n13556) );
  NAND2_X1 U12462 ( .A1(n13028), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15656) );
  NAND2_X1 U12463 ( .A1(n13359), .A2(n13358), .ZN(n20184) );
  AND2_X1 U12464 ( .A1(n13040), .A2(n13039), .ZN(n20174) );
  OR2_X1 U12465 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NAND2_X1 U12466 ( .A1(n10620), .A2(n16528), .ZN(n15745) );
  OR2_X1 U12467 ( .A1(n19613), .A2(n20019), .ZN(n19631) );
  INV_X1 U12468 ( .A(n19608), .ZN(n19630) );
  INV_X1 U12469 ( .A(n19676), .ZN(n19694) );
  AND2_X1 U12470 ( .A1(n19763), .A2(n19944), .ZN(n19747) );
  INV_X1 U12471 ( .A(n19783), .ZN(n19772) );
  NAND2_X1 U12472 ( .A1(n19794), .A2(n19793), .ZN(n19812) );
  AND2_X1 U12473 ( .A1(n19763), .A2(n20023), .ZN(n19811) );
  INV_X1 U12474 ( .A(n19826), .ZN(n19829) );
  NAND2_X1 U12475 ( .A1(n19864), .A2(n20162), .ZN(n19934) );
  OAI22_X1 U12476 ( .A1(n18409), .A2(n19560), .B1(n20421), .B2(n19562), .ZN(
        n19946) );
  INV_X1 U12477 ( .A(n20043), .ZN(n19988) );
  OAI22_X1 U12478 ( .A1(n19540), .A2(n19562), .B1(n19539), .B2(n19560), .ZN(
        n19992) );
  OAI21_X1 U12479 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n20006) );
  NOR2_X1 U12480 ( .A1(n19936), .A2(n19935), .ZN(n20004) );
  OAI22_X1 U12481 ( .A1(n19563), .A2(n19562), .B1(n19561), .B2(n19560), .ZN(
        n20005) );
  OAI22_X1 U12482 ( .A1(n14029), .A2(n19562), .B1(n14030), .B2(n19560), .ZN(
        n20040) );
  INV_X1 U12483 ( .A(n19995), .ZN(n20045) );
  OAI22_X1 U12484 ( .A1(n19546), .A2(n19560), .B1(n20462), .B2(n19562), .ZN(
        n20049) );
  NAND2_X1 U12485 ( .A1(n19864), .A2(n20023), .ZN(n20059) );
  INV_X1 U12486 ( .A(n20059), .ZN(n20066) );
  INV_X1 U12487 ( .A(n19106), .ZN(n16551) );
  INV_X1 U12488 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n20079) );
  INV_X1 U12489 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n12466) );
  AND3_X1 U12490 ( .A1(n20083), .A2(n20146), .A3(n20084), .ZN(n20224) );
  NAND2_X1 U12491 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20083), .ZN(n20230) );
  INV_X1 U12492 ( .A(n10165), .ZN(n16732) );
  NOR2_X1 U12493 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16920), .ZN(n16905) );
  NOR4_X1 U12494 ( .A1(n17120), .A2(n18980), .A3(n18977), .A4(n16960), .ZN(
        n16942) );
  INV_X1 U12495 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17914) );
  INV_X1 U12496 ( .A(n17028), .ZN(n17048) );
  NAND2_X1 U12497 ( .A1(n9828), .A2(n10033), .ZN(n19032) );
  NAND2_X1 U12498 ( .A1(n17101), .A2(n19037), .ZN(n10033) );
  INV_X1 U12499 ( .A(n17116), .ZN(n17091) );
  NAND2_X1 U12500 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17130), .ZN(n17116) );
  OAI211_X1 U12501 ( .C1(n18925), .C2(n18926), .A(n17057), .B(n19097), .ZN(
        n17130) );
  NOR2_X1 U12502 ( .A1(n16851), .A2(n17193), .ZN(n17198) );
  INV_X1 U12503 ( .A(n17437), .ZN(n17459) );
  OR2_X1 U12504 ( .A1(n17607), .A2(n17468), .ZN(n10191) );
  NAND2_X1 U12505 ( .A1(n17469), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17466) );
  NOR2_X1 U12506 ( .A1(n17475), .A2(n17675), .ZN(n17469) );
  AND2_X1 U12507 ( .A1(n17493), .A2(n9973), .ZN(n17478) );
  NAND2_X1 U12508 ( .A1(n17493), .A2(n9874), .ZN(n17484) );
  NOR2_X1 U12509 ( .A1(n18449), .A2(n17496), .ZN(n17493) );
  NAND2_X1 U12510 ( .A1(n17493), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17492) );
  NOR2_X1 U12511 ( .A1(n17534), .A2(n10195), .ZN(n17497) );
  NAND2_X1 U12512 ( .A1(n17497), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17496) );
  NOR2_X1 U12513 ( .A1(n17656), .A2(n17522), .ZN(n17517) );
  NOR3_X1 U12514 ( .A1(n18449), .A2(n17534), .A3(n17652), .ZN(n17526) );
  NAND2_X1 U12515 ( .A1(n17535), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17534) );
  NAND4_X1 U12516 ( .A1(n17576), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .A4(n17462), .ZN(n17539) );
  NOR2_X1 U12517 ( .A1(n17571), .A2(n17695), .ZN(n17576) );
  INV_X1 U12518 ( .A(n16619), .ZN(n17578) );
  OR2_X1 U12519 ( .A1(n10048), .A2(n15754), .ZN(n15756) );
  AND4_X1 U12520 ( .A1(n10411), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10295) );
  NOR2_X1 U12521 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  NOR2_X1 U12522 ( .A1(n17683), .A2(n17594), .ZN(n17600) );
  INV_X1 U12523 ( .A(n17605), .ZN(n17601) );
  NOR2_X1 U12524 ( .A1(n17603), .A2(n17681), .ZN(n17602) );
  INV_X1 U12525 ( .A(n17607), .ZN(n17573) );
  NOR2_X1 U12526 ( .A1(n18893), .A2(n17596), .ZN(n17605) );
  NOR2_X1 U12527 ( .A1(n19084), .A2(n17709), .ZN(n17669) );
  OAI211_X1 U12528 ( .C1(n19084), .C2(n19085), .A(n9877), .B(n17648), .ZN(
        n17702) );
  BUF_X1 U12529 ( .A(n17702), .Z(n17709) );
  CLKBUF_X1 U12530 ( .A(n17669), .Z(n17710) );
  INV_X1 U12531 ( .A(n16764), .ZN(n17045) );
  AND2_X1 U12532 ( .A1(n18083), .A2(n10176), .ZN(n17826) );
  AOI21_X1 U12533 ( .B1(n17805), .B2(n17982), .A(n17803), .ZN(n10176) );
  INV_X1 U12534 ( .A(n17929), .ZN(n17884) );
  NOR2_X2 U12535 ( .A1(n19042), .A2(n18078), .ZN(n17929) );
  INV_X1 U12536 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18054) );
  INV_X1 U12537 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18071) );
  INV_X1 U12538 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19042) );
  NOR2_X1 U12539 ( .A1(n10031), .A2(n15863), .ZN(n16565) );
  INV_X1 U12540 ( .A(n10089), .ZN(n17721) );
  NAND2_X1 U12541 ( .A1(n17780), .A2(n15860), .ZN(n17771) );
  INV_X1 U12542 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18177) );
  AND2_X1 U12543 ( .A1(n10175), .A2(n10173), .ZN(n18383) );
  INV_X1 U12544 ( .A(n18090), .ZN(n18307) );
  AND3_X1 U12545 ( .A1(n15857), .A2(n15856), .A3(n15855), .ZN(n17860) );
  NAND2_X1 U12546 ( .A1(n10169), .A2(n10175), .ZN(n18309) );
  NOR2_X1 U12547 ( .A1(n18874), .A2(n10172), .ZN(n10169) );
  INV_X1 U12548 ( .A(n10047), .ZN(n17938) );
  NAND2_X1 U12549 ( .A1(n18391), .A2(n16619), .ZN(n18299) );
  INV_X1 U12550 ( .A(n18299), .ZN(n18315) );
  INV_X1 U12551 ( .A(n10083), .ZN(n10082) );
  AND2_X1 U12552 ( .A1(n18188), .A2(n18357), .ZN(n18324) );
  INV_X1 U12553 ( .A(n18392), .ZN(n18328) );
  NOR2_X1 U12554 ( .A1(n10170), .A2(n18392), .ZN(n18322) );
  NOR2_X1 U12555 ( .A1(n18052), .A2(n15818), .ZN(n18041) );
  INV_X1 U12556 ( .A(n18371), .ZN(n18384) );
  INV_X1 U12557 ( .A(n18322), .ZN(n18395) );
  INV_X1 U12558 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18903) );
  INV_X1 U12559 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U12560 ( .A1(n18896), .A2(n13107), .B1(n9820), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19057) );
  OAI21_X1 U12561 ( .B1(n18872), .B2(n10034), .A(n18873), .ZN(n19036) );
  INV_X1 U12562 ( .A(n17101), .ZN(n10034) );
  INV_X1 U12563 ( .A(n19060), .ZN(n19062) );
  OAI211_X1 U12564 ( .C1(n19078), .C2(n18901), .A(n18410), .B(n15741), .ZN(
        n19060) );
  INV_X1 U12565 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18415) );
  INV_X1 U12566 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18435) );
  INV_X1 U12567 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18441) );
  INV_X1 U12568 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18454) );
  INV_X1 U12569 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18813) );
  NOR2_X1 U12570 ( .A1(n18925), .A2(n18177), .ZN(n18920) );
  NAND2_X1 U12571 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19042), .ZN(n18925) );
  AND2_X1 U12572 ( .A1(n18915), .A2(n18914), .ZN(n10019) );
  NAND2_X1 U12573 ( .A1(n18950), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19093) );
  AND2_X2 U12574 ( .A1(n12345), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20415)
         );
  CLKBUF_X1 U12575 ( .A(n16718), .Z(n16717) );
  NAND2_X1 U12576 ( .A1(n14685), .A2(n13719), .ZN(n12333) );
  NAND2_X1 U12577 ( .A1(n19429), .A2(n10266), .ZN(n10265) );
  AOI21_X1 U12578 ( .B1(n14394), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n9844), .ZN(n10250) );
  OAI21_X1 U12579 ( .B1(n15370), .B2(n15640), .A(n10248), .ZN(n10247) );
  NAND2_X1 U12580 ( .A1(n9919), .A2(n10006), .ZN(P2_U3029) );
  NAND2_X1 U12581 ( .A1(n15523), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10006) );
  AOI21_X1 U12582 ( .B1(n10097), .B2(n17076), .A(n9908), .ZN(n16782) );
  XNOR2_X1 U12583 ( .A(n16775), .B(n10098), .ZN(n10097) );
  OAI21_X1 U12584 ( .B1(n10193), .B2(n10192), .A(n10190), .ZN(P3_U2705) );
  AND2_X1 U12585 ( .A1(n17467), .A2(n10191), .ZN(n10190) );
  OAI21_X1 U12586 ( .B1(n17469), .B2(P3_EAX_REG_30__SCAN_IN), .A(n17596), .ZN(
        n10192) );
  INV_X1 U12587 ( .A(n17466), .ZN(n10193) );
  OAI21_X1 U12588 ( .B1(n16593), .B2(n17978), .A(n10303), .ZN(P3_U2801) );
  NOR3_X1 U12589 ( .A1(n10307), .A2(n10305), .A3(n10304), .ZN(n10303) );
  AND2_X1 U12590 ( .A1(n16594), .A2(n10306), .ZN(n10305) );
  NAND2_X1 U12591 ( .A1(n10087), .A2(n9854), .ZN(P3_U2802) );
  NAND2_X1 U12592 ( .A1(n17723), .A2(n17722), .ZN(n10088) );
  NAND2_X1 U12593 ( .A1(n17807), .A2(n10149), .ZN(P3_U2808) );
  AOI21_X1 U12594 ( .B1(n17808), .B2(n18159), .A(n10150), .ZN(n10149) );
  INV_X1 U12595 ( .A(n15772), .ZN(n15787) );
  INV_X1 U12596 ( .A(n11949), .ZN(n11268) );
  INV_X2 U12597 ( .A(n11268), .ZN(n11648) );
  INV_X1 U12598 ( .A(n17360), .ZN(n17344) );
  NAND2_X2 U12599 ( .A1(n9898), .A2(n12468), .ZN(n12473) );
  NOR3_X1 U12600 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14395), .ZN(n9844) );
  AND4_X1 U12601 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9845)
         );
  OR3_X1 U12602 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n13111), .ZN(n10408) );
  INV_X2 U12603 ( .A(n14110), .ZN(n14183) );
  AND2_X1 U12604 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15834), .ZN(
        n15835) );
  AND4_X1 U12605 ( .A1(n11088), .A2(n11090), .A3(n11089), .A4(n9985), .ZN(
        n9847) );
  INV_X1 U12606 ( .A(n11027), .ZN(n10904) );
  INV_X1 U12607 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14995) );
  AND4_X1 U12608 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n9848) );
  INV_X1 U12609 ( .A(n12581), .ZN(n12624) );
  INV_X1 U12610 ( .A(n15224), .ZN(n10370) );
  AND2_X1 U12611 ( .A1(n9884), .A2(n15449), .ZN(n9849) );
  OR3_X1 U12612 ( .A1(n14488), .A2(n12317), .A3(n10330), .ZN(n9850) );
  AND2_X1 U12613 ( .A1(n10221), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9851) );
  AND2_X1 U12614 ( .A1(n13369), .A2(n11128), .ZN(n9852) );
  AND2_X1 U12615 ( .A1(n10100), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9853) );
  AND3_X1 U12616 ( .A1(n17728), .A2(n9924), .A3(n10085), .ZN(n9854) );
  AND2_X1 U12617 ( .A1(n10073), .A2(n10072), .ZN(n9856) );
  AND2_X1 U12618 ( .A1(n9916), .A2(n10715), .ZN(n9857) );
  AND2_X1 U12619 ( .A1(n11234), .A2(n11232), .ZN(n9858) );
  NOR2_X1 U12620 ( .A1(n10354), .A2(n16398), .ZN(n9859) );
  AND2_X1 U12621 ( .A1(n10096), .A2(n17735), .ZN(n9860) );
  AND3_X1 U12622 ( .A1(n10618), .A2(n20217), .A3(n9922), .ZN(n9861) );
  AND2_X1 U12623 ( .A1(n20588), .A2(n10062), .ZN(n9862) );
  OR2_X1 U12624 ( .A1(n20423), .A2(n20440), .ZN(n12217) );
  AND2_X1 U12625 ( .A1(n10256), .A2(n11157), .ZN(n9863) );
  AND2_X1 U12626 ( .A1(n10301), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9864) );
  AND4_X1 U12627 ( .A1(n10231), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9865) );
  AND2_X1 U12628 ( .A1(n10090), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9866) );
  AND2_X1 U12629 ( .A1(n10224), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9867) );
  AND2_X1 U12630 ( .A1(n10227), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9868) );
  AND2_X1 U12631 ( .A1(n15864), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9869) );
  AND2_X1 U12632 ( .A1(n9866), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U12633 ( .A1(n9959), .A2(n12837), .ZN(n9871) );
  AND2_X1 U12634 ( .A1(n14275), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9872) );
  AND2_X1 U12635 ( .A1(n10080), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9873) );
  AND2_X1 U12636 ( .A1(n10196), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n9874) );
  AND2_X1 U12637 ( .A1(n10374), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9875) );
  NOR2_X1 U12638 ( .A1(n18879), .A2(n13112), .ZN(n13142) );
  INV_X1 U12639 ( .A(n13132), .ZN(n15793) );
  NOR2_X1 U12640 ( .A1(n15729), .A2(n10166), .ZN(n9877) );
  NAND2_X1 U12641 ( .A1(n13979), .A2(n10315), .ZN(n14038) );
  OR3_X1 U12642 ( .A1(n14597), .A2(n10336), .A3(n14535), .ZN(n9878) );
  INV_X1 U12643 ( .A(n17978), .ZN(n17989) );
  OR2_X1 U12644 ( .A1(n14105), .A2(n10204), .ZN(n9879) );
  NOR2_X1 U12645 ( .A1(n15885), .A2(n18883), .ZN(n18894) );
  INV_X1 U12646 ( .A(n10170), .ZN(n18868) );
  NAND2_X1 U12647 ( .A1(n10171), .A2(n10175), .ZN(n10170) );
  NAND2_X1 U12648 ( .A1(n13979), .A2(n13978), .ZN(n13977) );
  AND2_X1 U12649 ( .A1(n15254), .A2(n10376), .ZN(n9880) );
  NOR2_X1 U12650 ( .A1(n18936), .A2(n18055), .ZN(n17858) );
  AND2_X1 U12651 ( .A1(n17493), .A2(n10196), .ZN(n9881) );
  AND2_X1 U12652 ( .A1(n11324), .A2(n11323), .ZN(n9882) );
  AND2_X1 U12653 ( .A1(n12944), .A2(n10309), .ZN(n9883) );
  OR3_X1 U12654 ( .A1(n16346), .A2(n14110), .A3(n15437), .ZN(n9884) );
  INV_X1 U12655 ( .A(n15848), .ZN(n10072) );
  NOR2_X1 U12656 ( .A1(n15631), .A2(n15632), .ZN(n15614) );
  AND4_X1 U12657 ( .A1(n11243), .A2(n11242), .A3(n11241), .A4(n11240), .ZN(
        n9886) );
  OR2_X1 U12658 ( .A1(n15597), .A2(n15598), .ZN(n9887) );
  AND2_X1 U12659 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n9888) );
  AND2_X1 U12660 ( .A1(n10014), .A2(n9861), .ZN(n9889) );
  OR2_X1 U12661 ( .A1(n11112), .A2(n12833), .ZN(n9890) );
  INV_X1 U12662 ( .A(n15246), .ZN(n14240) );
  AND2_X1 U12663 ( .A1(n15065), .A2(n15064), .ZN(n9891) );
  INV_X1 U12664 ( .A(n15448), .ZN(n10353) );
  AND3_X1 U12665 ( .A1(n15369), .A2(n15368), .A3(n15367), .ZN(n9892) );
  AND2_X1 U12666 ( .A1(n10134), .A2(n10391), .ZN(n9893) );
  OR2_X1 U12667 ( .A1(n14465), .A2(n10319), .ZN(n9894) );
  AND2_X1 U12668 ( .A1(n19057), .A2(n18898), .ZN(n9896) );
  INV_X1 U12669 ( .A(n15820), .ZN(n10040) );
  OR2_X1 U12670 ( .A1(n14210), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9897) );
  AND2_X1 U12671 ( .A1(n14204), .A2(n12569), .ZN(n9898) );
  NAND2_X2 U12672 ( .A1(n10186), .A2(n14223), .ZN(n15637) );
  NAND2_X2 U12673 ( .A1(n10540), .A2(n10539), .ZN(n19554) );
  AND3_X1 U12674 ( .A1(n15530), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n14160), .ZN(n9899) );
  AND2_X1 U12675 ( .A1(n10355), .A2(n9859), .ZN(n9900) );
  NOR2_X1 U12676 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n15852), .ZN(
        n9901) );
  BUF_X1 U12677 ( .A(n14204), .Z(n19547) );
  INV_X1 U12678 ( .A(n13347), .ZN(n13350) );
  OAI21_X1 U12679 ( .B1(n10119), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10117), 
        .ZN(n13347) );
  OR2_X1 U12680 ( .A1(n12402), .A2(n19554), .ZN(n9902) );
  AND3_X1 U12681 ( .A1(n10251), .A2(n14403), .A3(n10250), .ZN(n9903) );
  AND2_X1 U12682 ( .A1(n15162), .A2(n15151), .ZN(n15142) );
  AND2_X1 U12683 ( .A1(n10074), .A2(n10040), .ZN(n9904) );
  NOR2_X1 U12684 ( .A1(n15056), .A2(n15055), .ZN(n9905) );
  AND2_X1 U12685 ( .A1(n13915), .A2(n10182), .ZN(n9906) );
  INV_X1 U12686 ( .A(n10015), .ZN(n15528) );
  OAI21_X1 U12687 ( .B1(n15515), .B2(n15514), .A(n15521), .ZN(n10015) );
  AND2_X1 U12688 ( .A1(n13818), .A2(n13862), .ZN(n9907) );
  INV_X1 U12689 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20218) );
  OR2_X1 U12690 ( .A1(n16778), .A2(n16779), .ZN(n9908) );
  AND2_X1 U12691 ( .A1(n13754), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9909) );
  AND2_X1 U12692 ( .A1(n14805), .A2(n16217), .ZN(n9910) );
  AND2_X1 U12693 ( .A1(n10636), .A2(n10635), .ZN(n9911) );
  AND2_X1 U12694 ( .A1(n15041), .A2(n15036), .ZN(n14255) );
  AND2_X1 U12695 ( .A1(n15860), .A2(n15920), .ZN(n9912) );
  AND2_X1 U12696 ( .A1(n10378), .A2(n13403), .ZN(n9913) );
  AND2_X1 U12697 ( .A1(n10632), .A2(n10631), .ZN(n9914) );
  OR2_X1 U12698 ( .A1(n10498), .A2(n10497), .ZN(n9915) );
  NAND2_X1 U12699 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9916) );
  NAND2_X1 U12700 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n9917) );
  NAND2_X1 U12701 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n9918) );
  AND2_X1 U12702 ( .A1(n10011), .A2(n10007), .ZN(n9919) );
  AND2_X1 U12703 ( .A1(n10076), .A2(n10075), .ZN(n9920) );
  INV_X1 U12704 ( .A(n15835), .ZN(n10073) );
  AND2_X1 U12705 ( .A1(n20423), .A2(n10311), .ZN(n9921) );
  AND2_X1 U12706 ( .A1(n10604), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9922) );
  AND2_X1 U12707 ( .A1(n10144), .A2(n10143), .ZN(n9923) );
  INV_X1 U12708 ( .A(n17577), .ZN(n18449) );
  NOR2_X1 U12709 ( .A1(n17724), .A2(n10086), .ZN(n9924) );
  INV_X2 U12710 ( .A(n14336), .ZN(n14334) );
  OR2_X1 U12711 ( .A1(n16591), .A2(n16592), .ZN(n9925) );
  AND2_X1 U12712 ( .A1(n9853), .A2(n10099), .ZN(n9926) );
  INV_X1 U12713 ( .A(n14330), .ZN(n10399) );
  NAND2_X1 U12714 ( .A1(n9859), .A2(n15599), .ZN(n9927) );
  NOR2_X1 U12715 ( .A1(n20710), .A2(n20429), .ZN(n9928) );
  AND2_X1 U12716 ( .A1(n15112), .A2(n13993), .ZN(n13992) );
  NOR2_X1 U12717 ( .A1(n13721), .A2(n10252), .ZN(n9929) );
  NOR2_X1 U12718 ( .A1(n13933), .A2(n13934), .ZN(n13932) );
  INV_X1 U12719 ( .A(n15264), .ZN(n10203) );
  AND2_X1 U12720 ( .A1(n12364), .A2(n10221), .ZN(n9930) );
  OR2_X1 U12721 ( .A1(n16081), .A2(n14678), .ZN(n9931) );
  AND2_X1 U12722 ( .A1(n10611), .A2(n10612), .ZN(n11111) );
  OR2_X1 U12723 ( .A1(n13721), .A2(n13722), .ZN(n9932) );
  NOR2_X1 U12724 ( .A1(n16467), .A2(n10243), .ZN(n9933) );
  OR2_X1 U12725 ( .A1(n15565), .A2(n10238), .ZN(n14019) );
  INV_X1 U12726 ( .A(n16070), .ZN(n10402) );
  AND2_X1 U12727 ( .A1(n15089), .A2(n15099), .ZN(n9934) );
  OR3_X1 U12728 ( .A1(n13735), .A2(n12273), .A3(n13734), .ZN(n9935) );
  OR3_X1 U12729 ( .A1(n13735), .A2(n12273), .A3(n10333), .ZN(n9936) );
  NOR2_X1 U12730 ( .A1(n15565), .A2(n10235), .ZN(n14023) );
  AND2_X1 U12731 ( .A1(n15855), .A2(n18203), .ZN(n9937) );
  OR2_X1 U12732 ( .A1(n14334), .A2(n14866), .ZN(n9938) );
  NOR2_X1 U12733 ( .A1(n15565), .A2(n10237), .ZN(n9939) );
  INV_X1 U12734 ( .A(n20588), .ZN(n10122) );
  INV_X1 U12735 ( .A(n10045), .ZN(n17924) );
  NAND2_X1 U12736 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  AND2_X1 U12737 ( .A1(n11596), .A2(n11546), .ZN(n9940) );
  AND2_X1 U12738 ( .A1(n10082), .A2(n17902), .ZN(n9941) );
  AND2_X1 U12739 ( .A1(n10116), .A2(n10121), .ZN(n9942) );
  INV_X1 U12740 ( .A(n10334), .ZN(n14588) );
  NOR2_X1 U12741 ( .A1(n14597), .A2(n10336), .ZN(n10334) );
  OR2_X1 U12742 ( .A1(n14334), .A2(n14348), .ZN(n9943) );
  AND2_X1 U12743 ( .A1(n13992), .A2(n10257), .ZN(n15067) );
  OR2_X1 U12744 ( .A1(n14096), .A2(n14204), .ZN(n14194) );
  AND2_X1 U12745 ( .A1(n10257), .A2(n15068), .ZN(n9944) );
  AND2_X1 U12746 ( .A1(n13544), .A2(n13513), .ZN(n9945) );
  INV_X1 U12747 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16407) );
  INV_X1 U12748 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19295) );
  AND2_X1 U12749 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n9946) );
  NOR2_X1 U12750 ( .A1(n19081), .A2(n15888), .ZN(n18890) );
  INV_X1 U12751 ( .A(n18890), .ZN(n10174) );
  INV_X1 U12752 ( .A(n15640), .ZN(n16492) );
  INV_X1 U12753 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21026) );
  NOR2_X1 U12754 ( .A1(n14093), .A2(n10717), .ZN(n13091) );
  AND2_X1 U12755 ( .A1(n15935), .A2(n10227), .ZN(n9947) );
  AND2_X1 U12756 ( .A1(n15940), .A2(n10224), .ZN(n9948) );
  AND2_X1 U12757 ( .A1(n15177), .A2(n15438), .ZN(n9949) );
  AND2_X1 U12758 ( .A1(n9949), .A2(n10241), .ZN(n9950) );
  AND2_X1 U12759 ( .A1(n14256), .A2(n15018), .ZN(n9951) );
  OR2_X1 U12760 ( .A1(n14208), .A2(n12459), .ZN(n9952) );
  NAND2_X1 U12761 ( .A1(n9847), .A2(n9987), .ZN(n13782) );
  INV_X1 U12762 ( .A(n13481), .ZN(n14994) );
  AND2_X1 U12763 ( .A1(n10210), .A2(n10208), .ZN(n9953) );
  NOR2_X1 U12764 ( .A1(n18026), .A2(n15822), .ZN(n9954) );
  OR2_X1 U12765 ( .A1(n14208), .A2(n14126), .ZN(n9955) );
  INV_X1 U12766 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10062) );
  AND2_X1 U12767 ( .A1(n11118), .A2(n11117), .ZN(n9956) );
  NOR2_X1 U12768 ( .A1(n14093), .A2(n10284), .ZN(n9957) );
  INV_X1 U12769 ( .A(n10269), .ZN(n10268) );
  NOR2_X1 U12770 ( .A1(n11051), .A2(n10270), .ZN(n10269) );
  NAND2_X1 U12771 ( .A1(n10941), .A2(n10940), .ZN(n9958) );
  AND2_X1 U12772 ( .A1(n12523), .A2(n13555), .ZN(n9959) );
  INV_X1 U12773 ( .A(n10316), .ZN(n10315) );
  NAND2_X1 U12774 ( .A1(n11763), .A2(n10317), .ZN(n10316) );
  OR2_X1 U12775 ( .A1(n10267), .A2(n10269), .ZN(n9960) );
  AND2_X1 U12776 ( .A1(n9960), .A2(n19429), .ZN(n9961) );
  NOR2_X1 U12777 ( .A1(n18041), .A2(n18040), .ZN(n9962) );
  AND2_X1 U12778 ( .A1(n9950), .A2(n10240), .ZN(n9963) );
  AND2_X1 U12779 ( .A1(n9951), .A2(n14226), .ZN(n9964) );
  INV_X1 U12780 ( .A(n11011), .ZN(n10263) );
  NOR2_X4 U12781 ( .A1(n13107), .A2(n10032), .ZN(n9965) );
  AND2_X1 U12782 ( .A1(n17927), .A2(n10100), .ZN(n9966) );
  AND2_X1 U12783 ( .A1(n17747), .A2(n10090), .ZN(n9967) );
  INV_X1 U12784 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10207) );
  OR2_X1 U12785 ( .A1(n16566), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9968) );
  OR2_X1 U12786 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9969) );
  AND2_X1 U12787 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .ZN(n9970) );
  INV_X1 U12788 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10091) );
  INV_X1 U12789 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10208) );
  INV_X1 U12790 ( .A(n13343), .ZN(n10283) );
  AND2_X1 U12791 ( .A1(n10187), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9971) );
  AND2_X1 U12792 ( .A1(n14355), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9972) );
  AND2_X1 U12793 ( .A1(n9874), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9973) );
  INV_X1 U12794 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n10197) );
  INV_X1 U12795 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10198) );
  INV_X1 U12796 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U12797 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9974) );
  INV_X1 U12798 ( .A(n9832), .ZN(n9975) );
  NAND3_X1 U12799 ( .A1(n19058), .A2(n18923), .A3(n18177), .ZN(n18388) );
  OAI22_X1 U12800 ( .A1(n18164), .A2(n17978), .B1(n18995), .B2(n18388), .ZN(
        n10154) );
  AOI22_X2 U12801 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19559), .ZN(n20060) );
  INV_X1 U12802 ( .A(n21024), .ZN(n9976) );
  INV_X1 U12803 ( .A(n9976), .ZN(n9977) );
  INV_X1 U12804 ( .A(n20914), .ZN(n9978) );
  INV_X1 U12805 ( .A(n9978), .ZN(n9979) );
  INV_X1 U12806 ( .A(n20929), .ZN(n9980) );
  INV_X1 U12807 ( .A(n9980), .ZN(n9981) );
  INV_X1 U12808 ( .A(n20902), .ZN(n9982) );
  INV_X1 U12809 ( .A(n9982), .ZN(n9983) );
  AOI22_X2 U12810 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20476), .B1(DATAI_22_), 
        .B2(n20477), .ZN(n20922) );
  AOI22_X2 U12811 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19559), .ZN(n20038) );
  AOI22_X2 U12812 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20476), .B1(DATAI_18_), 
        .B2(n20477), .ZN(n20906) );
  NOR2_X1 U12813 ( .A1(n20417), .A2(n20416), .ZN(n20476) );
  NOR2_X1 U12814 ( .A1(n20415), .A2(n20417), .ZN(n20477) );
  NOR4_X4 U12815 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n19042), .ZN(n17076) );
  INV_X1 U12816 ( .A(n11091), .ZN(n9987) );
  NOR2_X4 U12817 ( .A1(n9990), .A2(n9989), .ZN(n13926) );
  AND2_X2 U12818 ( .A1(n14112), .A2(n9993), .ZN(n14161) );
  NAND2_X2 U12820 ( .A1(n15246), .A2(n14241), .ZN(n14249) );
  OAI21_X2 U12821 ( .B1(n10352), .B2(n9995), .A(n9884), .ZN(n10351) );
  NAND3_X1 U12822 ( .A1(n10000), .A2(n10268), .A3(n9999), .ZN(n15117) );
  NAND2_X1 U12823 ( .A1(n15022), .A2(n10267), .ZN(n9999) );
  OR2_X2 U12824 ( .A1(n15022), .A2(n10270), .ZN(n10000) );
  XNOR2_X2 U12825 ( .A(n10692), .B(n11129), .ZN(n19509) );
  NOR2_X2 U12826 ( .A1(n13653), .A2(n13958), .ZN(n13725) );
  XNOR2_X2 U12827 ( .A(n10969), .B(n10965), .ZN(n15049) );
  AND3_X2 U12828 ( .A1(n10276), .A2(n10278), .A3(n9958), .ZN(n10969) );
  NAND2_X1 U12829 ( .A1(n13434), .A2(n13433), .ZN(n13432) );
  NAND2_X2 U12830 ( .A1(n10004), .A2(n14087), .ZN(n14093) );
  INV_X2 U12831 ( .A(n12402), .ZN(n14204) );
  NAND3_X1 U12832 ( .A1(n10714), .A2(n19541), .A3(n10005), .ZN(n10634) );
  AOI21_X2 U12833 ( .B1(n10262), .B2(n9855), .A(n15026), .ZN(n15034) );
  OAI211_X2 U12834 ( .C1(n13880), .C2(n13911), .A(n13879), .B(n13878), .ZN(
        n13881) );
  OAI21_X2 U12835 ( .B1(n10604), .B2(n20217), .A(n12581), .ZN(n13026) );
  NAND2_X1 U12836 ( .A1(n10557), .A2(n16502), .ZN(n10012) );
  NAND2_X1 U12837 ( .A1(n10562), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10013) );
  INV_X1 U12838 ( .A(n12614), .ZN(n10014) );
  NAND3_X1 U12839 ( .A1(n13783), .A2(n13782), .A3(n13818), .ZN(n13863) );
  NAND2_X1 U12840 ( .A1(n13822), .A2(n13863), .ZN(n13869) );
  NAND3_X1 U12841 ( .A1(n18913), .A2(n18912), .A3(n19075), .ZN(n10021) );
  NAND3_X1 U12842 ( .A1(n15721), .A2(n15716), .A3(n15720), .ZN(n15737) );
  INV_X2 U12843 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13107) );
  NOR2_X1 U12844 ( .A1(n15986), .A2(n10031), .ZN(n15987) );
  NAND3_X1 U12845 ( .A1(n10039), .A2(n10038), .A3(n10036), .ZN(n18027) );
  NAND4_X1 U12846 ( .A1(n10039), .A2(n10038), .A3(n9864), .A4(n10036), .ZN(
        n10041) );
  NAND2_X2 U12847 ( .A1(n10300), .A2(n10041), .ZN(n18016) );
  NAND3_X1 U12848 ( .A1(n15755), .A2(n10050), .A3(n10049), .ZN(n10048) );
  NAND4_X1 U12849 ( .A1(n10055), .A2(n15753), .A3(n10054), .A4(n10053), .ZN(
        n10052) );
  NAND2_X2 U12850 ( .A1(n11556), .A2(n11555), .ZN(n11586) );
  AND2_X2 U12851 ( .A1(n11226), .A2(n10058), .ZN(n11400) );
  AND2_X2 U12852 ( .A1(n11227), .A2(n10058), .ZN(n11399) );
  OAI21_X1 U12853 ( .B1(n10108), .B2(n11366), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11384) );
  NAND2_X1 U12854 ( .A1(n11366), .A2(n10061), .ZN(n10059) );
  NAND2_X1 U12855 ( .A1(n10108), .A2(n10061), .ZN(n10060) );
  AND2_X2 U12856 ( .A1(n10064), .A2(n10140), .ZN(n14714) );
  INV_X1 U12857 ( .A(n14724), .ZN(n10064) );
  NAND2_X2 U12858 ( .A1(n13769), .A2(n13768), .ZN(n14336) );
  INV_X1 U12859 ( .A(n18016), .ZN(n10068) );
  NAND3_X1 U12860 ( .A1(n10070), .A2(n10071), .A3(n10069), .ZN(n17994) );
  INV_X1 U12861 ( .A(n15849), .ZN(n17869) );
  NAND2_X1 U12862 ( .A1(n10077), .A2(n17756), .ZN(n17745) );
  INV_X1 U12863 ( .A(n17902), .ZN(n18271) );
  NAND3_X1 U12864 ( .A1(n10089), .A2(n17989), .A3(n10088), .ZN(n10087) );
  AOI21_X1 U12865 ( .B1(n16816), .B2(n17735), .A(n9840), .ZN(n16796) );
  NAND2_X1 U12866 ( .A1(n10093), .A2(n10092), .ZN(n16795) );
  NAND2_X1 U12867 ( .A1(n16816), .A2(n10094), .ZN(n10093) );
  INV_X1 U12868 ( .A(n10096), .ZN(n16805) );
  AND2_X1 U12869 ( .A1(n17916), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10102) );
  AND2_X1 U12870 ( .A1(n13394), .A2(n12806), .ZN(n10103) );
  MUX2_X1 U12871 ( .A(n12806), .B(n10104), .S(n12965), .Z(n11303) );
  NAND2_X1 U12872 ( .A1(n20471), .A2(n20463), .ZN(n10104) );
  AND2_X2 U12873 ( .A1(n11354), .A2(n20463), .ZN(n12806) );
  NAND2_X1 U12874 ( .A1(n11576), .A2(n20463), .ZN(n11360) );
  NAND2_X2 U12875 ( .A1(n9886), .A2(n9848), .ZN(n20463) );
  NAND3_X1 U12876 ( .A1(n10106), .A2(n11365), .A3(n10105), .ZN(n11367) );
  NAND4_X1 U12877 ( .A1(n9913), .A2(n11363), .A3(n11362), .A4(n10109), .ZN(
        n10108) );
  NAND2_X2 U12878 ( .A1(n10110), .A2(n9883), .ZN(n11366) );
  INV_X1 U12879 ( .A(n12942), .ZN(n10110) );
  NAND2_X1 U12880 ( .A1(n10118), .A2(n9862), .ZN(n10113) );
  INV_X1 U12881 ( .A(n10112), .ZN(n10111) );
  OAI21_X1 U12882 ( .B1(n10114), .B2(n11391), .A(n11511), .ZN(n10112) );
  NAND2_X1 U12883 ( .A1(n10115), .A2(n20588), .ZN(n10121) );
  INV_X1 U12884 ( .A(n11391), .ZN(n10115) );
  NAND3_X1 U12885 ( .A1(n13679), .A2(n13680), .A3(n13752), .ZN(n10388) );
  OAI21_X1 U12886 ( .B1(n10397), .B2(n10128), .A(n16081), .ZN(n10124) );
  OR2_X2 U12887 ( .A1(n10396), .A2(n10125), .ZN(n10130) );
  INV_X1 U12888 ( .A(n10397), .ZN(n10125) );
  INV_X1 U12889 ( .A(n9893), .ZN(n10132) );
  NAND2_X1 U12890 ( .A1(n10127), .A2(n10126), .ZN(n14760) );
  NAND3_X1 U12891 ( .A1(n9893), .A2(n10129), .A3(n10130), .ZN(n10126) );
  NAND3_X1 U12892 ( .A1(n10131), .A2(n14783), .A3(n10130), .ZN(n14768) );
  NAND2_X1 U12893 ( .A1(n10136), .A2(n10133), .ZN(n10134) );
  OR2_X2 U12894 ( .A1(n10139), .A2(n14679), .ZN(n10138) );
  NOR2_X2 U12895 ( .A1(n14714), .A2(n9943), .ZN(n14679) );
  AND2_X2 U12896 ( .A1(n14714), .A2(n14680), .ZN(n10139) );
  NAND2_X1 U12897 ( .A1(n13864), .A2(n13917), .ZN(n13868) );
  NOR2_X1 U12898 ( .A1(n12563), .A2(n12581), .ZN(n10612) );
  NAND2_X1 U12899 ( .A1(n14103), .A2(n9923), .ZN(n10142) );
  NAND2_X2 U12900 ( .A1(n16733), .A2(n9968), .ZN(n18083) );
  NAND4_X1 U12901 ( .A1(n13510), .A2(n13509), .A3(n13507), .A4(n13508), .ZN(
        n10177) );
  NAND4_X1 U12902 ( .A1(n13540), .A2(n13539), .A3(n13537), .A4(n13538), .ZN(
        n10178) );
  NAND2_X1 U12903 ( .A1(n10601), .A2(n16502), .ZN(n10180) );
  NAND2_X1 U12904 ( .A1(n10179), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10181) );
  NAND4_X1 U12905 ( .A1(n10597), .A2(n10600), .A3(n10598), .A4(n10599), .ZN(
        n10179) );
  NAND2_X2 U12906 ( .A1(n10181), .A2(n10180), .ZN(n10604) );
  NAND2_X1 U12907 ( .A1(n10618), .A2(n12467), .ZN(n13943) );
  INV_X1 U12908 ( .A(n14217), .ZN(n10184) );
  NAND2_X1 U12909 ( .A1(n13916), .A2(n13915), .ZN(n14219) );
  NAND2_X1 U12910 ( .A1(n15454), .A2(n10189), .ZN(n15280) );
  AND2_X2 U12911 ( .A1(n15454), .A2(n10187), .ZN(n15254) );
  INV_X2 U12912 ( .A(n17377), .ZN(n15837) );
  NAND3_X1 U12913 ( .A1(n9845), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .ZN(n10195) );
  AND2_X1 U12914 ( .A1(n9877), .A2(n18416), .ZN(n10200) );
  INV_X1 U12915 ( .A(n15885), .ZN(n10201) );
  INV_X1 U12916 ( .A(n10213), .ZN(n14181) );
  AND2_X2 U12917 ( .A1(n10212), .A2(n10209), .ZN(n14185) );
  NAND3_X1 U12918 ( .A1(n10361), .A2(n9897), .A3(n10359), .ZN(n10358) );
  NAND2_X1 U12919 ( .A1(n10360), .A2(n10370), .ZN(n10359) );
  NAND2_X1 U12920 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10230) );
  INV_X1 U12921 ( .A(n12359), .ZN(n10231) );
  NAND3_X1 U12922 ( .A1(n10231), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12360) );
  AND2_X2 U12923 ( .A1(n15176), .A2(n9963), .ZN(n15162) );
  NAND3_X1 U12924 ( .A1(n10633), .A2(n12564), .A3(n12614), .ZN(n10636) );
  NAND3_X1 U12925 ( .A1(n10254), .A2(n14008), .A3(n10253), .ZN(n10252) );
  INV_X1 U12926 ( .A(n13983), .ZN(n10255) );
  NAND2_X1 U12927 ( .A1(n14255), .A2(n9951), .ZN(n15017) );
  NAND2_X1 U12928 ( .A1(n14255), .A2(n9964), .ZN(n14234) );
  AND2_X1 U12929 ( .A1(n14255), .A2(n14256), .ZN(n15019) );
  NAND2_X1 U12930 ( .A1(n15022), .A2(n9961), .ZN(n10264) );
  OAI211_X1 U12931 ( .C1(n15022), .C2(n10265), .A(n10264), .B(n10271), .ZN(
        P2_U2889) );
  NAND2_X1 U12932 ( .A1(n13009), .A2(n13010), .ZN(n10275) );
  NAND2_X1 U12933 ( .A1(n15065), .A2(n10277), .ZN(n10276) );
  INV_X2 U12934 ( .A(n17415), .ZN(n13106) );
  NAND2_X2 U12935 ( .A1(n17859), .A2(n17951), .ZN(n17780) );
  NOR2_X1 U12936 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  INV_X1 U12937 ( .A(n15776), .ZN(n10289) );
  NAND4_X1 U12938 ( .A1(n10295), .A2(n10291), .A3(n10290), .A4(n10294), .ZN(
        n17597) );
  NAND2_X1 U12939 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10294) );
  NAND2_X1 U12940 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U12941 ( .A1(n15822), .A2(n10301), .ZN(n10300) );
  OR2_X2 U12942 ( .A1(n15854), .A2(n15863), .ZN(n17966) );
  INV_X1 U12943 ( .A(n17993), .ZN(n10302) );
  NAND3_X1 U12944 ( .A1(n16600), .A2(n9925), .A3(n16602), .ZN(n10304) );
  OAI22_X2 U12945 ( .A1(n12871), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13329), 
        .B2(n11492), .ZN(n11412) );
  INV_X1 U12946 ( .A(n12737), .ZN(n10312) );
  NAND4_X1 U12947 ( .A1(n10312), .A2(n9921), .A3(n11352), .A4(n13632), .ZN(
        n10309) );
  NAND3_X1 U12948 ( .A1(n13631), .A2(n12239), .A3(n10310), .ZN(n12944) );
  NAND4_X1 U12949 ( .A1(n10312), .A2(n13632), .A3(n11352), .A4(n20423), .ZN(
        n15971) );
  AND2_X2 U12950 ( .A1(n13979), .A2(n10314), .ZN(n14074) );
  OR2_X2 U12951 ( .A1(n14465), .A2(n10321), .ZN(n14440) );
  AND2_X2 U12952 ( .A1(n14576), .A2(n10323), .ZN(n14478) );
  NOR2_X2 U12953 ( .A1(n13099), .A2(n13098), .ZN(n13379) );
  NOR3_X4 U12954 ( .A1(n13735), .A2(n12273), .A3(n10332), .ZN(n14060) );
  INV_X1 U12955 ( .A(n14543), .ZN(n10338) );
  NAND2_X1 U12956 ( .A1(n10624), .A2(n10339), .ZN(n10625) );
  NAND2_X1 U12957 ( .A1(n12612), .A2(n10339), .ZN(n12613) );
  XNOR2_X2 U12958 ( .A(n13581), .B(n13580), .ZN(n13583) );
  AND3_X1 U12959 ( .A1(n10611), .A2(n10612), .A3(n9946), .ZN(n10414) );
  NAND2_X1 U12960 ( .A1(n13576), .A2(n13575), .ZN(n10343) );
  NAND2_X1 U12961 ( .A1(n10340), .A2(n10344), .ZN(n16448) );
  NAND3_X1 U12962 ( .A1(n10343), .A2(n13577), .A3(n10342), .ZN(n10340) );
  NAND3_X1 U12963 ( .A1(n13863), .A2(n13822), .A3(n14110), .ZN(n10341) );
  NAND2_X1 U12964 ( .A1(n16448), .A2(n16447), .ZN(n13830) );
  NOR2_X1 U12965 ( .A1(n9849), .A2(n15278), .ZN(n10348) );
  NAND3_X1 U12966 ( .A1(n10350), .A2(n10351), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10349) );
  INV_X1 U12967 ( .A(n15451), .ZN(n10350) );
  NAND2_X1 U12968 ( .A1(n14240), .A2(n10369), .ZN(n10363) );
  INV_X1 U12969 ( .A(n14250), .ZN(n10372) );
  NAND4_X1 U12970 ( .A1(n9819), .A2(n10605), .A3(n20217), .A4(n10628), .ZN(
        n12367) );
  XNOR2_X1 U12971 ( .A(n12983), .B(n12981), .ZN(n12970) );
  AND2_X1 U12972 ( .A1(n12878), .A2(n10378), .ZN(n12238) );
  MUX2_X1 U12973 ( .A(n11473), .B(n11474), .S(n11354), .Z(n11476) );
  OAI22_X1 U12974 ( .A1(n12944), .A2(n10380), .B1(n15971), .B2(n20440), .ZN(
        n12945) );
  NAND3_X1 U12975 ( .A1(n11417), .A2(n20890), .A3(n10062), .ZN(n11435) );
  NAND2_X1 U12976 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  NAND2_X1 U12977 ( .A1(n20366), .A2(n13670), .ZN(n10387) );
  NAND2_X1 U12978 ( .A1(n20366), .A2(n13670), .ZN(n10385) );
  OAI21_X1 U12979 ( .B1(n20366), .B2(n13670), .A(n13664), .ZN(n10386) );
  AND2_X2 U12980 ( .A1(n14335), .A2(n10398), .ZN(n10397) );
  NAND2_X1 U12981 ( .A1(n14478), .A2(n14480), .ZN(n14479) );
  NAND2_X1 U12982 ( .A1(n11668), .A2(n11667), .ZN(n13712) );
  NAND2_X1 U12983 ( .A1(n10403), .A2(n11584), .ZN(n12974) );
  NAND2_X1 U12984 ( .A1(n17906), .A2(n10410), .ZN(n17870) );
  NAND2_X1 U12985 ( .A1(n13103), .A2(n13102), .ZN(n13101) );
  NAND2_X1 U12986 ( .A1(n14595), .A2(n14594), .ZN(n14542) );
  CLKBUF_X1 U12987 ( .A(n13596), .Z(n13638) );
  INV_X1 U12988 ( .A(n13596), .ZN(n11668) );
  INV_X1 U12989 ( .A(n13382), .ZN(n11611) );
  NAND2_X1 U12990 ( .A1(n11611), .A2(n11610), .ZN(n13608) );
  OAI21_X1 U12991 ( .B1(n12986), .B2(n11762), .A(n11561), .ZN(n11562) );
  OR2_X1 U12992 ( .A1(n12986), .A2(n13350), .ZN(n20934) );
  OR2_X1 U12993 ( .A1(n12986), .A2(n13347), .ZN(n20686) );
  AND2_X1 U12994 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20190), .ZN(
        n11070) );
  AND2_X2 U12995 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15664) );
  AOI21_X1 U12996 ( .B1(n14414), .B2(n14411), .A(n14410), .ZN(n14412) );
  NAND2_X1 U12997 ( .A1(n15861), .A2(n15921), .ZN(n15859) );
  CLKBUF_X1 U12998 ( .A(n12642), .Z(n12908) );
  OR2_X1 U12999 ( .A1(n15852), .A2(n17993), .ZN(n15853) );
  INV_X4 U13000 ( .A(n10408), .ZN(n17412) );
  INV_X1 U13001 ( .A(n14343), .ZN(n11356) );
  OR2_X2 U13002 ( .A1(n13480), .A2(n13495), .ZN(n19977) );
  INV_X1 U13003 ( .A(n12962), .ZN(n11564) );
  NAND2_X1 U13004 ( .A1(n14760), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14712) );
  NAND2_X1 U13005 ( .A1(n13911), .A2(n13868), .ZN(n13878) );
  OR2_X1 U13006 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12178) );
  INV_X1 U13007 ( .A(n12178), .ZN(n12145) );
  NOR2_X1 U13008 ( .A1(n13997), .A2(n13998), .ZN(n10404) );
  OR2_X1 U13009 ( .A1(n10969), .A2(n10968), .ZN(n10405) );
  AND2_X1 U13010 ( .A1(n10986), .A2(n10418), .ZN(n10406) );
  AND4_X1 U13011 ( .A1(n10603), .A2(n16528), .A3(n10602), .A4(n10714), .ZN(
        n10407) );
  NAND2_X1 U13012 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10409) );
  AND3_X1 U13013 ( .A1(n18267), .A2(n17903), .A3(n18231), .ZN(n10410) );
  OR2_X1 U13014 ( .A1(n9885), .A2(n17262), .ZN(n10411) );
  AND2_X1 U13015 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10412) );
  OR2_X1 U13016 ( .A1(n12606), .A2(n20218), .ZN(n10413) );
  AND3_X1 U13017 ( .A1(n11253), .A2(n11252), .A3(n11251), .ZN(n10415) );
  INV_X1 U13018 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13670) );
  NAND2_X1 U13019 ( .A1(n10894), .A2(n16502), .ZN(n10416) );
  OR2_X1 U13020 ( .A1(n10541), .A2(n13469), .ZN(n10417) );
  INV_X1 U13021 ( .A(n12470), .ZN(n12503) );
  NOR2_X1 U13022 ( .A1(n17578), .A2(n16621), .ZN(n15851) );
  INV_X1 U13023 ( .A(n17951), .ZN(n15863) );
  AND3_X1 U13024 ( .A1(n11007), .A2(n11008), .A3(n10983), .ZN(n10418) );
  INV_X1 U13025 ( .A(n15802), .ZN(n17608) );
  OR2_X2 U13026 ( .A1(n19037), .A2(n13108), .ZN(n10419) );
  AND2_X1 U13027 ( .A1(n17459), .A2(n18449), .ZN(n17456) );
  OR3_X1 U13028 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17798), .ZN(n10420) );
  NAND2_X1 U13029 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10421) );
  INV_X1 U13030 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20083) );
  INV_X1 U13031 ( .A(n17596), .ZN(n17516) );
  INV_X1 U13032 ( .A(n12504), .ZN(n12517) );
  INV_X1 U13033 ( .A(n17858), .ZN(n17823) );
  NAND2_X1 U13034 ( .A1(n21026), .A2(n20422), .ZN(n20593) );
  INV_X2 U13035 ( .A(n13719), .ZN(n14610) );
  NOR2_X1 U13036 ( .A1(n14600), .A2(n14381), .ZN(n13719) );
  INV_X2 U13037 ( .A(n13047), .ZN(n20361) );
  AND2_X1 U13038 ( .A1(n12232), .A2(n12212), .ZN(n12220) );
  INV_X1 U13039 ( .A(n11061), .ZN(n10498) );
  INV_X1 U13040 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13478) );
  INV_X1 U13041 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13487) );
  INV_X1 U13042 ( .A(n12202), .ZN(n12200) );
  INV_X1 U13043 ( .A(n11545), .ZN(n11546) );
  OAI22_X1 U13044 ( .A1(n11027), .A2(n10590), .B1(n11028), .B2(n10589), .ZN(
        n10591) );
  NAND2_X1 U13045 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10454) );
  AND2_X1 U13046 ( .A1(n20889), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12197) );
  INV_X1 U13047 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11966) );
  OR2_X1 U13048 ( .A1(n11540), .A2(n11539), .ZN(n13759) );
  AND2_X1 U13049 ( .A1(n11527), .A2(n11526), .ZN(n11544) );
  INV_X1 U13050 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11230) );
  AND4_X1 U13051 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12456) );
  NAND2_X1 U13052 ( .A1(n10605), .A2(n9839), .ZN(n10606) );
  OAI21_X1 U13053 ( .B1(n12568), .B2(n10714), .A(n12569), .ZN(n10623) );
  OR2_X1 U13054 ( .A1(n13189), .A2(n15713), .ZN(n13185) );
  NOR2_X1 U13055 ( .A1(n20478), .A2(n21028), .ZN(n11578) );
  NOR2_X1 U13056 ( .A1(n11408), .A2(n11407), .ZN(n13329) );
  OR2_X1 U13057 ( .A1(n11624), .A2(n11623), .ZN(n13758) );
  INV_X1 U13058 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11214) );
  NOR2_X1 U13059 ( .A1(n11938), .A2(n12066), .ZN(n11215) );
  OR2_X1 U13060 ( .A1(n12436), .A2(n12435), .ZN(n13858) );
  OR2_X1 U13061 ( .A1(n10982), .A2(n10984), .ZN(n11007) );
  AND2_X1 U13062 ( .A1(n15075), .A2(n10874), .ZN(n10885) );
  NAND2_X1 U13063 ( .A1(n11082), .A2(n11081), .ZN(n11105) );
  NAND2_X1 U13064 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10479) );
  OAI21_X1 U13065 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19055), .A(
        n13185), .ZN(n13191) );
  OR2_X1 U13066 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20414), .ZN(
        n12230) );
  AND4_X1 U13067 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(
        n11324) );
  OR2_X1 U13068 ( .A1(n12119), .A2(n14696), .ZN(n12120) );
  NOR2_X1 U13069 ( .A1(n11982), .A2(n14763), .ZN(n11983) );
  INV_X1 U13070 ( .A(n11578), .ZN(n11633) );
  INV_X1 U13071 ( .A(n13639), .ZN(n11667) );
  AND3_X1 U13072 ( .A1(n13767), .A2(n13766), .A3(n13771), .ZN(n13768) );
  OR2_X1 U13073 ( .A1(n11509), .A2(n11508), .ZN(n13673) );
  AND4_X1 U13074 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11233) );
  INV_X1 U13075 ( .A(n12847), .ZN(n12723) );
  AND2_X1 U13076 ( .A1(n10885), .A2(n13962), .ZN(n10886) );
  AND2_X1 U13077 ( .A1(n12506), .A2(n12505), .ZN(n12512) );
  OR2_X2 U13078 ( .A1(n13480), .A2(n13496), .ZN(n19938) );
  INV_X1 U13079 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17397) );
  NOR2_X1 U13080 ( .A1(n9885), .A2(n17397), .ZN(n15761) );
  NAND2_X1 U13081 ( .A1(n15863), .A2(n18091), .ZN(n15865) );
  AND2_X1 U13082 ( .A1(n12231), .A2(n12230), .ZN(n12648) );
  INV_X1 U13083 ( .A(n11921), .ZN(n11922) );
  AND2_X1 U13084 ( .A1(n12271), .A2(n12270), .ZN(n13734) );
  NAND2_X1 U13085 ( .A1(n12318), .A2(n11356), .ZN(n12252) );
  NOR2_X1 U13086 ( .A1(n11938), .A2(n11963), .ZN(n11313) );
  NOR2_X1 U13087 ( .A1(n11938), .A2(n11332), .ZN(n11333) );
  OR2_X1 U13088 ( .A1(n12120), .A2(n14433), .ZN(n13397) );
  OR2_X1 U13089 ( .A1(n14368), .A2(n21026), .ZN(n12148) );
  INV_X1 U13090 ( .A(n12178), .ZN(n13391) );
  AND2_X1 U13091 ( .A1(n11764), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U13092 ( .A1(n11576), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U13093 ( .A1(n11647), .A2(n11646), .ZN(n13597) );
  INV_X1 U13094 ( .A(n16068), .ZN(n14327) );
  OR2_X1 U13095 ( .A1(n14958), .A2(n16180), .ZN(n13005) );
  INV_X1 U13096 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20839) );
  AND3_X1 U13097 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21026), .A3(n20422), 
        .ZN(n20479) );
  NAND2_X1 U13098 ( .A1(n11102), .A2(n11101), .ZN(n12589) );
  AND2_X1 U13099 ( .A1(n20218), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n10699) );
  NOR2_X1 U13100 ( .A1(n15465), .A2(n15471), .ZN(n15459) );
  OR2_X1 U13101 ( .A1(n14173), .A2(n15590), .ZN(n15581) );
  AND2_X1 U13102 ( .A1(n14274), .A2(n14273), .ZN(n15568) );
  INV_X1 U13103 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13547) );
  NAND2_X1 U13104 ( .A1(n10682), .A2(n12466), .ZN(n10704) );
  INV_X1 U13105 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17414) );
  AOI21_X1 U13106 ( .B1(n17318), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n15761), .ZN(n15762) );
  INV_X1 U13107 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17143) );
  NAND2_X1 U13108 ( .A1(n10422), .A2(n15865), .ZN(n15866) );
  NOR2_X1 U13109 ( .A1(n15863), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17853) );
  OR2_X1 U13110 ( .A1(n17588), .A2(n15897), .ZN(n15895) );
  INV_X1 U13111 ( .A(n18421), .ZN(n15728) );
  INV_X2 U13112 ( .A(n14343), .ZN(n12327) );
  INV_X1 U13113 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16029) );
  NAND2_X1 U13114 ( .A1(n11669), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11702) );
  AND2_X1 U13115 ( .A1(n12283), .A2(n12282), .ZN(n14606) );
  OR2_X1 U13116 ( .A1(n16018), .A2(n12178), .ZN(n11926) );
  AND2_X1 U13117 ( .A1(n20478), .A2(n20471), .ZN(n13631) );
  INV_X1 U13118 ( .A(n14377), .ZN(n12184) );
  NAND2_X1 U13119 ( .A1(n12036), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12087) );
  NOR2_X1 U13120 ( .A1(n11841), .A2(n16029), .ZN(n11878) );
  NOR2_X1 U13121 ( .A1(n11757), .A2(n11725), .ZN(n11764) );
  NOR2_X1 U13122 ( .A1(n11702), .A2(n11701), .ZN(n11706) );
  AND4_X1 U13123 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n13639) );
  AND2_X1 U13124 ( .A1(n11587), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11549) );
  OR2_X1 U13125 ( .A1(n20370), .A2(n12794), .ZN(n14824) );
  NAND2_X1 U13126 ( .A1(n12954), .A2(n12951), .ZN(n20398) );
  AND2_X1 U13127 ( .A1(n13693), .A2(n13692), .ZN(n14939) );
  INV_X1 U13128 ( .A(n20513), .ZN(n20420) );
  AND2_X1 U13129 ( .A1(n20930), .A2(n20427), .ZN(n20771) );
  INV_X1 U13130 ( .A(n20477), .ZN(n20468) );
  OR2_X1 U13131 ( .A1(n20934), .A2(n20813), .ZN(n20976) );
  AND2_X1 U13132 ( .A1(n12589), .A2(n12372), .ZN(n16529) );
  AND2_X1 U13133 ( .A1(n12462), .A2(n12461), .ZN(n14118) );
  OR3_X1 U13134 ( .A1(n12463), .A2(n9838), .A3(n16260), .ZN(n19328) );
  NOR2_X1 U13135 ( .A1(n13612), .A2(n13952), .ZN(n10774) );
  NAND2_X1 U13136 ( .A1(n16534), .A2(n13018), .ZN(n13025) );
  INV_X1 U13137 ( .A(n10921), .ZN(n15076) );
  OR2_X1 U13138 ( .A1(n10851), .A2(n13988), .ZN(n13989) );
  OAI21_X1 U13139 ( .B1(n12356), .B2(n12355), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12357) );
  OR3_X1 U13140 ( .A1(n15426), .A2(n15401), .A3(n15278), .ZN(n15379) );
  OR2_X1 U13141 ( .A1(n15493), .A2(n14276), .ZN(n15471) );
  INV_X1 U13142 ( .A(n19310), .ZN(n19294) );
  OAI21_X1 U13143 ( .B1(n13561), .B2(n15512), .A(n13560), .ZN(n14274) );
  OR2_X1 U13144 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  AND2_X1 U13145 ( .A1(n19583), .A2(n19582), .ZN(n19763) );
  AND2_X1 U13146 ( .A1(n20174), .A2(n19667), .ZN(n19944) );
  INV_X1 U13147 ( .A(n19944), .ZN(n19935) );
  OR2_X1 U13148 ( .A1(n19583), .A2(n20194), .ZN(n19936) );
  INV_X1 U13149 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20013) );
  NAND2_X1 U13150 ( .A1(n15874), .A2(n15875), .ZN(n18865) );
  INV_X1 U13151 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17055) );
  INV_X1 U13152 ( .A(n17115), .ZN(n17126) );
  INV_X1 U13153 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15691) );
  OAI21_X1 U13154 ( .B1(n15888), .B2(n18869), .A(n13200), .ZN(n16000) );
  INV_X1 U13155 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17932) );
  NOR2_X1 U13156 ( .A1(n15895), .A2(n17584), .ZN(n18012) );
  NOR2_X1 U13157 ( .A1(n18358), .A2(n18053), .ZN(n18052) );
  INV_X1 U13158 ( .A(n18864), .ZN(n16556) );
  NOR2_X1 U13159 ( .A1(n18075), .A2(n18082), .ZN(n18074) );
  NOR2_X1 U13160 ( .A1(n15971), .A2(n20235), .ZN(n12650) );
  NOR2_X1 U13161 ( .A1(n13404), .A2(n13394), .ZN(n13413) );
  AND2_X1 U13162 ( .A1(n20277), .A2(n13399), .ZN(n20292) );
  OAI22_X1 U13163 ( .A1(n14842), .A2(n14613), .B1(n21192), .B2(n14612), .ZN(
        n12331) );
  NAND2_X1 U13164 ( .A1(n14506), .A2(n14500), .ZN(n14499) );
  INV_X1 U13165 ( .A(n14613), .ZN(n14601) );
  INV_X1 U13166 ( .A(n13043), .ZN(n14316) );
  NAND2_X1 U13167 ( .A1(n11707), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11757) );
  AND2_X1 U13168 ( .A1(n14824), .A2(n12960), .ZN(n16094) );
  AND2_X1 U13169 ( .A1(n15965), .A2(n13627), .ZN(n20370) );
  AND2_X1 U13170 ( .A1(n14934), .A2(n14346), .ZN(n14919) );
  NOR2_X1 U13171 ( .A1(n16126), .A2(n14354), .ZN(n14934) );
  NAND2_X1 U13172 ( .A1(n13696), .A2(n20398), .ZN(n16234) );
  AND2_X1 U13173 ( .A1(n12954), .A2(n12950), .ZN(n14958) );
  INV_X1 U13174 ( .A(n20398), .ZN(n16180) );
  INV_X1 U13175 ( .A(n14939), .ZN(n20395) );
  AND2_X1 U13176 ( .A1(n12954), .A2(n14373), .ZN(n14956) );
  OAI22_X1 U13178 ( .A1(n20436), .A2(n20435), .B1(n20774), .B2(n20590), .ZN(
        n20483) );
  OAI22_X1 U13179 ( .A1(n20521), .A2(n20520), .B1(n20774), .B2(n20648), .ZN(
        n20544) );
  OR2_X1 U13180 ( .A1(n20419), .A2(n20418), .ZN(n20555) );
  INV_X1 U13181 ( .A(n20596), .ZN(n20613) );
  OR2_X1 U13182 ( .A1(n13316), .A2(n20420), .ZN(n20838) );
  OAI22_X1 U13183 ( .A1(n20650), .A2(n20649), .B1(n20648), .B2(n20930), .ZN(
        n20673) );
  NAND2_X1 U13184 ( .A1(n13316), .A2(n20420), .ZN(n20813) );
  OAI211_X1 U13185 ( .C1(n20731), .C2(n20847), .A(n20771), .B(n20715), .ZN(
        n20733) );
  OAI22_X1 U13186 ( .A1(n20776), .A2(n20775), .B1(n20774), .B2(n20931), .ZN(
        n20800) );
  AND2_X1 U13187 ( .A1(n20419), .A2(n12986), .ZN(n20815) );
  INV_X1 U13188 ( .A(n20894), .ZN(n20925) );
  INV_X1 U13189 ( .A(n21023), .ZN(n20958) );
  NOR2_X1 U13190 ( .A1(n21028), .A2(n21025), .ZN(n13321) );
  INV_X1 U13191 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20232) );
  INV_X1 U13192 ( .A(n19328), .ZN(n19346) );
  AND2_X1 U13193 ( .A1(n13951), .A2(n13950), .ZN(n14018) );
  NAND2_X1 U13194 ( .A1(n16259), .A2(n12375), .ZN(n19325) );
  AND2_X1 U13195 ( .A1(n16501), .A2(n12632), .ZN(n19333) );
  OR2_X1 U13196 ( .A1(n10862), .A2(n10861), .ZN(n15082) );
  AND2_X1 U13197 ( .A1(n19368), .A2(n13971), .ZN(n19362) );
  OR2_X1 U13198 ( .A1(n13997), .A2(n13941), .ZN(n15108) );
  INV_X1 U13199 ( .A(n19389), .ZN(n19396) );
  NOR2_X1 U13200 ( .A1(n15655), .A2(n13365), .ZN(n19582) );
  INV_X1 U13201 ( .A(n12659), .ZN(n19486) );
  AND2_X1 U13202 ( .A1(n19514), .A2(n20183), .ZN(n19510) );
  OR2_X1 U13203 ( .A1(n15430), .A2(n14271), .ZN(n15419) );
  NOR2_X1 U13204 ( .A1(n15636), .A2(n16460), .ZN(n16392) );
  INV_X1 U13205 ( .A(n16477), .ZN(n16490) );
  INV_X1 U13206 ( .A(n19509), .ZN(n13468) );
  NAND2_X1 U13207 ( .A1(n15512), .A2(n15519), .ZN(n15517) );
  AND2_X1 U13208 ( .A1(n19763), .A2(n20162), .ZN(n19693) );
  AND2_X1 U13209 ( .A1(n19725), .A2(n19944), .ZN(n19717) );
  AND2_X1 U13210 ( .A1(n19733), .A2(n19729), .ZN(n19751) );
  AND2_X1 U13211 ( .A1(n19583), .A2(n20194), .ZN(n19725) );
  NOR2_X1 U13212 ( .A1(n20174), .A2(n20184), .ZN(n19584) );
  AND2_X1 U13213 ( .A1(n19864), .A2(n19584), .ZN(n19859) );
  INV_X1 U13214 ( .A(n19863), .ZN(n19894) );
  NOR2_X1 U13215 ( .A1(n20174), .A2(n19667), .ZN(n20162) );
  NOR2_X2 U13216 ( .A1(n19969), .A2(n19935), .ZN(n19958) );
  NOR2_X1 U13217 ( .A1(n19969), .A2(n19968), .ZN(n20056) );
  NAND2_X1 U13218 ( .A1(n18920), .A2(n18865), .ZN(n17609) );
  INV_X1 U13219 ( .A(n17067), .ZN(n19097) );
  OR2_X1 U13220 ( .A1(n16787), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16774) );
  NOR2_X1 U13221 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16897), .ZN(n16883) );
  NOR2_X1 U13222 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16943), .ZN(n16925) );
  NOR2_X1 U13223 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16963), .ZN(n16949) );
  NOR2_X1 U13224 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16996), .ZN(n16995) );
  NOR2_X1 U13225 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17061), .ZN(n17040) );
  NAND2_X1 U13226 ( .A1(n18914), .A2(n16749), .ZN(n17120) );
  NOR4_X1 U13227 ( .A1(n17274), .A2(n17278), .A3(n17437), .A4(n17279), .ZN(
        n17260) );
  NAND3_X1 U13228 ( .A1(n18412), .A2(n16000), .A3(n16557), .ZN(n17437) );
  OAI211_X1 U13229 ( .C1(n9828), .C2(n18446), .A(n15833), .B(n15832), .ZN(
        n18008) );
  INV_X1 U13230 ( .A(n17646), .ZN(n17611) );
  NOR2_X1 U13231 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18411), .ZN(n18765) );
  INV_X1 U13232 ( .A(n18086), .ZN(n18076) );
  INV_X1 U13233 ( .A(n18148), .ZN(n18190) );
  INV_X1 U13234 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18290) );
  OAI211_X1 U13235 ( .C1(n16556), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        n15883) );
  NOR2_X1 U13236 ( .A1(n18863), .A2(n18392), .ZN(n18391) );
  NOR2_X1 U13237 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19031), .ZN(
        n19056) );
  INV_X1 U13238 ( .A(n18794), .ZN(n18767) );
  CLKBUF_X1 U13239 ( .A(n18515), .Z(n18511) );
  INV_X1 U13240 ( .A(n18519), .ZN(n18582) );
  INV_X1 U13241 ( .A(n18587), .ZN(n18663) );
  INV_X1 U13242 ( .A(n18669), .ZN(n18733) );
  INV_X1 U13243 ( .A(n18691), .ZN(n18757) );
  INV_X1 U13244 ( .A(n19085), .ZN(n18938) );
  NAND2_X1 U13245 ( .A1(n13620), .A2(n12650), .ZN(n12867) );
  INV_X1 U13246 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21220) );
  NAND2_X1 U13247 ( .A1(n13413), .A2(n13412), .ZN(n20313) );
  INV_X1 U13248 ( .A(n20292), .ZN(n16051) );
  OR2_X1 U13249 ( .A1(n20279), .A2(n13738), .ZN(n16055) );
  INV_X1 U13250 ( .A(n20264), .ZN(n20324) );
  INV_X1 U13251 ( .A(n12331), .ZN(n12332) );
  INV_X1 U13252 ( .A(n14788), .ZN(n14662) );
  OR2_X1 U13253 ( .A1(n14052), .A2(n14051), .ZN(n16091) );
  AND2_X1 U13254 ( .A1(n13628), .A2(n13627), .ZN(n14647) );
  OR2_X1 U13255 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16248), .ZN(n20326) );
  INV_X1 U13256 ( .A(n20328), .ZN(n20349) );
  NOR2_X1 U13257 ( .A1(n12867), .A2(n12866), .ZN(n13047) );
  OR2_X1 U13258 ( .A1(n20361), .A2(n20440), .ZN(n14320) );
  INV_X1 U13259 ( .A(n16094), .ZN(n20374) );
  INV_X1 U13260 ( .A(n20405), .ZN(n20387) );
  INV_X1 U13261 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20414) );
  OR2_X1 U13262 ( .A1(n20555), .A2(n20838), .ZN(n20506) );
  OR2_X1 U13263 ( .A1(n20555), .A2(n20742), .ZN(n20548) );
  OR2_X1 U13264 ( .A1(n20555), .A2(n20933), .ZN(n20582) );
  OR2_X1 U13265 ( .A1(n20686), .A2(n20838), .ZN(n20642) );
  OR2_X1 U13266 ( .A1(n20686), .A2(n20742), .ZN(n20677) );
  OR2_X1 U13267 ( .A1(n20686), .A2(n20813), .ZN(n20700) );
  NAND2_X1 U13268 ( .A1(n20815), .A2(n20709), .ZN(n20762) );
  NAND2_X1 U13269 ( .A1(n20815), .A2(n20763), .ZN(n20829) );
  NAND2_X1 U13270 ( .A1(n20815), .A2(n20814), .ZN(n20886) );
  NAND2_X1 U13271 ( .A1(n20888), .A2(n20887), .ZN(n20962) );
  INV_X1 U13272 ( .A(n20907), .ZN(n20997) );
  INV_X1 U13273 ( .A(n21030), .ZN(n21094) );
  NOR2_X1 U13274 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20232), .ZN(n21064) );
  INV_X1 U13275 ( .A(n21076), .ZN(n21082) );
  INV_X1 U13276 ( .A(n21064), .ZN(n21115) );
  NAND2_X1 U13277 ( .A1(n12706), .A2(n16551), .ZN(n19108) );
  INV_X1 U13278 ( .A(n19333), .ZN(n19340) );
  INV_X1 U13279 ( .A(n19290), .ZN(n19349) );
  INV_X1 U13280 ( .A(n15110), .ZN(n15106) );
  INV_X1 U13281 ( .A(n19429), .ZN(n19366) );
  AND2_X1 U13282 ( .A1(n19366), .A2(n19365), .ZN(n19389) );
  AND2_X1 U13283 ( .A1(n19370), .A2(n19369), .ZN(n19434) );
  NAND2_X1 U13284 ( .A1(n12749), .A2(n12748), .ZN(n19437) );
  NAND2_X1 U13285 ( .A1(n12747), .A2(n20224), .ZN(n19476) );
  NAND2_X1 U13286 ( .A1(n12638), .A2(n9838), .ZN(n12745) );
  INV_X1 U13287 ( .A(n16449), .ZN(n19501) );
  INV_X1 U13288 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16385) );
  INV_X1 U13289 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19273) );
  NAND2_X1 U13290 ( .A1(n12708), .A2(n9833), .ZN(n19493) );
  INV_X1 U13291 ( .A(n16493), .ZN(n16457) );
  INV_X1 U13292 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16517) );
  NAND2_X1 U13293 ( .A1(n19584), .A2(n19725), .ZN(n19604) );
  NAND2_X1 U13294 ( .A1(n19725), .A2(n20162), .ZN(n19666) );
  INV_X1 U13295 ( .A(n19717), .ZN(n19724) );
  INV_X1 U13296 ( .A(n19747), .ZN(n19755) );
  NAND2_X1 U13297 ( .A1(n20023), .A2(n19725), .ZN(n19783) );
  INV_X1 U13298 ( .A(n19811), .ZN(n19805) );
  NAND2_X1 U13299 ( .A1(n19835), .A2(n19584), .ZN(n19826) );
  NAND2_X1 U13300 ( .A1(n19835), .A2(n20162), .ZN(n19863) );
  INV_X1 U13301 ( .A(n20030), .ZN(n19914) );
  INV_X1 U13302 ( .A(n20049), .ZN(n19926) );
  INV_X1 U13303 ( .A(n20040), .ZN(n19991) );
  INV_X1 U13304 ( .A(n20004), .ZN(n20001) );
  INV_X1 U13305 ( .A(n19992), .ZN(n20048) );
  INV_X1 U13306 ( .A(n20056), .ZN(n20070) );
  INV_X1 U13307 ( .A(n20161), .ZN(n20081) );
  CLKBUF_X1 U13308 ( .A(n20151), .Z(n20145) );
  INV_X1 U13309 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19083) );
  INV_X1 U13310 ( .A(n17081), .ZN(n17127) );
  AND2_X1 U13311 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17198), .ZN(n17192) );
  NOR2_X1 U13312 ( .A1(n16986), .A2(n17389), .ZN(n17375) );
  NOR2_X1 U13313 ( .A1(n17543), .A2(n17565), .ZN(n17564) );
  NAND2_X1 U13314 ( .A1(n18893), .A2(n17460), .ZN(n17607) );
  NAND2_X1 U13315 ( .A1(n17611), .A2(n18412), .ZN(n17627) );
  NAND2_X1 U13316 ( .A1(n17648), .A2(n17610), .ZN(n17646) );
  NAND2_X1 U13317 ( .A1(n18076), .A2(n16619), .ZN(n17978) );
  OR2_X1 U13318 ( .A1(n18166), .A2(n18165), .ZN(n18186) );
  INV_X1 U13319 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18267) );
  OAI21_X2 U13320 ( .B1(n15884), .B2(n15883), .A(n18920), .ZN(n18392) );
  INV_X1 U13321 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18898) );
  INV_X1 U13322 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18429) );
  INV_X1 U13323 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18446) );
  INV_X1 U13324 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18626) );
  INV_X1 U13325 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18646) );
  INV_X1 U13326 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18654) );
  INV_X1 U13327 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18667) );
  INV_X1 U13328 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18806) );
  INV_X1 U13329 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18827) );
  INV_X1 U13330 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18923) );
  INV_X1 U13331 ( .A(n19027), .ZN(n18937) );
  INV_X1 U13332 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18950) );
  NOR2_X1 U13333 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12358), .ZN(n16718)
         );
  NAND2_X1 U13334 ( .A1(n12333), .A2(n12332), .ZN(P1_U2842) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10945) );
  OR2_X1 U13336 ( .A1(n10541), .A2(n10945), .ZN(n10426) );
  INV_X2 U13337 ( .A(n9895), .ZN(n10894) );
  NAND2_X1 U13338 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13339 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10424) );
  NAND2_X2 U13340 ( .A1(n11072), .A2(n15664), .ZN(n11028) );
  NAND2_X1 U13341 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10423) );
  NAND4_X1 U13342 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10438) );
  INV_X1 U13343 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10427) );
  AND2_X4 U13344 ( .A1(n10429), .A2(n10428), .ZN(n11061) );
  INV_X1 U13345 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10430) );
  INV_X1 U13346 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10432) );
  OR2_X1 U13347 ( .A1(n11037), .A2(n10432), .ZN(n10435) );
  AND3_X4 U13348 ( .A1(n15665), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10889) );
  NAND2_X1 U13349 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10434) );
  INV_X1 U13350 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10946) );
  OR2_X1 U13351 ( .A1(n11036), .A2(n10946), .ZN(n10433) );
  NAND4_X1 U13352 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10437) );
  INV_X1 U13353 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10954) );
  OR2_X1 U13354 ( .A1(n10541), .A2(n10954), .ZN(n10442) );
  NAND2_X1 U13355 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10441) );
  NAND2_X1 U13356 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U13357 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10439) );
  NAND4_X1 U13358 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10450) );
  INV_X1 U13359 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10443) );
  INV_X1 U13360 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10444) );
  OR2_X1 U13361 ( .A1(n11037), .A2(n10444), .ZN(n10447) );
  NAND2_X1 U13362 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10446) );
  INV_X1 U13363 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10955) );
  OR2_X1 U13364 ( .A1(n11036), .A2(n10955), .ZN(n10445) );
  NAND4_X1 U13365 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  NOR2_X1 U13366 ( .A1(n10450), .A2(n10449), .ZN(n10567) );
  MUX2_X2 U13367 ( .A(n10576), .B(n10567), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10618) );
  INV_X2 U13368 ( .A(n9895), .ZN(n15672) );
  NAND2_X1 U13369 ( .A1(n15672), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13370 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13371 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10451) );
  NAND4_X1 U13372 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10459) );
  INV_X1 U13373 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U13374 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10456) );
  NAND4_X1 U13375 ( .A1(n10421), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10458) );
  NOR2_X1 U13376 ( .A1(n10459), .A2(n10458), .ZN(n10563) );
  NAND2_X1 U13377 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13378 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13379 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10460) );
  NAND4_X1 U13380 ( .A1(n10417), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10468) );
  NAND2_X1 U13381 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10466) );
  INV_X1 U13382 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13499) );
  NAND2_X1 U13383 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10464) );
  NAND4_X1 U13384 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  NOR2_X1 U13385 ( .A1(n10468), .A2(n10467), .ZN(n10583) );
  INV_X1 U13386 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13387 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13388 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13389 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10471) );
  NAND4_X1 U13390 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10481) );
  INV_X1 U13391 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10475) );
  OR2_X1 U13392 ( .A1(n11037), .A2(n10475), .ZN(n10478) );
  NAND2_X1 U13393 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10477) );
  INV_X1 U13394 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10989) );
  OR2_X1 U13395 ( .A1(n11036), .A2(n10989), .ZN(n10476) );
  NAND4_X1 U13396 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10480) );
  NOR2_X1 U13397 ( .A1(n10481), .A2(n10480), .ZN(n10574) );
  INV_X1 U13398 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U13399 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10484) );
  NAND2_X1 U13400 ( .A1(n9827), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10483) );
  NAND2_X1 U13401 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10482) );
  NAND4_X1 U13402 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10491) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10486) );
  OR2_X1 U13404 ( .A1(n11037), .A2(n10486), .ZN(n10489) );
  NAND2_X1 U13405 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10488) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10998) );
  OR2_X1 U13407 ( .A1(n11036), .A2(n10998), .ZN(n10487) );
  NAND4_X1 U13408 ( .A1(n9917), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10490) );
  NOR2_X1 U13409 ( .A1(n10491), .A2(n10490), .ZN(n10564) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13411 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13412 ( .A1(n9827), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10494) );
  INV_X4 U13413 ( .A(n11028), .ZN(n11058) );
  NAND2_X1 U13414 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10493) );
  NAND4_X1 U13415 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10505) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10497) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10499) );
  OR2_X1 U13418 ( .A1(n11037), .A2(n10499), .ZN(n10503) );
  NAND2_X1 U13419 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10502) );
  INV_X1 U13420 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10500) );
  OR2_X1 U13421 ( .A1(n11036), .A2(n10500), .ZN(n10501) );
  NAND4_X1 U13422 ( .A1(n9915), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10504) );
  NAND2_X1 U13423 ( .A1(n10566), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10519) );
  INV_X1 U13424 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U13425 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13426 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10508) );
  NAND2_X1 U13427 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10507) );
  NAND4_X1 U13428 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10517) );
  INV_X1 U13429 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10511) );
  OR2_X1 U13430 ( .A1(n11037), .A2(n10511), .ZN(n10515) );
  NAND2_X1 U13431 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10514) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10512) );
  OR2_X1 U13433 ( .A1(n11036), .A2(n10512), .ZN(n10513) );
  NAND4_X1 U13434 ( .A1(n9918), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10516) );
  NAND2_X1 U13435 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13436 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13437 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10520) );
  NAND4_X1 U13438 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10528) );
  NAND2_X1 U13439 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10525) );
  NAND4_X1 U13440 ( .A1(n10409), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10527) );
  NAND2_X1 U13441 ( .A1(n10579), .A2(n16502), .ZN(n10540) );
  NAND2_X1 U13442 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10531) );
  NAND2_X1 U13443 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13444 ( .A1(n11058), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10529) );
  NAND4_X1 U13445 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10538) );
  NAND2_X1 U13446 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U13447 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10534) );
  NAND4_X1 U13448 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10537) );
  NAND2_X1 U13449 ( .A1(n10565), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10539) );
  AOI22_X1 U13450 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13451 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10544) );
  INV_X2 U13452 ( .A(n11027), .ZN(n11020) );
  AOI22_X1 U13453 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10543) );
  NAND4_X1 U13454 ( .A1(n10545), .A2(n10544), .A3(n10543), .A4(n10542), .ZN(
        n10571) );
  NAND2_X1 U13455 ( .A1(n10571), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10551) );
  AOI22_X1 U13456 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13457 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13458 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13459 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n10889), .ZN(n10546) );
  NAND4_X1 U13460 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10578) );
  NAND2_X1 U13461 ( .A1(n10578), .A2(n16502), .ZN(n10550) );
  INV_X1 U13462 ( .A(n12402), .ZN(n10552) );
  AOI22_X1 U13463 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13464 ( .A1(n15672), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13465 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13466 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10553) );
  NAND4_X1 U13467 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10557) );
  AOI22_X1 U13468 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13469 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13470 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13471 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10558) );
  NAND4_X1 U13472 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n10562) );
  NAND3_X1 U13473 ( .A1(n10564), .A2(n10563), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10573) );
  INV_X1 U13474 ( .A(n10565), .ZN(n10570) );
  INV_X1 U13475 ( .A(n10566), .ZN(n10569) );
  INV_X1 U13476 ( .A(n10567), .ZN(n10568) );
  NAND4_X1 U13477 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  INV_X1 U13478 ( .A(n10574), .ZN(n10575) );
  NOR2_X1 U13479 ( .A1(n10575), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10586) );
  INV_X1 U13480 ( .A(n10576), .ZN(n10577) );
  AND2_X1 U13481 ( .A1(n10578), .A2(n10577), .ZN(n10585) );
  INV_X1 U13482 ( .A(n10579), .ZN(n10582) );
  INV_X1 U13483 ( .A(n10580), .ZN(n10581) );
  AND2_X1 U13484 ( .A1(n10582), .A2(n10581), .ZN(n10584) );
  NAND4_X1 U13485 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10587) );
  AOI22_X1 U13486 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10596) );
  INV_X1 U13487 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10590) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10589) );
  INV_X1 U13489 ( .A(n10591), .ZN(n10593) );
  AOI22_X1 U13490 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10592) );
  AND2_X1 U13491 ( .A1(n10593), .A2(n10592), .ZN(n10595) );
  AOI22_X1 U13492 ( .A1(n10723), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10594) );
  NAND3_X1 U13493 ( .A1(n10596), .A2(n10595), .A3(n10594), .ZN(n10601) );
  AOI22_X1 U13494 ( .A1(n10718), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13495 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13496 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13497 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10723), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10597) );
  INV_X1 U13498 ( .A(n13943), .ZN(n10602) );
  NAND2_X1 U13499 ( .A1(n10646), .A2(n9838), .ZN(n10610) );
  NAND3_X1 U13500 ( .A1(n13026), .A2(n12568), .A3(n12569), .ZN(n10609) );
  NAND2_X1 U13501 ( .A1(n10607), .A2(n10619), .ZN(n10608) );
  NOR2_X2 U13502 ( .A1(n10609), .A2(n10608), .ZN(n11108) );
  NAND2_X1 U13503 ( .A1(n11108), .A2(n12607), .ZN(n10662) );
  NAND2_X1 U13504 ( .A1(n10610), .A2(n10662), .ZN(n12626) );
  NAND2_X2 U13505 ( .A1(n12626), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11112) );
  INV_X1 U13506 ( .A(n10634), .ZN(n10611) );
  INV_X1 U13507 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14996) );
  NOR2_X1 U13508 ( .A1(n10688), .A2(n16528), .ZN(n10613) );
  NAND2_X1 U13509 ( .A1(n11113), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10615) );
  NAND2_X1 U13510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10614) );
  OAI211_X1 U13511 ( .C1(n11196), .C2(n14996), .A(n10615), .B(n10614), .ZN(
        n10616) );
  INV_X1 U13512 ( .A(n10616), .ZN(n10617) );
  NAND2_X1 U13513 ( .A1(n10714), .A2(n12402), .ZN(n10626) );
  NAND3_X1 U13514 ( .A1(n10619), .A2(n10618), .A3(n10626), .ZN(n10622) );
  NAND3_X1 U13515 ( .A1(n10634), .A2(n9838), .A3(n12507), .ZN(n10653) );
  NAND2_X1 U13516 ( .A1(n10653), .A2(n16528), .ZN(n10624) );
  NAND2_X1 U13517 ( .A1(n10625), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10632) );
  INV_X1 U13518 ( .A(n12575), .ZN(n12579) );
  INV_X1 U13519 ( .A(n10626), .ZN(n10627) );
  NAND3_X1 U13520 ( .A1(n10628), .A2(n9819), .A3(n10627), .ZN(n16527) );
  INV_X1 U13521 ( .A(n10618), .ZN(n10629) );
  NOR2_X1 U13522 ( .A1(n9838), .A2(n10629), .ZN(n10630) );
  NAND2_X1 U13523 ( .A1(n16527), .A2(n10630), .ZN(n11109) );
  NAND2_X1 U13524 ( .A1(n20217), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20222) );
  INV_X1 U13525 ( .A(n20222), .ZN(n12748) );
  NAND3_X1 U13526 ( .A1(n12579), .A2(n11109), .A3(n12748), .ZN(n10631) );
  NAND2_X1 U13527 ( .A1(n12507), .A2(n9902), .ZN(n12565) );
  NAND2_X1 U13528 ( .A1(n12565), .A2(n19541), .ZN(n12564) );
  NAND2_X1 U13529 ( .A1(n12507), .A2(n12568), .ZN(n12566) );
  AND2_X1 U13530 ( .A1(n12566), .A2(n12569), .ZN(n10633) );
  NAND2_X1 U13531 ( .A1(n12624), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10659) );
  NOR2_X1 U13532 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16499) );
  AND2_X1 U13533 ( .A1(n16499), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10637) );
  INV_X1 U13534 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12833) );
  INV_X1 U13535 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13536 ( .A1(n11113), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10639) );
  NAND2_X1 U13537 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10638) );
  OAI211_X1 U13538 ( .C1(n11196), .C2(n10640), .A(n10639), .B(n10638), .ZN(
        n10641) );
  INV_X1 U13539 ( .A(n10641), .ZN(n10642) );
  INV_X1 U13540 ( .A(n10691), .ZN(n11130) );
  OAI21_X1 U13541 ( .B1(n20181), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20079), 
        .ZN(n10643) );
  NAND2_X1 U13542 ( .A1(n11130), .A2(n11131), .ZN(n10673) );
  INV_X1 U13543 ( .A(n10673), .ZN(n10644) );
  NOR2_X1 U13544 ( .A1(n11134), .A2(n10644), .ZN(n10681) );
  INV_X1 U13545 ( .A(n11131), .ZN(n10645) );
  NAND2_X1 U13546 ( .A1(n10691), .A2(n10645), .ZN(n10675) );
  AND2_X1 U13547 ( .A1(n11134), .A2(n10675), .ZN(n10680) );
  NAND2_X1 U13548 ( .A1(n10661), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10648) );
  AOI22_X1 U13549 ( .A1(n10646), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16499), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10647) );
  INV_X1 U13550 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15660) );
  INV_X1 U13551 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12391) );
  NAND2_X1 U13552 ( .A1(n11113), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U13553 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10649) );
  OAI211_X1 U13554 ( .C1(n11196), .C2(n12391), .A(n10650), .B(n10649), .ZN(
        n10651) );
  INV_X1 U13555 ( .A(n10651), .ZN(n10652) );
  OAI21_X2 U13556 ( .B1(n11112), .B2(n15660), .A(n10652), .ZN(n10668) );
  XNOR2_X2 U13557 ( .A(n10669), .B(n10668), .ZN(n10696) );
  INV_X1 U13558 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15654) );
  NAND2_X1 U13559 ( .A1(n9911), .A2(n10653), .ZN(n12606) );
  INV_X1 U13560 ( .A(n16499), .ZN(n10663) );
  NAND2_X1 U13561 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U13562 ( .A1(n10663), .A2(n10654), .ZN(n10655) );
  AOI21_X1 U13563 ( .B1(n11113), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10655), .ZN(
        n10656) );
  NAND2_X1 U13564 ( .A1(n10656), .A2(n9914), .ZN(n10657) );
  NOR2_X1 U13565 ( .A1(n10659), .A2(n12563), .ZN(n10660) );
  INV_X1 U13566 ( .A(n10662), .ZN(n10665) );
  NOR2_X1 U13567 ( .A1(n10663), .A2(n20199), .ZN(n10664) );
  NAND2_X1 U13568 ( .A1(n10696), .A2(n10703), .ZN(n10672) );
  INV_X1 U13569 ( .A(n10668), .ZN(n10670) );
  NAND2_X1 U13570 ( .A1(n10670), .A2(n10669), .ZN(n10671) );
  NAND2_X2 U13571 ( .A1(n10672), .A2(n10671), .ZN(n11129) );
  NAND2_X1 U13572 ( .A1(n11134), .A2(n10673), .ZN(n10674) );
  INV_X1 U13573 ( .A(n11134), .ZN(n10676) );
  AND2_X1 U13574 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13575 ( .A1(n11129), .A2(n10677), .ZN(n10678) );
  OAI211_X2 U13576 ( .C1(n10681), .C2(n10680), .A(n10679), .B(n10678), .ZN(
        n13481) );
  BUF_X1 U13577 ( .A(n13481), .Z(n13011) );
  NAND2_X1 U13578 ( .A1(n10714), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U13579 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20012) );
  INV_X1 U13580 ( .A(n20012), .ZN(n10683) );
  NAND2_X1 U13581 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10683), .ZN(
        n10693) );
  INV_X1 U13582 ( .A(n10693), .ZN(n10684) );
  NAND2_X1 U13583 ( .A1(n10684), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20020) );
  INV_X1 U13584 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U13585 ( .A1(n10685), .A2(n10693), .ZN(n10686) );
  AND3_X1 U13586 ( .A1(n20020), .A2(n20169), .A3(n10686), .ZN(n19898) );
  AOI21_X1 U13587 ( .B1(n10704), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19898), .ZN(n10687) );
  OAI21_X2 U13588 ( .B1(n13011), .B2(n12716), .A(n10687), .ZN(n10716) );
  NOR2_X1 U13589 ( .A1(n10688), .A2(n13469), .ZN(n10689) );
  OR2_X1 U13590 ( .A1(n10716), .A2(n10689), .ZN(n10690) );
  NAND2_X1 U13591 ( .A1(n10716), .A2(n10689), .ZN(n14089) );
  AND2_X2 U13592 ( .A1(n10690), .A2(n14089), .ZN(n13010) );
  XNOR2_X1 U13593 ( .A(n10691), .B(n11131), .ZN(n10692) );
  NAND2_X1 U13594 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19865) );
  NAND2_X1 U13595 ( .A1(n19865), .A2(n20181), .ZN(n10694) );
  AND2_X1 U13596 ( .A1(n10694), .A2(n10693), .ZN(n19668) );
  AOI22_X1 U13597 ( .A1(n10704), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20169), .B2(n19668), .ZN(n10695) );
  NAND2_X1 U13598 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13599 ( .A1(n10704), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10697) );
  NAND2_X1 U13600 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20190), .ZN(
        n19574) );
  NAND2_X1 U13601 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20199), .ZN(
        n19836) );
  NAND2_X1 U13602 ( .A1(n19574), .A2(n19836), .ZN(n19669) );
  NAND2_X1 U13603 ( .A1(n20169), .A2(n19669), .ZN(n19839) );
  NAND2_X1 U13604 ( .A1(n10697), .A2(n19839), .ZN(n10698) );
  AOI22_X1 U13605 ( .A1(n10704), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20169), .B2(n20199), .ZN(n10705) );
  NAND2_X1 U13606 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10707) );
  INV_X1 U13607 ( .A(n15655), .ZN(n10708) );
  NAND2_X1 U13608 ( .A1(n10708), .A2(n10707), .ZN(n10709) );
  INV_X1 U13609 ( .A(n10710), .ZN(n10711) );
  NAND2_X1 U13610 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  NAND2_X1 U13611 ( .A1(n10714), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10715) );
  NOR2_X1 U13612 ( .A1(n10688), .A2(n10988), .ZN(n14087) );
  NAND2_X1 U13613 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10717) );
  AND2_X2 U13614 ( .A1(n11061), .A2(n16502), .ZN(n12489) );
  AND2_X2 U13615 ( .A1(n11057), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12477) );
  AOI22_X1 U13616 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13617 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10721) );
  INV_X2 U13618 ( .A(n10416), .ZN(n12482) );
  AOI22_X1 U13619 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13620 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13621 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10731) );
  AND2_X2 U13622 ( .A1(n10889), .A2(n16502), .ZN(n12490) );
  AOI22_X1 U13623 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13624 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10728) );
  AND2_X1 U13625 ( .A1(n10724), .A2(n16502), .ZN(n10780) );
  AOI22_X1 U13626 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10727) );
  AND2_X1 U13627 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10725) );
  AND2_X1 U13628 ( .A1(n13012), .A2(n10725), .ZN(n12491) );
  AOI22_X1 U13629 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10726) );
  NAND4_X1 U13630 ( .A1(n10729), .A2(n10728), .A3(n10727), .A4(n10726), .ZN(
        n10730) );
  NOR2_X1 U13631 ( .A1(n10731), .A2(n10730), .ZN(n13343) );
  AOI22_X1 U13632 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13633 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13635 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10733) );
  NAND4_X1 U13636 ( .A1(n10736), .A2(n10735), .A3(n10734), .A4(n10733), .ZN(
        n10742) );
  AOI22_X1 U13637 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13638 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13639 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13640 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12491), .ZN(n10737) );
  NAND4_X1 U13641 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(
        n10741) );
  NOR2_X1 U13642 ( .A1(n10742), .A2(n10741), .ZN(n13372) );
  AOI22_X1 U13643 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13644 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13645 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12479), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13646 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12480), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13647 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10753) );
  AOI22_X1 U13648 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11087), .B1(
        n10747), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13649 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13650 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12490), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13651 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12491), .ZN(n10748) );
  NAND4_X1 U13652 ( .A1(n10751), .A2(n10750), .A3(n10749), .A4(n10748), .ZN(
        n10752) );
  INV_X1 U13653 ( .A(n13432), .ZN(n10775) );
  AOI22_X1 U13654 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13655 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13656 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12481), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13657 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10754) );
  NAND4_X1 U13658 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10763) );
  AOI22_X1 U13659 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13660 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13661 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13662 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12491), .ZN(n10758) );
  NAND4_X1 U13663 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10762) );
  OR2_X1 U13664 ( .A1(n10763), .A2(n10762), .ZN(n12469) );
  INV_X1 U13665 ( .A(n12469), .ZN(n13612) );
  AOI22_X1 U13666 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12416), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13667 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13668 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12479), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13669 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12480), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10764) );
  NAND4_X1 U13670 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(
        n10773) );
  AOI22_X1 U13671 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11087), .B1(
        n10747), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13672 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13673 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13674 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12491), .ZN(n10768) );
  NAND4_X1 U13675 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10772) );
  NOR2_X1 U13676 ( .A1(n10773), .A2(n10772), .ZN(n13952) );
  AOI22_X1 U13677 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13678 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10778) );
  INV_X1 U13679 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13680 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13681 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10776) );
  NAND4_X1 U13682 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10786) );
  AOI22_X1 U13683 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13684 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13685 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13686 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10781) );
  NAND4_X1 U13687 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10785) );
  NOR2_X1 U13688 ( .A1(n10786), .A2(n10785), .ZN(n13958) );
  AOI22_X1 U13689 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13690 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13691 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13692 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10787) );
  NAND4_X1 U13693 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(
        n10798) );
  AOI22_X1 U13694 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13695 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13696 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10794) );
  INV_X1 U13697 ( .A(n12488), .ZN(n12560) );
  INV_X1 U13698 ( .A(n12487), .ZN(n10813) );
  INV_X1 U13699 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13799) );
  OAI22_X1 U13700 ( .A1(n10791), .A2(n12560), .B1(n10813), .B2(n13799), .ZN(
        n10792) );
  INV_X1 U13701 ( .A(n10792), .ZN(n10793) );
  NAND4_X1 U13702 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10797) );
  OR2_X1 U13703 ( .A1(n10798), .A2(n10797), .ZN(n15087) );
  AOI22_X1 U13704 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13705 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13706 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13707 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10799) );
  NAND4_X1 U13708 ( .A1(n10802), .A2(n10801), .A3(n10800), .A4(n10799), .ZN(
        n10808) );
  AOI22_X1 U13709 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13710 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13712 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12491), .ZN(n10803) );
  NAND4_X1 U13713 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10807) );
  OR2_X1 U13714 ( .A1(n10808), .A2(n10807), .ZN(n15097) );
  INV_X1 U13715 ( .A(n15097), .ZN(n10852) );
  AOI22_X1 U13716 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13717 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13718 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13719 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10809) );
  NAND4_X1 U13720 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10820) );
  AOI22_X1 U13721 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13722 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13723 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12491), .ZN(n10816) );
  INV_X1 U13724 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13491) );
  OAI22_X1 U13725 ( .A1(n13469), .A2(n12560), .B1(n10813), .B2(n13491), .ZN(
        n10814) );
  INV_X1 U13726 ( .A(n10814), .ZN(n10815) );
  NAND4_X1 U13727 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10819) );
  OR2_X1 U13728 ( .A1(n10820), .A2(n10819), .ZN(n13991) );
  INV_X1 U13729 ( .A(n13991), .ZN(n10851) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13731 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13732 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13733 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10821) );
  NAND4_X1 U13734 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10830) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13736 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13737 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13738 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12491), .ZN(n10825) );
  NAND4_X1 U13739 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  NOR2_X1 U13740 ( .A1(n10830), .A2(n10829), .ZN(n15109) );
  AOI22_X1 U13741 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13742 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13743 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13744 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10831) );
  NAND4_X1 U13745 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n10840) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13747 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13749 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12491), .ZN(n10835) );
  NAND4_X1 U13750 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10839) );
  NOR2_X1 U13751 ( .A1(n10840), .A2(n10839), .ZN(n13940) );
  AOI22_X1 U13752 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13753 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13754 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13755 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10841) );
  NAND4_X1 U13756 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        n10850) );
  AOI22_X1 U13757 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13758 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13759 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13760 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10845) );
  NAND4_X1 U13761 ( .A1(n10848), .A2(n10847), .A3(n10846), .A4(n10845), .ZN(
        n10849) );
  NOR2_X1 U13762 ( .A1(n10850), .A2(n10849), .ZN(n13998) );
  OR2_X1 U13763 ( .A1(n13940), .A2(n13998), .ZN(n13941) );
  OR2_X1 U13764 ( .A1(n15109), .A2(n13941), .ZN(n13988) );
  NOR2_X1 U13765 ( .A1(n10852), .A2(n13989), .ZN(n15084) );
  AND2_X1 U13766 ( .A1(n15087), .A2(n15084), .ZN(n10863) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13768 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13769 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10853) );
  NAND4_X1 U13771 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10862) );
  AOI22_X1 U13772 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13773 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13774 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13775 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12491), .ZN(n10857) );
  NAND4_X1 U13776 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12477), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13778 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10864) );
  NAND4_X1 U13781 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10873) );
  AOI22_X1 U13782 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13783 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13784 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13785 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12491), .ZN(n10868) );
  NAND4_X1 U13786 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10872) );
  NOR2_X1 U13787 ( .A1(n10873), .A2(n10872), .ZN(n15077) );
  INV_X1 U13788 ( .A(n15077), .ZN(n10874) );
  AOI22_X1 U13789 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12416), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13790 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10732), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13792 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12480), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10875) );
  NAND4_X1 U13793 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10884) );
  AOI22_X1 U13794 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10747), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13795 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12488), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13797 ( .A1(n12487), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12491), .ZN(n10879) );
  NAND4_X1 U13798 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n10883) );
  INV_X1 U13799 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10888) );
  INV_X1 U13800 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10887) );
  OAI22_X1 U13801 ( .A1(n10900), .A2(n10888), .B1(n9837), .B2(n10887), .ZN(
        n10893) );
  INV_X1 U13802 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10891) );
  INV_X1 U13803 ( .A(n10889), .ZN(n11035) );
  INV_X1 U13804 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10890) );
  OAI22_X1 U13805 ( .A1(n9836), .A2(n10891), .B1(n11035), .B2(n10890), .ZN(
        n10892) );
  NOR2_X1 U13806 ( .A1(n10893), .A2(n10892), .ZN(n10897) );
  AOI22_X1 U13807 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13808 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10895) );
  XNOR2_X1 U13809 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11054) );
  NAND4_X1 U13810 ( .A1(n10897), .A2(n10896), .A3(n10895), .A4(n11054), .ZN(
        n10909) );
  INV_X1 U13811 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10899) );
  INV_X1 U13812 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10898) );
  OAI22_X1 U13813 ( .A1(n10900), .A2(n10899), .B1(n9837), .B2(n10898), .ZN(
        n10903) );
  INV_X1 U13814 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10901) );
  INV_X1 U13815 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13466) );
  OAI22_X1 U13816 ( .A1(n9836), .A2(n10901), .B1(n11035), .B2(n13466), .ZN(
        n10902) );
  NOR2_X1 U13817 ( .A1(n10903), .A2(n10902), .ZN(n10907) );
  INV_X1 U13818 ( .A(n11054), .ZN(n11062) );
  AOI22_X1 U13819 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13820 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10905) );
  NAND4_X1 U13821 ( .A1(n10907), .A2(n11062), .A3(n10906), .A4(n10905), .ZN(
        n10908) );
  AND2_X1 U13822 ( .A1(n10909), .A2(n10908), .ZN(n10935) );
  NAND2_X1 U13823 ( .A1(n9833), .A2(n10935), .ZN(n10920) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12489), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13825 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13826 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10732), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12480), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10910) );
  NAND4_X1 U13828 ( .A1(n10913), .A2(n10912), .A3(n10911), .A4(n10910), .ZN(
        n10919) );
  AOI22_X1 U13829 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11087), .B1(
        n10747), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13830 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13831 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10780), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13832 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12491), .ZN(n10914) );
  NAND4_X1 U13833 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  OR2_X1 U13834 ( .A1(n10919), .A2(n10918), .ZN(n10936) );
  XNOR2_X1 U13835 ( .A(n10920), .B(n10936), .ZN(n10940) );
  INV_X1 U13836 ( .A(n10935), .ZN(n10939) );
  NOR2_X1 U13837 ( .A1(n9833), .A2(n10939), .ZN(n15064) );
  INV_X1 U13838 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13520) );
  INV_X1 U13839 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13533) );
  OAI22_X1 U13840 ( .A1(n10900), .A2(n13520), .B1(n9837), .B2(n13533), .ZN(
        n10924) );
  INV_X1 U13841 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13530) );
  OAI22_X1 U13842 ( .A1(n9836), .A2(n10590), .B1(n11035), .B2(n13530), .ZN(
        n10923) );
  NOR2_X1 U13843 ( .A1(n10924), .A2(n10923), .ZN(n10927) );
  AOI22_X1 U13844 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13845 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10925) );
  NAND4_X1 U13846 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n11054), .ZN(
        n10934) );
  INV_X1 U13847 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13516) );
  INV_X1 U13848 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13514) );
  OAI22_X1 U13849 ( .A1(n10900), .A2(n13516), .B1(n9837), .B2(n13514), .ZN(
        n10929) );
  INV_X1 U13850 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13527) );
  INV_X1 U13851 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13532) );
  OAI22_X1 U13852 ( .A1(n9836), .A2(n13527), .B1(n11035), .B2(n13532), .ZN(
        n10928) );
  NOR2_X1 U13853 ( .A1(n10929), .A2(n10928), .ZN(n10932) );
  AOI22_X1 U13854 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13855 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10930) );
  NAND4_X1 U13856 ( .A1(n10932), .A2(n11062), .A3(n10931), .A4(n10930), .ZN(
        n10933) );
  NAND2_X1 U13857 ( .A1(n10934), .A2(n10933), .ZN(n10942) );
  NAND2_X1 U13858 ( .A1(n10936), .A2(n10935), .ZN(n10943) );
  XOR2_X1 U13859 ( .A(n10942), .B(n10943), .Z(n10937) );
  NAND2_X1 U13860 ( .A1(n10937), .A2(n11008), .ZN(n15055) );
  INV_X1 U13861 ( .A(n10942), .ZN(n10938) );
  NAND2_X1 U13862 ( .A1(n9839), .A2(n10938), .ZN(n15058) );
  NOR2_X1 U13863 ( .A1(n15058), .A2(n10939), .ZN(n10941) );
  NOR2_X1 U13864 ( .A1(n10943), .A2(n10942), .ZN(n10964) );
  INV_X1 U13865 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10944) );
  OAI22_X1 U13866 ( .A1(n10900), .A2(n10945), .B1(n9837), .B2(n10944), .ZN(
        n10949) );
  INV_X1 U13867 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10947) );
  OAI22_X1 U13868 ( .A1(n9836), .A2(n10947), .B1(n11035), .B2(n10946), .ZN(
        n10948) );
  NOR2_X1 U13869 ( .A1(n10949), .A2(n10948), .ZN(n10952) );
  AOI22_X1 U13870 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13871 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10950) );
  NAND4_X1 U13872 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n11054), .ZN(
        n10963) );
  INV_X1 U13873 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10953) );
  OAI22_X1 U13874 ( .A1(n10900), .A2(n10954), .B1(n9837), .B2(n10953), .ZN(
        n10958) );
  INV_X1 U13875 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10956) );
  OAI22_X1 U13876 ( .A1(n9836), .A2(n10956), .B1(n11035), .B2(n10955), .ZN(
        n10957) );
  NOR2_X1 U13877 ( .A1(n10958), .A2(n10957), .ZN(n10961) );
  AOI22_X1 U13878 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13879 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10959) );
  NAND4_X1 U13880 ( .A1(n10961), .A2(n11062), .A3(n10960), .A4(n10959), .ZN(
        n10962) );
  AND2_X1 U13881 ( .A1(n10963), .A2(n10962), .ZN(n10966) );
  NAND2_X1 U13882 ( .A1(n10964), .A2(n10966), .ZN(n10982) );
  OAI211_X1 U13883 ( .C1(n10964), .C2(n10966), .A(n11008), .B(n10982), .ZN(
        n10968) );
  INV_X1 U13884 ( .A(n10968), .ZN(n10965) );
  INV_X1 U13885 ( .A(n10966), .ZN(n10967) );
  NOR2_X1 U13886 ( .A1(n9833), .A2(n10967), .ZN(n15048) );
  OAI22_X1 U13887 ( .A1(n10900), .A2(n13469), .B1(n9837), .B2(n13491), .ZN(
        n10971) );
  INV_X1 U13888 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13503) );
  OAI22_X1 U13889 ( .A1(n9836), .A2(n13503), .B1(n11035), .B2(n13498), .ZN(
        n10970) );
  NOR2_X1 U13890 ( .A1(n10971), .A2(n10970), .ZN(n10974) );
  AOI22_X1 U13891 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13892 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U13893 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n11054), .ZN(
        n10981) );
  INV_X1 U13894 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13472) );
  OAI22_X1 U13895 ( .A1(n10900), .A2(n13478), .B1(n9837), .B2(n13472), .ZN(
        n10976) );
  INV_X1 U13896 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13484) );
  OAI22_X1 U13897 ( .A1(n9836), .A2(n13484), .B1(n11035), .B2(n13487), .ZN(
        n10975) );
  NOR2_X1 U13898 ( .A1(n10976), .A2(n10975), .ZN(n10979) );
  AOI22_X1 U13899 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13900 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10977) );
  NAND4_X1 U13901 ( .A1(n10979), .A2(n11062), .A3(n10978), .A4(n10977), .ZN(
        n10980) );
  NAND2_X1 U13902 ( .A1(n10981), .A2(n10980), .ZN(n10984) );
  NAND2_X1 U13903 ( .A1(n10982), .A2(n10984), .ZN(n10983) );
  XNOR2_X2 U13904 ( .A(n10986), .B(n10418), .ZN(n15044) );
  INV_X1 U13905 ( .A(n10984), .ZN(n10985) );
  NAND2_X1 U13906 ( .A1(n9839), .A2(n10985), .ZN(n15043) );
  INV_X1 U13907 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10987) );
  OAI22_X1 U13908 ( .A1(n10900), .A2(n10988), .B1(n9837), .B2(n10987), .ZN(
        n10992) );
  INV_X1 U13909 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10990) );
  OAI22_X1 U13910 ( .A1(n9836), .A2(n10990), .B1(n11035), .B2(n10989), .ZN(
        n10991) );
  NOR2_X1 U13911 ( .A1(n10992), .A2(n10991), .ZN(n10995) );
  AOI22_X1 U13912 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13913 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U13914 ( .A1(n10995), .A2(n10994), .A3(n10993), .A4(n11054), .ZN(
        n11006) );
  INV_X1 U13915 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10996) );
  OAI22_X1 U13916 ( .A1(n10900), .A2(n10997), .B1(n9837), .B2(n10996), .ZN(
        n11001) );
  INV_X1 U13917 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10999) );
  OAI22_X1 U13918 ( .A1(n9836), .A2(n10999), .B1(n11035), .B2(n10998), .ZN(
        n11000) );
  NOR2_X1 U13919 ( .A1(n11001), .A2(n11000), .ZN(n11004) );
  AOI22_X1 U13920 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U13921 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11002) );
  NAND4_X1 U13922 ( .A1(n11004), .A2(n11062), .A3(n11003), .A4(n11002), .ZN(
        n11005) );
  NAND2_X1 U13923 ( .A1(n11006), .A2(n11005), .ZN(n11012) );
  INV_X1 U13924 ( .A(n11012), .ZN(n11010) );
  INV_X1 U13925 ( .A(n11007), .ZN(n11009) );
  OR2_X1 U13926 ( .A1(n11007), .A2(n11012), .ZN(n11045) );
  OAI211_X1 U13927 ( .C1(n11010), .C2(n11009), .A(n11045), .B(n11008), .ZN(
        n11011) );
  NOR2_X1 U13928 ( .A1(n9833), .A2(n11012), .ZN(n15033) );
  NAND2_X1 U13929 ( .A1(n15034), .A2(n15033), .ZN(n15032) );
  INV_X1 U13930 ( .A(n15026), .ZN(n11026) );
  OAI22_X1 U13931 ( .A1(n10900), .A2(n10791), .B1(n9837), .B2(n13799), .ZN(
        n11014) );
  INV_X1 U13932 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13806) );
  INV_X1 U13933 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13785) );
  OAI22_X1 U13934 ( .A1(n9836), .A2(n13806), .B1(n11035), .B2(n13785), .ZN(
        n11013) );
  NOR2_X1 U13935 ( .A1(n11014), .A2(n11013), .ZN(n11017) );
  AOI22_X1 U13936 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U13937 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11015) );
  NAND4_X1 U13938 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11054), .ZN(
        n11025) );
  INV_X1 U13939 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13789) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13797) );
  OAI22_X1 U13941 ( .A1(n10900), .A2(n13789), .B1(n9837), .B2(n13797), .ZN(
        n11019) );
  INV_X1 U13942 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13803) );
  INV_X1 U13943 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13792) );
  OAI22_X1 U13944 ( .A1(n9836), .A2(n13803), .B1(n11035), .B2(n13792), .ZN(
        n11018) );
  NOR2_X1 U13945 ( .A1(n11019), .A2(n11018), .ZN(n11023) );
  AOI22_X1 U13946 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15672), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U13947 ( .A1(n10904), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11021) );
  NAND4_X1 U13948 ( .A1(n11023), .A2(n11062), .A3(n11022), .A4(n11021), .ZN(
        n11024) );
  NAND2_X1 U13949 ( .A1(n11025), .A2(n11024), .ZN(n11046) );
  OAI22_X1 U13950 ( .A1(n10900), .A2(n13844), .B1(n11027), .B2(n13837), .ZN(
        n11031) );
  INV_X1 U13951 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11029) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13834) );
  OAI22_X1 U13953 ( .A1(n11029), .A2(n11028), .B1(n9895), .B2(n13834), .ZN(
        n11030) );
  NOR2_X1 U13954 ( .A1(n11031), .A2(n11030), .ZN(n11034) );
  AOI22_X1 U13955 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11032) );
  NAND4_X1 U13956 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11054), .ZN(
        n11044) );
  OAI22_X1 U13957 ( .A1(n10900), .A2(n13840), .B1(n11035), .B2(n13831), .ZN(
        n11039) );
  INV_X1 U13958 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13839) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13833) );
  OAI22_X1 U13960 ( .A1(n9836), .A2(n13839), .B1(n9837), .B2(n13833), .ZN(
        n11038) );
  NOR2_X1 U13961 ( .A1(n11039), .A2(n11038), .ZN(n11042) );
  AOI22_X1 U13962 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U13963 ( .A1(n15672), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U13964 ( .A1(n11042), .A2(n11062), .A3(n11041), .A4(n11040), .ZN(
        n11043) );
  NAND2_X1 U13965 ( .A1(n11044), .A2(n11043), .ZN(n11049) );
  INV_X1 U13966 ( .A(n11045), .ZN(n15025) );
  INV_X1 U13967 ( .A(n11046), .ZN(n15027) );
  AND2_X1 U13968 ( .A1(n9833), .A2(n15027), .ZN(n11047) );
  NAND2_X1 U13969 ( .A1(n15025), .A2(n11047), .ZN(n11048) );
  NOR2_X1 U13970 ( .A1(n11048), .A2(n11049), .ZN(n11050) );
  AOI21_X1 U13971 ( .B1(n11049), .B2(n11048), .A(n11050), .ZN(n15020) );
  INV_X1 U13972 ( .A(n11050), .ZN(n11051) );
  AOI22_X1 U13973 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U13974 ( .A1(n15672), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9834), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U13975 ( .A1(n11053), .A2(n11052), .ZN(n11068) );
  AOI22_X1 U13976 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11056) );
  NAND3_X1 U13977 ( .A1(n11056), .A2(n11055), .A3(n11054), .ZN(n11067) );
  AOI22_X1 U13978 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10904), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13979 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11058), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11059) );
  NAND2_X1 U13980 ( .A1(n11060), .A2(n11059), .ZN(n11066) );
  AOI22_X1 U13981 ( .A1(n11061), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10724), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11064) );
  NAND3_X1 U13982 ( .A1(n11064), .A2(n11063), .A3(n11062), .ZN(n11065) );
  OAI22_X1 U13983 ( .A1(n11068), .A2(n11067), .B1(n11066), .B2(n11065), .ZN(
        n11069) );
  NAND2_X1 U13984 ( .A1(n20222), .A2(n9833), .ZN(n11074) );
  MUX2_X1 U13985 ( .A(n20190), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12583) );
  INV_X1 U13986 ( .A(n11075), .ZN(n11071) );
  NAND2_X1 U13987 ( .A1(n11072), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11094) );
  OAI21_X1 U13988 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n11072), .A(
        n11094), .ZN(n11073) );
  XNOR2_X1 U13989 ( .A(n11093), .B(n11073), .ZN(n12389) );
  MUX2_X1 U13990 ( .A(n12581), .B(n11074), .S(n12389), .Z(n11082) );
  OAI21_X1 U13991 ( .B1(n20199), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11075), .ZN(n12559) );
  INV_X1 U13992 ( .A(n12559), .ZN(n12582) );
  XNOR2_X1 U13993 ( .A(n12583), .B(n11075), .ZN(n12371) );
  OAI21_X1 U13994 ( .B1(n9833), .B2(n12582), .A(n12371), .ZN(n11076) );
  OAI21_X1 U13995 ( .B1(n12389), .B2(n9833), .A(n11076), .ZN(n11077) );
  NAND2_X1 U13996 ( .A1(n11077), .A2(n16528), .ZN(n11080) );
  NAND2_X1 U13997 ( .A1(n12582), .A2(n12583), .ZN(n11078) );
  NAND2_X1 U13998 ( .A1(n12624), .A2(n11078), .ZN(n11079) );
  NAND2_X1 U13999 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  AOI22_X1 U14000 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12489), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14001 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14002 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12481), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14003 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10732), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U14004 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11091) );
  AOI22_X1 U14005 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14006 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14007 ( .A1(n11087), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12491), .ZN(n11088) );
  NAND2_X1 U14008 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20181), .ZN(
        n11092) );
  NAND2_X1 U14009 ( .A1(n11093), .A2(n11092), .ZN(n11095) );
  NAND2_X1 U14010 ( .A1(n11095), .A2(n11094), .ZN(n11097) );
  MUX2_X1 U14011 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n10685), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11096) );
  OAI22_X1 U14012 ( .A1(n11097), .A2(n11096), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16502), .ZN(n11100) );
  XNOR2_X1 U14013 ( .A(n11097), .B(n11096), .ZN(n12369) );
  INV_X1 U14014 ( .A(n12369), .ZN(n12414) );
  NAND2_X1 U14015 ( .A1(n12587), .A2(n12414), .ZN(n11104) );
  NAND3_X1 U14016 ( .A1(n11105), .A2(n12368), .A3(n12414), .ZN(n11098) );
  NAND2_X1 U14017 ( .A1(n11098), .A2(n12624), .ZN(n11103) );
  AND2_X1 U14018 ( .A1(n16517), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11099) );
  OR2_X1 U14019 ( .A1(n11100), .A2(n11099), .ZN(n11102) );
  INV_X1 U14020 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15748) );
  NAND2_X1 U14021 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15748), .ZN(
        n11101) );
  OAI211_X1 U14022 ( .C1(n11105), .C2(n11104), .A(n11103), .B(n12589), .ZN(
        n11106) );
  MUX2_X1 U14023 ( .A(n11106), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20218), .Z(n12597) );
  INV_X1 U14024 ( .A(n13028), .ZN(n16534) );
  INV_X1 U14025 ( .A(n11109), .ZN(n11110) );
  AND2_X1 U14026 ( .A1(n11108), .A2(n11110), .ZN(n13018) );
  INV_X1 U14027 ( .A(n11111), .ZN(n13014) );
  NAND2_X1 U14028 ( .A1(n20079), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20078) );
  AOI21_X4 U14029 ( .B1(n13025), .B2(n13014), .A(n19106), .ZN(n15104) );
  NAND2_X1 U14030 ( .A1(n15117), .A2(n15110), .ZN(n11207) );
  INV_X1 U14031 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15549) );
  OR2_X1 U14032 ( .A1(n14232), .A2(n15549), .ZN(n11118) );
  INV_X1 U14033 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U14034 ( .A1(n14227), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11115) );
  NAND2_X1 U14035 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11114) );
  OAI211_X1 U14036 ( .C1(n11196), .C2(n14125), .A(n11115), .B(n11114), .ZN(
        n11116) );
  INV_X1 U14037 ( .A(n11116), .ZN(n11117) );
  INV_X1 U14038 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11119) );
  OR2_X1 U14039 ( .A1(n14232), .A2(n11119), .ZN(n11125) );
  INV_X1 U14040 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U14041 ( .A1(n14227), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14042 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11120) );
  OAI211_X1 U14043 ( .C1(n11196), .C2(n11122), .A(n11121), .B(n11120), .ZN(
        n11123) );
  INV_X1 U14044 ( .A(n11123), .ZN(n11124) );
  NAND2_X1 U14045 ( .A1(n11125), .A2(n11124), .ZN(n12547) );
  INV_X1 U14046 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16470) );
  AOI22_X1 U14047 ( .A1(n14227), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14048 ( .A1(n14228), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11126) );
  OAI211_X1 U14049 ( .C1(n14232), .C2(n16470), .A(n11127), .B(n11126), .ZN(
        n11128) );
  INV_X1 U14050 ( .A(n11128), .ZN(n13342) );
  NAND2_X1 U14051 ( .A1(n11133), .A2(n11132), .ZN(n11135) );
  NAND2_X1 U14052 ( .A1(n11135), .A2(n11134), .ZN(n11140) );
  INV_X1 U14053 ( .A(n11136), .ZN(n11138) );
  NAND2_X1 U14054 ( .A1(n11138), .A2(n11137), .ZN(n11139) );
  INV_X1 U14055 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16480) );
  OR2_X1 U14056 ( .A1(n14232), .A2(n16480), .ZN(n11145) );
  INV_X1 U14057 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U14058 ( .A1(n14227), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11142) );
  NAND2_X1 U14059 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11141) );
  OAI211_X1 U14060 ( .C1(n11196), .C2(n14094), .A(n11142), .B(n11141), .ZN(
        n11143) );
  INV_X1 U14061 ( .A(n11143), .ZN(n11144) );
  INV_X1 U14062 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U14063 ( .A1(n14227), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14064 ( .A1(n14228), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11146) );
  OAI211_X1 U14065 ( .C1(n14232), .C2(n16497), .A(n11147), .B(n11146), .ZN(
        n14083) );
  NAND2_X1 U14066 ( .A1(n14082), .A2(n14083), .ZN(n14081) );
  INV_X1 U14067 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U14068 ( .A1(n14227), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11149) );
  NAND2_X1 U14069 ( .A1(n14228), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11148) );
  OAI211_X1 U14070 ( .C1(n14232), .C2(n13890), .A(n11149), .B(n11148), .ZN(
        n11150) );
  INV_X1 U14071 ( .A(n11150), .ZN(n13094) );
  NOR2_X2 U14072 ( .A1(n14081), .A2(n13094), .ZN(n13368) );
  INV_X1 U14073 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12458) );
  INV_X1 U14074 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13927) );
  OR2_X1 U14075 ( .A1(n14232), .A2(n13927), .ZN(n11152) );
  AOI22_X1 U14076 ( .A1(n14227), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11151) );
  OAI211_X1 U14077 ( .C1(n11196), .C2(n12458), .A(n11152), .B(n11151), .ZN(
        n13369) );
  INV_X1 U14078 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15643) );
  OR2_X1 U14079 ( .A1(n14232), .A2(n15643), .ZN(n11154) );
  AOI22_X1 U14080 ( .A1(n14227), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11153) );
  OAI211_X1 U14081 ( .C1(n10207), .C2(n11196), .A(n11154), .B(n11153), .ZN(
        n13375) );
  INV_X1 U14082 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U14083 ( .A1(n14227), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11156) );
  NAND2_X1 U14084 ( .A1(n14228), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11155) );
  OAI211_X1 U14085 ( .C1(n14232), .C2(n15622), .A(n11156), .B(n11155), .ZN(
        n11157) );
  INV_X1 U14086 ( .A(n11157), .ZN(n13437) );
  INV_X1 U14087 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11160) );
  INV_X1 U14088 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15589) );
  OR2_X1 U14089 ( .A1(n14232), .A2(n15589), .ZN(n11159) );
  AOI22_X1 U14090 ( .A1(n14227), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11158) );
  OAI211_X1 U14091 ( .C1(n11160), .C2(n11196), .A(n11159), .B(n11158), .ZN(
        n13609) );
  INV_X1 U14092 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14121) );
  INV_X1 U14093 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15590) );
  OR2_X1 U14094 ( .A1(n14232), .A2(n15590), .ZN(n11162) );
  AOI22_X1 U14095 ( .A1(n14227), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11161) );
  OAI211_X1 U14096 ( .C1(n14121), .C2(n11196), .A(n11162), .B(n11161), .ZN(
        n13654) );
  INV_X1 U14097 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15563) );
  OR2_X1 U14098 ( .A1(n14232), .A2(n15563), .ZN(n11168) );
  INV_X1 U14099 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14100 ( .A1(n14227), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U14101 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11163) );
  OAI211_X1 U14102 ( .C1(n11196), .C2(n11165), .A(n11164), .B(n11163), .ZN(
        n11166) );
  INV_X1 U14103 ( .A(n11166), .ZN(n11167) );
  INV_X1 U14104 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14145) );
  INV_X1 U14105 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15529) );
  OR2_X1 U14106 ( .A1(n14232), .A2(n15529), .ZN(n11170) );
  AOI22_X1 U14107 ( .A1(n14227), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11169) );
  OAI211_X1 U14108 ( .C1(n11196), .C2(n14145), .A(n11170), .B(n11169), .ZN(
        n14008) );
  INV_X1 U14109 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n14155) );
  INV_X1 U14110 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14160) );
  OR2_X1 U14111 ( .A1(n14232), .A2(n14160), .ZN(n11172) );
  AOI22_X1 U14112 ( .A1(n14227), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11171) );
  OAI211_X1 U14113 ( .C1(n11196), .C2(n14155), .A(n11172), .B(n11171), .ZN(
        n13983) );
  INV_X1 U14114 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11175) );
  INV_X1 U14115 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14137) );
  OR2_X1 U14116 ( .A1(n14232), .A2(n14137), .ZN(n11174) );
  AOI22_X1 U14117 ( .A1(n14227), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11173) );
  OAI211_X1 U14118 ( .C1(n11196), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n15111) );
  INV_X1 U14119 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n14138) );
  INV_X1 U14120 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15478) );
  OR2_X1 U14121 ( .A1(n14232), .A2(n15478), .ZN(n11177) );
  AOI22_X1 U14122 ( .A1(n14227), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11176) );
  OAI211_X1 U14123 ( .C1(n11196), .C2(n14138), .A(n11177), .B(n11176), .ZN(
        n13993) );
  INV_X1 U14124 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14129) );
  INV_X1 U14125 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15479) );
  OR2_X1 U14126 ( .A1(n14232), .A2(n15479), .ZN(n11179) );
  AOI22_X1 U14127 ( .A1(n14227), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11178) );
  OAI211_X1 U14128 ( .C1(n11196), .C2(n14129), .A(n11179), .B(n11178), .ZN(
        n15099) );
  INV_X1 U14129 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14130) );
  INV_X1 U14130 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15465) );
  OR2_X1 U14131 ( .A1(n14232), .A2(n15465), .ZN(n11181) );
  AOI22_X1 U14132 ( .A1(n14227), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11180) );
  OAI211_X1 U14133 ( .C1(n11196), .C2(n14130), .A(n11181), .B(n11180), .ZN(
        n15089) );
  INV_X1 U14134 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n14180) );
  INV_X1 U14135 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15458) );
  OR2_X1 U14136 ( .A1(n14232), .A2(n15458), .ZN(n11183) );
  AOI22_X1 U14137 ( .A1(n14227), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11182) );
  OAI211_X1 U14138 ( .C1(n11196), .C2(n14180), .A(n11183), .B(n11182), .ZN(
        n15078) );
  INV_X1 U14139 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15074) );
  INV_X1 U14140 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15437) );
  OR2_X1 U14141 ( .A1(n14232), .A2(n15437), .ZN(n11185) );
  AOI22_X1 U14142 ( .A1(n14227), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11184) );
  OAI211_X1 U14143 ( .C1(n11196), .C2(n15074), .A(n11185), .B(n11184), .ZN(
        n15068) );
  INV_X1 U14144 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15278) );
  OR2_X1 U14145 ( .A1(n14232), .A2(n15278), .ZN(n11187) );
  AOI22_X1 U14146 ( .A1(n14227), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11186) );
  OAI211_X1 U14147 ( .C1(n11196), .C2(n10208), .A(n11187), .B(n11186), .ZN(
        n15059) );
  INV_X1 U14148 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11190) );
  INV_X1 U14149 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14199) );
  OR2_X1 U14150 ( .A1(n14232), .A2(n14199), .ZN(n11189) );
  AOI22_X1 U14151 ( .A1(n14227), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11188) );
  OAI211_X1 U14152 ( .C1(n11196), .C2(n11190), .A(n11189), .B(n11188), .ZN(
        n15050) );
  INV_X1 U14153 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16310) );
  INV_X1 U14154 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15255) );
  OR2_X1 U14155 ( .A1(n14232), .A2(n15255), .ZN(n11192) );
  AOI22_X1 U14156 ( .A1(n14227), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11191) );
  OAI211_X1 U14157 ( .C1(n11196), .C2(n16310), .A(n11192), .B(n11191), .ZN(
        n15039) );
  INV_X1 U14158 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11195) );
  INV_X1 U14159 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14392) );
  OR2_X1 U14160 ( .A1(n14232), .A2(n14392), .ZN(n11194) );
  AOI22_X1 U14161 ( .A1(n14227), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11193) );
  OAI211_X1 U14162 ( .C1(n11196), .C2(n11195), .A(n11194), .B(n11193), .ZN(
        n15036) );
  INV_X1 U14163 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11199) );
  INV_X1 U14164 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15381) );
  OR2_X1 U14165 ( .A1(n14232), .A2(n15381), .ZN(n11198) );
  AOI22_X1 U14166 ( .A1(n14227), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11197) );
  OAI211_X1 U14167 ( .C1(n11196), .C2(n11199), .A(n11198), .B(n11197), .ZN(
        n14256) );
  INV_X1 U14168 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U14169 ( .A1(n14227), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11201) );
  NAND2_X1 U14170 ( .A1(n14228), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11200) );
  OAI211_X1 U14171 ( .C1(n14232), .C2(n15382), .A(n11201), .B(n11200), .ZN(
        n15018) );
  INV_X1 U14172 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14207) );
  INV_X1 U14173 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15367) );
  OR2_X1 U14174 ( .A1(n14232), .A2(n15367), .ZN(n11203) );
  AOI22_X1 U14175 ( .A1(n14227), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11202) );
  OAI211_X1 U14176 ( .C1(n11196), .C2(n14207), .A(n11203), .B(n11202), .ZN(
        n14226) );
  XNOR2_X1 U14177 ( .A(n15017), .B(n14226), .ZN(n16269) );
  INV_X1 U14178 ( .A(n16269), .ZN(n15370) );
  NAND2_X1 U14179 ( .A1(n9831), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11204) );
  OAI21_X1 U14180 ( .B1(n15370), .B2(n9831), .A(n11204), .ZN(n11205) );
  INV_X1 U14181 ( .A(n11205), .ZN(n11206) );
  NAND2_X1 U14182 ( .A1(n11207), .A2(n11206), .ZN(P2_U2857) );
  NAND2_X1 U14183 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11213) );
  AND2_X2 U14184 ( .A1(n11209), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13292) );
  AND2_X4 U14185 ( .A1(n11227), .A2(n13292), .ZN(n12166) );
  NAND2_X1 U14186 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11212) );
  NOR2_X4 U14187 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14971) );
  NAND2_X1 U14188 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11211) );
  NAND2_X1 U14189 ( .A1(n9823), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11210) );
  NAND4_X1 U14190 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11216) );
  AND2_X2 U14191 ( .A1(n13295), .A2(n14971), .ZN(n11427) );
  NAND2_X1 U14192 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14193 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14194 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11218) );
  NAND2_X1 U14195 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11217) );
  AND2_X2 U14196 ( .A1(n13292), .A2(n14971), .ZN(n11308) );
  NAND2_X1 U14197 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11225) );
  INV_X2 U14198 ( .A(n12128), .ZN(n11928) );
  NAND2_X1 U14199 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14200 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14201 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14202 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11229) );
  AND2_X4 U14203 ( .A1(n13295), .A2(n11227), .ZN(n11494) );
  NAND2_X1 U14204 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11228) );
  OAI211_X1 U14205 ( .C1(n12163), .C2(n11230), .A(n11229), .B(n11228), .ZN(
        n11231) );
  INV_X1 U14206 ( .A(n11231), .ZN(n11232) );
  INV_X1 U14207 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U14208 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U14209 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11236) );
  OAI211_X1 U14210 ( .C1(n12163), .C2(n11238), .A(n11237), .B(n11236), .ZN(
        n11239) );
  INV_X1 U14211 ( .A(n11239), .ZN(n11243) );
  AOI22_X1 U14212 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14213 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11241) );
  INV_X2 U14214 ( .A(n11938), .ZN(n11444) );
  NAND2_X1 U14215 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11240) );
  AOI22_X1 U14216 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14217 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14218 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14219 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14220 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U14221 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11252) );
  INV_X1 U14222 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U14223 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11249) );
  NAND2_X1 U14224 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11248) );
  OAI211_X1 U14225 ( .C1(n12163), .C2(n12127), .A(n11249), .B(n11248), .ZN(
        n11250) );
  INV_X1 U14226 ( .A(n11250), .ZN(n11251) );
  AOI22_X1 U14227 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14228 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14229 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14230 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11258) );
  AND3_X2 U14231 ( .A1(n10415), .A2(n11259), .A3(n11258), .ZN(n11576) );
  INV_X1 U14232 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14233 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11261) );
  NAND2_X1 U14234 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11260) );
  OAI211_X1 U14235 ( .C1(n12163), .C2(n11262), .A(n11261), .B(n11260), .ZN(
        n11263) );
  INV_X1 U14236 ( .A(n11263), .ZN(n11267) );
  AOI22_X1 U14237 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14238 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U14239 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11264) );
  NAND4_X1 U14240 ( .A1(n11267), .A2(n11266), .A3(n11265), .A4(n11264), .ZN(
        n11274) );
  INV_X2 U14241 ( .A(n12018), .ZN(n12165) );
  AOI22_X1 U14242 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14243 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11271) );
  INV_X2 U14244 ( .A(n11268), .ZN(n12105) );
  AOI22_X1 U14245 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14246 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U14247 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11273) );
  INV_X1 U14248 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11277) );
  NAND2_X1 U14249 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14250 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11275) );
  OAI211_X1 U14251 ( .C1(n12163), .C2(n11277), .A(n11276), .B(n11275), .ZN(
        n11278) );
  INV_X1 U14252 ( .A(n11278), .ZN(n11282) );
  AOI22_X1 U14253 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14254 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11280) );
  NAND2_X1 U14255 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11279) );
  NAND4_X1 U14256 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11288) );
  AOI22_X1 U14257 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14258 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14259 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14260 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11283) );
  NAND4_X1 U14261 ( .A1(n11286), .A2(n11285), .A3(n11284), .A4(n11283), .ZN(
        n11287) );
  NAND2_X1 U14262 ( .A1(n11354), .A2(n11576), .ZN(n11351) );
  INV_X1 U14263 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U14264 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14265 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11289) );
  OAI211_X1 U14266 ( .C1(n11729), .C2(n11950), .A(n11290), .B(n11289), .ZN(
        n11291) );
  INV_X1 U14267 ( .A(n11291), .ZN(n11295) );
  AOI22_X1 U14268 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14269 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U14270 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11292) );
  NAND4_X1 U14271 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11301) );
  AOI22_X1 U14272 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11401), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14273 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14274 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14275 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11296) );
  NAND4_X1 U14276 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n11300) );
  OR2_X2 U14277 ( .A1(n11301), .A2(n11300), .ZN(n20478) );
  NAND2_X1 U14278 ( .A1(n11351), .A2(n20478), .ZN(n11359) );
  NAND2_X1 U14279 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U14280 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14281 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11305) );
  NAND2_X1 U14282 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14283 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11312) );
  NAND2_X1 U14284 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14285 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14286 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11309) );
  NAND4_X1 U14287 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n11314) );
  NAND2_X1 U14288 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U14289 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11317) );
  NAND2_X1 U14290 ( .A1(n9823), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14291 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11315) );
  NAND2_X1 U14292 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U14293 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11320) );
  OAI211_X1 U14294 ( .C1(n13298), .C2(n11966), .A(n11321), .B(n11320), .ZN(
        n11322) );
  INV_X1 U14295 ( .A(n11322), .ZN(n11323) );
  NAND3_X4 U14296 ( .A1(n11326), .A2(n11325), .A3(n9882), .ZN(n20423) );
  INV_X1 U14297 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11327) );
  NAND2_X1 U14298 ( .A1(n11401), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14299 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14300 ( .A1(n9823), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11328) );
  NAND4_X1 U14301 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11334) );
  NAND2_X1 U14302 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14303 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14304 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14305 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14306 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14307 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14308 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11340) );
  NAND2_X1 U14309 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11339) );
  INV_X1 U14310 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11345) );
  NAND2_X1 U14311 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14312 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11343) );
  OAI211_X1 U14313 ( .C1(n12163), .C2(n11345), .A(n11344), .B(n11343), .ZN(
        n11346) );
  INV_X1 U14314 ( .A(n11346), .ZN(n11347) );
  NAND4_X4 U14315 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n20440) );
  NAND2_X1 U14316 ( .A1(n12642), .A2(n12868), .ZN(n12887) );
  NAND2_X1 U14317 ( .A1(n12965), .A2(n20452), .ZN(n12737) );
  INV_X1 U14318 ( .A(n11351), .ZN(n11352) );
  NAND2_X1 U14319 ( .A1(n12904), .A2(n12254), .ZN(n11353) );
  NAND2_X1 U14320 ( .A1(n12887), .A2(n11353), .ZN(n12942) );
  XNOR2_X1 U14321 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12733) );
  NOR2_X2 U14322 ( .A1(n20452), .A2(n20446), .ZN(n12892) );
  AND2_X4 U14323 ( .A1(n20452), .A2(n20440), .ZN(n14343) );
  NAND2_X1 U14324 ( .A1(n12806), .A2(n14343), .ZN(n12949) );
  NAND2_X1 U14325 ( .A1(n20423), .A2(n20446), .ZN(n12877) );
  OAI211_X1 U14326 ( .C1(n11354), .C2(n21104), .A(n12949), .B(n12877), .ZN(
        n11375) );
  INV_X1 U14327 ( .A(n20452), .ZN(n11355) );
  OAI21_X1 U14328 ( .B1(n12872), .B2(n12892), .A(n13394), .ZN(n11363) );
  NAND2_X1 U14329 ( .A1(n12806), .A2(n11576), .ZN(n11358) );
  NAND2_X1 U14330 ( .A1(n12218), .A2(n20471), .ZN(n11357) );
  AND2_X1 U14331 ( .A1(n11357), .A2(n20478), .ZN(n11373) );
  NAND2_X1 U14332 ( .A1(n12879), .A2(n11354), .ZN(n12876) );
  INV_X1 U14333 ( .A(n11359), .ZN(n11361) );
  NAND2_X1 U14334 ( .A1(n12876), .A2(n14368), .ZN(n11362) );
  NAND2_X1 U14335 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11386) );
  OAI21_X1 U14336 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11386), .ZN(n20768) );
  OR2_X1 U14337 ( .A1(n15976), .A2(n20839), .ZN(n11379) );
  OAI21_X1 U14338 ( .B1(n12795), .B2(n20768), .A(n11379), .ZN(n11364) );
  INV_X1 U14339 ( .A(n11364), .ZN(n11365) );
  MUX2_X1 U14340 ( .A(n15976), .B(n12795), .S(n20889), .Z(n11368) );
  INV_X1 U14341 ( .A(n11369), .ZN(n11370) );
  OAI21_X1 U14342 ( .B1(n13400), .B2(n11370), .A(n12872), .ZN(n11378) );
  INV_X1 U14343 ( .A(n16242), .ZN(n14987) );
  NOR2_X1 U14344 ( .A1(n14987), .A2(n21026), .ZN(n11371) );
  AND2_X1 U14345 ( .A1(n13403), .A2(n11371), .ZN(n11372) );
  NAND2_X1 U14346 ( .A1(n12892), .A2(n11576), .ZN(n12947) );
  OAI211_X1 U14347 ( .C1(n11373), .C2(n21104), .A(n11372), .B(n12947), .ZN(
        n11374) );
  NOR2_X1 U14348 ( .A1(n11375), .A2(n11374), .ZN(n11377) );
  NAND3_X1 U14349 ( .A1(n12876), .A2(n20440), .A3(n14368), .ZN(n11376) );
  NAND3_X1 U14350 ( .A1(n11378), .A2(n11377), .A3(n11376), .ZN(n11436) );
  INV_X1 U14351 ( .A(n11379), .ZN(n11382) );
  INV_X1 U14352 ( .A(n11380), .ZN(n11381) );
  OAI21_X1 U14353 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11382), .A(
        n11381), .ZN(n11383) );
  INV_X1 U14354 ( .A(n12795), .ZN(n11388) );
  INV_X1 U14355 ( .A(n11386), .ZN(n11385) );
  NAND2_X1 U14356 ( .A1(n11385), .A2(n20764), .ZN(n20805) );
  NAND2_X1 U14357 ( .A1(n11386), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U14358 ( .A1(n20805), .A2(n11387), .ZN(n20433) );
  NAND2_X1 U14359 ( .A1(n11388), .A2(n20433), .ZN(n11389) );
  INV_X1 U14360 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14361 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11393) );
  NAND2_X1 U14362 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11392) );
  OAI211_X1 U14363 ( .C1(n11729), .C2(n11409), .A(n11393), .B(n11392), .ZN(
        n11394) );
  INV_X1 U14364 ( .A(n11394), .ZN(n11398) );
  AOI22_X1 U14365 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14366 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11396) );
  NAND2_X1 U14367 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11395) );
  NAND4_X1 U14368 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11408) );
  INV_X1 U14369 ( .A(n11399), .ZN(n11503) );
  AOI22_X1 U14370 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11406) );
  INV_X1 U14371 ( .A(n11400), .ZN(n11418) );
  AOI22_X1 U14372 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14373 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11404) );
  INV_X1 U14374 ( .A(n11401), .ZN(n12015) );
  INV_X2 U14375 ( .A(n12015), .ZN(n12138) );
  INV_X1 U14376 ( .A(n11402), .ZN(n11449) );
  AOI22_X1 U14377 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14378 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  OAI22_X1 U14379 ( .A1(n12226), .A2(n11409), .B1(n11493), .B2(n13329), .ZN(
        n11410) );
  INV_X1 U14380 ( .A(n11410), .ZN(n11411) );
  XNOR2_X2 U14381 ( .A(n11412), .B(n11411), .ZN(n11556) );
  INV_X1 U14382 ( .A(n11413), .ZN(n20551) );
  INV_X1 U14383 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11478) );
  NAND2_X1 U14384 ( .A1(n12136), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11420) );
  NAND2_X1 U14385 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11419) );
  OAI211_X1 U14386 ( .C1(n11729), .C2(n11478), .A(n11420), .B(n11419), .ZN(
        n11421) );
  INV_X1 U14387 ( .A(n11421), .ZN(n11426) );
  AOI22_X1 U14388 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14389 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14390 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11423) );
  NAND4_X1 U14391 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11433) );
  BUF_X1 U14392 ( .A(n11427), .Z(n11910) );
  AOI22_X1 U14393 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11900), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14394 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11430) );
  INV_X1 U14395 ( .A(n12166), .ZN(n12130) );
  AOI22_X1 U14396 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14397 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11428) );
  NAND4_X1 U14398 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11432) );
  NAND2_X1 U14399 ( .A1(n13767), .A2(n12963), .ZN(n11434) );
  INV_X1 U14400 ( .A(n11436), .ZN(n11437) );
  XNOR2_X2 U14401 ( .A(n11438), .B(n11437), .ZN(n14370) );
  INV_X1 U14402 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11442) );
  NAND2_X1 U14403 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U14405 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11440) );
  OAI211_X1 U14406 ( .C1(n11729), .C2(n11442), .A(n11441), .B(n11440), .ZN(
        n11443) );
  INV_X1 U14407 ( .A(n11443), .ZN(n11448) );
  AOI22_X1 U14408 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14409 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14411 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11445) );
  NAND4_X1 U14412 ( .A1(n11448), .A2(n11447), .A3(n11446), .A4(n11445), .ZN(
        n11455) );
  AOI22_X1 U14413 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14414 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14415 ( .A1(n11648), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14416 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11450) );
  NAND4_X1 U14417 ( .A1(n11453), .A2(n11452), .A3(n11451), .A4(n11450), .ZN(
        n11454) );
  INV_X1 U14418 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U14419 ( .A1(n11456), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U14420 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11457) );
  OAI211_X1 U14421 ( .C1(n11729), .C2(n11459), .A(n11458), .B(n11457), .ZN(
        n11460) );
  INV_X1 U14422 ( .A(n11460), .ZN(n11465) );
  AOI22_X1 U14423 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14424 ( .A1(n11308), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11463) );
  NAND2_X1 U14425 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11462) );
  NAND4_X1 U14426 ( .A1(n11465), .A2(n11464), .A3(n11463), .A4(n11462), .ZN(
        n11471) );
  AOI22_X1 U14427 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14428 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14429 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14430 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11466) );
  NAND4_X1 U14431 ( .A1(n11469), .A2(n11468), .A3(n11467), .A4(n11466), .ZN(
        n11470) );
  XNOR2_X1 U14432 ( .A(n13771), .B(n12964), .ZN(n11472) );
  NOR2_X1 U14433 ( .A1(n11472), .A2(n11492), .ZN(n11571) );
  INV_X1 U14434 ( .A(n13771), .ZN(n11474) );
  NAND2_X1 U14435 ( .A1(n20423), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11473) );
  AOI21_X1 U14436 ( .B1(n13394), .B2(n12964), .A(n21026), .ZN(n11475) );
  NAND2_X1 U14437 ( .A1(n11476), .A2(n11475), .ZN(n11573) );
  AOI22_X1 U14438 ( .A1(n11571), .A2(n11573), .B1(n13767), .B2(n13771), .ZN(
        n11477) );
  NAND2_X1 U14439 ( .A1(n11575), .A2(n11477), .ZN(n11483) );
  OR2_X1 U14440 ( .A1(n12226), .A2(n11478), .ZN(n11481) );
  INV_X1 U14441 ( .A(n11493), .ZN(n11479) );
  NAND2_X1 U14442 ( .A1(n11479), .A2(n12963), .ZN(n11480) );
  OAI211_X1 U14443 ( .C1(n11492), .C2(n13771), .A(n11481), .B(n11480), .ZN(
        n11482) );
  NAND2_X1 U14444 ( .A1(n11483), .A2(n11482), .ZN(n11484) );
  AOI21_X2 U14445 ( .B1(n12962), .B2(n11563), .A(n11486), .ZN(n11555) );
  NOR3_X1 U14446 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20764), .A3(
        n20839), .ZN(n20685) );
  NAND2_X1 U14447 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20685), .ZN(
        n20678) );
  NAND2_X1 U14448 ( .A1(n20804), .A2(n20678), .ZN(n11488) );
  NAND3_X1 U14449 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20971) );
  INV_X1 U14450 ( .A(n20971), .ZN(n11487) );
  NAND2_X1 U14451 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11487), .ZN(
        n20966) );
  NAND2_X1 U14452 ( .A1(n11488), .A2(n20966), .ZN(n20425) );
  OAI22_X1 U14453 ( .A1(n12795), .A2(n20425), .B1(n15976), .B2(n20804), .ZN(
        n11489) );
  INV_X1 U14454 ( .A(n11489), .ZN(n11490) );
  INV_X1 U14455 ( .A(n12226), .ZN(n11510) );
  INV_X1 U14456 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14457 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14458 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11495) );
  OAI211_X1 U14459 ( .C1(n11729), .C2(n11497), .A(n11496), .B(n11495), .ZN(
        n11498) );
  INV_X1 U14460 ( .A(n11498), .ZN(n11502) );
  AOI22_X1 U14461 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14462 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14463 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11499) );
  NAND4_X1 U14464 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11509) );
  AOI22_X1 U14465 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14466 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14467 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14468 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U14469 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11508) );
  AOI22_X1 U14470 ( .A1(n11510), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12232), .B2(n13673), .ZN(n11511) );
  INV_X1 U14471 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14472 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U14473 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11512) );
  OAI211_X1 U14474 ( .C1(n11729), .C2(n11525), .A(n11513), .B(n11512), .ZN(
        n11514) );
  INV_X1 U14475 ( .A(n11514), .ZN(n11518) );
  INV_X1 U14476 ( .A(n12155), .ZN(n11905) );
  AOI22_X1 U14477 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11905), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14478 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12166), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14479 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11515) );
  NAND4_X1 U14480 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(
        n11524) );
  AOI22_X1 U14481 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n9821), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14482 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12076), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14483 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14484 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11519) );
  NAND4_X1 U14485 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11523) );
  NAND2_X1 U14486 ( .A1(n12232), .A2(n13672), .ZN(n11527) );
  OR2_X1 U14487 ( .A1(n12226), .A2(n11525), .ZN(n11526) );
  NAND2_X1 U14488 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14489 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11528) );
  OAI211_X1 U14490 ( .C1(n11729), .C2(n11541), .A(n11529), .B(n11528), .ZN(
        n11530) );
  INV_X1 U14491 ( .A(n11530), .ZN(n11534) );
  AOI22_X1 U14492 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14493 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14494 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11531) );
  NAND4_X1 U14495 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11540) );
  AOI22_X1 U14496 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14497 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14498 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14499 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14500 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11539) );
  NAND2_X1 U14501 ( .A1(n12232), .A2(n13759), .ZN(n11543) );
  INV_X1 U14502 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11541) );
  OR2_X1 U14503 ( .A1(n12226), .A2(n11541), .ZN(n11542) );
  OAI21_X1 U14504 ( .B1(n11597), .B2(n11544), .A(n11545), .ZN(n11547) );
  INV_X1 U14505 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14506 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11588) );
  INV_X1 U14507 ( .A(n11588), .ZN(n11548) );
  INV_X1 U14508 ( .A(n11627), .ZN(n11629) );
  INV_X1 U14509 ( .A(n11549), .ZN(n11606) );
  INV_X1 U14510 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14511 ( .A1(n11606), .A2(n11550), .ZN(n11551) );
  NAND2_X1 U14512 ( .A1(n11629), .A2(n11551), .ZN(n20305) );
  AOI22_X1 U14513 ( .A1(n20305), .A2(n12145), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14514 ( .B1(n11633), .B2(n11553), .A(n11552), .ZN(n11554) );
  AOI21_X1 U14515 ( .B1(n13671), .B2(n11796), .A(n11554), .ZN(n13382) );
  NAND2_X1 U14516 ( .A1(n13631), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11601) );
  XNOR2_X1 U14517 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13421) );
  AOI21_X1 U14518 ( .B1(n13391), .B2(n13421), .A(n14378), .ZN(n11559) );
  NAND2_X1 U14519 ( .A1(n12180), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11558) );
  OAI211_X1 U14520 ( .C1(n11601), .C2(n11208), .A(n11559), .B(n11558), .ZN(
        n11560) );
  INV_X1 U14521 ( .A(n11560), .ZN(n11561) );
  NAND2_X1 U14522 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11585) );
  XNOR2_X2 U14523 ( .A(n11565), .B(n11564), .ZN(n13316) );
  NAND2_X1 U14524 ( .A1(n13316), .A2(n11796), .ZN(n11570) );
  INV_X1 U14525 ( .A(n11601), .ZN(n11566) );
  NAND2_X1 U14526 ( .A1(n11566), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11568) );
  AOI22_X1 U14527 ( .A1(n12180), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21028), .ZN(n11567) );
  AND2_X1 U14528 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  NAND2_X1 U14529 ( .A1(n11570), .A2(n11569), .ZN(n12860) );
  INV_X1 U14530 ( .A(n11571), .ZN(n11572) );
  XNOR2_X1 U14531 ( .A(n11573), .B(n11572), .ZN(n11574) );
  NAND2_X1 U14532 ( .A1(n20513), .A2(n11576), .ZN(n11577) );
  NAND2_X1 U14533 ( .A1(n11577), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U14534 ( .A1(n11578), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U14535 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11579) );
  OAI211_X1 U14536 ( .C1(n11601), .C2(n15948), .A(n11580), .B(n11579), .ZN(
        n11581) );
  AOI21_X1 U14537 ( .B1(n14370), .B2(n11796), .A(n11581), .ZN(n12797) );
  OR2_X1 U14538 ( .A1(n12798), .A2(n12797), .ZN(n12800) );
  INV_X1 U14539 ( .A(n12797), .ZN(n11582) );
  OR2_X1 U14540 ( .A1(n11582), .A2(n12178), .ZN(n11583) );
  NAND2_X1 U14541 ( .A1(n12800), .A2(n11583), .ZN(n12859) );
  NAND2_X1 U14542 ( .A1(n12860), .A2(n12859), .ZN(n12973) );
  NAND2_X1 U14543 ( .A1(n20419), .A2(n11796), .ZN(n11595) );
  INV_X1 U14544 ( .A(n11587), .ZN(n11604) );
  INV_X1 U14545 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11589) );
  NAND2_X1 U14546 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  NAND2_X1 U14547 ( .A1(n11604), .A2(n11590), .ZN(n13443) );
  AOI22_X1 U14548 ( .A1(n13443), .A2(n12145), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14549 ( .A1(n12180), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11591) );
  OAI211_X1 U14550 ( .C1(n11601), .C2(n11214), .A(n11592), .B(n11591), .ZN(
        n11593) );
  INV_X1 U14551 ( .A(n11593), .ZN(n11594) );
  NAND2_X1 U14552 ( .A1(n11595), .A2(n11594), .ZN(n13102) );
  XNOR2_X1 U14553 ( .A(n11597), .B(n11596), .ZN(n13669) );
  INV_X1 U14554 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14555 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U14556 ( .A1(n12180), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11598) );
  OAI211_X1 U14557 ( .C1(n11601), .C2(n11600), .A(n11599), .B(n11598), .ZN(
        n11602) );
  NAND2_X1 U14558 ( .A1(n11602), .A2(n12178), .ZN(n11608) );
  INV_X1 U14559 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14560 ( .A1(n11604), .A2(n11603), .ZN(n11605) );
  NAND2_X1 U14561 ( .A1(n11606), .A2(n11605), .ZN(n20373) );
  NAND2_X1 U14562 ( .A1(n20373), .A2(n12145), .ZN(n11607) );
  NAND2_X1 U14563 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  INV_X1 U14564 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U14565 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U14566 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11612) );
  OAI211_X1 U14567 ( .C1(n11729), .C2(n12124), .A(n11613), .B(n11612), .ZN(
        n11614) );
  INV_X1 U14568 ( .A(n11614), .ZN(n11618) );
  AOI22_X1 U14569 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14570 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14571 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11615) );
  NAND4_X1 U14572 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11624) );
  AOI22_X1 U14573 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14574 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14575 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14576 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11619) );
  NAND4_X1 U14577 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11623) );
  NAND2_X1 U14578 ( .A1(n12232), .A2(n13758), .ZN(n11626) );
  OR2_X1 U14579 ( .A1(n12226), .A2(n12124), .ZN(n11625) );
  XNOR2_X1 U14580 ( .A(n11635), .B(n11636), .ZN(n13683) );
  INV_X1 U14581 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11632) );
  INV_X1 U14582 ( .A(n11639), .ZN(n11641) );
  INV_X1 U14583 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14584 ( .A1(n11629), .A2(n11628), .ZN(n11630) );
  NAND2_X1 U14585 ( .A1(n11641), .A2(n11630), .ZN(n20296) );
  AOI22_X1 U14586 ( .A1(n20296), .A2(n12145), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11631) );
  OAI21_X1 U14587 ( .B1(n11633), .B2(n11632), .A(n11631), .ZN(n11634) );
  NOR2_X2 U14588 ( .A1(n13608), .A2(n13606), .ZN(n13598) );
  NAND2_X1 U14589 ( .A1(n12232), .A2(n13771), .ZN(n11637) );
  OAI21_X1 U14590 ( .B1(n11442), .B2(n12226), .A(n11637), .ZN(n11638) );
  XNOR2_X1 U14591 ( .A(n13769), .B(n11638), .ZN(n13755) );
  NAND2_X1 U14592 ( .A1(n13755), .A2(n11796), .ZN(n11647) );
  INV_X1 U14593 ( .A(n11669), .ZN(n11643) );
  INV_X1 U14594 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14595 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  NAND2_X1 U14596 ( .A1(n11643), .A2(n11642), .ZN(n20284) );
  AOI22_X1 U14597 ( .A1(n20284), .A2(n12145), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U14598 ( .A1(n12180), .A2(P1_EAX_REG_7__SCAN_IN), .ZN(n11644) );
  AND2_X1 U14599 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  NAND2_X1 U14600 ( .A1(n13598), .A2(n13597), .ZN(n13596) );
  AOI22_X1 U14601 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14602 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14603 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11648), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14604 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11649) );
  NAND4_X1 U14605 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11662) );
  INV_X1 U14606 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U14607 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11654) );
  NAND2_X1 U14608 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11653) );
  OAI211_X1 U14609 ( .C1(n11729), .C2(n11655), .A(n11654), .B(n11653), .ZN(
        n11656) );
  INV_X1 U14610 ( .A(n11656), .ZN(n11660) );
  AOI22_X1 U14611 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14612 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U14613 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11657) );
  NAND4_X1 U14614 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11661) );
  OAI21_X1 U14615 ( .B1(n11662), .B2(n11661), .A(n11796), .ZN(n11666) );
  NAND2_X1 U14616 ( .A1(n12180), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11665) );
  XNOR2_X1 U14617 ( .A(n11669), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13777) );
  NAND2_X1 U14618 ( .A1(n13777), .A2(n12145), .ZN(n11664) );
  NAND2_X1 U14619 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11663) );
  XNOR2_X1 U14620 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11702), .ZN(
        n20263) );
  INV_X1 U14621 ( .A(n20263), .ZN(n13908) );
  AOI22_X1 U14622 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14623 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14624 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14625 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11670) );
  NAND4_X1 U14626 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11683) );
  INV_X1 U14627 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14628 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11675) );
  NAND2_X1 U14629 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11674) );
  OAI211_X1 U14630 ( .C1(n11729), .C2(n11676), .A(n11675), .B(n11674), .ZN(
        n11677) );
  INV_X1 U14631 ( .A(n11677), .ZN(n11681) );
  AOI22_X1 U14632 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14633 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U14634 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11678) );
  NAND4_X1 U14635 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11682) );
  OAI21_X1 U14636 ( .B1(n11683), .B2(n11682), .A(n11796), .ZN(n11686) );
  NAND2_X1 U14637 ( .A1(n12180), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11685) );
  NAND2_X1 U14638 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11684) );
  NAND3_X1 U14639 ( .A1(n11686), .A2(n11685), .A3(n11684), .ZN(n11687) );
  INV_X1 U14640 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U14641 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14642 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11688) );
  OAI211_X1 U14643 ( .C1(n11729), .C2(n12016), .A(n11689), .B(n11688), .ZN(
        n11690) );
  INV_X1 U14644 ( .A(n11690), .ZN(n11694) );
  AOI22_X1 U14645 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14646 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14647 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11691) );
  NAND4_X1 U14648 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11700) );
  AOI22_X1 U14649 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14650 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14651 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14652 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14653 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  NOR2_X1 U14654 ( .A1(n11700), .A2(n11699), .ZN(n11705) );
  XNOR2_X1 U14655 ( .A(n11706), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14837) );
  NAND2_X1 U14656 ( .A1(n14837), .A2(n12145), .ZN(n11704) );
  AOI22_X1 U14657 ( .A1(n12180), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n14378), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11703) );
  OAI211_X1 U14658 ( .C1(n11705), .C2(n11762), .A(n11704), .B(n11703), .ZN(
        n13730) );
  NAND2_X1 U14659 ( .A1(n12180), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11709) );
  OAI21_X1 U14660 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11707), .A(
        n11757), .ZN(n16103) );
  AOI22_X1 U14661 ( .A1(n13391), .A2(n16103), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14662 ( .A1(n11709), .A2(n11708), .ZN(n13978) );
  INV_X1 U14663 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14664 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11711) );
  NAND2_X1 U14665 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11710) );
  OAI211_X1 U14666 ( .C1(n11729), .C2(n11712), .A(n11711), .B(n11710), .ZN(
        n11713) );
  INV_X1 U14667 ( .A(n11713), .ZN(n11717) );
  AOI22_X1 U14668 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14669 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14670 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11714) );
  NAND4_X1 U14671 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11723) );
  AOI22_X1 U14672 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14673 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14674 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14675 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11718) );
  NAND4_X1 U14676 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11722) );
  OR2_X1 U14677 ( .A1(n11723), .A2(n11722), .ZN(n11724) );
  XOR2_X1 U14678 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11764), .Z(
        n14826) );
  INV_X1 U14679 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11728) );
  NAND2_X1 U14680 ( .A1(n12136), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14681 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11726) );
  OAI211_X1 U14682 ( .C1(n11729), .C2(n11728), .A(n11727), .B(n11726), .ZN(
        n11730) );
  INV_X1 U14683 ( .A(n11730), .ZN(n11734) );
  AOI22_X1 U14684 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14685 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14686 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11731) );
  NAND4_X1 U14687 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n11740) );
  AOI22_X1 U14688 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14689 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14690 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14691 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11735) );
  NAND4_X1 U14692 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11739) );
  OR2_X1 U14693 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  AOI22_X1 U14694 ( .A1(n11796), .A2(n11741), .B1(n14378), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U14695 ( .A1(n12180), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11742) );
  OAI211_X1 U14696 ( .C1(n14826), .C2(n12178), .A(n11743), .B(n11742), .ZN(
        n14039) );
  INV_X1 U14697 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U14698 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14699 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11744) );
  OAI211_X1 U14700 ( .C1(n13298), .C2(n12068), .A(n11745), .B(n11744), .ZN(
        n11746) );
  INV_X1 U14701 ( .A(n11746), .ZN(n11750) );
  AOI22_X1 U14702 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14703 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14704 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11747) );
  NAND4_X1 U14705 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11756) );
  AOI22_X1 U14706 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14707 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14708 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12076), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14709 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U14710 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11755) );
  NOR2_X1 U14711 ( .A1(n11756), .A2(n11755), .ZN(n11761) );
  XNOR2_X1 U14712 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11757), .ZN(
        n16093) );
  INV_X1 U14713 ( .A(n16093), .ZN(n11758) );
  AOI22_X1 U14714 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13391), .B2(n11758), .ZN(n11760) );
  NAND2_X1 U14715 ( .A1(n12180), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11759) );
  OAI211_X1 U14716 ( .C1(n11762), .C2(n11761), .A(n11760), .B(n11759), .ZN(
        n14049) );
  XOR2_X1 U14717 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11804), .Z(
        n16084) );
  INV_X1 U14718 ( .A(n16084), .ZN(n11782) );
  AOI22_X1 U14719 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U14720 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14721 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14722 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11765) );
  NAND4_X1 U14723 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11777) );
  INV_X1 U14724 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U14725 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U14726 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11769) );
  OAI211_X1 U14727 ( .C1(n13298), .C2(n12157), .A(n11770), .B(n11769), .ZN(
        n11771) );
  INV_X1 U14728 ( .A(n11771), .ZN(n11775) );
  AOI22_X1 U14729 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14730 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14731 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11772) );
  NAND4_X1 U14732 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11776) );
  OAI21_X1 U14733 ( .B1(n11777), .B2(n11776), .A(n11796), .ZN(n11780) );
  NAND2_X1 U14734 ( .A1(n12180), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U14735 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11778) );
  NAND3_X1 U14736 ( .A1(n11780), .A2(n11779), .A3(n11778), .ZN(n11781) );
  AOI21_X1 U14737 ( .B1(n11782), .B2(n12145), .A(n11781), .ZN(n14078) );
  XNOR2_X1 U14738 ( .A(n11783), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14809) );
  AOI22_X1 U14739 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14740 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14741 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14742 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14743 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11798) );
  INV_X1 U14744 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U14745 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U14746 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11788) );
  OAI211_X1 U14747 ( .C1(n13298), .C2(n11790), .A(n11789), .B(n11788), .ZN(
        n11791) );
  INV_X1 U14748 ( .A(n11791), .ZN(n11795) );
  AOI22_X1 U14749 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14750 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U14751 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11792) );
  NAND4_X1 U14752 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11797) );
  OAI21_X1 U14753 ( .B1(n11798), .B2(n11797), .A(n11796), .ZN(n11801) );
  NAND2_X1 U14754 ( .A1(n12180), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11800) );
  NAND2_X1 U14755 ( .A1(n14378), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11799) );
  NAND3_X1 U14756 ( .A1(n11801), .A2(n11800), .A3(n11799), .ZN(n11802) );
  AOI21_X1 U14757 ( .B1(n14809), .B2(n12145), .A(n11802), .ZN(n14055) );
  OR2_X1 U14758 ( .A1(n14078), .A2(n14055), .ZN(n11803) );
  INV_X1 U14759 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11805) );
  XNOR2_X1 U14760 ( .A(n11824), .B(n11805), .ZN(n14560) );
  NAND2_X1 U14761 ( .A1(n14560), .A2(n12145), .ZN(n11822) );
  NAND2_X1 U14762 ( .A1(n12148), .A2(n12178), .ZN(n11944) );
  AOI22_X1 U14763 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14764 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14765 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14766 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11806) );
  NAND4_X1 U14767 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11817) );
  AOI22_X1 U14768 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14769 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11812) );
  AOI21_X1 U14770 ( .B1(n9823), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13391), .ZN(n11811) );
  NAND2_X1 U14771 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11810) );
  NAND4_X1 U14772 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n11816) );
  INV_X1 U14773 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11964) );
  INV_X1 U14774 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11814) );
  OAI22_X1 U14775 ( .A1(n13298), .A2(n11964), .B1(n11938), .B2(n11814), .ZN(
        n11815) );
  OR3_X1 U14776 ( .A1(n11817), .A2(n11816), .A3(n11815), .ZN(n11818) );
  NAND2_X1 U14777 ( .A1(n11944), .A2(n11818), .ZN(n11820) );
  AOI22_X1 U14778 ( .A1(n12180), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21028), .ZN(n11819) );
  NAND2_X1 U14779 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  NAND2_X1 U14780 ( .A1(n11822), .A2(n11821), .ZN(n14554) );
  INV_X1 U14781 ( .A(n14554), .ZN(n11823) );
  AND2_X2 U14782 ( .A1(n14074), .A2(n11823), .ZN(n14595) );
  XNOR2_X1 U14783 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11841), .ZN(
        n16076) );
  AOI22_X1 U14784 ( .A1(n12180), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14378), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14785 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14786 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14787 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14788 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U14789 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11838) );
  INV_X1 U14790 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14791 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U14792 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11829) );
  OAI211_X1 U14793 ( .C1(n13298), .C2(n11831), .A(n11830), .B(n11829), .ZN(
        n11832) );
  INV_X1 U14794 ( .A(n11832), .ZN(n11836) );
  AOI22_X1 U14795 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14796 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U14797 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11833) );
  NAND4_X1 U14798 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11837) );
  OAI21_X1 U14799 ( .B1(n11838), .B2(n11837), .A(n12175), .ZN(n11839) );
  OAI211_X1 U14800 ( .C1(n16076), .C2(n12178), .A(n11840), .B(n11839), .ZN(
        n14594) );
  INV_X1 U14801 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11842) );
  XNOR2_X1 U14802 ( .A(n11878), .B(n11842), .ZN(n14545) );
  NAND2_X1 U14803 ( .A1(n14545), .A2(n12145), .ZN(n11859) );
  AOI22_X1 U14804 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14805 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14806 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14807 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U14808 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11854) );
  AOI22_X1 U14809 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14810 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11849) );
  AOI21_X1 U14811 ( .B1(n12076), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n12145), .ZN(n11848) );
  NAND2_X1 U14812 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11847) );
  NAND4_X1 U14813 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11853) );
  INV_X1 U14814 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12013) );
  INV_X1 U14815 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11851) );
  OAI22_X1 U14816 ( .A1(n13298), .A2(n12013), .B1(n11938), .B2(n11851), .ZN(
        n11852) );
  OR3_X1 U14817 ( .A1(n11854), .A2(n11853), .A3(n11852), .ZN(n11855) );
  NAND2_X1 U14818 ( .A1(n11944), .A2(n11855), .ZN(n11857) );
  AOI22_X1 U14819 ( .A1(n12180), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21028), .ZN(n11856) );
  NAND2_X1 U14820 ( .A1(n11857), .A2(n11856), .ZN(n11858) );
  NAND2_X1 U14821 ( .A1(n11859), .A2(n11858), .ZN(n14583) );
  INV_X1 U14822 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U14823 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11861) );
  NAND2_X1 U14824 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11860) );
  OAI211_X1 U14825 ( .C1(n13298), .C2(n11862), .A(n11861), .B(n11860), .ZN(
        n11863) );
  INV_X1 U14826 ( .A(n11863), .ZN(n11867) );
  AOI22_X1 U14827 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14828 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14829 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11864) );
  NAND4_X1 U14830 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11873) );
  AOI22_X1 U14831 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14832 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14833 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14834 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U14835 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  NOR2_X1 U14836 ( .A1(n11873), .A2(n11872), .ZN(n11877) );
  OAI21_X1 U14837 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21220), .A(
        n21028), .ZN(n11874) );
  INV_X1 U14838 ( .A(n11874), .ZN(n11875) );
  AOI21_X1 U14839 ( .B1(n12180), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11875), .ZN(
        n11876) );
  OAI21_X1 U14840 ( .B1(n12148), .B2(n11877), .A(n11876), .ZN(n11881) );
  OAI21_X1 U14841 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11879), .A(
        n11921), .ZN(n16067) );
  OR2_X1 U14842 ( .A1(n12178), .A2(n16067), .ZN(n11880) );
  NAND2_X1 U14843 ( .A1(n11881), .A2(n11880), .ZN(n14586) );
  NOR2_X2 U14844 ( .A1(n14542), .A2(n11882), .ZN(n14532) );
  AOI22_X1 U14845 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12138), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14846 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14847 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11399), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14848 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9821), .B1(n9823), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U14849 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11895) );
  AOI22_X1 U14850 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14851 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12166), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11889) );
  AOI21_X1 U14852 ( .B1(n12076), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12145), .ZN(n11888) );
  NAND2_X1 U14853 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11887) );
  NAND4_X1 U14854 ( .A1(n11890), .A2(n11889), .A3(n11888), .A4(n11887), .ZN(
        n11894) );
  INV_X1 U14855 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11892) );
  INV_X1 U14856 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11891) );
  OAI22_X1 U14857 ( .A1(n11892), .A2(n13298), .B1(n11938), .B2(n11891), .ZN(
        n11893) );
  OR3_X1 U14858 ( .A1(n11895), .A2(n11894), .A3(n11893), .ZN(n11896) );
  NAND2_X1 U14859 ( .A1(n11944), .A2(n11896), .ZN(n11899) );
  AOI22_X1 U14860 ( .A1(n12180), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21028), .ZN(n11898) );
  XNOR2_X1 U14861 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11921), .ZN(
        n14779) );
  AND2_X1 U14862 ( .A1(n13391), .A2(n14779), .ZN(n11897) );
  AOI21_X1 U14863 ( .B1(n11899), .B2(n11898), .A(n11897), .ZN(n14533) );
  AND2_X2 U14864 ( .A1(n14532), .A2(n14533), .ZN(n14576) );
  INV_X1 U14865 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U14866 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11902) );
  NAND2_X1 U14867 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11901) );
  OAI211_X1 U14868 ( .C1(n13298), .C2(n11903), .A(n11902), .B(n11901), .ZN(
        n11904) );
  INV_X1 U14869 ( .A(n11904), .ZN(n11909) );
  AOI22_X1 U14870 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14871 ( .A1(n11905), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U14872 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11906) );
  NAND4_X1 U14873 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11916) );
  AOI22_X1 U14874 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14875 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14876 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14877 ( .A1(n11962), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11911) );
  NAND4_X1 U14878 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n11915) );
  NOR2_X1 U14879 ( .A1(n11916), .A2(n11915), .ZN(n11920) );
  OAI21_X1 U14880 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21220), .A(
        n21028), .ZN(n11917) );
  INV_X1 U14881 ( .A(n11917), .ZN(n11918) );
  AOI21_X1 U14882 ( .B1(n12180), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11918), .ZN(
        n11919) );
  OAI21_X1 U14883 ( .B1(n12148), .B2(n11920), .A(n11919), .ZN(n11927) );
  INV_X1 U14884 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16010) );
  INV_X1 U14885 ( .A(n11923), .ZN(n11924) );
  NAND2_X1 U14886 ( .A1(n16010), .A2(n11924), .ZN(n11925) );
  NAND2_X1 U14887 ( .A1(n11982), .A2(n11925), .ZN(n16018) );
  AOI22_X1 U14888 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14889 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14890 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14891 ( .A1(n12136), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11929) );
  NAND4_X1 U14892 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11942) );
  AOI22_X1 U14893 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12166), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14894 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12105), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11935) );
  AOI21_X1 U14895 ( .B1(n11905), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12145), .ZN(n11934) );
  NAND2_X1 U14896 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11933) );
  NAND4_X1 U14897 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n11941) );
  INV_X1 U14898 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11939) );
  INV_X1 U14899 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11937) );
  OAI22_X1 U14900 ( .A1(n13298), .A2(n11939), .B1(n11938), .B2(n11937), .ZN(
        n11940) );
  OR3_X1 U14901 ( .A1(n11942), .A2(n11941), .A3(n11940), .ZN(n11943) );
  NAND2_X1 U14902 ( .A1(n11944), .A2(n11943), .ZN(n11946) );
  AOI22_X1 U14903 ( .A1(n12180), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21028), .ZN(n11945) );
  NAND2_X1 U14904 ( .A1(n11946), .A2(n11945), .ZN(n11948) );
  XNOR2_X1 U14905 ( .A(n11982), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14765) );
  NAND2_X1 U14906 ( .A1(n14765), .A2(n12145), .ZN(n11947) );
  NAND2_X1 U14907 ( .A1(n11948), .A2(n11947), .ZN(n14521) );
  INV_X1 U14908 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11955) );
  INV_X1 U14909 ( .A(n11949), .ZN(n12126) );
  INV_X1 U14910 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12162) );
  OAI22_X1 U14911 ( .A1(n12126), .A2(n12162), .B1(n9824), .B2(n11950), .ZN(
        n11952) );
  INV_X1 U14912 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12154) );
  OAI22_X1 U14913 ( .A1(n12018), .A2(n12154), .B1(n11503), .B2(n12157), .ZN(
        n11951) );
  AOI211_X1 U14914 ( .C1(n11461), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n11952), .B(n11951), .ZN(n11954) );
  AOI22_X1 U14915 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11953) );
  OAI211_X1 U14916 ( .C1(n12163), .C2(n11955), .A(n11954), .B(n11953), .ZN(
        n11961) );
  AOI22_X1 U14917 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U14918 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U14919 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U14920 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U14921 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  NOR2_X1 U14922 ( .A1(n11961), .A2(n11960), .ZN(n11988) );
  INV_X1 U14923 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11971) );
  OAI22_X1 U14924 ( .A1(n11503), .A2(n11964), .B1(n11449), .B2(n11963), .ZN(
        n11968) );
  INV_X1 U14925 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11965) );
  OAI22_X1 U14926 ( .A1(n12128), .A2(n11966), .B1(n12126), .B2(n11965), .ZN(
        n11967) );
  AOI211_X1 U14927 ( .C1(n11461), .C2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n11968), .B(n11967), .ZN(n11970) );
  AOI22_X1 U14928 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12165), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11969) );
  OAI211_X1 U14929 ( .C1(n12163), .C2(n11971), .A(n11970), .B(n11969), .ZN(
        n11977) );
  AOI22_X1 U14930 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U14931 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9821), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14932 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U14933 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11972) );
  NAND4_X1 U14934 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n11976) );
  NOR2_X1 U14935 ( .A1(n11977), .A2(n11976), .ZN(n11989) );
  XNOR2_X1 U14936 ( .A(n11988), .B(n11989), .ZN(n11981) );
  NAND2_X1 U14937 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U14938 ( .A1(n12178), .A2(n11978), .ZN(n11979) );
  AOI21_X1 U14939 ( .B1(n12180), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11979), .ZN(
        n11980) );
  OAI21_X1 U14940 ( .B1(n12148), .B2(n11981), .A(n11980), .ZN(n11987) );
  INV_X1 U14941 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14763) );
  INV_X1 U14942 ( .A(n11983), .ZN(n11984) );
  INV_X1 U14943 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14510) );
  NAND2_X1 U14944 ( .A1(n11984), .A2(n14510), .ZN(n11985) );
  NAND2_X1 U14945 ( .A1(n12034), .A2(n11985), .ZN(n14755) );
  NAND2_X1 U14946 ( .A1(n11987), .A2(n11986), .ZN(n14509) );
  NOR2_X1 U14947 ( .A1(n11989), .A2(n11988), .ZN(n12012) );
  INV_X1 U14948 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11992) );
  NAND2_X1 U14949 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U14950 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11990) );
  OAI211_X1 U14951 ( .C1(n12163), .C2(n11992), .A(n11991), .B(n11990), .ZN(
        n11993) );
  INV_X1 U14952 ( .A(n11993), .ZN(n11997) );
  AOI22_X1 U14953 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U14954 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U14955 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11994) );
  NAND4_X1 U14956 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n12003) );
  AOI22_X1 U14957 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U14958 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U14959 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U14960 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U14961 ( .A1(n12001), .A2(n12000), .A3(n11999), .A4(n11998), .ZN(
        n12002) );
  OR2_X1 U14962 ( .A1(n12003), .A2(n12002), .ZN(n12011) );
  INV_X1 U14963 ( .A(n12011), .ZN(n12004) );
  XNOR2_X1 U14964 ( .A(n12012), .B(n12004), .ZN(n12005) );
  NAND2_X1 U14965 ( .A1(n12005), .A2(n12175), .ZN(n12010) );
  NAND2_X1 U14966 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U14967 ( .A1(n12178), .A2(n12006), .ZN(n12007) );
  AOI21_X1 U14968 ( .B1(n12180), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12007), .ZN(
        n12009) );
  XNOR2_X1 U14969 ( .A(n12034), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14747) );
  AOI21_X1 U14970 ( .B1(n12010), .B2(n12009), .A(n12008), .ZN(n14494) );
  NAND2_X1 U14971 ( .A1(n12012), .A2(n12011), .ZN(n12042) );
  INV_X1 U14972 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12023) );
  INV_X1 U14973 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12014) );
  OAI22_X1 U14974 ( .A1(n12015), .A2(n12014), .B1(n11503), .B2(n12013), .ZN(
        n12020) );
  INV_X1 U14975 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12017) );
  OAI22_X1 U14976 ( .A1(n12018), .A2(n12017), .B1(n11418), .B2(n12016), .ZN(
        n12019) );
  AOI211_X1 U14977 ( .C1(n11461), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n12020), .B(n12019), .ZN(n12022) );
  AOI22_X1 U14978 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11439), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12021) );
  OAI211_X1 U14979 ( .C1(n12163), .C2(n12023), .A(n12022), .B(n12021), .ZN(
        n12029) );
  AOI22_X1 U14980 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U14981 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11905), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U14982 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U14983 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12024) );
  NAND4_X1 U14984 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12028) );
  NOR2_X1 U14985 ( .A1(n12029), .A2(n12028), .ZN(n12043) );
  XNOR2_X1 U14986 ( .A(n12042), .B(n12043), .ZN(n12033) );
  NAND2_X1 U14987 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12030) );
  NAND2_X1 U14988 ( .A1(n12178), .A2(n12030), .ZN(n12031) );
  AOI21_X1 U14989 ( .B1(n12180), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12031), .ZN(
        n12032) );
  OAI21_X1 U14990 ( .B1(n12033), .B2(n12148), .A(n12032), .ZN(n12041) );
  INV_X1 U14991 ( .A(n12034), .ZN(n12035) );
  INV_X1 U14992 ( .A(n12036), .ZN(n12038) );
  INV_X1 U14993 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12037) );
  NAND2_X1 U14994 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  NAND2_X1 U14995 ( .A1(n12087), .A2(n12039), .ZN(n14738) );
  NOR2_X1 U14996 ( .A1(n12043), .A2(n12042), .ZN(n12065) );
  INV_X1 U14997 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U14998 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12045) );
  NAND2_X1 U14999 ( .A1(n11439), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12044) );
  OAI211_X1 U15000 ( .C1(n12163), .C2(n12046), .A(n12045), .B(n12044), .ZN(
        n12047) );
  INV_X1 U15001 ( .A(n12047), .ZN(n12051) );
  AOI22_X1 U15002 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15003 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U15004 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12048) );
  NAND4_X1 U15005 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12057) );
  AOI22_X1 U15006 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15007 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15008 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15009 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11456), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12052) );
  NAND4_X1 U15010 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(
        n12056) );
  OR2_X1 U15011 ( .A1(n12057), .A2(n12056), .ZN(n12064) );
  XNOR2_X1 U15012 ( .A(n12065), .B(n12064), .ZN(n12061) );
  NAND2_X1 U15013 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12058) );
  NAND2_X1 U15014 ( .A1(n12178), .A2(n12058), .ZN(n12059) );
  AOI21_X1 U15015 ( .B1(n12180), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12059), .ZN(
        n12060) );
  OAI21_X1 U15016 ( .B1(n12061), .B2(n12148), .A(n12060), .ZN(n12063) );
  XNOR2_X1 U15017 ( .A(n12087), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14729) );
  NAND2_X1 U15018 ( .A1(n14729), .A2(n12145), .ZN(n12062) );
  NAND2_X1 U15019 ( .A1(n12063), .A2(n12062), .ZN(n14464) );
  OR2_X2 U15020 ( .A1(n14479), .A2(n14464), .ZN(n14465) );
  NAND2_X1 U15021 ( .A1(n12065), .A2(n12064), .ZN(n12095) );
  INV_X1 U15022 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12075) );
  INV_X1 U15023 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12067) );
  OAI22_X1 U15024 ( .A1(n12067), .A2(n12126), .B1(n11449), .B2(n12066), .ZN(
        n12072) );
  INV_X1 U15025 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12069) );
  OAI22_X1 U15026 ( .A1(n12070), .A2(n12069), .B1(n11418), .B2(n12068), .ZN(
        n12071) );
  AOI211_X1 U15027 ( .C1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .C2(n11461), .A(
        n12072), .B(n12071), .ZN(n12074) );
  AOI22_X1 U15028 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11494), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12073) );
  OAI211_X1 U15029 ( .C1(n12075), .C2(n13298), .A(n12074), .B(n12073), .ZN(
        n12082) );
  AOI22_X1 U15030 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12076), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15031 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12166), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15032 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11962), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15033 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15034 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12081) );
  NOR2_X1 U15035 ( .A1(n12082), .A2(n12081), .ZN(n12096) );
  XNOR2_X1 U15036 ( .A(n12095), .B(n12096), .ZN(n12086) );
  NAND2_X1 U15037 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12083) );
  NAND2_X1 U15038 ( .A1(n12178), .A2(n12083), .ZN(n12084) );
  AOI21_X1 U15039 ( .B1(n12180), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12084), .ZN(
        n12085) );
  OAI21_X1 U15040 ( .B1(n12086), .B2(n12148), .A(n12085), .ZN(n12094) );
  INV_X1 U15041 ( .A(n12087), .ZN(n12088) );
  INV_X1 U15042 ( .A(n12089), .ZN(n12091) );
  INV_X1 U15043 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12090) );
  NAND2_X1 U15044 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U15045 ( .A1(n12119), .A2(n12092), .ZN(n14718) );
  OR2_X1 U15046 ( .A1(n14718), .A2(n12178), .ZN(n12093) );
  NAND2_X1 U15047 ( .A1(n12094), .A2(n12093), .ZN(n14455) );
  NOR2_X1 U15048 ( .A1(n12096), .A2(n12095), .ZN(n12123) );
  INV_X1 U15049 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12099) );
  NAND2_X1 U15050 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12098) );
  NAND2_X1 U15051 ( .A1(n11494), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12097) );
  OAI211_X1 U15052 ( .C1(n12163), .C2(n12099), .A(n12098), .B(n12097), .ZN(
        n12100) );
  INV_X1 U15053 ( .A(n12100), .ZN(n12104) );
  AOI22_X1 U15054 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15055 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U15056 ( .A1(n11444), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12101) );
  NAND4_X1 U15057 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12111) );
  AOI22_X1 U15058 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15059 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15060 ( .A1(n12105), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9823), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15061 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12106) );
  NAND4_X1 U15062 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  OR2_X1 U15063 ( .A1(n12111), .A2(n12110), .ZN(n12122) );
  INV_X1 U15064 ( .A(n12122), .ZN(n12112) );
  XNOR2_X1 U15065 ( .A(n12123), .B(n12112), .ZN(n12113) );
  NAND2_X1 U15066 ( .A1(n12113), .A2(n12175), .ZN(n12118) );
  NAND2_X1 U15067 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12114) );
  NAND2_X1 U15068 ( .A1(n12178), .A2(n12114), .ZN(n12115) );
  AOI21_X1 U15069 ( .B1(n12180), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12115), .ZN(
        n12117) );
  XNOR2_X1 U15070 ( .A(n12119), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14698) );
  AOI21_X1 U15071 ( .B1(n12118), .B2(n12117), .A(n12116), .ZN(n14441) );
  INV_X1 U15072 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14696) );
  INV_X1 U15073 ( .A(n12120), .ZN(n12121) );
  INV_X1 U15074 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U15075 ( .B1(n12121), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13397), .ZN(n14692) );
  NAND2_X1 U15076 ( .A1(n12123), .A2(n12122), .ZN(n12151) );
  INV_X1 U15077 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12135) );
  INV_X1 U15078 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12125) );
  OAI22_X1 U15079 ( .A1(n12126), .A2(n12125), .B1(n9824), .B2(n12124), .ZN(
        n12132) );
  INV_X1 U15080 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12129) );
  OAI22_X1 U15081 ( .A1(n12130), .A2(n12129), .B1(n12128), .B2(n12127), .ZN(
        n12131) );
  AOI211_X1 U15082 ( .C1(n11444), .C2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12132), .B(n12131), .ZN(n12134) );
  AOI22_X1 U15083 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11494), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12133) );
  OAI211_X1 U15084 ( .C1(n12163), .C2(n12135), .A(n12134), .B(n12133), .ZN(
        n12144) );
  AOI22_X1 U15085 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11308), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15086 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15087 ( .A1(n9821), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15088 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12139) );
  NAND4_X1 U15089 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12143) );
  NOR2_X1 U15090 ( .A1(n12144), .A2(n12143), .ZN(n12152) );
  XNOR2_X1 U15091 ( .A(n12151), .B(n12152), .ZN(n12149) );
  AOI21_X1 U15092 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21028), .A(
        n12145), .ZN(n12147) );
  NAND2_X1 U15093 ( .A1(n12180), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12146) );
  OAI211_X1 U15094 ( .C1(n12149), .C2(n12148), .A(n12147), .B(n12146), .ZN(
        n12150) );
  OAI21_X1 U15095 ( .B1(n12178), .B2(n14692), .A(n12150), .ZN(n14430) );
  NOR2_X1 U15096 ( .A1(n12152), .A2(n12151), .ZN(n12174) );
  OAI22_X1 U15097 ( .A1(n12155), .A2(n12154), .B1(n9824), .B2(n11442), .ZN(
        n12159) );
  INV_X1 U15098 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12156) );
  OAI22_X1 U15099 ( .A1(n11418), .A2(n12157), .B1(n11449), .B2(n12156), .ZN(
        n12158) );
  AOI211_X1 U15100 ( .C1(n11444), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n12159), .B(n12158), .ZN(n12161) );
  AOI22_X1 U15101 ( .A1(n11427), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11494), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12160) );
  OAI211_X1 U15102 ( .C1(n12163), .C2(n12162), .A(n12161), .B(n12160), .ZN(
        n12172) );
  AOI22_X1 U15103 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15104 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11399), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15105 ( .A1(n12165), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12137), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15106 ( .A1(n12166), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15107 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  NOR2_X1 U15108 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  XNOR2_X1 U15109 ( .A(n12174), .B(n12173), .ZN(n12176) );
  NAND2_X1 U15110 ( .A1(n12176), .A2(n12175), .ZN(n12183) );
  NAND2_X1 U15111 ( .A1(n21028), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12177) );
  NAND2_X1 U15112 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  AOI21_X1 U15113 ( .B1(n12180), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12179), .ZN(
        n12182) );
  XNOR2_X1 U15114 ( .A(n13397), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14681) );
  AOI21_X1 U15115 ( .B1(n12183), .B2(n12182), .A(n12181), .ZN(n14377) );
  XNOR2_X1 U15116 ( .A(n14429), .B(n12184), .ZN(n14685) );
  XNOR2_X1 U15117 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U15118 ( .A1(n12197), .A2(n12198), .ZN(n12186) );
  NAND2_X1 U15119 ( .A1(n20839), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12185) );
  NAND2_X1 U15120 ( .A1(n12186), .A2(n12185), .ZN(n12210) );
  XNOR2_X1 U15121 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12209) );
  NAND2_X1 U15122 ( .A1(n12210), .A2(n12209), .ZN(n12188) );
  NAND2_X1 U15123 ( .A1(n20764), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12187) );
  NAND2_X1 U15124 ( .A1(n12188), .A2(n12187), .ZN(n12192) );
  XNOR2_X1 U15125 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15126 ( .A1(n12192), .A2(n12191), .ZN(n12190) );
  NAND2_X1 U15127 ( .A1(n20804), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12189) );
  NAND2_X1 U15128 ( .A1(n12190), .A2(n12189), .ZN(n12229) );
  NAND2_X1 U15129 ( .A1(n20440), .A2(n20463), .ZN(n13756) );
  XNOR2_X1 U15130 ( .A(n12192), .B(n12191), .ZN(n12643) );
  NAND2_X1 U15131 ( .A1(n13403), .A2(n20463), .ZN(n12193) );
  NAND2_X1 U15132 ( .A1(n12193), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U15133 ( .A1(n13767), .A2(n20440), .ZN(n12194) );
  NOR3_X1 U15134 ( .A1(n12200), .A2(n12868), .A3(n12196), .ZN(n12224) );
  AOI21_X1 U15135 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n15948), .A(
        n12197), .ZN(n12203) );
  NAND2_X1 U15136 ( .A1(n12232), .A2(n12203), .ZN(n12206) );
  INV_X1 U15137 ( .A(n12235), .ZN(n12205) );
  XNOR2_X1 U15138 ( .A(n12198), .B(n12197), .ZN(n12645) );
  INV_X1 U15139 ( .A(n12645), .ZN(n12201) );
  NOR2_X1 U15140 ( .A1(n12226), .A2(n12201), .ZN(n12199) );
  NOR2_X1 U15141 ( .A1(n12200), .A2(n12199), .ZN(n12207) );
  AOI21_X1 U15142 ( .B1(n12202), .B2(n20440), .A(n12201), .ZN(n12208) );
  NAND2_X1 U15143 ( .A1(n12218), .A2(n20423), .ZN(n12211) );
  OAI211_X1 U15144 ( .C1(n13767), .C2(n12868), .A(n12211), .B(n13403), .ZN(
        n12204) );
  AOI222_X1 U15145 ( .A1(n12206), .A2(n12205), .B1(n12207), .B2(n12208), .C1(
        n12204), .C2(n12203), .ZN(n12216) );
  NOR2_X1 U15146 ( .A1(n12208), .A2(n12207), .ZN(n12215) );
  XNOR2_X1 U15147 ( .A(n12210), .B(n12209), .ZN(n12644) );
  INV_X1 U15148 ( .A(n12644), .ZN(n12212) );
  INV_X1 U15149 ( .A(n12211), .ZN(n12213) );
  OAI22_X1 U15150 ( .A1(n12213), .A2(n20440), .B1(n12212), .B2(n12226), .ZN(
        n12214) );
  OAI22_X1 U15151 ( .A1(n12216), .A2(n12215), .B1(n12220), .B2(n12214), .ZN(
        n12222) );
  OAI21_X1 U15152 ( .B1(n12218), .B2(n20440), .A(n12217), .ZN(n12219) );
  NAND2_X1 U15153 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  AOI22_X1 U15154 ( .A1(n12222), .A2(n12221), .B1(n12226), .B2(n12643), .ZN(
        n12223) );
  AOI211_X1 U15155 ( .C1(n12235), .C2(n12643), .A(n12224), .B(n12223), .ZN(
        n12225) );
  AOI21_X1 U15156 ( .B1(n12646), .B2(n12226), .A(n12225), .ZN(n12227) );
  AOI21_X1 U15157 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21026), .A(
        n12227), .ZN(n12234) );
  NOR2_X1 U15158 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11600), .ZN(
        n12228) );
  NAND2_X1 U15159 ( .A1(n12648), .A2(n12232), .ZN(n12233) );
  NAND2_X1 U15160 ( .A1(n12234), .A2(n12233), .ZN(n12237) );
  NAND2_X1 U15161 ( .A1(n12235), .A2(n12648), .ZN(n12236) );
  NAND2_X4 U15162 ( .A1(n12237), .A2(n12236), .ZN(n13620) );
  NOR2_X1 U15163 ( .A1(n14368), .A2(n12868), .ZN(n12928) );
  INV_X1 U15164 ( .A(n12806), .ZN(n12786) );
  INV_X1 U15165 ( .A(n13403), .ZN(n12807) );
  NAND2_X1 U15166 ( .A1(n12786), .A2(n12807), .ZN(n12878) );
  NAND2_X1 U15167 ( .A1(n12928), .A2(n12238), .ZN(n12740) );
  INV_X1 U15168 ( .A(n20478), .ZN(n14381) );
  AND3_X1 U15169 ( .A1(n11354), .A2(n14381), .A3(n20471), .ZN(n13621) );
  NAND3_X1 U15170 ( .A1(n12239), .A2(n13619), .A3(n13621), .ZN(n12240) );
  INV_X1 U15171 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20397) );
  NAND2_X1 U15172 ( .A1(n12318), .A2(n20397), .ZN(n12243) );
  INV_X1 U15173 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21272) );
  NAND2_X1 U15174 ( .A1(n12254), .A2(n21272), .ZN(n12242) );
  NAND3_X1 U15175 ( .A1(n12243), .A2(n12327), .A3(n12242), .ZN(n12245) );
  NAND2_X1 U15176 ( .A1(n14343), .A2(n21272), .ZN(n12244) );
  NAND2_X1 U15177 ( .A1(n12245), .A2(n12244), .ZN(n12247) );
  NAND2_X1 U15178 ( .A1(n12318), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12246) );
  OAI21_X1 U15179 ( .B1(n14343), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12246), .ZN(
        n12858) );
  XNOR2_X1 U15180 ( .A(n12247), .B(n12858), .ZN(n12862) );
  NAND2_X1 U15181 ( .A1(n12862), .A2(n13619), .ZN(n12863) );
  INV_X1 U15182 ( .A(n12247), .ZN(n12248) );
  NAND2_X1 U15183 ( .A1(n12248), .A2(n12858), .ZN(n12249) );
  NAND2_X1 U15184 ( .A1(n12863), .A2(n12249), .ZN(n12976) );
  INV_X1 U15185 ( .A(n12318), .ZN(n12312) );
  MUX2_X1 U15186 ( .A(n14343), .B(n12312), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12251) );
  INV_X1 U15187 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20411) );
  NOR2_X1 U15188 ( .A1(n13619), .A2(n20411), .ZN(n12250) );
  NOR2_X1 U15189 ( .A1(n12251), .A2(n12250), .ZN(n12975) );
  OR2_X2 U15190 ( .A1(n12976), .A2(n12975), .ZN(n13099) );
  MUX2_X1 U15191 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12253) );
  OAI21_X1 U15192 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14341), .A(
        n12253), .ZN(n13098) );
  MUX2_X1 U15193 ( .A(n12327), .B(n12318), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12256) );
  INV_X1 U15194 ( .A(n12254), .ZN(n14340) );
  NAND2_X1 U15195 ( .A1(n14340), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12255) );
  NAND2_X1 U15196 ( .A1(n12256), .A2(n12255), .ZN(n13378) );
  INV_X1 U15197 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16239) );
  INV_X1 U15198 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21450) );
  NAND2_X1 U15199 ( .A1(n13619), .A2(n21450), .ZN(n12257) );
  OAI211_X1 U15200 ( .C1(n14343), .C2(n16239), .A(n12257), .B(n12318), .ZN(
        n12258) );
  OAI21_X1 U15201 ( .B1(n12315), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12258), .ZN(
        n13386) );
  MUX2_X1 U15202 ( .A(n14343), .B(n12312), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12261) );
  INV_X1 U15203 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12259) );
  NOR2_X1 U15204 ( .A1(n13619), .A2(n12259), .ZN(n12260) );
  NOR2_X1 U15205 ( .A1(n12261), .A2(n12260), .ZN(n13602) );
  INV_X1 U15206 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16231) );
  INV_X1 U15207 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21337) );
  NAND2_X1 U15208 ( .A1(n13619), .A2(n21337), .ZN(n12262) );
  OAI211_X1 U15209 ( .C1(n14343), .C2(n16231), .A(n12262), .B(n12318), .ZN(
        n12263) );
  OAI21_X1 U15210 ( .B1(n12315), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12263), .ZN(
        n13600) );
  NOR2_X2 U15211 ( .A1(n13605), .A2(n13600), .ZN(n13645) );
  MUX2_X1 U15212 ( .A(n12327), .B(n12318), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12265) );
  NAND2_X1 U15213 ( .A1(n14340), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12264) );
  NAND2_X1 U15214 ( .A1(n12265), .A2(n12264), .ZN(n13644) );
  NAND2_X1 U15215 ( .A1(n13645), .A2(n13644), .ZN(n13715) );
  INV_X1 U15216 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16217) );
  INV_X1 U15217 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U15218 ( .A1(n13619), .A2(n13717), .ZN(n12266) );
  OAI211_X1 U15219 ( .C1(n14343), .C2(n16217), .A(n12266), .B(n12318), .ZN(
        n12267) );
  OAI21_X1 U15220 ( .B1(n12315), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12267), .ZN(
        n13714) );
  OR2_X2 U15221 ( .A1(n13715), .A2(n13714), .ZN(n13735) );
  NAND2_X1 U15222 ( .A1(n12318), .A2(n16207), .ZN(n12269) );
  INV_X1 U15223 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21507) );
  NAND2_X1 U15224 ( .A1(n13619), .A2(n21507), .ZN(n12268) );
  NAND3_X1 U15225 ( .A1(n12269), .A2(n12327), .A3(n12268), .ZN(n12271) );
  NAND2_X1 U15226 ( .A1(n14343), .A2(n21507), .ZN(n12270) );
  MUX2_X1 U15227 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12272) );
  OAI21_X1 U15228 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14341), .A(
        n12272), .ZN(n12273) );
  INV_X1 U15229 ( .A(n12273), .ZN(n14013) );
  MUX2_X1 U15230 ( .A(n14343), .B(n12312), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12275) );
  INV_X1 U15231 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14818) );
  NOR2_X1 U15232 ( .A1(n13619), .A2(n14818), .ZN(n12274) );
  NOR2_X1 U15233 ( .A1(n12275), .A2(n12274), .ZN(n14070) );
  MUX2_X1 U15234 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12276) );
  OAI21_X1 U15235 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14341), .A(
        n12276), .ZN(n14040) );
  INV_X1 U15236 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14331) );
  NAND2_X1 U15237 ( .A1(n12318), .A2(n14331), .ZN(n12278) );
  INV_X1 U15238 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15239 ( .A1(n13619), .A2(n12279), .ZN(n12277) );
  NAND3_X1 U15240 ( .A1(n12278), .A2(n12327), .A3(n12277), .ZN(n12281) );
  NAND2_X1 U15241 ( .A1(n14343), .A2(n12279), .ZN(n12280) );
  NAND2_X1 U15242 ( .A1(n12281), .A2(n12280), .ZN(n14059) );
  MUX2_X1 U15243 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12283) );
  INV_X1 U15244 ( .A(n14341), .ZN(n12309) );
  INV_X1 U15245 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16159) );
  NAND2_X1 U15246 ( .A1(n12309), .A2(n16159), .ZN(n12282) );
  INV_X1 U15247 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16156) );
  NAND2_X1 U15248 ( .A1(n12318), .A2(n16156), .ZN(n12285) );
  INV_X1 U15249 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U15250 ( .A1(n13619), .A2(n14603), .ZN(n12284) );
  NAND3_X1 U15251 ( .A1(n12285), .A2(n12327), .A3(n12284), .ZN(n12287) );
  NAND2_X1 U15252 ( .A1(n14343), .A2(n14603), .ZN(n12286) );
  AND2_X1 U15253 ( .A1(n12287), .A2(n12286), .ZN(n14558) );
  OR2_X2 U15254 ( .A1(n14609), .A2(n14558), .ZN(n14597) );
  INV_X1 U15255 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16141) );
  INV_X1 U15256 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21485) );
  NAND2_X1 U15257 ( .A1(n13619), .A2(n21485), .ZN(n12288) );
  OAI211_X1 U15258 ( .C1(n14343), .C2(n16141), .A(n12288), .B(n12318), .ZN(
        n12289) );
  OAI21_X1 U15259 ( .B1(n12315), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12289), .ZN(
        n14596) );
  MUX2_X1 U15260 ( .A(n12327), .B(n12318), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12291) );
  NAND2_X1 U15261 ( .A1(n14340), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12290) );
  NAND2_X1 U15262 ( .A1(n12291), .A2(n12290), .ZN(n14543) );
  MUX2_X1 U15263 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12292) );
  OAI21_X1 U15264 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14341), .A(
        n12292), .ZN(n14590) );
  INV_X1 U15265 ( .A(n14590), .ZN(n12293) );
  MUX2_X1 U15266 ( .A(n14343), .B(n12312), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12295) );
  INV_X1 U15267 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14950) );
  NOR2_X1 U15268 ( .A1(n13619), .A2(n14950), .ZN(n12294) );
  NOR2_X1 U15269 ( .A1(n12295), .A2(n12294), .ZN(n14535) );
  MUX2_X1 U15270 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12296) );
  OAI21_X1 U15271 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14341), .A(
        n12296), .ZN(n14577) );
  OR2_X2 U15272 ( .A1(n9878), .A2(n14577), .ZN(n14579) );
  INV_X1 U15273 ( .A(n12315), .ZN(n12297) );
  INV_X1 U15274 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21336) );
  NAND2_X1 U15275 ( .A1(n12297), .A2(n21336), .ZN(n12300) );
  INV_X1 U15276 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14918) );
  NAND2_X1 U15277 ( .A1(n13619), .A2(n21336), .ZN(n12298) );
  OAI211_X1 U15278 ( .C1(n14343), .C2(n14918), .A(n12298), .B(n12318), .ZN(
        n12299) );
  AND2_X1 U15279 ( .A1(n12300), .A2(n12299), .ZN(n14504) );
  MUX2_X1 U15280 ( .A(n12327), .B(n12318), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12302) );
  NAND2_X1 U15281 ( .A1(n14340), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U15282 ( .A1(n12302), .A2(n12301), .ZN(n14522) );
  NAND2_X1 U15283 ( .A1(n14504), .A2(n14522), .ZN(n12303) );
  NOR2_X2 U15284 ( .A1(n14579), .A2(n12303), .ZN(n14506) );
  INV_X1 U15285 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14909) );
  NAND2_X1 U15286 ( .A1(n12318), .A2(n14909), .ZN(n12305) );
  INV_X1 U15287 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21479) );
  NAND2_X1 U15288 ( .A1(n13619), .A2(n21479), .ZN(n12304) );
  NAND3_X1 U15289 ( .A1(n12305), .A2(n12327), .A3(n12304), .ZN(n12307) );
  NAND2_X1 U15290 ( .A1(n14343), .A2(n21479), .ZN(n12306) );
  NAND2_X1 U15291 ( .A1(n12307), .A2(n12306), .ZN(n14500) );
  MUX2_X1 U15292 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12311) );
  INV_X1 U15293 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U15294 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  NAND2_X1 U15295 ( .A1(n12311), .A2(n12310), .ZN(n14487) );
  OR2_X2 U15296 ( .A1(n14499), .A2(n14487), .ZN(n14488) );
  MUX2_X1 U15297 ( .A(n14343), .B(n12312), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12314) );
  INV_X1 U15298 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14888) );
  NOR2_X1 U15299 ( .A1(n13619), .A2(n14888), .ZN(n12313) );
  NOR2_X1 U15300 ( .A1(n12314), .A2(n12313), .ZN(n14473) );
  MUX2_X1 U15301 ( .A(n12315), .B(n12327), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12316) );
  OAI21_X1 U15302 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14341), .A(
        n12316), .ZN(n12317) );
  INV_X1 U15303 ( .A(n12317), .ZN(n14451) );
  INV_X1 U15304 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U15305 ( .A1(n12318), .A2(n14862), .ZN(n12320) );
  INV_X1 U15306 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U15307 ( .A1(n13619), .A2(n14571), .ZN(n12319) );
  NAND3_X1 U15308 ( .A1(n12320), .A2(n12327), .A3(n12319), .ZN(n12322) );
  NAND2_X1 U15309 ( .A1(n14343), .A2(n14571), .ZN(n12321) );
  NAND2_X1 U15310 ( .A1(n12322), .A2(n12321), .ZN(n14442) );
  OR2_X1 U15311 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12324) );
  INV_X1 U15312 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U15313 ( .A1(n13619), .A2(n12323), .ZN(n12325) );
  NAND2_X1 U15314 ( .A1(n12324), .A2(n12325), .ZN(n12326) );
  MUX2_X1 U15315 ( .A(n12326), .B(n12325), .S(n14343), .Z(n14432) );
  OAI22_X1 U15316 ( .A1(n14431), .A2(n12327), .B1(n12326), .B2(n9850), .ZN(
        n12330) );
  NAND2_X1 U15317 ( .A1(n14341), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12329) );
  NAND2_X1 U15318 ( .A1(n14340), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12328) );
  NAND2_X1 U15319 ( .A1(n12329), .A2(n12328), .ZN(n14342) );
  XNOR2_X1 U15320 ( .A(n12330), .B(n14342), .ZN(n14842) );
  OR2_X2 U15321 ( .A1(n14600), .A2(n20478), .ZN(n14613) );
  INV_X1 U15322 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21192) );
  NOR2_X1 U15323 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12335) );
  NOR4_X1 U15324 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12334) );
  NAND4_X1 U15325 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12335), .A4(n12334), .ZN(n12358) );
  NOR4_X1 U15326 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12339) );
  NOR4_X1 U15327 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12338) );
  NOR4_X1 U15328 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12337) );
  NOR4_X1 U15329 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12336) );
  AND4_X1 U15330 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12344) );
  NOR4_X1 U15331 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12342) );
  NOR4_X1 U15332 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12341) );
  NOR4_X1 U15333 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12340) );
  INV_X1 U15334 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21046) );
  AND4_X1 U15335 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n21046), .ZN(
        n12343) );
  NAND2_X1 U15336 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  INV_X1 U15337 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21223) );
  INV_X1 U15338 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21465) );
  NOR4_X1 U15339 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21223), .A4(n21465), .ZN(n12347) );
  NOR4_X1 U15340 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12346)
         );
  NAND3_X1 U15341 ( .A1(n20415), .A2(n12347), .A3(n12346), .ZN(U214) );
  NOR4_X1 U15342 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12351) );
  NOR4_X1 U15343 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12350) );
  NOR4_X1 U15344 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12349) );
  NOR4_X1 U15345 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15346 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12356) );
  NOR4_X1 U15347 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12354) );
  NOR4_X1 U15348 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12353) );
  NOR4_X1 U15349 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12352) );
  INV_X1 U15350 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20102) );
  NAND4_X1 U15351 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n20102), .ZN(
        n12355) );
  NOR2_X1 U15352 ( .A1(n15125), .A2(n12358), .ZN(n16633) );
  NAND2_X1 U15353 ( .A1(n16633), .A2(U214), .ZN(U212) );
  AOI21_X1 U15354 ( .B1(n16407), .B2(n12365), .A(n15938), .ZN(n16391) );
  AOI21_X1 U15355 ( .B1(n19252), .B2(n12363), .A(n9930), .ZN(n19256) );
  AOI21_X1 U15356 ( .B1(n19273), .B2(n12362), .A(n12364), .ZN(n19277) );
  AOI21_X1 U15357 ( .B1(n19295), .B2(n12360), .A(n9865), .ZN(n19301) );
  AOI21_X1 U15358 ( .B1(n14995), .B2(n12359), .A(n12361), .ZN(n14992) );
  OAI22_X1 U15359 ( .A1(n20218), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19359) );
  INV_X1 U15360 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19334) );
  OAI22_X1 U15361 ( .A1(n20218), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19334), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15659) );
  AND2_X1 U15362 ( .A1(n19359), .A2(n15659), .ZN(n15011) );
  OAI21_X1 U15363 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12359), .ZN(n19502) );
  NAND2_X1 U15364 ( .A1(n15011), .A2(n19502), .ZN(n14990) );
  NOR2_X1 U15365 ( .A1(n14992), .A2(n14990), .ZN(n19314) );
  OAI21_X1 U15366 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12361), .A(
        n12360), .ZN(n19499) );
  NAND2_X1 U15367 ( .A1(n19314), .A2(n19499), .ZN(n19299) );
  NOR2_X1 U15368 ( .A1(n19301), .A2(n19299), .ZN(n19282) );
  OAI21_X1 U15369 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9865), .A(
        n12362), .ZN(n19283) );
  NAND2_X1 U15370 ( .A1(n19282), .A2(n19283), .ZN(n19275) );
  NOR2_X1 U15371 ( .A1(n19277), .A2(n19275), .ZN(n19264) );
  OAI21_X1 U15372 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12364), .A(
        n12363), .ZN(n19265) );
  NAND2_X1 U15373 ( .A1(n19264), .A2(n19265), .ZN(n19254) );
  NOR2_X1 U15374 ( .A1(n19256), .A2(n19254), .ZN(n19243) );
  OAI21_X1 U15375 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9930), .A(
        n12365), .ZN(n19244) );
  NAND2_X1 U15376 ( .A1(n19243), .A2(n19244), .ZN(n12366) );
  NOR2_X1 U15377 ( .A1(n16391), .A2(n12366), .ZN(n19233) );
  INV_X1 U15378 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14231) );
  INV_X1 U15379 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16321) );
  INV_X1 U15380 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16345) );
  INV_X1 U15381 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n19127) );
  INV_X1 U15382 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15332) );
  INV_X1 U15383 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15350) );
  INV_X1 U15384 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U15385 ( .A1(n19303), .A2(n15010), .ZN(n19358) );
  AOI211_X1 U15386 ( .C1(n16391), .C2(n12366), .A(n19233), .B(n19358), .ZN(
        n12556) );
  INV_X1 U15387 ( .A(n12368), .ZN(n12370) );
  NOR3_X1 U15388 ( .A1(n12370), .A2(n12389), .A3(n12369), .ZN(n12557) );
  NAND2_X1 U15389 ( .A1(n12371), .A2(n12557), .ZN(n12372) );
  INV_X1 U15390 ( .A(n12632), .ZN(n12373) );
  INV_X2 U15391 ( .A(n20230), .ZN(n20148) );
  NAND2_X2 U15392 ( .A1(n20148), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20146) );
  NOR2_X1 U15393 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20091) );
  INV_X1 U15394 ( .A(n20091), .ZN(n20084) );
  NAND2_X1 U15395 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20216) );
  NAND2_X1 U15396 ( .A1(n20224), .A2(n20216), .ZN(n12594) );
  NOR2_X1 U15397 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12594), .ZN(n12464) );
  OR2_X1 U15398 ( .A1(n12745), .A2(n12464), .ZN(n16259) );
  INV_X1 U15399 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n12714) );
  NAND2_X1 U15400 ( .A1(n12714), .A2(n20216), .ZN(n12374) );
  NAND2_X1 U15401 ( .A1(n12638), .A2(n12374), .ZN(n12463) );
  OR2_X1 U15402 ( .A1(n12463), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12375) );
  AND2_X1 U15403 ( .A1(n12376), .A2(n12632), .ZN(n20214) );
  NAND2_X1 U15404 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20013), .ZN(n20075) );
  NOR2_X1 U15405 ( .A1(n20078), .A2(n20075), .ZN(n16542) );
  AND2_X2 U15406 ( .A1(n20169), .A2(n16499), .ZN(n19310) );
  OR2_X1 U15407 ( .A1(n19310), .A2(n19303), .ZN(n12377) );
  OR2_X1 U15408 ( .A1(n16542), .A2(n12377), .ZN(n12378) );
  NOR2_X2 U15409 ( .A1(n19323), .A2(n12466), .ZN(n19324) );
  OAI22_X1 U15410 ( .A1(n19343), .A2(n11122), .B1(n16407), .B2(n19353), .ZN(
        n12555) );
  INV_X1 U15411 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20112) );
  AOI22_X1 U15412 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12416), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15413 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15414 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12481), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15415 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10732), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15416 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12388) );
  AOI22_X1 U15417 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15418 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15419 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15420 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12491), .ZN(n12383) );
  NAND4_X1 U15421 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12387) );
  INV_X1 U15422 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12390) );
  NAND2_X1 U15423 ( .A1(n12391), .A2(n12390), .ZN(n12403) );
  AOI22_X1 U15424 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12416), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15425 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15426 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12479), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15427 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10732), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12392) );
  NAND4_X1 U15428 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12401) );
  AOI22_X1 U15429 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12490), .B1(
        n12488), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15430 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15431 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10780), .B1(
        n10747), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15432 ( .A1(n12487), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12491), .ZN(n12396) );
  NAND4_X1 U15433 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  MUX2_X1 U15434 ( .A(n12403), .B(n12723), .S(n14208), .Z(n12827) );
  AOI22_X1 U15435 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12416), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15436 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12481), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15437 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12479), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15438 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10732), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12404) );
  NAND4_X1 U15439 ( .A1(n12407), .A2(n12406), .A3(n12405), .A4(n12404), .ZN(
        n12413) );
  AOI22_X1 U15440 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15441 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15442 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15443 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12491), .ZN(n12408) );
  NAND4_X1 U15444 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12412) );
  MUX2_X1 U15445 ( .A(n13511), .B(n12414), .S(n12581), .Z(n12586) );
  MUX2_X1 U15446 ( .A(n12586), .B(n14996), .S(n19547), .Z(n13545) );
  INV_X1 U15447 ( .A(n12587), .ZN(n12415) );
  MUX2_X1 U15448 ( .A(n12415), .B(P2_EBX_REG_4__SCAN_IN), .S(n19547), .Z(
        n13578) );
  NOR2_X2 U15449 ( .A1(n13579), .A2(n13578), .ZN(n13824) );
  INV_X1 U15450 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U15451 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15452 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15453 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15454 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12417) );
  NAND4_X1 U15455 ( .A1(n12420), .A2(n12419), .A3(n12418), .A4(n12417), .ZN(
        n12426) );
  AOI22_X1 U15456 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15457 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15458 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15459 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15460 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12425) );
  MUX2_X1 U15461 ( .A(n14084), .B(n13814), .S(n14208), .Z(n13823) );
  INV_X1 U15462 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U15463 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12478), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15464 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15465 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12481), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15466 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12482), .B1(
        n10732), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12427) );
  NAND4_X1 U15467 ( .A1(n12430), .A2(n12429), .A3(n12428), .A4(n12427), .ZN(
        n12436) );
  AOI22_X1 U15468 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12488), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15469 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15470 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12490), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15471 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12491), .ZN(n12431) );
  NAND4_X1 U15472 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12435) );
  MUX2_X1 U15473 ( .A(n13097), .B(n13858), .S(n14208), .Z(n13865) );
  NAND2_X1 U15474 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12440) );
  NAND2_X1 U15475 ( .A1(n12477), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12439) );
  NAND2_X1 U15476 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12438) );
  NAND2_X1 U15477 ( .A1(n12479), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12437) );
  NAND2_X1 U15478 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12444) );
  NAND2_X1 U15479 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12443) );
  NAND2_X1 U15480 ( .A1(n12487), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12442) );
  NAND2_X1 U15481 ( .A1(n12491), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12441) );
  NAND2_X1 U15482 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12448) );
  NAND2_X1 U15483 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12447) );
  NAND2_X1 U15484 ( .A1(n11087), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12446) );
  NAND2_X1 U15485 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12445) );
  NAND2_X1 U15486 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12452) );
  NAND2_X1 U15487 ( .A1(n12480), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12451) );
  NAND2_X1 U15488 ( .A1(n12482), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12450) );
  NAND2_X1 U15489 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12449) );
  NAND4_X1 U15490 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12457) );
  MUX2_X1 U15491 ( .A(n12458), .B(n12457), .S(n14208), .Z(n13924) );
  INV_X1 U15492 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12459) );
  INV_X1 U15493 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U15494 ( .A1(n14204), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12460) );
  OR2_X1 U15495 ( .A1(n14109), .A2(n12460), .ZN(n12462) );
  INV_X1 U15496 ( .A(n14112), .ZN(n12461) );
  INV_X1 U15497 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16260) );
  AND2_X1 U15498 ( .A1(n9839), .A2(n20217), .ZN(n12591) );
  AND2_X1 U15499 ( .A1(n12591), .A2(n12464), .ZN(n12465) );
  AND2_X1 U15500 ( .A1(n12575), .A2(n12465), .ZN(n16501) );
  AND2_X2 U15501 ( .A1(n12468), .A2(n14208), .ZN(n13966) );
  AOI22_X1 U15502 ( .A1(n14399), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n13966), 
        .B2(n12469), .ZN(n12472) );
  AND2_X1 U15503 ( .A1(n19565), .A2(n12466), .ZN(n12470) );
  AND2_X2 U15504 ( .A1(n9833), .A2(n12466), .ZN(n12504) );
  AOI22_X1 U15505 ( .A1(n14398), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12471) );
  INV_X2 U15506 ( .A(n12503), .ZN(n14398) );
  AOI222_X1 U15507 ( .A1(n14399), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n14398), 
        .B2(P2_EAX_REG_7__SCAN_IN), .C1(n12504), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13933) );
  INV_X1 U15508 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15509 ( .A1(n14398), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12504), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U15510 ( .A1(n13966), .A2(n13814), .ZN(n12474) );
  OAI211_X1 U15511 ( .C1(n12473), .C2(n12476), .A(n12475), .B(n12474), .ZN(
        n16482) );
  AOI22_X1 U15512 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12477), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15513 ( .A1(n12416), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15514 ( .A1(n12481), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12480), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15515 ( .A1(n10732), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12482), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12483) );
  NAND4_X1 U15516 ( .A1(n12486), .A2(n12485), .A3(n12484), .A4(n12483), .ZN(
        n12497) );
  AOI22_X1 U15517 ( .A1(n12488), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12487), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15518 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15519 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11087), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15520 ( .A1(n10747), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12491), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12492) );
  NAND4_X1 U15521 ( .A1(n12495), .A2(n12494), .A3(n12493), .A4(n12492), .ZN(
        n12496) );
  NAND2_X1 U15522 ( .A1(n13966), .A2(n12722), .ZN(n12499) );
  INV_X1 U15523 ( .A(n12507), .ZN(n13949) );
  NAND2_X1 U15524 ( .A1(n13949), .A2(n9841), .ZN(n12515) );
  NAND2_X1 U15525 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12498) );
  NAND4_X1 U15526 ( .A1(n12499), .A2(n12503), .A3(n12515), .A4(n12498), .ZN(
        n12622) );
  INV_X1 U15527 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19341) );
  AOI21_X1 U15528 ( .B1(n9833), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U15529 ( .A1(n19565), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12500) );
  AND2_X1 U15530 ( .A1(n12501), .A2(n12500), .ZN(n12502) );
  NAND2_X1 U15531 ( .A1(n12622), .A2(n12621), .ZN(n12511) );
  NAND2_X1 U15532 ( .A1(n14399), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15533 ( .A1(n12470), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9842), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12505) );
  XNOR2_X1 U15534 ( .A(n12511), .B(n12512), .ZN(n12780) );
  NAND2_X1 U15535 ( .A1(n12507), .A2(n12569), .ZN(n12508) );
  MUX2_X1 U15536 ( .A(n12508), .B(n20190), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12510) );
  NAND2_X1 U15537 ( .A1(n13966), .A2(n12847), .ZN(n12509) );
  NAND2_X1 U15538 ( .A1(n12510), .A2(n12509), .ZN(n12779) );
  NAND2_X1 U15539 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND2_X1 U15540 ( .A1(n12782), .A2(n12513), .ZN(n12521) );
  NAND2_X1 U15541 ( .A1(n13966), .A2(n12514), .ZN(n12516) );
  OAI211_X1 U15542 ( .C1(n12466), .C2(n20181), .A(n12516), .B(n12515), .ZN(
        n12520) );
  XNOR2_X1 U15543 ( .A(n12521), .B(n12520), .ZN(n12836) );
  NAND2_X1 U15544 ( .A1(n14399), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15545 ( .A1(n14398), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12504), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12518) );
  AND2_X1 U15546 ( .A1(n12519), .A2(n12518), .ZN(n12835) );
  INV_X1 U15547 ( .A(n12520), .ZN(n12522) );
  NAND2_X1 U15548 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  INV_X1 U15549 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13568) );
  NOR2_X1 U15550 ( .A1(n10685), .A2(n12466), .ZN(n12524) );
  AOI21_X1 U15551 ( .B1(n12504), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12524), .ZN(n12526) );
  NAND2_X1 U15552 ( .A1(n14398), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12525) );
  AND2_X1 U15553 ( .A1(n12526), .A2(n12525), .ZN(n12528) );
  NAND2_X1 U15554 ( .A1(n13966), .A2(n13511), .ZN(n12527) );
  OAI211_X1 U15555 ( .C1(n12473), .C2(n13568), .A(n12528), .B(n12527), .ZN(
        n13555) );
  INV_X1 U15556 ( .A(n13555), .ZN(n12529) );
  INV_X1 U15557 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15558 ( .A1(n14398), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12504), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U15559 ( .A1(n13966), .A2(n13782), .ZN(n12530) );
  OAI211_X1 U15560 ( .C1(n12473), .C2(n12532), .A(n12531), .B(n12530), .ZN(
        n13591) );
  NAND2_X1 U15561 ( .A1(n16482), .A2(n16481), .ZN(n16484) );
  NAND2_X1 U15562 ( .A1(n13966), .A2(n13858), .ZN(n12533) );
  INV_X1 U15563 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U15564 ( .A1(n14398), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12504), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12534) );
  OAI21_X1 U15565 ( .B1(n12473), .B2(n12535), .A(n12534), .ZN(n13892) );
  AOI21_X1 U15566 ( .B1(n13966), .B2(n14183), .A(n13895), .ZN(n13934) );
  INV_X1 U15567 ( .A(n13966), .ZN(n13959) );
  AOI22_X1 U15568 ( .A1(n14398), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12504), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U15569 ( .A1(n14399), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12536) );
  OAI211_X1 U15570 ( .C1(n13959), .C2(n13343), .A(n12537), .B(n12536), .ZN(
        n16468) );
  NOR2_X1 U15571 ( .A1(n12517), .A2(n15643), .ZN(n12540) );
  INV_X1 U15572 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12538) );
  OAI22_X1 U15573 ( .A1(n13959), .A2(n13372), .B1(n12538), .B2(n12473), .ZN(
        n12539) );
  AOI211_X1 U15574 ( .C1(P2_EAX_REG_9__SCAN_IN), .C2(n14398), .A(n12540), .B(
        n12539), .ZN(n15639) );
  INV_X1 U15575 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15576 ( .A1(n14398), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15577 ( .A1(n13966), .A2(n13433), .ZN(n12541) );
  OAI211_X1 U15578 ( .C1(n12473), .C2(n12543), .A(n12542), .B(n12541), .ZN(
        n15623) );
  AOI21_X1 U15579 ( .B1(n12544), .B2(n15624), .A(n9933), .ZN(n19380) );
  AOI22_X1 U15580 ( .A1(n14118), .A2(n19346), .B1(n19333), .B2(n19380), .ZN(
        n12545) );
  OAI211_X1 U15581 ( .C1(n20112), .C2(n19342), .A(n12545), .B(n19294), .ZN(
        n12554) );
  INV_X1 U15582 ( .A(n12546), .ZN(n13610) );
  INV_X1 U15583 ( .A(n12547), .ZN(n12549) );
  INV_X1 U15584 ( .A(n13435), .ZN(n12548) );
  NAND2_X1 U15585 ( .A1(n12549), .A2(n12548), .ZN(n12550) );
  NAND2_X1 U15586 ( .A1(n13610), .A2(n12550), .ZN(n16401) );
  AND2_X1 U15587 ( .A1(n9833), .A2(n20216), .ZN(n12551) );
  INV_X1 U15588 ( .A(n16391), .ZN(n12552) );
  INV_X1 U15589 ( .A(n19335), .ZN(n19352) );
  OAI22_X1 U15590 ( .A1(n16401), .A2(n19349), .B1(n12552), .B2(n19352), .ZN(
        n12553) );
  OR4_X1 U15591 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        P2_U2844) );
  INV_X1 U15592 ( .A(n12557), .ZN(n12558) );
  OAI21_X1 U15593 ( .B1(n12559), .B2(n12558), .A(n16529), .ZN(n12561) );
  AOI21_X1 U15594 ( .B1(n13012), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16522) );
  AOI21_X1 U15595 ( .B1(n12560), .B2(n16522), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n20192) );
  MUX2_X1 U15596 ( .A(n12561), .B(n20192), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20205) );
  INV_X1 U15597 ( .A(n20205), .ZN(n16544) );
  NOR2_X1 U15598 ( .A1(n16527), .A2(n9838), .ZN(n12562) );
  NAND2_X1 U15599 ( .A1(n16544), .A2(n12562), .ZN(n12602) );
  AND2_X1 U15600 ( .A1(n12564), .A2(n12563), .ZN(n12574) );
  OAI21_X1 U15601 ( .B1(n12565), .B2(n19565), .A(n12591), .ZN(n12610) );
  NAND2_X1 U15602 ( .A1(n12566), .A2(n10618), .ZN(n12567) );
  NAND2_X1 U15603 ( .A1(n12567), .A2(n15745), .ZN(n12573) );
  NAND2_X1 U15604 ( .A1(n9838), .A2(n12568), .ZN(n12604) );
  NAND2_X1 U15605 ( .A1(n12604), .A2(n16528), .ZN(n12570) );
  NAND2_X1 U15606 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  NAND2_X1 U15607 ( .A1(n12571), .A2(n10618), .ZN(n12572) );
  NAND4_X1 U15608 ( .A1(n12574), .A2(n12610), .A3(n12573), .A4(n12572), .ZN(
        n12605) );
  INV_X1 U15609 ( .A(n12605), .ZN(n12577) );
  INV_X1 U15610 ( .A(n12594), .ZN(n16519) );
  NAND3_X1 U15611 ( .A1(n12575), .A2(n16529), .A3(n16519), .ZN(n12576) );
  NAND2_X1 U15612 ( .A1(n12577), .A2(n12576), .ZN(n13023) );
  NAND3_X1 U15613 ( .A1(n16529), .A2(n13943), .A3(n20216), .ZN(n12578) );
  AOI21_X1 U15614 ( .B1(n12579), .B2(n9833), .A(n12578), .ZN(n12580) );
  NOR2_X1 U15615 ( .A1(n13023), .A2(n12580), .ZN(n12593) );
  MUX2_X1 U15616 ( .A(n12722), .B(n12582), .S(n12581), .Z(n12623) );
  NAND2_X1 U15617 ( .A1(n12623), .A2(n12583), .ZN(n12585) );
  NAND2_X1 U15618 ( .A1(n12585), .A2(n12584), .ZN(n12588) );
  NAND3_X1 U15619 ( .A1(n12588), .A2(n12587), .A3(n12586), .ZN(n12590) );
  AND2_X1 U15620 ( .A1(n12590), .A2(n12589), .ZN(n20201) );
  INV_X1 U15621 ( .A(n12591), .ZN(n12592) );
  NOR2_X1 U15622 ( .A1(n16527), .A2(n12592), .ZN(n20203) );
  NAND2_X1 U15623 ( .A1(n20201), .A2(n20203), .ZN(n12704) );
  AND2_X1 U15624 ( .A1(n12593), .A2(n12704), .ZN(n12601) );
  NAND2_X1 U15625 ( .A1(n13028), .A2(n9833), .ZN(n13030) );
  INV_X1 U15626 ( .A(n13030), .ZN(n12596) );
  NOR2_X1 U15627 ( .A1(n10618), .A2(n12594), .ZN(n12595) );
  NAND2_X1 U15628 ( .A1(n12596), .A2(n12595), .ZN(n12600) );
  AOI21_X1 U15629 ( .B1(n12597), .B2(n16528), .A(n19541), .ZN(n12598) );
  NAND2_X1 U15630 ( .A1(n13030), .A2(n12598), .ZN(n12599) );
  NAND4_X1 U15631 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12603) );
  NAND2_X1 U15632 ( .A1(n12627), .A2(n16533), .ZN(n15512) );
  NAND2_X1 U15633 ( .A1(n12606), .A2(n13026), .ZN(n12608) );
  NAND2_X1 U15634 ( .A1(n12608), .A2(n12607), .ZN(n12617) );
  NAND2_X1 U15635 ( .A1(n12609), .A2(n9833), .ZN(n15649) );
  NAND2_X1 U15636 ( .A1(n15649), .A2(n12610), .ZN(n12615) );
  OAI22_X1 U15637 ( .A1(n13026), .A2(n19541), .B1(n10618), .B2(n16528), .ZN(
        n12611) );
  INV_X1 U15638 ( .A(n12611), .ZN(n12612) );
  AOI21_X1 U15639 ( .B1(n12615), .B2(n12614), .A(n12613), .ZN(n12616) );
  NAND2_X1 U15640 ( .A1(n12617), .A2(n12616), .ZN(n15652) );
  OR2_X1 U15641 ( .A1(n15652), .A2(n11111), .ZN(n12618) );
  NAND2_X1 U15642 ( .A1(n12627), .A2(n12618), .ZN(n15519) );
  NOR2_X1 U15643 ( .A1(n12627), .A2(n19310), .ZN(n13562) );
  MUX2_X1 U15644 ( .A(n15517), .B(n13562), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n12631) );
  AND2_X1 U15645 ( .A1(n9839), .A2(n12722), .ZN(n12848) );
  INV_X1 U15646 ( .A(n12848), .ZN(n12619) );
  NAND2_X1 U15647 ( .A1(n12619), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12842) );
  OAI21_X1 U15648 ( .B1(n12619), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12842), .ZN(n12711) );
  INV_X1 U15649 ( .A(n12376), .ZN(n16530) );
  INV_X1 U15650 ( .A(n13018), .ZN(n16531) );
  OAI21_X1 U15651 ( .B1(n9839), .B2(n16530), .A(n16531), .ZN(n12620) );
  OAI21_X1 U15652 ( .B1(n12622), .B2(n12621), .A(n12511), .ZN(n19398) );
  OAI22_X1 U15653 ( .A1(n16457), .A2(n12711), .B1(n16469), .B2(n19398), .ZN(
        n12630) );
  MUX2_X1 U15654 ( .A(n12623), .B(P2_EBX_REG_0__SCAN_IN), .S(n19547), .Z(
        n19347) );
  NAND2_X1 U15655 ( .A1(n19347), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12824) );
  OAI21_X1 U15656 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19347), .A(
        n12824), .ZN(n12709) );
  INV_X1 U15657 ( .A(n16527), .ZN(n12625) );
  NAND2_X1 U15658 ( .A1(n12625), .A2(n12624), .ZN(n12705) );
  INV_X1 U15659 ( .A(n12705), .ZN(n20204) );
  NAND2_X1 U15660 ( .A1(n12627), .A2(n12626), .ZN(n15640) );
  INV_X1 U15661 ( .A(n19350), .ZN(n15653) );
  NAND2_X1 U15662 ( .A1(n16492), .A2(n15653), .ZN(n12628) );
  NAND2_X1 U15663 ( .A1(n19310), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12710) );
  OAI211_X1 U15664 ( .C1(n12709), .C2(n16477), .A(n12628), .B(n12710), .ZN(
        n12629) );
  OR3_X1 U15665 ( .A1(n12631), .A2(n12630), .A3(n12629), .ZN(P2_U3046) );
  INV_X1 U15666 ( .A(n15745), .ZN(n16524) );
  AND2_X1 U15667 ( .A1(n12632), .A2(n16524), .ZN(n19356) );
  INV_X1 U15668 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12634) );
  INV_X1 U15669 ( .A(n12638), .ZN(n12633) );
  NAND2_X1 U15670 ( .A1(n20169), .A2(n20079), .ZN(n19103) );
  OAI211_X1 U15671 ( .C1(n19356), .C2(n12634), .A(n12633), .B(n19103), .ZN(
        P2_U2814) );
  INV_X1 U15672 ( .A(n13026), .ZN(n12637) );
  INV_X1 U15673 ( .A(n19103), .ZN(n12635) );
  NOR4_X1 U15674 ( .A1(n12638), .A2(n19356), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .A4(n12635), .ZN(n12636) );
  AOI21_X1 U15675 ( .B1(n20214), .B2(n12637), .A(n12636), .ZN(P2_U3612) );
  INV_X1 U15676 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12641) );
  INV_X1 U15677 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12640) );
  OAI21_X1 U15678 ( .B1(n9838), .B2(n20216), .A(n12638), .ZN(n19483) );
  INV_X1 U15679 ( .A(n19483), .ZN(n12659) );
  INV_X1 U15680 ( .A(n19481), .ZN(n12639) );
  AOI22_X1 U15681 ( .A1(n13971), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15125), .ZN(n19371) );
  OAI222_X1 U15682 ( .A1(n12745), .A2(n12641), .B1(n12640), .B2(n12659), .C1(
        n12639), .C2(n19371), .ZN(P2_U2982) );
  NOR4_X1 U15683 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12647) );
  NOR2_X1 U15684 ( .A1(n12648), .A2(n12647), .ZN(n12917) );
  AND2_X1 U15685 ( .A1(n12917), .A2(n13627), .ZN(n12649) );
  NAND2_X1 U15686 ( .A1(n12908), .A2(n12649), .ZN(n12701) );
  INV_X1 U15687 ( .A(n12701), .ZN(n12651) );
  INV_X1 U15688 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21324) );
  INV_X1 U15689 ( .A(n13627), .ZN(n20235) );
  NOR2_X2 U15690 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20842) );
  NAND2_X1 U15691 ( .A1(n20842), .A2(n21025), .ZN(n20238) );
  OAI211_X1 U15692 ( .C1(n12651), .C2(n21324), .A(n12867), .B(n20238), .ZN(
        P1_U2801) );
  INV_X2 U15693 ( .A(n12745), .ZN(n19487) );
  AOI22_X1 U15694 ( .A1(n19487), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19483), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15695 ( .A1(n13971), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15125), .ZN(n19531) );
  INV_X1 U15696 ( .A(n19531), .ZN(n15210) );
  NAND2_X1 U15697 ( .A1(n19481), .A2(n15210), .ZN(n12697) );
  NAND2_X1 U15698 ( .A1(n12652), .A2(n12697), .ZN(P2_U2954) );
  AOI22_X1 U15699 ( .A1(n19487), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n19483), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15700 ( .A1(n13971), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15125), .ZN(n19535) );
  INV_X1 U15701 ( .A(n19535), .ZN(n14026) );
  NAND2_X1 U15702 ( .A1(n19481), .A2(n14026), .ZN(n12668) );
  NAND2_X1 U15703 ( .A1(n12653), .A2(n12668), .ZN(P2_U2970) );
  AOI22_X1 U15704 ( .A1(n19487), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n19483), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15705 ( .A1(n13971), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n15125), .ZN(n19377) );
  INV_X1 U15706 ( .A(n19377), .ZN(n15137) );
  NAND2_X1 U15707 ( .A1(n19481), .A2(n15137), .ZN(n12682) );
  NAND2_X1 U15708 ( .A1(n12654), .A2(n12682), .ZN(P2_U2964) );
  AOI22_X1 U15709 ( .A1(n19487), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n19483), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15710 ( .A1(n13971), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15125), .ZN(n19435) );
  INV_X1 U15711 ( .A(n19435), .ZN(n14002) );
  NAND2_X1 U15712 ( .A1(n19481), .A2(n14002), .ZN(n12692) );
  NAND2_X1 U15713 ( .A1(n12655), .A2(n12692), .ZN(P2_U2967) );
  AOI22_X1 U15714 ( .A1(n19487), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n19483), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15715 ( .A1(n13971), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15125), .ZN(n19526) );
  INV_X1 U15716 ( .A(n19526), .ZN(n13972) );
  NAND2_X1 U15717 ( .A1(n19481), .A2(n13972), .ZN(n12670) );
  NAND2_X1 U15718 ( .A1(n12656), .A2(n12670), .ZN(P2_U2968) );
  INV_X1 U15719 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19456) );
  NAND2_X1 U15720 ( .A1(n15125), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12658) );
  INV_X1 U15721 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16666) );
  OR2_X1 U15722 ( .A1(n15125), .A2(n16666), .ZN(n12657) );
  NAND2_X1 U15723 ( .A1(n12658), .A2(n12657), .ZN(n19385) );
  NAND2_X1 U15724 ( .A1(n19481), .A2(n19385), .ZN(n12667) );
  NAND2_X1 U15725 ( .A1(n19486), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12660) );
  OAI211_X1 U15726 ( .C1(n19456), .C2(n12745), .A(n12667), .B(n12660), .ZN(
        P2_U2976) );
  INV_X1 U15727 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19452) );
  NAND2_X1 U15728 ( .A1(n15125), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12662) );
  INV_X1 U15729 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16662) );
  OR2_X1 U15730 ( .A1(n15125), .A2(n16662), .ZN(n12661) );
  NAND2_X1 U15731 ( .A1(n12662), .A2(n12661), .ZN(n19379) );
  NAND2_X1 U15732 ( .A1(n19481), .A2(n19379), .ZN(n12665) );
  NAND2_X1 U15733 ( .A1(n19486), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12663) );
  OAI211_X1 U15734 ( .C1(n19452), .C2(n12745), .A(n12665), .B(n12663), .ZN(
        P2_U2978) );
  INV_X1 U15735 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U15736 ( .A1(n19486), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12664) );
  OAI211_X1 U15737 ( .C1(n12753), .C2(n12745), .A(n12665), .B(n12664), .ZN(
        P2_U2963) );
  INV_X1 U15738 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U15739 ( .A1(n19486), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12666) );
  OAI211_X1 U15740 ( .C1(n12767), .C2(n12745), .A(n12667), .B(n12666), .ZN(
        P2_U2961) );
  AOI22_X1 U15741 ( .A1(n19487), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n12669) );
  NAND2_X1 U15742 ( .A1(n12669), .A2(n12668), .ZN(P2_U2955) );
  AOI22_X1 U15743 ( .A1(n19487), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n12671) );
  NAND2_X1 U15744 ( .A1(n12671), .A2(n12670), .ZN(P2_U2953) );
  AOI22_X1 U15745 ( .A1(n19487), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15746 ( .A1(n13971), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15125), .ZN(n19542) );
  INV_X1 U15747 ( .A(n19542), .ZN(n15202) );
  NAND2_X1 U15748 ( .A1(n19481), .A2(n15202), .ZN(n12688) );
  NAND2_X1 U15749 ( .A1(n12672), .A2(n12688), .ZN(P2_U2971) );
  AOI22_X1 U15750 ( .A1(n19487), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15751 ( .A1(n13971), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15125), .ZN(n19555) );
  INV_X1 U15752 ( .A(n19555), .ZN(n15179) );
  NAND2_X1 U15753 ( .A1(n19481), .A2(n15179), .ZN(n12694) );
  NAND2_X1 U15754 ( .A1(n12673), .A2(n12694), .ZN(P2_U2958) );
  AOI22_X1 U15755 ( .A1(n19487), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n12677) );
  INV_X1 U15756 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n12674) );
  OR2_X1 U15757 ( .A1(n15125), .A2(n12674), .ZN(n12676) );
  NAND2_X1 U15758 ( .A1(n15125), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12675) );
  AND2_X1 U15759 ( .A1(n12676), .A2(n12675), .ZN(n19388) );
  INV_X1 U15760 ( .A(n19388), .ZN(n15170) );
  NAND2_X1 U15761 ( .A1(n19481), .A2(n15170), .ZN(n12686) );
  NAND2_X1 U15762 ( .A1(n12677), .A2(n12686), .ZN(P2_U2975) );
  AOI22_X1 U15763 ( .A1(n19487), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15764 ( .A1(n13971), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15125), .ZN(n19549) );
  INV_X1 U15765 ( .A(n19549), .ZN(n15187) );
  NAND2_X1 U15766 ( .A1(n19481), .A2(n15187), .ZN(n12684) );
  NAND2_X1 U15767 ( .A1(n12678), .A2(n12684), .ZN(P2_U2972) );
  AOI22_X1 U15768 ( .A1(n19487), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12681) );
  INV_X1 U15769 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16664) );
  OR2_X1 U15770 ( .A1(n15125), .A2(n16664), .ZN(n12680) );
  NAND2_X1 U15771 ( .A1(n15125), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12679) );
  AND2_X1 U15772 ( .A1(n12680), .A2(n12679), .ZN(n19382) );
  INV_X1 U15773 ( .A(n19382), .ZN(n15153) );
  NAND2_X1 U15774 ( .A1(n19481), .A2(n15153), .ZN(n12690) );
  NAND2_X1 U15775 ( .A1(n12681), .A2(n12690), .ZN(P2_U2977) );
  AOI22_X1 U15776 ( .A1(n19487), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U15777 ( .A1(n12683), .A2(n12682), .ZN(P2_U2979) );
  AOI22_X1 U15778 ( .A1(n19487), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15779 ( .A1(n12685), .A2(n12684), .ZN(P2_U2957) );
  AOI22_X1 U15780 ( .A1(n19487), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U15781 ( .A1(n12687), .A2(n12686), .ZN(P2_U2960) );
  AOI22_X1 U15782 ( .A1(n19487), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12689) );
  NAND2_X1 U15783 ( .A1(n12689), .A2(n12688), .ZN(P2_U2956) );
  AOI22_X1 U15784 ( .A1(n19487), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U15785 ( .A1(n12691), .A2(n12690), .ZN(P2_U2962) );
  AOI22_X1 U15786 ( .A1(n19487), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U15787 ( .A1(n12693), .A2(n12692), .ZN(P2_U2952) );
  AOI22_X1 U15788 ( .A1(n19487), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n12695) );
  NAND2_X1 U15789 ( .A1(n12695), .A2(n12694), .ZN(P2_U2973) );
  AOI22_X1 U15790 ( .A1(n19487), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n12696) );
  OAI22_X1 U15791 ( .A1(n15125), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13971), .ZN(n19567) );
  INV_X1 U15792 ( .A(n19567), .ZN(n16355) );
  NAND2_X1 U15793 ( .A1(n19481), .A2(n16355), .ZN(n12699) );
  NAND2_X1 U15794 ( .A1(n12696), .A2(n12699), .ZN(P2_U2974) );
  AOI22_X1 U15795 ( .A1(n19487), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U15796 ( .A1(n12698), .A2(n12697), .ZN(P2_U2969) );
  AOI22_X1 U15797 ( .A1(n19487), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15798 ( .A1(n12700), .A2(n12699), .ZN(P2_U2959) );
  INV_X1 U15799 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21221) );
  AND2_X1 U15800 ( .A1(n20238), .A2(n21221), .ZN(n12703) );
  OAI21_X1 U15801 ( .B1(n13400), .B2(n14343), .A(n21108), .ZN(n12702) );
  OAI21_X1 U15802 ( .B1(n12703), .B2(n21108), .A(n12702), .ZN(P1_U3487) );
  OAI21_X1 U15803 ( .B1(n20205), .B2(n12705), .A(n12704), .ZN(n12706) );
  NOR2_X1 U15804 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20163) );
  OR2_X1 U15805 ( .A1(n20169), .A2(n20163), .ZN(n20182) );
  NAND2_X1 U15806 ( .A1(n20182), .A2(n20218), .ZN(n12707) );
  AND2_X1 U15807 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20183) );
  INV_X1 U15808 ( .A(n19108), .ZN(n12708) );
  INV_X1 U15809 ( .A(n12709), .ZN(n12713) );
  NOR2_X2 U15810 ( .A1(n19108), .A2(n9833), .ZN(n16449) );
  OAI21_X1 U15811 ( .B1(n19501), .B2(n12711), .A(n12710), .ZN(n12712) );
  AOI21_X1 U15812 ( .B1(n19504), .B2(n12713), .A(n12712), .ZN(n12718) );
  NAND2_X1 U15813 ( .A1(n12714), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U15814 ( .A1(n12716), .A2(n12715), .ZN(n12721) );
  OAI21_X1 U15815 ( .B1(n19490), .B2(n12721), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12717) );
  OAI211_X1 U15816 ( .C1(n16438), .C2(n19350), .A(n12718), .B(n12717), .ZN(
        P2_U3014) );
  INV_X1 U15817 ( .A(n13479), .ZN(n19330) );
  NAND3_X1 U15818 ( .A1(n14204), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15819 ( .A1(n12827), .A2(n12719), .ZN(n19329) );
  NAND2_X1 U15820 ( .A1(n12824), .A2(n19329), .ZN(n12825) );
  OAI21_X1 U15821 ( .B1(n12824), .B2(n19329), .A(n12825), .ZN(n12720) );
  XNOR2_X1 U15822 ( .A(n12720), .B(n15660), .ZN(n12777) );
  OAI22_X1 U15823 ( .A1(n12777), .A2(n19493), .B1(n19503), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12728) );
  INV_X1 U15824 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20099) );
  AND2_X1 U15825 ( .A1(n19310), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12774) );
  NOR2_X1 U15826 ( .A1(n19514), .A2(n19334), .ZN(n12727) );
  XNOR2_X1 U15827 ( .A(n12723), .B(n12722), .ZN(n12843) );
  XNOR2_X1 U15828 ( .A(n12842), .B(n12843), .ZN(n12724) );
  OR2_X1 U15829 ( .A1(n12724), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12725) );
  NAND2_X1 U15830 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12724), .ZN(
        n12845) );
  AND2_X1 U15831 ( .A1(n12725), .A2(n12845), .ZN(n12783) );
  AND2_X1 U15832 ( .A1(n16449), .A2(n12783), .ZN(n12726) );
  NOR4_X1 U15833 ( .A1(n12728), .A2(n12774), .A3(n12727), .A4(n12726), .ZN(
        n12729) );
  OAI21_X1 U15834 ( .B1(n19330), .B2(n16438), .A(n12729), .ZN(P2_U3013) );
  OR2_X1 U15835 ( .A1(n13620), .A2(n13400), .ZN(n12732) );
  NAND2_X1 U15836 ( .A1(n12908), .A2(n12917), .ZN(n12730) );
  NAND2_X1 U15837 ( .A1(n12730), .A2(n15971), .ZN(n12731) );
  AND2_X1 U15838 ( .A1(n12732), .A2(n12731), .ZN(n20234) );
  NOR2_X1 U15839 ( .A1(n12733), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15996) );
  INV_X1 U15840 ( .A(n15996), .ZN(n12929) );
  NAND2_X1 U15841 ( .A1(n12217), .A2(n12929), .ZN(n12734) );
  NAND2_X1 U15842 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21110) );
  OAI21_X1 U15843 ( .B1(n12734), .B2(n13619), .A(n21110), .ZN(n21107) );
  NAND2_X1 U15844 ( .A1(n20234), .A2(n21107), .ZN(n15962) );
  AND2_X1 U15845 ( .A1(n15962), .A2(n13627), .ZN(n20243) );
  INV_X1 U15846 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21252) );
  INV_X1 U15847 ( .A(n12908), .ZN(n12735) );
  OAI22_X1 U15848 ( .A1(n13620), .A2(n15971), .B1(n12917), .B2(n12735), .ZN(
        n12743) );
  INV_X1 U15849 ( .A(n12736), .ZN(n12873) );
  AOI21_X1 U15850 ( .B1(n13394), .B2(n12873), .A(n12737), .ZN(n12738) );
  NAND2_X1 U15851 ( .A1(n12879), .A2(n12738), .ZN(n12906) );
  NOR2_X1 U15852 ( .A1(n12806), .A2(n13400), .ZN(n12739) );
  OR2_X1 U15853 ( .A1(n12906), .A2(n12739), .ZN(n12940) );
  INV_X1 U15854 ( .A(n12740), .ZN(n12951) );
  NAND2_X1 U15855 ( .A1(n13620), .A2(n12951), .ZN(n12741) );
  OAI21_X1 U15856 ( .B1(n13620), .B2(n12940), .A(n12741), .ZN(n12742) );
  OR2_X1 U15857 ( .A1(n12743), .A2(n12742), .ZN(n15963) );
  NAND2_X1 U15858 ( .A1(n20243), .A2(n15963), .ZN(n12744) );
  OAI21_X1 U15859 ( .B1(n20243), .B2(n21252), .A(n12744), .ZN(P1_U3484) );
  INV_X1 U15860 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15861 ( .A1(n16524), .A2(n16551), .ZN(n12746) );
  OAI21_X1 U15862 ( .B1(n13030), .B2(n12746), .A(n12745), .ZN(n12747) );
  INV_X1 U15863 ( .A(n19476), .ZN(n12749) );
  NAND2_X1 U15864 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20191) );
  OR2_X1 U15865 ( .A1(n20191), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20211) );
  INV_X2 U15866 ( .A(n20211), .ZN(n19474) );
  AOI22_X1 U15867 ( .A1(n19474), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U15868 ( .B1(n12751), .B2(n19437), .A(n12750), .ZN(P2_U2929) );
  AOI22_X1 U15869 ( .A1(n19474), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U15870 ( .B1(n12753), .B2(n19437), .A(n12752), .ZN(P2_U2924) );
  INV_X1 U15871 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15872 ( .A1(n19474), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12754) );
  OAI21_X1 U15873 ( .B1(n12755), .B2(n19437), .A(n12754), .ZN(P2_U2933) );
  INV_X1 U15874 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15875 ( .A1(n19474), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12756) );
  OAI21_X1 U15876 ( .B1(n12757), .B2(n19437), .A(n12756), .ZN(P2_U2934) );
  INV_X1 U15877 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15878 ( .A1(n19474), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12758) );
  OAI21_X1 U15879 ( .B1(n12759), .B2(n19437), .A(n12758), .ZN(P2_U2935) );
  INV_X1 U15880 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15881 ( .A1(n19474), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12760) );
  OAI21_X1 U15882 ( .B1(n12761), .B2(n19437), .A(n12760), .ZN(P2_U2927) );
  INV_X1 U15883 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15884 ( .A1(n19474), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12762) );
  OAI21_X1 U15885 ( .B1(n12763), .B2(n19437), .A(n12762), .ZN(P2_U2923) );
  INV_X1 U15886 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15887 ( .A1(n19474), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12764) );
  OAI21_X1 U15888 ( .B1(n12765), .B2(n19437), .A(n12764), .ZN(P2_U2928) );
  AOI22_X1 U15889 ( .A1(n19474), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12766) );
  OAI21_X1 U15890 ( .B1(n12767), .B2(n19437), .A(n12766), .ZN(P2_U2926) );
  INV_X1 U15891 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15892 ( .A1(n19474), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12768) );
  OAI21_X1 U15893 ( .B1(n12769), .B2(n19437), .A(n12768), .ZN(P2_U2925) );
  INV_X1 U15894 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U15895 ( .A1(n19474), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12770) );
  OAI21_X1 U15896 ( .B1(n15189), .B2(n19437), .A(n12770), .ZN(P2_U2930) );
  INV_X1 U15897 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U15898 ( .A1(n19474), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12771) );
  OAI21_X1 U15899 ( .B1(n14028), .B2(n19437), .A(n12771), .ZN(P2_U2932) );
  INV_X1 U15900 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15901 ( .A1(n19474), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12772) );
  OAI21_X1 U15902 ( .B1(n12773), .B2(n19437), .A(n12772), .ZN(P2_U2931) );
  AOI21_X1 U15903 ( .B1(n13562), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12774), .ZN(n12776) );
  NAND2_X1 U15904 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12840) );
  OAI211_X1 U15905 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15517), .B(n12840), .ZN(n12775) );
  OAI211_X1 U15906 ( .C1(n12777), .C2(n16477), .A(n12776), .B(n12775), .ZN(
        n12778) );
  INV_X1 U15907 ( .A(n12778), .ZN(n12785) );
  NAND2_X1 U15908 ( .A1(n12780), .A2(n12779), .ZN(n12781) );
  NAND2_X1 U15909 ( .A1(n12782), .A2(n12781), .ZN(n20188) );
  AOI22_X1 U15910 ( .A1(n16493), .A2(n12783), .B1(n16485), .B2(n20188), .ZN(
        n12784) );
  OAI211_X1 U15911 ( .C1(n19330), .C2(n15640), .A(n12785), .B(n12784), .ZN(
        P2_U3045) );
  NOR2_X1 U15912 ( .A1(n12906), .A2(n12786), .ZN(n12787) );
  OR2_X1 U15913 ( .A1(n20513), .A2(n13756), .ZN(n12790) );
  NAND2_X1 U15914 ( .A1(n13394), .A2(n20452), .ZN(n12987) );
  OAI21_X1 U15915 ( .B1(n21104), .B2(n12964), .A(n12987), .ZN(n12788) );
  INV_X1 U15916 ( .A(n12788), .ZN(n12789) );
  NAND2_X1 U15917 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  OAI21_X1 U15918 ( .B1(n12791), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12981), .ZN(n12957) );
  NAND2_X1 U15919 ( .A1(n21026), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12793) );
  NAND2_X1 U15920 ( .A1(n21220), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12792) );
  AND2_X1 U15921 ( .A1(n12793), .A2(n12792), .ZN(n12959) );
  INV_X1 U15922 ( .A(n20842), .ZN(n20967) );
  NAND2_X1 U15923 ( .A1(n20967), .A2(n12795), .ZN(n21109) );
  AND2_X1 U15924 ( .A1(n21109), .A2(n21026), .ZN(n12794) );
  NAND2_X1 U15925 ( .A1(n12959), .A2(n14824), .ZN(n12804) );
  INV_X1 U15926 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n12796) );
  OR2_X1 U15927 ( .A1(n16210), .A2(n12796), .ZN(n12952) );
  INV_X1 U15928 ( .A(n12952), .ZN(n12803) );
  NAND2_X1 U15929 ( .A1(n12798), .A2(n12797), .ZN(n12799) );
  AND2_X1 U15930 ( .A1(n12800), .A2(n12799), .ZN(n13417) );
  INV_X1 U15931 ( .A(n13417), .ZN(n13707) );
  NAND3_X1 U15932 ( .A1(n21026), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16247) );
  INV_X1 U15933 ( .A(n16247), .ZN(n12801) );
  NOR2_X1 U15934 ( .A1(n13707), .A2(n20417), .ZN(n12802) );
  AOI211_X1 U15935 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12804), .A(
        n12803), .B(n12802), .ZN(n12805) );
  OAI21_X1 U15936 ( .B1(n20242), .B2(n12957), .A(n12805), .ZN(P1_U2999) );
  INV_X1 U15937 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21478) );
  NAND2_X1 U15938 ( .A1(n12868), .A2(n15996), .ZN(n15970) );
  NAND2_X1 U15939 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  AND2_X1 U15940 ( .A1(n14373), .A2(n15996), .ZN(n12809) );
  NAND2_X1 U15941 ( .A1(n13620), .A2(n12809), .ZN(n12920) );
  NAND2_X1 U15942 ( .A1(n20328), .A2(n20423), .ZN(n13090) );
  INV_X1 U15943 ( .A(n13321), .ZN(n16248) );
  INV_X2 U15944 ( .A(n20326), .ZN(n21111) );
  NOR2_X4 U15945 ( .A1(n20328), .A2(n21111), .ZN(n15999) );
  AOI22_X1 U15946 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U15947 ( .B1(n21478), .B2(n13090), .A(n12810), .ZN(P1_U2912) );
  INV_X1 U15948 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15949 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12811) );
  OAI21_X1 U15950 ( .B1(n12812), .B2(n13090), .A(n12811), .ZN(P1_U2920) );
  INV_X1 U15951 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21466) );
  AOI22_X1 U15952 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12813) );
  OAI21_X1 U15953 ( .B1(n21466), .B2(n13090), .A(n12813), .ZN(P1_U2911) );
  INV_X1 U15954 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15955 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12814) );
  OAI21_X1 U15956 ( .B1(n12815), .B2(n13090), .A(n12814), .ZN(P1_U2914) );
  INV_X1 U15957 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U15958 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12816) );
  OAI21_X1 U15959 ( .B1(n14654), .B2(n13090), .A(n12816), .ZN(P1_U2917) );
  INV_X1 U15960 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21484) );
  AOI22_X1 U15961 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12817) );
  OAI21_X1 U15962 ( .B1(n21484), .B2(n13090), .A(n12817), .ZN(P1_U2909) );
  INV_X1 U15963 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21459) );
  AOI22_X1 U15964 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12818) );
  OAI21_X1 U15965 ( .B1(n21459), .B2(n13090), .A(n12818), .ZN(P1_U2908) );
  INV_X1 U15966 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21226) );
  AOI22_X1 U15967 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12819) );
  OAI21_X1 U15968 ( .B1(n21226), .B2(n13090), .A(n12819), .ZN(P1_U2915) );
  INV_X1 U15969 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15970 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U15971 ( .B1(n12821), .B2(n13090), .A(n12820), .ZN(P1_U2919) );
  INV_X1 U15972 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U15973 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12822) );
  OAI21_X1 U15974 ( .B1(n12823), .B2(n13090), .A(n12822), .ZN(P1_U2918) );
  INV_X1 U15975 ( .A(n13562), .ZN(n12834) );
  NOR2_X1 U15976 ( .A1(n12824), .A2(n19329), .ZN(n12826) );
  OAI21_X1 U15977 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12826), .A(
        n12825), .ZN(n12831) );
  INV_X1 U15978 ( .A(n12827), .ZN(n12828) );
  XNOR2_X1 U15979 ( .A(n12829), .B(n12828), .ZN(n15004) );
  XNOR2_X1 U15980 ( .A(n15004), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12830) );
  OR2_X1 U15981 ( .A1(n12831), .A2(n12830), .ZN(n19506) );
  NAND2_X1 U15982 ( .A1(n12831), .A2(n12830), .ZN(n19505) );
  NAND3_X1 U15983 ( .A1(n19506), .A2(n16490), .A3(n19505), .ZN(n12832) );
  NAND2_X1 U15984 ( .A1(n19310), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19511) );
  OAI211_X1 U15985 ( .C1(n12834), .C2(n12833), .A(n12832), .B(n19511), .ZN(
        n12855) );
  OR2_X1 U15986 ( .A1(n12836), .A2(n12835), .ZN(n12838) );
  NAND2_X1 U15987 ( .A1(n12838), .A2(n12837), .ZN(n20179) );
  INV_X1 U15988 ( .A(n20179), .ZN(n12841) );
  INV_X1 U15989 ( .A(n12840), .ZN(n12839) );
  NAND2_X1 U15990 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12839), .ZN(
        n13564) );
  NAND2_X1 U15991 ( .A1(n12833), .A2(n12840), .ZN(n14264) );
  NAND2_X1 U15992 ( .A1(n13564), .A2(n14264), .ZN(n12851) );
  OAI22_X1 U15993 ( .A1(n16469), .A2(n12841), .B1(n12851), .B2(n15519), .ZN(
        n12854) );
  INV_X1 U15994 ( .A(n12842), .ZN(n12844) );
  NAND2_X1 U15995 ( .A1(n12844), .A2(n12843), .ZN(n12846) );
  NAND2_X1 U15996 ( .A1(n12846), .A2(n12845), .ZN(n13552) );
  XNOR2_X1 U15997 ( .A(n12833), .B(n13552), .ZN(n12850) );
  AND2_X1 U15998 ( .A1(n12848), .A2(n12847), .ZN(n13541) );
  XOR2_X1 U15999 ( .A(n13542), .B(n13541), .Z(n12849) );
  NAND2_X1 U16000 ( .A1(n12850), .A2(n12849), .ZN(n13554) );
  OAI21_X1 U16001 ( .B1(n12850), .B2(n12849), .A(n13554), .ZN(n19500) );
  INV_X1 U16002 ( .A(n12851), .ZN(n12852) );
  OAI22_X1 U16003 ( .A1(n16457), .A2(n19500), .B1(n12852), .B2(n15512), .ZN(
        n12853) );
  NOR3_X1 U16004 ( .A1(n12855), .A2(n12854), .A3(n12853), .ZN(n12856) );
  OAI21_X1 U16005 ( .B1(n13468), .B2(n15640), .A(n12856), .ZN(P2_U3044) );
  INV_X1 U16006 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n21314) );
  OR2_X1 U16007 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12857) );
  NAND2_X1 U16008 ( .A1(n12858), .A2(n12857), .ZN(n13414) );
  OAI222_X1 U16009 ( .A1(n13707), .A2(n14610), .B1(n21314), .B2(n14612), .C1(
        n13414), .C2(n14613), .ZN(P1_U2872) );
  OR2_X1 U16010 ( .A1(n12860), .A2(n12859), .ZN(n12861) );
  NAND2_X1 U16011 ( .A1(n12973), .A2(n12861), .ZN(n13709) );
  OR2_X1 U16012 ( .A1(n12862), .A2(n13619), .ZN(n12864) );
  AND2_X1 U16013 ( .A1(n12864), .A2(n12863), .ZN(n12998) );
  INV_X1 U16014 ( .A(n12998), .ZN(n13426) );
  AOI22_X1 U16015 ( .A1(n14601), .A2(n13426), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14600), .ZN(n12865) );
  OAI21_X1 U16016 ( .B1(n14610), .B2(n13709), .A(n12865), .ZN(P1_U2871) );
  INV_X1 U16017 ( .A(n21110), .ZN(n15997) );
  AND2_X1 U16018 ( .A1(n21104), .A2(n15997), .ZN(n12866) );
  INV_X1 U16019 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14079) );
  INV_X1 U16020 ( .A(DATAI_15_), .ZN(n12870) );
  INV_X1 U16021 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12869) );
  MUX2_X1 U16022 ( .A(n12870), .B(n12869), .S(n20415), .Z(n14080) );
  INV_X1 U16023 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20327) );
  OAI222_X1 U16024 ( .A1(n14320), .A2(n14079), .B1(n13043), .B2(n14080), .C1(
        n13047), .C2(n20327), .ZN(P1_U2967) );
  NAND2_X1 U16025 ( .A1(n12872), .A2(n13400), .ZN(n12883) );
  NAND2_X1 U16026 ( .A1(n12873), .A2(n20423), .ZN(n12874) );
  NAND2_X1 U16027 ( .A1(n12874), .A2(n21104), .ZN(n12875) );
  NAND2_X1 U16028 ( .A1(n12876), .A2(n12875), .ZN(n12909) );
  INV_X1 U16029 ( .A(n12892), .ZN(n13300) );
  NAND2_X1 U16030 ( .A1(n12879), .A2(n13300), .ZN(n12880) );
  NAND2_X1 U16031 ( .A1(n12880), .A2(n20440), .ZN(n12881) );
  NAND4_X1 U16032 ( .A1(n12883), .A2(n12909), .A3(n12882), .A4(n12881), .ZN(
        n12946) );
  INV_X1 U16033 ( .A(n13622), .ZN(n12885) );
  INV_X1 U16034 ( .A(n12904), .ZN(n12884) );
  NAND3_X1 U16035 ( .A1(n12885), .A2(n12884), .A3(n12949), .ZN(n12886) );
  NOR2_X1 U16036 ( .A1(n12946), .A2(n12886), .ZN(n12889) );
  AND2_X1 U16037 ( .A1(n12889), .A2(n12888), .ZN(n14975) );
  OR2_X1 U16038 ( .A1(n20845), .A2(n14975), .ZN(n12901) );
  INV_X1 U16039 ( .A(n14975), .ZN(n14369) );
  INV_X1 U16040 ( .A(n13299), .ZN(n12891) );
  INV_X1 U16041 ( .A(n13291), .ZN(n14978) );
  NAND2_X1 U16042 ( .A1(n14978), .A2(n11208), .ZN(n12890) );
  NAND2_X1 U16043 ( .A1(n12891), .A2(n12890), .ZN(n12895) );
  INV_X1 U16044 ( .A(n12895), .ZN(n12903) );
  NAND2_X1 U16045 ( .A1(n12892), .A2(n12903), .ZN(n12898) );
  NAND2_X1 U16046 ( .A1(n14373), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12894) );
  NAND2_X1 U16047 ( .A1(n14373), .A2(n12893), .ZN(n14974) );
  MUX2_X1 U16048 ( .A(n12894), .B(n14974), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12897) );
  NOR2_X1 U16049 ( .A1(n12906), .A2(n12217), .ZN(n12916) );
  OR2_X1 U16050 ( .A1(n12951), .A2(n12916), .ZN(n13293) );
  NAND2_X1 U16051 ( .A1(n13293), .A2(n12895), .ZN(n12896) );
  OAI211_X1 U16052 ( .C1(n14369), .C2(n12898), .A(n12897), .B(n12896), .ZN(
        n12899) );
  INV_X1 U16053 ( .A(n12899), .ZN(n12900) );
  NAND2_X1 U16054 ( .A1(n12901), .A2(n12900), .ZN(n13306) );
  INV_X1 U16055 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13691) );
  NOR2_X1 U16056 ( .A1(n21025), .A2(n13691), .ZN(n14371) );
  INV_X1 U16057 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16058 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20397), .B2(n12902), .ZN(
        n14982) );
  INV_X1 U16059 ( .A(n14986), .ZN(n14976) );
  AOI222_X1 U16060 ( .A1(n13306), .A2(n16242), .B1(n14371), .B2(n14982), .C1(
        n14976), .C2(n12903), .ZN(n12924) );
  AND2_X1 U16061 ( .A1(n12904), .A2(n21110), .ZN(n13618) );
  OR2_X1 U16062 ( .A1(n13619), .A2(n15996), .ZN(n12905) );
  NAND2_X1 U16063 ( .A1(n13618), .A2(n12905), .ZN(n12933) );
  INV_X1 U16064 ( .A(n12933), .ZN(n12913) );
  INV_X1 U16065 ( .A(n12906), .ZN(n12907) );
  OR2_X1 U16066 ( .A1(n12908), .A2(n12907), .ZN(n12910) );
  NAND2_X1 U16067 ( .A1(n12910), .A2(n12909), .ZN(n12927) );
  INV_X1 U16068 ( .A(n12927), .ZN(n12911) );
  OAI21_X1 U16069 ( .B1(n20446), .B2(n13403), .A(n12911), .ZN(n12912) );
  AOI21_X1 U16070 ( .B1(n13620), .B2(n12913), .A(n12912), .ZN(n12915) );
  AND2_X1 U16071 ( .A1(n12915), .A2(n12914), .ZN(n12923) );
  NAND2_X1 U16072 ( .A1(n13620), .A2(n12916), .ZN(n12919) );
  NAND2_X1 U16073 ( .A1(n12917), .A2(n21110), .ZN(n12930) );
  OR2_X1 U16074 ( .A1(n12888), .A2(n12930), .ZN(n12918) );
  NAND2_X1 U16075 ( .A1(n12919), .A2(n12918), .ZN(n13626) );
  INV_X1 U16076 ( .A(n13626), .ZN(n12922) );
  OR2_X1 U16077 ( .A1(n12920), .A2(n15997), .ZN(n12921) );
  NAND2_X1 U16078 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13321), .ZN(n16252) );
  INV_X1 U16079 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21311) );
  OAI22_X1 U16080 ( .A1(n15949), .A2(n20235), .B1(n16252), .B2(n21311), .ZN(
        n16243) );
  AOI21_X1 U16081 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21026), .A(n16243), 
        .ZN(n14375) );
  INV_X1 U16082 ( .A(n14375), .ZN(n16245) );
  MUX2_X1 U16083 ( .A(n11209), .B(n12924), .S(n16245), .Z(n12926) );
  INV_X1 U16084 ( .A(n12926), .ZN(P1_U3472) );
  INV_X1 U16085 ( .A(n13620), .ZN(n15980) );
  AOI21_X1 U16086 ( .B1(n15980), .B2(n12928), .A(n12927), .ZN(n12938) );
  NAND2_X1 U16087 ( .A1(n20440), .A2(n12929), .ZN(n12932) );
  INV_X1 U16088 ( .A(n12930), .ZN(n12931) );
  NAND2_X1 U16089 ( .A1(n12932), .A2(n12931), .ZN(n12936) );
  INV_X1 U16090 ( .A(n13631), .ZN(n13629) );
  NAND3_X1 U16091 ( .A1(n12933), .A2(n20423), .A3(n13629), .ZN(n12934) );
  NAND2_X1 U16092 ( .A1(n13620), .A2(n12934), .ZN(n12935) );
  MUX2_X1 U16093 ( .A(n12936), .B(n12935), .S(n12965), .Z(n12937) );
  NAND2_X1 U16094 ( .A1(n12938), .A2(n12937), .ZN(n12939) );
  OAI21_X1 U16095 ( .B1(n12944), .B2(n11354), .A(n12940), .ZN(n12941) );
  OR2_X1 U16096 ( .A1(n12942), .A2(n12941), .ZN(n12943) );
  INV_X1 U16097 ( .A(n12946), .ZN(n12948) );
  OAI211_X1 U16098 ( .C1(n12949), .C2(n20423), .A(n12948), .B(n12947), .ZN(
        n12950) );
  NAND2_X1 U16099 ( .A1(n13691), .A2(n13005), .ZN(n13000) );
  OAI211_X1 U16100 ( .C1(n16211), .C2(n13414), .A(n13000), .B(n12952), .ZN(
        n12953) );
  INV_X1 U16101 ( .A(n12953), .ZN(n12956) );
  INV_X2 U16102 ( .A(n16210), .ZN(n20380) );
  NOR2_X1 U16103 ( .A1(n20380), .A2(n12954), .ZN(n12999) );
  OAI21_X1 U16104 ( .B1(n14956), .B2(n12999), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12955) );
  OAI211_X1 U16105 ( .C1(n20387), .C2(n12957), .A(n12956), .B(n12955), .ZN(
        P1_U3031) );
  INV_X1 U16106 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n12958) );
  NOR2_X1 U16107 ( .A1(n16210), .A2(n12958), .ZN(n13002) );
  INV_X1 U16108 ( .A(n12959), .ZN(n12960) );
  NOR2_X1 U16109 ( .A1(n20374), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12961) );
  AOI211_X1 U16110 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13002), .B(n12961), .ZN(n12972) );
  NAND2_X1 U16111 ( .A1(n12962), .A2(n20440), .ZN(n12969) );
  NAND2_X1 U16112 ( .A1(n12963), .A2(n12964), .ZN(n13330) );
  OAI21_X1 U16113 ( .B1(n12964), .B2(n12963), .A(n13330), .ZN(n12966) );
  OAI211_X1 U16114 ( .C1(n12966), .C2(n21104), .A(n12965), .B(n20463), .ZN(
        n12967) );
  INV_X1 U16115 ( .A(n12967), .ZN(n12968) );
  INV_X1 U16116 ( .A(n12985), .ZN(n12997) );
  NOR2_X1 U16117 ( .A1(n12970), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12996) );
  OR3_X1 U16118 ( .A1(n12997), .A2(n12996), .A3(n20242), .ZN(n12971) );
  OAI211_X1 U16119 ( .C1(n13709), .C2(n20417), .A(n12972), .B(n12971), .ZN(
        P1_U2998) );
  OAI21_X1 U16120 ( .B1(n10403), .B2(n11584), .A(n12974), .ZN(n13701) );
  INV_X1 U16121 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21233) );
  NAND2_X1 U16122 ( .A1(n12976), .A2(n12975), .ZN(n12977) );
  AND2_X1 U16123 ( .A1(n13099), .A2(n12977), .ZN(n20403) );
  INV_X1 U16124 ( .A(n20403), .ZN(n12978) );
  OAI222_X1 U16125 ( .A1(n13701), .A2(n14610), .B1(n14612), .B2(n21233), .C1(
        n12978), .C2(n14613), .ZN(P1_U2870) );
  INV_X1 U16126 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n12979) );
  NOR2_X1 U16127 ( .A1(n16210), .A2(n12979), .ZN(n20402) );
  NOR2_X1 U16128 ( .A1(n20374), .A2(n13421), .ZN(n12980) );
  AOI211_X1 U16129 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20402), .B(n12980), .ZN(n12995) );
  INV_X1 U16130 ( .A(n12981), .ZN(n12982) );
  NAND2_X1 U16131 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  XNOR2_X1 U16132 ( .A(n13326), .B(n20411), .ZN(n12992) );
  OR2_X1 U16133 ( .A1(n12986), .A2(n13756), .ZN(n12991) );
  XNOR2_X1 U16134 ( .A(n13330), .B(n13329), .ZN(n12989) );
  INV_X1 U16135 ( .A(n21104), .ZN(n13772) );
  INV_X1 U16136 ( .A(n12987), .ZN(n12988) );
  AOI21_X1 U16137 ( .B1(n12989), .B2(n13772), .A(n12988), .ZN(n12990) );
  NAND2_X1 U16138 ( .A1(n12991), .A2(n12990), .ZN(n12993) );
  OR2_X1 U16139 ( .A1(n12992), .A2(n12993), .ZN(n20406) );
  NAND2_X1 U16140 ( .A1(n12993), .A2(n12992), .ZN(n13328) );
  NAND3_X1 U16141 ( .A1(n20406), .A2(n13328), .A3(n20370), .ZN(n12994) );
  OAI211_X1 U16142 ( .C1(n20417), .C2(n13701), .A(n12995), .B(n12994), .ZN(
        P1_U2997) );
  NOR3_X1 U16143 ( .A1(n20387), .A2(n12997), .A3(n12996), .ZN(n13004) );
  NOR2_X1 U16144 ( .A1(n16211), .A2(n12998), .ZN(n13003) );
  INV_X1 U16145 ( .A(n12999), .ZN(n13692) );
  AOI21_X1 U16146 ( .B1(n13692), .B2(n13000), .A(n20397), .ZN(n13001) );
  NOR4_X1 U16147 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13008) );
  NAND2_X2 U16148 ( .A1(n13006), .A2(n13690), .ZN(n16219) );
  OAI211_X1 U16149 ( .C1(n14956), .C2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16219), .B(n20397), .ZN(n13007) );
  NAND2_X1 U16150 ( .A1(n13008), .A2(n13007), .ZN(P1_U3030) );
  INV_X1 U16151 ( .A(n19583), .ZN(n20167) );
  INV_X1 U16152 ( .A(n15656), .ZN(n16547) );
  INV_X1 U16153 ( .A(n15652), .ZN(n15682) );
  AND2_X1 U16154 ( .A1(n10646), .A2(n13012), .ZN(n13017) );
  NOR2_X1 U16155 ( .A1(n15664), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15673) );
  INV_X1 U16156 ( .A(n15673), .ZN(n15679) );
  INV_X1 U16157 ( .A(n13012), .ZN(n13013) );
  NAND2_X1 U16158 ( .A1(n10646), .A2(n13013), .ZN(n15674) );
  AOI21_X1 U16159 ( .B1(n10662), .B2(n13014), .A(n15672), .ZN(n15680) );
  INV_X1 U16160 ( .A(n15680), .ZN(n13015) );
  NAND3_X1 U16161 ( .A1(n15679), .A2(n15674), .A3(n13015), .ZN(n13016) );
  MUX2_X1 U16162 ( .A(n13017), .B(n13016), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13021) );
  NOR2_X1 U16163 ( .A1(n16533), .A2(n13018), .ZN(n15677) );
  OR2_X1 U16164 ( .A1(n15677), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13019) );
  AOI21_X1 U16165 ( .B1(n13019), .B2(n10416), .A(n15673), .ZN(n13020) );
  NOR2_X1 U16166 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  OAI21_X1 U16167 ( .B1(n13011), .B2(n15682), .A(n13022), .ZN(n16504) );
  AOI22_X1 U16168 ( .A1(n20167), .A2(n16547), .B1(n20163), .B2(n16504), .ZN(
        n13036) );
  NAND2_X1 U16169 ( .A1(n16524), .A2(n16519), .ZN(n13031) );
  INV_X1 U16170 ( .A(n13023), .ZN(n13024) );
  AND2_X1 U16171 ( .A1(n13025), .A2(n13024), .ZN(n13029) );
  AND2_X1 U16172 ( .A1(n13026), .A2(n20216), .ZN(n16521) );
  AND3_X1 U16173 ( .A1(n12376), .A2(n16529), .A3(n16521), .ZN(n13027) );
  AOI21_X1 U16174 ( .B1(n13028), .B2(n16533), .A(n13027), .ZN(n13947) );
  OAI211_X1 U16175 ( .C1(n13031), .C2(n13030), .A(n13029), .B(n13947), .ZN(
        n16505) );
  NAND2_X1 U16176 ( .A1(n16505), .A2(n16551), .ZN(n13034) );
  NOR2_X1 U16177 ( .A1(n20218), .A2(n20191), .ZN(n16554) );
  NOR2_X1 U16178 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12466), .ZN(n13032) );
  AOI21_X1 U16179 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16554), .A(n13032), .ZN(
        n13033) );
  NAND2_X1 U16180 ( .A1(n13034), .A2(n13033), .ZN(n15749) );
  INV_X1 U16181 ( .A(n15749), .ZN(n15686) );
  NAND2_X1 U16182 ( .A1(n15686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13035) );
  OAI21_X1 U16183 ( .B1(n13036), .B2(n15686), .A(n13035), .ZN(P2_U3596) );
  MUX2_X1 U16184 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n19509), .S(n15104), .Z(
        n13041) );
  AOI21_X1 U16185 ( .B1(n20174), .B2(n15110), .A(n13041), .ZN(n13042) );
  INV_X1 U16186 ( .A(n13042), .ZN(P2_U2885) );
  AOI22_X1 U16187 ( .A1(n20362), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20361), .ZN(n13046) );
  INV_X1 U16188 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16686) );
  NAND2_X1 U16189 ( .A1(n20415), .A2(n16686), .ZN(n13044) );
  OAI21_X1 U16190 ( .B1(n20415), .B2(DATAI_0_), .A(n13044), .ZN(n20431) );
  INV_X1 U16191 ( .A(n20431), .ZN(n13045) );
  NAND2_X1 U16192 ( .A1(n14316), .A2(n13045), .ZN(n13073) );
  NAND2_X1 U16193 ( .A1(n13046), .A2(n13073), .ZN(P1_U2952) );
  AOI22_X1 U16194 ( .A1(n20362), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20361), .ZN(n13050) );
  INV_X1 U16195 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16681) );
  NAND2_X1 U16196 ( .A1(n20415), .A2(n16681), .ZN(n13048) );
  OAI21_X1 U16197 ( .B1(n20415), .B2(DATAI_1_), .A(n13048), .ZN(n20442) );
  INV_X1 U16198 ( .A(n20442), .ZN(n13049) );
  NAND2_X1 U16199 ( .A1(n14316), .A2(n13049), .ZN(n13071) );
  NAND2_X1 U16200 ( .A1(n13050), .A2(n13071), .ZN(P1_U2953) );
  AOI22_X1 U16201 ( .A1(n20362), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20361), .ZN(n13053) );
  INV_X1 U16202 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16675) );
  NAND2_X1 U16203 ( .A1(n20415), .A2(n16675), .ZN(n13051) );
  OAI21_X1 U16204 ( .B1(n20415), .B2(DATAI_4_), .A(n13051), .ZN(n20459) );
  INV_X1 U16205 ( .A(n20459), .ZN(n13052) );
  NAND2_X1 U16206 ( .A1(n14316), .A2(n13052), .ZN(n13064) );
  NAND2_X1 U16207 ( .A1(n13053), .A2(n13064), .ZN(P1_U2956) );
  AOI22_X1 U16208 ( .A1(n20362), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20361), .ZN(n13057) );
  INV_X1 U16209 ( .A(n20415), .ZN(n20416) );
  NAND2_X1 U16210 ( .A1(n20416), .A2(DATAI_2_), .ZN(n13055) );
  NAND2_X1 U16211 ( .A1(n20415), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13054) );
  AND2_X1 U16212 ( .A1(n13055), .A2(n13054), .ZN(n20448) );
  INV_X1 U16213 ( .A(n20448), .ZN(n13056) );
  NAND2_X1 U16214 ( .A1(n14316), .A2(n13056), .ZN(n13069) );
  NAND2_X1 U16215 ( .A1(n13057), .A2(n13069), .ZN(P1_U2954) );
  AOI22_X1 U16216 ( .A1(n20362), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20361), .ZN(n13060) );
  INV_X1 U16217 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16671) );
  NAND2_X1 U16218 ( .A1(n20415), .A2(n16671), .ZN(n13058) );
  OAI21_X1 U16219 ( .B1(n20415), .B2(DATAI_6_), .A(n13058), .ZN(n20473) );
  INV_X1 U16220 ( .A(n20473), .ZN(n13059) );
  NAND2_X1 U16221 ( .A1(n14316), .A2(n13059), .ZN(n13081) );
  NAND2_X1 U16222 ( .A1(n13060), .A2(n13081), .ZN(P1_U2943) );
  AOI22_X1 U16223 ( .A1(n20362), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20361), .ZN(n13063) );
  INV_X1 U16224 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16673) );
  NAND2_X1 U16225 ( .A1(n20415), .A2(n16673), .ZN(n13061) );
  OAI21_X1 U16226 ( .B1(n20415), .B2(DATAI_5_), .A(n13061), .ZN(n20465) );
  INV_X1 U16227 ( .A(n20465), .ZN(n13062) );
  NAND2_X1 U16228 ( .A1(n14316), .A2(n13062), .ZN(n13079) );
  NAND2_X1 U16229 ( .A1(n13063), .A2(n13079), .ZN(P1_U2942) );
  AOI22_X1 U16230 ( .A1(n20362), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20361), .ZN(n13065) );
  NAND2_X1 U16231 ( .A1(n13065), .A2(n13064), .ZN(P1_U2941) );
  AOI22_X1 U16232 ( .A1(n20362), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20361), .ZN(n13068) );
  INV_X1 U16233 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16677) );
  NAND2_X1 U16234 ( .A1(n20415), .A2(n16677), .ZN(n13066) );
  OAI21_X1 U16235 ( .B1(n20415), .B2(DATAI_3_), .A(n13066), .ZN(n20454) );
  INV_X1 U16236 ( .A(n20454), .ZN(n13067) );
  NAND2_X1 U16237 ( .A1(n14316), .A2(n13067), .ZN(n13077) );
  NAND2_X1 U16238 ( .A1(n13068), .A2(n13077), .ZN(P1_U2940) );
  AOI22_X1 U16239 ( .A1(n20362), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20361), .ZN(n13070) );
  NAND2_X1 U16240 ( .A1(n13070), .A2(n13069), .ZN(P1_U2939) );
  AOI22_X1 U16241 ( .A1(n20362), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20361), .ZN(n13072) );
  NAND2_X1 U16242 ( .A1(n13072), .A2(n13071), .ZN(P1_U2938) );
  AOI22_X1 U16243 ( .A1(n20362), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20361), .ZN(n13074) );
  NAND2_X1 U16244 ( .A1(n13074), .A2(n13073), .ZN(P1_U2937) );
  AOI22_X1 U16245 ( .A1(n20362), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20361), .ZN(n13076) );
  INV_X1 U16246 ( .A(DATAI_7_), .ZN(n21203) );
  INV_X1 U16247 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16669) );
  MUX2_X1 U16248 ( .A(n21203), .B(n16669), .S(n20415), .Z(n20482) );
  INV_X1 U16249 ( .A(n20482), .ZN(n13075) );
  NAND2_X1 U16250 ( .A1(n14316), .A2(n13075), .ZN(n13083) );
  NAND2_X1 U16251 ( .A1(n13076), .A2(n13083), .ZN(P1_U2944) );
  AOI22_X1 U16252 ( .A1(n20362), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20361), .ZN(n13078) );
  NAND2_X1 U16253 ( .A1(n13078), .A2(n13077), .ZN(P1_U2955) );
  AOI22_X1 U16254 ( .A1(n20362), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20361), .ZN(n13080) );
  NAND2_X1 U16255 ( .A1(n13080), .A2(n13079), .ZN(P1_U2957) );
  AOI22_X1 U16256 ( .A1(n20362), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20361), .ZN(n13082) );
  NAND2_X1 U16257 ( .A1(n13082), .A2(n13081), .ZN(P1_U2958) );
  AOI22_X1 U16258 ( .A1(n20362), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20361), .ZN(n13084) );
  NAND2_X1 U16259 ( .A1(n13084), .A2(n13083), .ZN(P1_U2959) );
  INV_X1 U16260 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21475) );
  AOI22_X1 U16261 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21111), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15999), .ZN(n13085) );
  OAI21_X1 U16262 ( .B1(n21475), .B2(n13090), .A(n13085), .ZN(P1_U2906) );
  INV_X1 U16263 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16264 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13086) );
  OAI21_X1 U16265 ( .B1(n14314), .B2(n13090), .A(n13086), .ZN(P1_U2910) );
  INV_X1 U16266 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21323) );
  AOI22_X1 U16267 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13087) );
  OAI21_X1 U16268 ( .B1(n21323), .B2(n13090), .A(n13087), .ZN(P1_U2916) );
  INV_X1 U16269 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21238) );
  AOI22_X1 U16270 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13088) );
  OAI21_X1 U16271 ( .B1(n21238), .B2(n13090), .A(n13088), .ZN(P1_U2913) );
  INV_X1 U16272 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U16273 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13089) );
  OAI21_X1 U16274 ( .B1(n14307), .B2(n13090), .A(n13089), .ZN(P1_U2907) );
  NOR2_X1 U16275 ( .A1(n14093), .A2(n10791), .ZN(n13093) );
  INV_X1 U16276 ( .A(n13091), .ZN(n13092) );
  OAI211_X1 U16277 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13093), .A(
        n13092), .B(n15110), .ZN(n13096) );
  AOI21_X1 U16278 ( .B1(n13094), .B2(n14081), .A(n13368), .ZN(n19289) );
  NAND2_X1 U16279 ( .A1(n19289), .A2(n15104), .ZN(n13095) );
  OAI211_X1 U16280 ( .C1(n15104), .C2(n13097), .A(n13096), .B(n13095), .ZN(
        P2_U2881) );
  AND2_X1 U16281 ( .A1(n13099), .A2(n13098), .ZN(n13100) );
  NOR2_X1 U16282 ( .A1(n13379), .A2(n13100), .ZN(n20386) );
  INV_X1 U16283 ( .A(n20386), .ZN(n13104) );
  INV_X1 U16284 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21191) );
  OAI21_X1 U16285 ( .B1(n13103), .B2(n13102), .A(n13384), .ZN(n13710) );
  OAI222_X1 U16286 ( .A1(n13104), .A2(n14613), .B1(n14612), .B2(n21191), .C1(
        n13710), .C2(n14610), .ZN(P1_U2869) );
  AND2_X1 U16287 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17171) );
  AOI22_X1 U16288 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17398), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n9830), .ZN(n13105) );
  OAI21_X1 U16289 ( .B1(n18454), .B2(n17238), .A(n13105), .ZN(n13120) );
  AOI22_X1 U16290 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13106), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n9822), .ZN(n13118) );
  NOR2_X4 U16291 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13108), .ZN(
        n15772) );
  AOI22_X1 U16292 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n15772), .ZN(n13109) );
  OAI21_X1 U16293 ( .B1(n17298), .B2(n18667), .A(n13109), .ZN(n13116) );
  INV_X1 U16294 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18862) );
  INV_X2 U16295 ( .A(n9885), .ZN(n17281) );
  AOI22_X1 U16296 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17281), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n15837), .ZN(n13114) );
  AOI22_X1 U16297 ( .A1(n17360), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17359), .ZN(n13113) );
  OAI211_X1 U16298 ( .C1(n18862), .C2(n9828), .A(n13114), .B(n13113), .ZN(
        n13115) );
  AOI211_X1 U16299 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n13116), .B(n13115), .ZN(n13117) );
  OAI211_X1 U16300 ( .C1(n10408), .C2(n17143), .A(n13118), .B(n13117), .ZN(
        n13119) );
  AOI211_X4 U16301 ( .C1(n17363), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13120), .B(n13119), .ZN(n17577) );
  INV_X2 U16302 ( .A(n9876), .ZN(n17394) );
  AOI22_X1 U16303 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16304 ( .B1(n17238), .B2(n18415), .A(n13121), .ZN(n13130) );
  AOI22_X1 U16305 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16306 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13122) );
  OAI21_X1 U16307 ( .B1(n9828), .B2(n18806), .A(n13122), .ZN(n13126) );
  AOI22_X1 U16308 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16309 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13123) );
  OAI211_X1 U16310 ( .C1(n15793), .C2(n18646), .A(n13124), .B(n13123), .ZN(
        n13125) );
  AOI211_X1 U16311 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13126), .B(n13125), .ZN(n13127) );
  OAI211_X1 U16312 ( .C1(n15787), .C2(n17414), .A(n13128), .B(n13127), .ZN(
        n13129) );
  AOI22_X1 U16313 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U16314 ( .B1(n17328), .B2(n18626), .A(n13131), .ZN(n13141) );
  AOI22_X1 U16315 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13139) );
  INV_X1 U16316 ( .A(n13132), .ZN(n17298) );
  AOI22_X1 U16317 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13133) );
  OAI21_X1 U16318 ( .B1(n17298), .B2(n18654), .A(n13133), .ZN(n13137) );
  AOI22_X1 U16319 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16320 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17412), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13134) );
  OAI211_X1 U16321 ( .C1(n9828), .C2(n18827), .A(n13135), .B(n13134), .ZN(
        n13136) );
  AOI211_X1 U16322 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13137), .B(n13136), .ZN(n13138) );
  OAI211_X1 U16323 ( .C1(n17238), .C2(n18429), .A(n13139), .B(n13138), .ZN(
        n13140) );
  OAI22_X1 U16324 ( .A1(n10419), .A2(n15691), .B1(n9876), .B2(n15792), .ZN(
        n13152) );
  INV_X1 U16325 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U16326 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16327 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13143) );
  OAI21_X1 U16328 ( .B1(n17238), .B2(n18441), .A(n13143), .ZN(n13148) );
  AOI22_X1 U16329 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U16330 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U16331 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13144) );
  NAND3_X1 U16332 ( .A1(n13146), .A2(n13145), .A3(n13144), .ZN(n13147) );
  AOI211_X1 U16333 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n13148), .B(n13147), .ZN(n13149) );
  OAI211_X1 U16334 ( .C1(n13155), .C2(n17216), .A(n13150), .B(n13149), .ZN(
        n13151) );
  AOI22_X1 U16335 ( .A1(n17359), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13163) );
  INV_X1 U16336 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18820) );
  AOI22_X1 U16337 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U16338 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13153) );
  OAI211_X1 U16339 ( .C1(n9828), .C2(n18820), .A(n13154), .B(n13153), .ZN(
        n13161) );
  AOI22_X1 U16340 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U16341 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16342 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U16343 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13156) );
  NAND4_X1 U16344 ( .A1(n13159), .A2(n13158), .A3(n13157), .A4(n13156), .ZN(
        n13160) );
  NAND2_X1 U16345 ( .A1(n18437), .A2(n15728), .ZN(n15879) );
  AOI22_X1 U16346 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13164) );
  OAI21_X1 U16347 ( .B1(n17238), .B2(n18435), .A(n13164), .ZN(n13173) );
  INV_X1 U16348 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U16349 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13171) );
  INV_X1 U16350 ( .A(n17298), .ZN(n17311) );
  INV_X1 U16351 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U16352 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16353 ( .B1(n9846), .B2(n17349), .A(n13165), .ZN(n13169) );
  INV_X1 U16354 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18834) );
  AOI22_X1 U16355 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U16356 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13166) );
  OAI211_X1 U16357 ( .C1(n9828), .C2(n18834), .A(n13167), .B(n13166), .ZN(
        n13168) );
  AOI211_X1 U16358 ( .C1(n17311), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n13169), .B(n13168), .ZN(n13170) );
  OAI211_X1 U16359 ( .C1(n10408), .C2(n17234), .A(n13171), .B(n13170), .ZN(
        n13172) );
  AOI22_X1 U16360 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13183) );
  INV_X1 U16361 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18850) );
  AOI22_X1 U16362 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17412), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16363 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13174) );
  OAI211_X1 U16364 ( .C1(n9828), .C2(n18850), .A(n13175), .B(n13174), .ZN(
        n13181) );
  AOI22_X1 U16365 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16366 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16367 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13177) );
  NAND2_X1 U16368 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13176) );
  NAND4_X1 U16369 ( .A1(n13179), .A2(n13178), .A3(n13177), .A4(n13176), .ZN(
        n13180) );
  NAND2_X1 U16370 ( .A1(n18432), .A2(n17463), .ZN(n15735) );
  AOI22_X1 U16371 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18903), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13184), .ZN(n13190) );
  AOI22_X1 U16372 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18898), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19055), .ZN(n15714) );
  INV_X1 U16373 ( .A(n15714), .ZN(n13189) );
  NAND2_X1 U16374 ( .A1(n18897), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15713) );
  NAND2_X1 U16375 ( .A1(n13190), .A2(n13191), .ZN(n13186) );
  OAI22_X1 U16376 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18405), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13187), .ZN(n13192) );
  NOR2_X1 U16377 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18405), .ZN(
        n13188) );
  NAND2_X1 U16378 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13187), .ZN(
        n13193) );
  AOI22_X1 U16379 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13192), .B1(
        n13188), .B2(n13193), .ZN(n13198) );
  OAI21_X1 U16380 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18897), .A(
        n15713), .ZN(n15873) );
  NOR2_X1 U16381 ( .A1(n13189), .A2(n15873), .ZN(n13197) );
  XNOR2_X1 U16382 ( .A(n13191), .B(n13190), .ZN(n13196) );
  INV_X1 U16383 ( .A(n13198), .ZN(n13195) );
  AOI21_X1 U16384 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13193), .A(
        n13192), .ZN(n13194) );
  AOI21_X1 U16385 ( .B1(n13198), .B2(n13197), .A(n15874), .ZN(n13199) );
  NOR2_X1 U16386 ( .A1(n17463), .A2(n18437), .ZN(n15717) );
  NAND4_X1 U16387 ( .A1(n17577), .A2(n15728), .A3(n15716), .A4(n15717), .ZN(
        n13200) );
  AOI22_X1 U16388 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U16389 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13201) );
  OAI211_X1 U16390 ( .C1(n9828), .C2(n18813), .A(n13202), .B(n13201), .ZN(
        n13208) );
  AOI22_X1 U16391 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U16392 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16393 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16394 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13203) );
  NAND4_X1 U16395 ( .A1(n13206), .A2(n13205), .A3(n13204), .A4(n13203), .ZN(
        n13207) );
  NAND2_X1 U16396 ( .A1(n17577), .A2(n17459), .ZN(n17453) );
  INV_X2 U16397 ( .A(n17456), .ZN(n17451) );
  INV_X1 U16398 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16851) );
  INV_X1 U16399 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16875) );
  INV_X1 U16400 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17274) );
  INV_X1 U16401 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17278) );
  INV_X1 U16402 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17458) );
  INV_X1 U16403 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17452) );
  NOR2_X1 U16404 ( .A1(n17458), .A2(n17452), .ZN(n17447) );
  NAND4_X1 U16405 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n17447), .ZN(n17436) );
  NAND4_X1 U16406 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n17392) );
  NAND4_X1 U16407 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n13212)
         );
  NAND4_X1 U16408 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), .ZN(n13211)
         );
  OR4_X1 U16409 ( .A1(n17436), .A2(n17392), .A3(n13212), .A4(n13211), .ZN(
        n17279) );
  NAND2_X1 U16410 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17260), .ZN(n17258) );
  NOR2_X1 U16411 ( .A1(n18449), .A2(n17258), .ZN(n17244) );
  NAND2_X1 U16412 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17244), .ZN(n17230) );
  NOR2_X1 U16413 ( .A1(n16875), .A2(n17230), .ZN(n17199) );
  NAND2_X1 U16414 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17199), .ZN(n17193) );
  NAND2_X1 U16415 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17192), .ZN(n17177) );
  INV_X1 U16416 ( .A(n17177), .ZN(n17187) );
  NAND2_X1 U16417 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17187), .ZN(n17182) );
  NAND2_X1 U16418 ( .A1(n17451), .A2(n17182), .ZN(n13213) );
  OAI21_X1 U16419 ( .B1(n17171), .B2(n17453), .A(n13213), .ZN(n17172) );
  INV_X1 U16420 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U16421 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13214) );
  OAI21_X1 U16422 ( .B1(n17238), .B2(n17221), .A(n13214), .ZN(n13223) );
  INV_X1 U16423 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15700) );
  AOI22_X1 U16424 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U16425 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13215) );
  OAI21_X1 U16426 ( .B1(n15793), .B2(n15691), .A(n13215), .ZN(n13219) );
  INV_X1 U16427 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15798) );
  AOI22_X1 U16428 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U16429 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13216) );
  OAI211_X1 U16430 ( .C1(n9846), .C2(n15798), .A(n13217), .B(n13216), .ZN(
        n13218) );
  AOI211_X1 U16431 ( .C1(n9965), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13219), .B(n13218), .ZN(n13220) );
  OAI211_X1 U16432 ( .C1(n10408), .C2(n15700), .A(n13221), .B(n13220), .ZN(
        n13222) );
  AOI211_X1 U16433 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13223), .B(n13222), .ZN(n13286) );
  AOI22_X1 U16434 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13224) );
  OAI21_X1 U16435 ( .B1(n17396), .B2(n15752), .A(n13224), .ZN(n13233) );
  INV_X1 U16436 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U16437 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16438 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16439 ( .B1(n15787), .B2(n18654), .A(n13225), .ZN(n13229) );
  INV_X1 U16440 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U16441 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16442 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13226) );
  OAI211_X1 U16443 ( .C1(n9828), .C2(n17362), .A(n13227), .B(n13226), .ZN(
        n13228) );
  AOI211_X1 U16444 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n13229), .B(n13228), .ZN(n13230) );
  OAI211_X1 U16445 ( .C1(n10419), .C2(n17248), .A(n13231), .B(n13230), .ZN(
        n13232) );
  AOI211_X1 U16446 ( .C1(n13275), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n13233), .B(n13232), .ZN(n17180) );
  INV_X1 U16447 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18419) );
  AOI22_X1 U16448 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U16449 ( .B1(n9885), .B2(n18419), .A(n13234), .ZN(n13244) );
  INV_X1 U16450 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18649) );
  AOI22_X1 U16451 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13242) );
  INV_X1 U16452 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16453 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16454 ( .B1(n9846), .B2(n13236), .A(n13235), .ZN(n13240) );
  AOI22_X1 U16455 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16456 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U16457 ( .C1(n17298), .C2(n17397), .A(n13238), .B(n13237), .ZN(
        n13239) );
  AOI211_X1 U16458 ( .C1(n9965), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n13240), .B(n13239), .ZN(n13241) );
  OAI211_X1 U16459 ( .C1(n15787), .C2(n18649), .A(n13242), .B(n13241), .ZN(
        n13243) );
  AOI211_X1 U16460 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n13244), .B(n13243), .ZN(n17189) );
  AOI22_X1 U16461 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16462 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16463 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13245) );
  OAI211_X1 U16464 ( .C1(n9846), .C2(n17414), .A(n13246), .B(n13245), .ZN(
        n13252) );
  AOI22_X1 U16465 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16466 ( .A1(n17359), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U16467 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U16468 ( .A1(n9965), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13247) );
  NAND4_X1 U16469 ( .A1(n13250), .A2(n13249), .A3(n13248), .A4(n13247), .ZN(
        n13251) );
  AOI211_X1 U16470 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n13252), .B(n13251), .ZN(n13253) );
  OAI211_X1 U16471 ( .C1(n15787), .C2(n18646), .A(n13254), .B(n13253), .ZN(
        n17195) );
  AOI22_X1 U16472 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13264) );
  AOI22_X1 U16473 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n9830), .ZN(n13256) );
  AOI22_X1 U16474 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17417), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17398), .ZN(n13255) );
  OAI211_X1 U16475 ( .C1(n17143), .C2(n9828), .A(n13256), .B(n13255), .ZN(
        n13262) );
  AOI22_X1 U16476 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17359), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U16477 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n13106), .ZN(n13259) );
  AOI22_X1 U16478 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16479 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13257) );
  NAND4_X1 U16480 ( .A1(n13260), .A2(n13259), .A3(n13258), .A4(n13257), .ZN(
        n13261) );
  AOI211_X1 U16481 ( .C1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .C2(n17311), .A(
        n13262), .B(n13261), .ZN(n13263) );
  OAI211_X1 U16482 ( .C1(n10419), .C2(n18454), .A(n13264), .B(n13263), .ZN(
        n17196) );
  NAND2_X1 U16483 ( .A1(n17195), .A2(n17196), .ZN(n17194) );
  NOR2_X1 U16484 ( .A1(n17189), .A2(n17194), .ZN(n17188) );
  INV_X1 U16485 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18623) );
  AOI22_X1 U16486 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16487 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16488 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13265) );
  OAI211_X1 U16489 ( .C1(n15793), .C2(n17262), .A(n13266), .B(n13265), .ZN(
        n13272) );
  AOI22_X1 U16490 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U16491 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U16492 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16493 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13267) );
  NAND4_X1 U16494 ( .A1(n13270), .A2(n13269), .A3(n13268), .A4(n13267), .ZN(
        n13271) );
  AOI211_X1 U16495 ( .C1(n9965), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n13272), .B(n13271), .ZN(n13273) );
  OAI211_X1 U16496 ( .C1(n17344), .C2(n18623), .A(n13274), .B(n13273), .ZN(
        n17185) );
  NAND2_X1 U16497 ( .A1(n17188), .A2(n17185), .ZN(n17184) );
  NOR2_X1 U16498 ( .A1(n17180), .A2(n17184), .ZN(n17179) );
  AOI22_X1 U16499 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13285) );
  INV_X1 U16500 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U16501 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16502 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13276) );
  OAI211_X1 U16503 ( .C1(n9828), .C2(n17346), .A(n13277), .B(n13276), .ZN(
        n13283) );
  AOI22_X1 U16504 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16505 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16506 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U16507 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13278) );
  NAND4_X1 U16508 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13282) );
  AOI211_X1 U16509 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n13283), .B(n13282), .ZN(n13284) );
  OAI211_X1 U16510 ( .C1(n10419), .C2(n17349), .A(n13285), .B(n13284), .ZN(
        n17175) );
  NAND2_X1 U16511 ( .A1(n17179), .A2(n17175), .ZN(n17174) );
  NOR2_X1 U16512 ( .A1(n13286), .A2(n17174), .ZN(n17169) );
  AOI21_X1 U16513 ( .B1(n13286), .B2(n17174), .A(n17169), .ZN(n17474) );
  AOI22_X1 U16514 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17172), .B1(n17474), 
        .B2(n17456), .ZN(n13290) );
  INV_X1 U16515 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13288) );
  INV_X1 U16516 ( .A(n17182), .ZN(n13287) );
  NAND3_X1 U16517 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13288), .A3(n13287), 
        .ZN(n13289) );
  NAND2_X1 U16518 ( .A1(n13290), .A2(n13289), .ZN(P3_U2675) );
  NOR2_X1 U16519 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21025), .ZN(n13314) );
  INV_X1 U16520 ( .A(n20710), .ZN(n13305) );
  INV_X1 U16521 ( .A(n14974), .ZN(n13303) );
  AOI21_X1 U16522 ( .B1(n13295), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13292), .ZN(n13297) );
  INV_X1 U16523 ( .A(n14373), .ZN(n15947) );
  MUX2_X1 U16524 ( .A(n13292), .B(n11214), .S(n13291), .Z(n13294) );
  OAI21_X1 U16525 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13296) );
  OAI21_X1 U16526 ( .B1(n13297), .B2(n15947), .A(n13296), .ZN(n13302) );
  OAI21_X1 U16527 ( .B1(n13299), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13298), .ZN(n14985) );
  NOR3_X1 U16528 ( .A1(n14369), .A2(n13300), .A3(n14985), .ZN(n13301) );
  AOI211_X1 U16529 ( .C1(n13303), .C2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13302), .B(n13301), .ZN(n13304) );
  OAI21_X1 U16530 ( .B1(n13305), .B2(n14975), .A(n13304), .ZN(n14984) );
  MUX2_X1 U16531 ( .A(n14984), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15949), .Z(n15959) );
  AOI22_X1 U16532 ( .A1(n13314), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21025), .B2(n15959), .ZN(n13308) );
  MUX2_X1 U16533 ( .A(n13306), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15949), .Z(n15955) );
  AOI22_X1 U16534 ( .A1(n15955), .A2(n21025), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13314), .ZN(n13307) );
  OR2_X1 U16535 ( .A1(n13308), .A2(n13307), .ZN(n15961) );
  OR2_X1 U16536 ( .A1(n15961), .A2(n14971), .ZN(n13322) );
  OR2_X1 U16537 ( .A1(n13309), .A2(n10122), .ZN(n13310) );
  XNOR2_X1 U16538 ( .A(n13310), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20308) );
  INV_X1 U16539 ( .A(n20308), .ZN(n13311) );
  NOR2_X1 U16540 ( .A1(n13311), .A2(n12888), .ZN(n16241) );
  OAI21_X1 U16541 ( .B1(n15949), .B2(n16241), .A(n21025), .ZN(n13312) );
  AOI21_X1 U16542 ( .B1(n15949), .B2(n11600), .A(n13312), .ZN(n13313) );
  AOI21_X1 U16543 ( .B1(n13314), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13313), .ZN(n15968) );
  AND3_X1 U16544 ( .A1(n13322), .A2(n21311), .A3(n15968), .ZN(n13315) );
  NOR2_X1 U16545 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21105) );
  INV_X1 U16546 ( .A(n20593), .ZN(n20427) );
  INV_X1 U16547 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U16548 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20847), .ZN(n13351) );
  INV_X1 U16549 ( .A(n13351), .ZN(n14968) );
  NOR2_X1 U16550 ( .A1(n20845), .A2(n14968), .ZN(n13319) );
  NAND2_X1 U16551 ( .A1(n13316), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13349) );
  NAND2_X1 U16552 ( .A1(n13349), .A2(n20842), .ZN(n20808) );
  INV_X1 U16553 ( .A(n20808), .ZN(n20554) );
  NOR2_X1 U16554 ( .A1(n13349), .A2(n20967), .ZN(n13317) );
  MUX2_X1 U16555 ( .A(n20554), .B(n13317), .S(n12986), .Z(n13318) );
  OAI21_X1 U16556 ( .B1(n13319), .B2(n13318), .A(n20413), .ZN(n13320) );
  OAI21_X1 U16557 ( .B1(n20413), .B2(n20764), .A(n13320), .ZN(P1_U3476) );
  NAND3_X1 U16558 ( .A1(n13322), .A2(n15968), .A3(n13321), .ZN(n15982) );
  INV_X1 U16559 ( .A(n15982), .ZN(n13324) );
  INV_X1 U16560 ( .A(n14370), .ZN(n20552) );
  OAI22_X1 U16561 ( .A1(n20513), .A2(n20967), .B1(n20552), .B2(n14968), .ZN(
        n13323) );
  OAI21_X1 U16562 ( .B1(n13324), .B2(n13323), .A(n20413), .ZN(n13325) );
  OAI21_X1 U16563 ( .B1(n20413), .B2(n20889), .A(n13325), .ZN(P1_U3478) );
  NAND2_X1 U16564 ( .A1(n13326), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13327) );
  NAND2_X1 U16565 ( .A1(n13328), .A2(n13327), .ZN(n13663) );
  INV_X1 U16566 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20393) );
  XNOR2_X1 U16567 ( .A(n13663), .B(n20393), .ZN(n13336) );
  INV_X1 U16568 ( .A(n13756), .ZN(n13766) );
  NAND2_X1 U16569 ( .A1(n20419), .A2(n13766), .ZN(n13334) );
  NAND2_X1 U16570 ( .A1(n13330), .A2(n13329), .ZN(n13675) );
  INV_X1 U16571 ( .A(n13673), .ZN(n13331) );
  XNOR2_X1 U16572 ( .A(n13675), .B(n13331), .ZN(n13332) );
  NAND2_X1 U16573 ( .A1(n13332), .A2(n13772), .ZN(n13333) );
  NAND2_X1 U16574 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  NAND2_X1 U16575 ( .A1(n13336), .A2(n13335), .ZN(n13665) );
  OR2_X1 U16576 ( .A1(n13336), .A2(n13335), .ZN(n13337) );
  NAND2_X1 U16577 ( .A1(n13665), .A2(n13337), .ZN(n20388) );
  INV_X1 U16578 ( .A(n13710), .ZN(n13340) );
  INV_X1 U16579 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13444) );
  NOR2_X1 U16580 ( .A1(n16210), .A2(n13444), .ZN(n20385) );
  AOI21_X1 U16581 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20385), .ZN(n13338) );
  OAI21_X1 U16582 ( .B1(n20374), .B2(n13443), .A(n13338), .ZN(n13339) );
  AOI21_X1 U16583 ( .B1(n13340), .B2(n14411), .A(n13339), .ZN(n13341) );
  OAI21_X1 U16584 ( .B1(n20242), .B2(n20388), .A(n13341), .ZN(P1_U2996) );
  AOI21_X1 U16585 ( .B1(n13342), .B2(n13367), .A(n13374), .ZN(n19267) );
  INV_X1 U16586 ( .A(n19267), .ZN(n13346) );
  OAI211_X1 U16587 ( .C1(n9957), .C2(n10283), .A(n15110), .B(n13373), .ZN(
        n13345) );
  NAND2_X1 U16588 ( .A1(n9831), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13344) );
  OAI211_X1 U16589 ( .C1(n13346), .C2(n9831), .A(n13345), .B(n13344), .ZN(
        P2_U2879) );
  INV_X1 U16590 ( .A(n20413), .ZN(n13355) );
  OAI21_X1 U16591 ( .B1(n20815), .B2(n21220), .A(n20419), .ZN(n13348) );
  OAI21_X1 U16592 ( .B1(n20686), .B2(n13349), .A(n13348), .ZN(n13352) );
  INV_X1 U16593 ( .A(n13316), .ZN(n20972) );
  NOR3_X1 U16594 ( .A1(n20934), .A2(n20967), .A3(n21220), .ZN(n20970) );
  AOI222_X1 U16595 ( .A1(n13352), .A2(n20842), .B1(n20972), .B2(n20970), .C1(
        n20710), .C2(n13351), .ZN(n13354) );
  NAND2_X1 U16596 ( .A1(n13355), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13353) );
  OAI21_X1 U16597 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(P1_U3475) );
  MUX2_X1 U16598 ( .A(n12391), .B(n19330), .S(n15104), .Z(n13360) );
  OAI21_X1 U16599 ( .B1(n19667), .B2(n15106), .A(n13360), .ZN(P2_U2886) );
  NOR2_X1 U16600 ( .A1(n13481), .A2(n9831), .ZN(n13361) );
  AOI21_X1 U16601 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n9831), .A(n13361), .ZN(
        n13362) );
  OAI21_X1 U16602 ( .B1(n19583), .B2(n15106), .A(n13362), .ZN(P2_U2884) );
  AOI21_X1 U16603 ( .B1(n9833), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13363) );
  AND2_X1 U16604 ( .A1(n13364), .A2(n13363), .ZN(n13365) );
  MUX2_X1 U16605 ( .A(n12390), .B(n19350), .S(n15104), .Z(n13366) );
  OAI21_X1 U16606 ( .B1(n20194), .B2(n15106), .A(n13366), .ZN(P2_U2887) );
  XNOR2_X1 U16607 ( .A(n13091), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13371) );
  OAI21_X1 U16608 ( .B1(n13369), .B2(n13368), .A(n13367), .ZN(n19281) );
  MUX2_X1 U16609 ( .A(n12458), .B(n19281), .S(n15104), .Z(n13370) );
  OAI21_X1 U16610 ( .B1(n13371), .B2(n15106), .A(n13370), .ZN(P2_U2880) );
  XNOR2_X1 U16611 ( .A(n13373), .B(n13372), .ZN(n13377) );
  OAI21_X1 U16612 ( .B1(n13375), .B2(n13374), .A(n13436), .ZN(n19260) );
  MUX2_X1 U16613 ( .A(n10207), .B(n19260), .S(n15104), .Z(n13376) );
  OAI21_X1 U16614 ( .B1(n13377), .B2(n15106), .A(n13376), .ZN(P2_U2878) );
  OR2_X1 U16615 ( .A1(n13379), .A2(n13378), .ZN(n13380) );
  AND2_X1 U16616 ( .A1(n13387), .A2(n13380), .ZN(n20379) );
  INV_X1 U16617 ( .A(n20379), .ZN(n20312) );
  INV_X1 U16618 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21259) );
  INV_X1 U16619 ( .A(n13383), .ZN(n13381) );
  XNOR2_X1 U16620 ( .A(n13384), .B(n13381), .ZN(n20369) );
  INV_X1 U16621 ( .A(n20369), .ZN(n13635) );
  OAI222_X1 U16622 ( .A1(n14613), .A2(n20312), .B1(n14612), .B2(n21259), .C1(
        n14610), .C2(n13635), .ZN(P1_U2868) );
  OAI21_X1 U16623 ( .B1(n13384), .B2(n13383), .A(n13382), .ZN(n13385) );
  AND2_X1 U16624 ( .A1(n13385), .A2(n13608), .ZN(n20302) );
  INV_X1 U16625 ( .A(n20302), .ZN(n13708) );
  NAND2_X1 U16626 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  NAND2_X1 U16627 ( .A1(n13603), .A2(n13388), .ZN(n20299) );
  INV_X1 U16628 ( .A(n20299), .ZN(n16232) );
  AOI22_X1 U16629 ( .A1(n14601), .A2(n16232), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14600), .ZN(n13389) );
  OAI21_X1 U16630 ( .B1(n13708), .B2(n14610), .A(n13389), .ZN(P1_U2867) );
  NAND2_X1 U16631 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21105), .ZN(n15979) );
  AND2_X1 U16632 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21026), .ZN(n13390) );
  NAND2_X1 U16633 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  OAI21_X1 U16634 ( .B1(n15979), .B2(n21026), .A(n13392), .ZN(n13393) );
  OR2_X1 U16635 ( .A1(n20440), .A2(n15996), .ZN(n13395) );
  NAND2_X1 U16636 ( .A1(n21110), .A2(n21220), .ZN(n15972) );
  INV_X1 U16637 ( .A(n15972), .ZN(n13410) );
  NAND2_X1 U16638 ( .A1(n13395), .A2(n13410), .ZN(n13408) );
  INV_X1 U16639 ( .A(n13408), .ZN(n13396) );
  INV_X1 U16640 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14683) );
  NOR2_X1 U16641 ( .A1(n13397), .A2(n14683), .ZN(n13398) );
  XNOR2_X1 U16642 ( .A(n13398), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14409) );
  NOR2_X1 U16643 ( .A1(n14409), .A2(n21025), .ZN(n13399) );
  INV_X1 U16644 ( .A(n13404), .ZN(n13401) );
  NAND2_X1 U16645 ( .A1(n13401), .A2(n13400), .ZN(n13402) );
  NAND2_X1 U16646 ( .A1(n16051), .A2(n13402), .ZN(n20321) );
  NOR2_X1 U16647 ( .A1(n13404), .A2(n13403), .ZN(n20309) );
  NAND2_X1 U16648 ( .A1(n20309), .A2(n14370), .ZN(n13407) );
  AND2_X2 U16649 ( .A1(n20277), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20307) );
  AND2_X1 U16650 ( .A1(n14409), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16651 ( .B1(n20307), .B2(n20264), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13406) );
  NAND2_X1 U16652 ( .A1(n13407), .A2(n13406), .ZN(n13416) );
  NAND2_X1 U16653 ( .A1(n20440), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13411) );
  AND2_X1 U16654 ( .A1(n13408), .A2(n13411), .ZN(n13409) );
  NOR2_X1 U16655 ( .A1(n13411), .A2(n13410), .ZN(n13412) );
  OAI22_X1 U16656 ( .A1(n21314), .A2(n20297), .B1(n20313), .B2(n13414), .ZN(
        n13415) );
  AOI211_X1 U16657 ( .C1(n13417), .C2(n20321), .A(n13416), .B(n13415), .ZN(
        n13418) );
  OAI21_X1 U16658 ( .B1(n20279), .B2(n12796), .A(n13418), .ZN(P1_U2840) );
  INV_X1 U16659 ( .A(n20321), .ZN(n13449) );
  AOI22_X1 U16660 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n20315), .B1(n20288), .B2(
        n20403), .ZN(n13425) );
  XOR2_X1 U16661 ( .A(P1_REIP_REG_2__SCAN_IN), .B(P1_REIP_REG_1__SCAN_IN), .Z(
        n13423) );
  INV_X1 U16662 ( .A(n20845), .ZN(n20429) );
  NAND2_X1 U16663 ( .A1(n20309), .A2(n20429), .ZN(n13420) );
  INV_X1 U16664 ( .A(n20277), .ZN(n13640) );
  AOI22_X1 U16665 ( .A1(n20307), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13640), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13419) );
  OAI211_X1 U16666 ( .C1(n20324), .C2(n13421), .A(n13420), .B(n13419), .ZN(
        n13422) );
  AOI21_X1 U16667 ( .B1(n20270), .B2(n13423), .A(n13422), .ZN(n13424) );
  OAI211_X1 U16668 ( .C1(n13701), .C2(n13449), .A(n13425), .B(n13424), .ZN(
        P1_U2838) );
  AOI22_X1 U16669 ( .A1(n20288), .A2(n13426), .B1(n20315), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13431) );
  INV_X1 U16670 ( .A(n20932), .ZN(n20936) );
  NAND2_X1 U16671 ( .A1(n20309), .A2(n20936), .ZN(n13428) );
  AOI22_X1 U16672 ( .A1(n20307), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13640), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13427) );
  OAI211_X1 U16673 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20324), .A(
        n13428), .B(n13427), .ZN(n13429) );
  AOI21_X1 U16674 ( .B1(n20270), .B2(n12958), .A(n13429), .ZN(n13430) );
  OAI211_X1 U16675 ( .C1(n13449), .C2(n13709), .A(n13431), .B(n13430), .ZN(
        P1_U2839) );
  OAI211_X1 U16676 ( .C1(n13434), .C2(n13433), .A(n13613), .B(n15110), .ZN(
        n13439) );
  AOI21_X1 U16677 ( .B1(n13437), .B2(n13436), .A(n13435), .ZN(n19247) );
  NAND2_X1 U16678 ( .A1(n19247), .A2(n15104), .ZN(n13438) );
  OAI211_X1 U16679 ( .C1(n15104), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        P2_U2877) );
  OAI221_X1 U16680 ( .B1(n20318), .B2(P1_REIP_REG_2__SCAN_IN), .C1(n20318), 
        .C2(P1_REIP_REG_1__SCAN_IN), .A(n20277), .ZN(n13441) );
  AOI22_X1 U16681 ( .A1(n20307), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13441), .ZN(n13442) );
  OAI21_X1 U16682 ( .B1(n20324), .B2(n13443), .A(n13442), .ZN(n13446) );
  AND4_X1 U16683 ( .A1(n20270), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n13444), .ZN(n13445) );
  AOI211_X1 U16684 ( .C1(n20309), .C2(n20710), .A(n13446), .B(n13445), .ZN(
        n13448) );
  AOI22_X1 U16685 ( .A1(n20288), .A2(n20386), .B1(n20315), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13447) );
  OAI211_X1 U16686 ( .C1(n13449), .C2(n13710), .A(n13448), .B(n13447), .ZN(
        P1_U2837) );
  XNOR2_X1 U16687 ( .A(n13613), .B(n13612), .ZN(n13451) );
  MUX2_X1 U16688 ( .A(n11122), .B(n16401), .S(n15104), .Z(n13450) );
  OAI21_X1 U16689 ( .B1(n13451), .B2(n15106), .A(n13450), .ZN(P2_U2876) );
  INV_X1 U16690 ( .A(n19584), .ZN(n13452) );
  OR2_X1 U16691 ( .A1(n19583), .A2(n12714), .ZN(n19872) );
  OAI21_X1 U16692 ( .B1(n13452), .B2(n19872), .A(n20169), .ZN(n13461) );
  NAND2_X1 U16693 ( .A1(n20181), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19869) );
  OR2_X1 U16694 ( .A1(n19869), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19784) );
  INV_X1 U16695 ( .A(n19784), .ZN(n13457) );
  NOR2_X1 U16696 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16548) );
  INV_X1 U16697 ( .A(n16548), .ZN(n20215) );
  NAND2_X1 U16698 ( .A1(n20215), .A2(n20191), .ZN(n13453) );
  NOR2_X1 U16699 ( .A1(n13481), .A2(n19509), .ZN(n13454) );
  OR2_X1 U16700 ( .A1(n10696), .A2(n19350), .ZN(n13496) );
  INV_X1 U16701 ( .A(n13496), .ZN(n13490) );
  INV_X1 U16702 ( .A(n20169), .ZN(n19973) );
  NOR2_X1 U16703 ( .A1(n19574), .A2(n19869), .ZN(n19840) );
  INV_X1 U16704 ( .A(n19840), .ZN(n13455) );
  OAI211_X1 U16705 ( .C1(n13531), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19973), 
        .B(n13455), .ZN(n13456) );
  OAI211_X1 U16706 ( .C1(n13461), .C2(n13457), .A(n19975), .B(n13456), .ZN(
        n19831) );
  INV_X1 U16707 ( .A(n19831), .ZN(n13467) );
  INV_X1 U16708 ( .A(n13531), .ZN(n13459) );
  OAI21_X1 U16709 ( .B1(n13459), .B2(n19840), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13460) );
  OAI21_X1 U16710 ( .B1(n13461), .B2(n19784), .A(n13460), .ZN(n19830) );
  INV_X1 U16711 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18409) );
  INV_X1 U16712 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20421) );
  INV_X1 U16713 ( .A(n19946), .ZN(n20028) );
  AOI22_X1 U16714 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19559), .ZN(n19949) );
  INV_X1 U16715 ( .A(n19949), .ZN(n20025) );
  NOR2_X2 U16716 ( .A1(n16528), .A2(n19564), .ZN(n20016) );
  AOI22_X1 U16717 ( .A1(n20025), .A2(n19859), .B1(n20016), .B2(n19840), .ZN(
        n13463) );
  OAI21_X1 U16718 ( .B1(n20028), .B2(n19826), .A(n13463), .ZN(n13464) );
  AOI21_X1 U16719 ( .B1(n13458), .B2(n19830), .A(n13464), .ZN(n13465) );
  OAI21_X1 U16720 ( .B1(n13467), .B2(n13466), .A(n13465), .ZN(P2_U3120) );
  INV_X1 U16721 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13470) );
  INV_X1 U16722 ( .A(n13489), .ZN(n13471) );
  OAI22_X1 U16723 ( .A1(n13470), .A2(n19636), .B1(n19516), .B2(n13469), .ZN(
        n13475) );
  INV_X1 U16724 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13473) );
  OAI22_X1 U16725 ( .A1(n13473), .A2(n20011), .B1(n19938), .B2(n13472), .ZN(
        n13474) );
  NOR2_X1 U16726 ( .A1(n13475), .A2(n13474), .ZN(n13510) );
  INV_X1 U16727 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13477) );
  OAI22_X1 U16728 ( .A1(n13478), .A2(n19786), .B1(n19899), .B2(n13477), .ZN(
        n13486) );
  AND2_X1 U16729 ( .A1(n13479), .A2(n19350), .ZN(n13501) );
  INV_X1 U16730 ( .A(n13501), .ZN(n13495) );
  AND2_X2 U16731 ( .A1(n13481), .A2(n19509), .ZN(n13502) );
  INV_X1 U16732 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13483) );
  OAI22_X1 U16733 ( .A1(n19977), .A2(n13484), .B1(n13787), .B2(n13483), .ZN(
        n13485) );
  NOR2_X1 U16734 ( .A1(n13486), .A2(n13485), .ZN(n13509) );
  INV_X1 U16735 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13488) );
  OAI22_X1 U16736 ( .A1(n13488), .A2(n19868), .B1(n13531), .B2(n13487), .ZN(
        n13494) );
  INV_X1 U16737 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16738 ( .A1(n13502), .A2(n13489), .ZN(n19760) );
  NAND2_X1 U16739 ( .A1(n13502), .A2(n13490), .ZN(n19697) );
  OAI22_X1 U16740 ( .A1(n13492), .A2(n19760), .B1(n19697), .B2(n13491), .ZN(
        n13493) );
  NOR2_X1 U16741 ( .A1(n13494), .A2(n13493), .ZN(n13508) );
  OAI22_X1 U16742 ( .A1(n13499), .A2(n13805), .B1(n19572), .B2(n13498), .ZN(
        n13506) );
  NAND2_X1 U16743 ( .A1(n13502), .A2(n13501), .ZN(n19726) );
  OAI22_X1 U16744 ( .A1(n13784), .A2(n13504), .B1(n19726), .B2(n13503), .ZN(
        n13505) );
  NOR2_X1 U16745 ( .A1(n13506), .A2(n13505), .ZN(n13507) );
  INV_X1 U16746 ( .A(n13511), .ZN(n13512) );
  NAND2_X1 U16747 ( .A1(n13512), .A2(n9839), .ZN(n13513) );
  INV_X1 U16748 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13515) );
  OAI22_X1 U16749 ( .A1(n19786), .A2(n13516), .B1(n19726), .B2(n10590), .ZN(
        n13517) );
  NOR2_X1 U16750 ( .A1(n13518), .A2(n13517), .ZN(n13540) );
  INV_X1 U16751 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13519) );
  OAI22_X1 U16752 ( .A1(n13519), .A2(n19868), .B1(n19636), .B2(n10589), .ZN(
        n13523) );
  INV_X1 U16753 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13521) );
  OAI22_X1 U16754 ( .A1(n13521), .A2(n13784), .B1(n19516), .B2(n13520), .ZN(
        n13522) );
  NOR2_X1 U16755 ( .A1(n13523), .A2(n13522), .ZN(n13539) );
  INV_X1 U16756 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13525) );
  NAND2_X1 U16757 ( .A1(n19672), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13524) );
  OAI211_X1 U16758 ( .C1(n20011), .C2(n13525), .A(n13524), .B(n9833), .ZN(
        n13529) );
  INV_X1 U16759 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13526) );
  OAI22_X1 U16760 ( .A1(n19977), .A2(n13527), .B1(n19760), .B2(n13526), .ZN(
        n13528) );
  NOR2_X1 U16761 ( .A1(n13529), .A2(n13528), .ZN(n13538) );
  OAI22_X1 U16762 ( .A1(n13532), .A2(n13531), .B1(n19572), .B2(n13530), .ZN(
        n13536) );
  INV_X1 U16763 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13534) );
  OAI22_X1 U16764 ( .A1(n13805), .A2(n13534), .B1(n19697), .B2(n13533), .ZN(
        n13535) );
  NOR2_X1 U16765 ( .A1(n13536), .A2(n13535), .ZN(n13537) );
  INV_X1 U16766 ( .A(n13541), .ZN(n13543) );
  NAND2_X1 U16767 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  OAI21_X1 U16768 ( .B1(n13546), .B2(n13545), .A(n13579), .ZN(n15000) );
  NAND2_X1 U16769 ( .A1(n13549), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13576) );
  NAND2_X1 U16770 ( .A1(n13577), .A2(n13576), .ZN(n13551) );
  NAND2_X1 U16771 ( .A1(n15004), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13550) );
  AND2_X1 U16772 ( .A1(n19506), .A2(n13550), .ZN(n13575) );
  XNOR2_X1 U16773 ( .A(n13551), .B(n13575), .ZN(n13574) );
  NAND2_X1 U16774 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13552), .ZN(
        n13553) );
  NAND2_X1 U16775 ( .A1(n13554), .A2(n13553), .ZN(n13584) );
  XNOR2_X1 U16776 ( .A(n13584), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13582) );
  XOR2_X1 U16777 ( .A(n13583), .B(n13582), .Z(n13572) );
  XNOR2_X1 U16778 ( .A(n13556), .B(n13555), .ZN(n20166) );
  NOR2_X1 U16779 ( .A1(n13568), .A2(n19294), .ZN(n13557) );
  AOI21_X1 U16780 ( .B1(n16485), .B2(n20166), .A(n13557), .ZN(n13558) );
  OAI21_X1 U16781 ( .B1(n13011), .B2(n15640), .A(n13558), .ZN(n13566) );
  INV_X1 U16782 ( .A(n14264), .ZN(n13561) );
  INV_X1 U16783 ( .A(n15519), .ZN(n13563) );
  INV_X1 U16784 ( .A(n13564), .ZN(n13559) );
  NAND2_X1 U16785 ( .A1(n13563), .A2(n13559), .ZN(n13560) );
  AOI21_X1 U16786 ( .B1(n13564), .B2(n13563), .A(n13562), .ZN(n14263) );
  OAI21_X1 U16787 ( .B1(n15512), .B2(n14264), .A(n14263), .ZN(n13888) );
  MUX2_X1 U16788 ( .A(n14274), .B(n13888), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13565) );
  AOI211_X1 U16789 ( .C1(n13572), .C2(n16493), .A(n13566), .B(n13565), .ZN(
        n13567) );
  OAI21_X1 U16790 ( .B1(n13574), .B2(n16477), .A(n13567), .ZN(P2_U3043) );
  OAI22_X1 U16791 ( .A1(n19514), .A2(n14995), .B1(n13568), .B2(n19294), .ZN(
        n13569) );
  AOI21_X1 U16792 ( .B1(n16442), .B2(n14992), .A(n13569), .ZN(n13570) );
  OAI21_X1 U16793 ( .B1(n13011), .B2(n16438), .A(n13570), .ZN(n13571) );
  AOI21_X1 U16794 ( .B1(n13572), .B2(n16449), .A(n13571), .ZN(n13573) );
  OAI21_X1 U16795 ( .B1(n13574), .B2(n19493), .A(n13573), .ZN(P2_U3011) );
  XNOR2_X1 U16796 ( .A(n13579), .B(n13578), .ZN(n19308) );
  XNOR2_X1 U16797 ( .A(n19308), .B(n16480), .ZN(n13826) );
  XNOR2_X1 U16798 ( .A(n13827), .B(n13826), .ZN(n19494) );
  XNOR2_X1 U16799 ( .A(n13872), .B(n16480), .ZN(n13586) );
  NAND2_X1 U16800 ( .A1(n13584), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13585) );
  XNOR2_X1 U16801 ( .A(n13586), .B(n13871), .ZN(n19491) );
  NAND2_X1 U16802 ( .A1(n13588), .A2(n13587), .ZN(n13590) );
  INV_X1 U16803 ( .A(n14082), .ZN(n13589) );
  AND2_X1 U16804 ( .A1(n13590), .A2(n13589), .ZN(n19496) );
  INV_X1 U16805 ( .A(n19496), .ZN(n19311) );
  XNOR2_X1 U16806 ( .A(n13591), .B(n9871), .ZN(n19404) );
  INV_X1 U16807 ( .A(n19404), .ZN(n19399) );
  OAI22_X1 U16808 ( .A1(n19311), .A2(n15640), .B1(n19399), .B2(n16469), .ZN(
        n13594) );
  NAND2_X1 U16809 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14274), .ZN(
        n16479) );
  AOI21_X1 U16810 ( .B1(n13547), .B2(n15517), .A(n13888), .ZN(n16498) );
  NAND2_X1 U16811 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19310), .ZN(n13592) );
  OAI221_X1 U16812 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16479), .C1(
        n16480), .C2(n16498), .A(n13592), .ZN(n13593) );
  AOI211_X1 U16813 ( .C1(n19491), .C2(n16493), .A(n13594), .B(n13593), .ZN(
        n13595) );
  OAI21_X1 U16814 ( .B1(n19494), .B2(n16477), .A(n13595), .ZN(P2_U3042) );
  OR2_X1 U16815 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  AND2_X1 U16816 ( .A1(n13638), .A2(n13599), .ZN(n20281) );
  INV_X1 U16817 ( .A(n20281), .ZN(n13702) );
  AOI21_X1 U16818 ( .B1(n13600), .B2(n13605), .A(n13645), .ZN(n20269) );
  AOI22_X1 U16819 ( .A1(n14601), .A2(n20269), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14600), .ZN(n13601) );
  OAI21_X1 U16820 ( .B1(n13702), .B2(n14610), .A(n13601), .ZN(P1_U2865) );
  NAND2_X1 U16821 ( .A1(n13603), .A2(n13602), .ZN(n13604) );
  NAND2_X1 U16822 ( .A1(n13605), .A2(n13604), .ZN(n20285) );
  INV_X1 U16823 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21248) );
  INV_X1 U16824 ( .A(n13606), .ZN(n13607) );
  XNOR2_X1 U16825 ( .A(n13608), .B(n13607), .ZN(n20291) );
  INV_X1 U16826 ( .A(n20291), .ZN(n13634) );
  OAI222_X1 U16827 ( .A1(n20285), .A2(n14613), .B1(n14612), .B2(n21248), .C1(
        n14610), .C2(n13634), .ZN(P1_U2866) );
  INV_X1 U16828 ( .A(n13609), .ZN(n13611) );
  AOI21_X1 U16829 ( .B1(n13611), .B2(n13610), .A(n13655), .ZN(n19237) );
  INV_X1 U16830 ( .A(n19237), .ZN(n13617) );
  OAI21_X1 U16831 ( .B1(n13613), .B2(n13612), .A(n13952), .ZN(n13614) );
  NAND3_X1 U16832 ( .A1(n13614), .A2(n15110), .A3(n13653), .ZN(n13616) );
  NAND2_X1 U16833 ( .A1(n9831), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13615) );
  OAI211_X1 U16834 ( .C1(n13617), .C2(n9831), .A(n13616), .B(n13615), .ZN(
        P2_U2875) );
  NAND3_X1 U16835 ( .A1(n13620), .A2(n13619), .A3(n13618), .ZN(n13624) );
  NAND2_X1 U16836 ( .A1(n13622), .A2(n13621), .ZN(n13623) );
  NAND2_X1 U16837 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  NAND2_X1 U16838 ( .A1(n14674), .A2(n13632), .ZN(n14666) );
  NOR2_X1 U16839 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  OAI222_X1 U16840 ( .A1(n20473), .A2(n14676), .B1(n14672), .B2(n13634), .C1(
        n11632), .C2(n14647), .ZN(P1_U2898) );
  INV_X1 U16841 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20341) );
  OAI222_X1 U16842 ( .A1(n20459), .A2(n14676), .B1(n14672), .B2(n13635), .C1(
        n20341), .C2(n14647), .ZN(P1_U2900) );
  INV_X1 U16843 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21052) );
  INV_X1 U16844 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21265) );
  NAND3_X1 U16845 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n20317) );
  NOR2_X1 U16846 ( .A1(n21265), .A2(n20317), .ZN(n20276) );
  NAND4_X1 U16847 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20276), .A3(
        P1_REIP_REG_5__SCAN_IN), .A4(P1_REIP_REG_6__SCAN_IN), .ZN(n13647) );
  NOR2_X1 U16848 ( .A1(n21052), .A2(n13647), .ZN(n20257) );
  AND2_X1 U16849 ( .A1(n20277), .A2(n20257), .ZN(n13636) );
  OR2_X1 U16850 ( .A1(n20279), .A2(n13636), .ZN(n20268) );
  INV_X1 U16851 ( .A(n13712), .ZN(n13637) );
  AOI21_X1 U16852 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13779) );
  NAND2_X1 U16853 ( .A1(n13779), .A2(n20292), .ZN(n13652) );
  INV_X1 U16854 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21305) );
  NOR2_X2 U16855 ( .A1(n13640), .A2(n20238), .ZN(n20306) );
  AOI21_X1 U16856 ( .B1(n20307), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20306), .ZN(n13643) );
  INV_X1 U16857 ( .A(n13777), .ZN(n13641) );
  NAND2_X1 U16858 ( .A1(n20264), .A2(n13641), .ZN(n13642) );
  OAI211_X1 U16859 ( .C1(n20297), .C2(n21305), .A(n13643), .B(n13642), .ZN(
        n13650) );
  OR2_X1 U16860 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  AND2_X1 U16861 ( .A1(n13646), .A2(n13715), .ZN(n16221) );
  INV_X1 U16862 ( .A(n16221), .ZN(n13659) );
  OR3_X1 U16863 ( .A1(n20318), .A2(n13647), .A3(P1_REIP_REG_8__SCAN_IN), .ZN(
        n13648) );
  OAI21_X1 U16864 ( .B1(n13659), .B2(n20313), .A(n13648), .ZN(n13649) );
  NOR2_X1 U16865 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  OAI211_X1 U16866 ( .C1(n21052), .C2(n20268), .A(n13652), .B(n13651), .ZN(
        P1_U2832) );
  XNOR2_X1 U16867 ( .A(n13653), .B(n13958), .ZN(n13658) );
  OR2_X1 U16868 ( .A1(n13655), .A2(n13654), .ZN(n13656) );
  NAND2_X1 U16869 ( .A1(n13656), .A2(n13721), .ZN(n19229) );
  MUX2_X1 U16870 ( .A(n19229), .B(n14121), .S(n9831), .Z(n13657) );
  OAI21_X1 U16871 ( .B1(n13658), .B2(n15106), .A(n13657), .ZN(P2_U2874) );
  INV_X1 U16872 ( .A(n13779), .ZN(n13662) );
  OAI222_X1 U16873 ( .A1(n13662), .A2(n14610), .B1(n14612), .B2(n21305), .C1(
        n13659), .C2(n14613), .ZN(P1_U2864) );
  INV_X1 U16874 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13661) );
  NAND2_X1 U16875 ( .A1(n20415), .A2(n12674), .ZN(n13660) );
  OAI21_X1 U16876 ( .B1(n20415), .B2(DATAI_8_), .A(n13660), .ZN(n14635) );
  OAI222_X1 U16877 ( .A1(n13662), .A2(n14672), .B1(n13661), .B2(n14674), .C1(
        n14635), .C2(n14676), .ZN(P1_U2896) );
  NAND2_X1 U16878 ( .A1(n13663), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13664) );
  NAND2_X1 U16879 ( .A1(n13675), .A2(n13673), .ZN(n13666) );
  XNOR2_X1 U16880 ( .A(n13666), .B(n13672), .ZN(n13667) );
  AND2_X1 U16881 ( .A1(n13667), .A2(n13772), .ZN(n13668) );
  AOI21_X1 U16882 ( .B1(n13669), .B2(n13766), .A(n13668), .ZN(n20366) );
  AND2_X1 U16883 ( .A1(n13673), .A2(n13672), .ZN(n13674) );
  NAND2_X1 U16884 ( .A1(n13675), .A2(n13674), .ZN(n13684) );
  XNOR2_X1 U16885 ( .A(n13684), .B(n13759), .ZN(n13676) );
  NAND2_X1 U16886 ( .A1(n13676), .A2(n13772), .ZN(n13677) );
  NAND2_X1 U16887 ( .A1(n13678), .A2(n13677), .ZN(n13681) );
  XNOR2_X1 U16888 ( .A(n13681), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16117) );
  NAND2_X1 U16889 ( .A1(n13681), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13682) );
  NAND2_X1 U16890 ( .A1(n13683), .A2(n13766), .ZN(n13688) );
  INV_X1 U16891 ( .A(n13684), .ZN(n13761) );
  NAND2_X1 U16892 ( .A1(n13761), .A2(n13759), .ZN(n13685) );
  XNOR2_X1 U16893 ( .A(n13685), .B(n13758), .ZN(n13686) );
  NAND2_X1 U16894 ( .A1(n13686), .A2(n13772), .ZN(n13687) );
  NAND2_X1 U16895 ( .A1(n13688), .A2(n13687), .ZN(n13754) );
  XOR2_X1 U16896 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13754), .Z(
        n13689) );
  XNOR2_X1 U16897 ( .A(n13753), .B(n13689), .ZN(n16110) );
  NAND2_X1 U16898 ( .A1(n14958), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14942) );
  NAND2_X1 U16899 ( .A1(n14942), .A2(n13690), .ZN(n14903) );
  NAND2_X1 U16900 ( .A1(n14903), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20412) );
  NAND2_X1 U16901 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20381) );
  NOR2_X1 U16902 ( .A1(n20381), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16235) );
  INV_X1 U16903 ( .A(n16235), .ZN(n13694) );
  INV_X1 U16904 ( .A(n20396), .ZN(n16175) );
  AOI21_X1 U16905 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n16175), .ZN(n20377) );
  NOR2_X1 U16906 ( .A1(n16239), .A2(n20381), .ZN(n13695) );
  AOI21_X1 U16907 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16233) );
  NAND2_X1 U16908 ( .A1(n14958), .A2(n13691), .ZN(n13693) );
  AOI21_X1 U16909 ( .B1(n16180), .B2(n16233), .A(n20395), .ZN(n20375) );
  OAI21_X1 U16910 ( .B1(n13695), .B2(n20398), .A(n20375), .ZN(n16177) );
  OR2_X1 U16911 ( .A1(n20377), .A2(n16177), .ZN(n16199) );
  AOI21_X1 U16912 ( .B1(n20381), .B2(n20396), .A(n16199), .ZN(n16240) );
  OAI211_X1 U16913 ( .C1(n13696), .C2(n13694), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16240), .ZN(n16218) );
  INV_X1 U16914 ( .A(n13695), .ZN(n14351) );
  NOR2_X1 U16915 ( .A1(n16233), .A2(n14351), .ZN(n16197) );
  NAND2_X1 U16916 ( .A1(n16197), .A2(n16234), .ZN(n16222) );
  NAND2_X1 U16917 ( .A1(n12259), .A2(n16222), .ZN(n13699) );
  INV_X1 U16918 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13697) );
  OAI22_X1 U16919 ( .A1(n16211), .A2(n20285), .B1(n16210), .B2(n13697), .ZN(
        n13698) );
  AOI21_X1 U16920 ( .B1(n16218), .B2(n13699), .A(n13698), .ZN(n13700) );
  OAI21_X1 U16921 ( .B1(n20387), .B2(n16110), .A(n13700), .ZN(P1_U3025) );
  INV_X1 U16922 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20345) );
  OAI222_X1 U16923 ( .A1(n14672), .A2(n13701), .B1(n20448), .B2(n14676), .C1(
        n14674), .C2(n20345), .ZN(P1_U2902) );
  INV_X1 U16924 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20337) );
  OAI222_X1 U16925 ( .A1(n14672), .A2(n13702), .B1(n20482), .B2(n14676), .C1(
        n14674), .C2(n20337), .ZN(P1_U2897) );
  XNOR2_X1 U16926 ( .A(n15083), .B(n15082), .ZN(n13706) );
  INV_X1 U16927 ( .A(n14009), .ZN(n13704) );
  NAND2_X1 U16928 ( .A1(n9956), .A2(n9932), .ZN(n13703) );
  NAND2_X1 U16929 ( .A1(n13704), .A2(n13703), .ZN(n19203) );
  MUX2_X1 U16930 ( .A(n14125), .B(n19203), .S(n15104), .Z(n13705) );
  OAI21_X1 U16931 ( .B1(n13706), .B2(n15106), .A(n13705), .ZN(P2_U2872) );
  INV_X1 U16932 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20350) );
  OAI222_X1 U16933 ( .A1(n13707), .A2(n14672), .B1(n14647), .B2(n20350), .C1(
        n20431), .C2(n14676), .ZN(P1_U2904) );
  OAI222_X1 U16934 ( .A1(n13708), .A2(n14672), .B1(n14674), .B2(n11553), .C1(
        n20465), .C2(n14676), .ZN(P1_U2899) );
  INV_X1 U16935 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20347) );
  OAI222_X1 U16936 ( .A1(n13709), .A2(n14672), .B1(n14647), .B2(n20347), .C1(
        n20442), .C2(n14676), .ZN(P1_U2903) );
  INV_X1 U16937 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20343) );
  OAI222_X1 U16938 ( .A1(n13710), .A2(n14672), .B1(n14674), .B2(n20343), .C1(
        n20454), .C2(n14676), .ZN(P1_U2901) );
  AND2_X1 U16939 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  NOR2_X1 U16940 ( .A1(n13731), .A2(n13713), .ZN(n20265) );
  NAND2_X1 U16941 ( .A1(n13715), .A2(n13714), .ZN(n13716) );
  NAND2_X1 U16942 ( .A1(n13735), .A2(n13716), .ZN(n20258) );
  OAI22_X1 U16943 ( .A1(n20258), .A2(n14613), .B1(n14612), .B2(n13717), .ZN(
        n13718) );
  AOI21_X1 U16944 ( .B1(n20265), .B2(n13719), .A(n13718), .ZN(n13720) );
  INV_X1 U16945 ( .A(n13720), .ZN(P1_U2863) );
  NAND2_X1 U16946 ( .A1(n13722), .A2(n13721), .ZN(n13723) );
  AND2_X1 U16947 ( .A1(n13723), .A2(n9932), .ZN(n19214) );
  INV_X1 U16948 ( .A(n19214), .ZN(n15573) );
  INV_X1 U16949 ( .A(n15083), .ZN(n13724) );
  OAI211_X1 U16950 ( .C1(n13725), .C2(n13962), .A(n13724), .B(n15110), .ZN(
        n13727) );
  NAND2_X1 U16951 ( .A1(n9831), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13726) );
  OAI211_X1 U16952 ( .C1(n15573), .C2(n9831), .A(n13727), .B(n13726), .ZN(
        P2_U2873) );
  INV_X1 U16953 ( .A(n20265), .ZN(n13729) );
  INV_X1 U16954 ( .A(DATAI_9_), .ZN(n21343) );
  MUX2_X1 U16955 ( .A(n21343), .B(n16666), .S(n20415), .Z(n14631) );
  INV_X1 U16956 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13728) );
  OAI222_X1 U16957 ( .A1(n13729), .A2(n14672), .B1(n14631), .B2(n14676), .C1(
        n13728), .C2(n14647), .ZN(P1_U2895) );
  INV_X1 U16958 ( .A(n13730), .ZN(n13733) );
  INV_X1 U16959 ( .A(n13731), .ZN(n13732) );
  AOI21_X1 U16960 ( .B1(n13733), .B2(n13732), .A(n13979), .ZN(n14839) );
  INV_X1 U16961 ( .A(n14839), .ZN(n13751) );
  AND2_X1 U16962 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  NOR2_X1 U16963 ( .A1(n14014), .A2(n13736), .ZN(n13742) );
  AOI22_X1 U16964 ( .A1(n14601), .A2(n13742), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14600), .ZN(n13737) );
  OAI21_X1 U16965 ( .B1(n13751), .B2(n14610), .A(n13737), .ZN(P1_U2862) );
  INV_X1 U16966 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21054) );
  NAND2_X1 U16967 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20257), .ZN(n13743) );
  NOR2_X1 U16968 ( .A1(n21054), .A2(n13743), .ZN(n16044) );
  AND2_X1 U16969 ( .A1(n20277), .A2(n16044), .ZN(n13738) );
  NAND2_X1 U16970 ( .A1(n14839), .A2(n20292), .ZN(n13748) );
  AOI21_X1 U16971 ( .B1(n20307), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20306), .ZN(n13741) );
  INV_X1 U16972 ( .A(n14837), .ZN(n13739) );
  NAND2_X1 U16973 ( .A1(n20264), .A2(n13739), .ZN(n13740) );
  OAI211_X1 U16974 ( .C1(n20297), .C2(n21507), .A(n13741), .B(n13740), .ZN(
        n13746) );
  INV_X1 U16975 ( .A(n13742), .ZN(n16202) );
  OR3_X1 U16976 ( .A1(n20318), .A2(n13743), .A3(P1_REIP_REG_10__SCAN_IN), .ZN(
        n13744) );
  OAI21_X1 U16977 ( .B1(n16202), .B2(n20313), .A(n13744), .ZN(n13745) );
  NOR2_X1 U16978 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  OAI211_X1 U16979 ( .C1(n21054), .C2(n16055), .A(n13748), .B(n13747), .ZN(
        P1_U2830) );
  INV_X1 U16980 ( .A(DATAI_10_), .ZN(n13749) );
  MUX2_X1 U16981 ( .A(n13749), .B(n16664), .S(n20415), .Z(n14627) );
  INV_X1 U16982 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13750) );
  OAI222_X1 U16983 ( .A1(n14672), .A2(n13751), .B1(n14627), .B2(n14676), .C1(
        n13750), .C2(n14647), .ZN(P1_U2894) );
  INV_X1 U16984 ( .A(n13755), .ZN(n13757) );
  OR2_X1 U16985 ( .A1(n13757), .A2(n13756), .ZN(n13764) );
  AND2_X1 U16986 ( .A1(n13759), .A2(n13758), .ZN(n13760) );
  NAND2_X1 U16987 ( .A1(n13761), .A2(n13760), .ZN(n13770) );
  XNOR2_X1 U16988 ( .A(n13770), .B(n13771), .ZN(n13762) );
  NAND2_X1 U16989 ( .A1(n13762), .A2(n13772), .ZN(n13763) );
  NAND2_X1 U16990 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  OR2_X1 U16991 ( .A1(n13765), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16105) );
  NAND2_X1 U16992 ( .A1(n13765), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16104) );
  INV_X1 U16993 ( .A(n13770), .ZN(n13773) );
  NAND3_X1 U16994 ( .A1(n13773), .A2(n13772), .A3(n13771), .ZN(n13774) );
  NAND2_X1 U16995 ( .A1(n14805), .A2(n13774), .ZN(n13904) );
  XNOR2_X1 U16996 ( .A(n13904), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13775) );
  XNOR2_X1 U16997 ( .A(n13903), .B(n13775), .ZN(n16220) );
  INV_X1 U16998 ( .A(n16220), .ZN(n13781) );
  AOI22_X1 U16999 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13776) );
  OAI21_X1 U17000 ( .B1(n20374), .B2(n13777), .A(n13776), .ZN(n13778) );
  AOI21_X1 U17001 ( .B1(n13779), .B2(n14411), .A(n13778), .ZN(n13780) );
  OAI21_X1 U17002 ( .B1(n13781), .B2(n20242), .A(n13780), .ZN(P1_U2991) );
  INV_X1 U17003 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13786) );
  OAI22_X1 U17004 ( .A1(n13786), .A2(n13784), .B1(n19572), .B2(n13785), .ZN(
        n13791) );
  INV_X1 U17005 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13788) );
  OAI22_X1 U17006 ( .A1(n19786), .A2(n13789), .B1(n13787), .B2(n13788), .ZN(
        n13790) );
  NOR2_X1 U17007 ( .A1(n13791), .A2(n13790), .ZN(n13813) );
  OAI22_X1 U17008 ( .A1(n13792), .A2(n13531), .B1(n19516), .B2(n10791), .ZN(
        n13796) );
  INV_X1 U17009 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13794) );
  INV_X1 U17010 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13793) );
  OAI22_X1 U17011 ( .A1(n19868), .A2(n13794), .B1(n19760), .B2(n13793), .ZN(
        n13795) );
  NOR2_X1 U17012 ( .A1(n13796), .A2(n13795), .ZN(n13812) );
  INV_X1 U17013 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13798) );
  OAI22_X1 U17014 ( .A1(n13798), .A2(n19636), .B1(n19938), .B2(n13797), .ZN(
        n13802) );
  INV_X1 U17015 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13800) );
  OAI22_X1 U17016 ( .A1(n20011), .A2(n13800), .B1(n19697), .B2(n13799), .ZN(
        n13801) );
  NOR2_X1 U17017 ( .A1(n13802), .A2(n13801), .ZN(n13811) );
  INV_X1 U17018 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13804) );
  OAI22_X1 U17019 ( .A1(n13804), .A2(n19899), .B1(n19977), .B2(n13803), .ZN(
        n13809) );
  INV_X1 U17020 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13807) );
  OAI22_X1 U17021 ( .A1(n13805), .A2(n13807), .B1(n19726), .B2(n13806), .ZN(
        n13808) );
  NOR2_X1 U17022 ( .A1(n13809), .A2(n13808), .ZN(n13810) );
  NAND4_X1 U17023 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        n13817) );
  INV_X1 U17024 ( .A(n13814), .ZN(n13815) );
  NAND2_X1 U17025 ( .A1(n13815), .A2(n9838), .ZN(n13816) );
  NAND2_X1 U17026 ( .A1(n13817), .A2(n13816), .ZN(n13820) );
  NAND2_X1 U17027 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  NOR2_X1 U17028 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  OR2_X1 U17029 ( .A1(n13866), .A2(n13825), .ZN(n19296) );
  NAND2_X1 U17030 ( .A1(n13828), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13829) );
  NAND2_X1 U17031 ( .A1(n13830), .A2(n13829), .ZN(n13922) );
  INV_X1 U17032 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13832) );
  OAI22_X1 U17033 ( .A1(n13832), .A2(n19868), .B1(n13531), .B2(n13831), .ZN(
        n13836) );
  OAI22_X1 U17034 ( .A1(n13834), .A2(n19636), .B1(n19938), .B2(n13833), .ZN(
        n13835) );
  NOR2_X1 U17035 ( .A1(n13836), .A2(n13835), .ZN(n13857) );
  OAI22_X1 U17036 ( .A1(n13838), .A2(n13784), .B1(n13805), .B2(n13837), .ZN(
        n13842) );
  OAI22_X1 U17037 ( .A1(n13840), .A2(n19786), .B1(n19977), .B2(n13839), .ZN(
        n13841) );
  NOR2_X1 U17038 ( .A1(n13842), .A2(n13841), .ZN(n13856) );
  INV_X1 U17039 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13843) );
  OAI22_X1 U17040 ( .A1(n13844), .A2(n19516), .B1(n20011), .B2(n13843), .ZN(
        n13847) );
  INV_X1 U17041 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13845) );
  OAI22_X1 U17042 ( .A1(n13845), .A2(n19697), .B1(n19760), .B2(n11029), .ZN(
        n13846) );
  NOR2_X1 U17043 ( .A1(n13847), .A2(n13846), .ZN(n13855) );
  INV_X1 U17044 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13848) );
  OAI22_X1 U17045 ( .A1(n19572), .A2(n13849), .B1(n19726), .B2(n13848), .ZN(
        n13853) );
  INV_X1 U17046 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13850) );
  OAI22_X1 U17047 ( .A1(n19899), .A2(n13851), .B1(n13787), .B2(n13850), .ZN(
        n13852) );
  NOR2_X1 U17048 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  NAND4_X1 U17049 ( .A1(n13857), .A2(n13856), .A3(n13855), .A4(n13854), .ZN(
        n13861) );
  INV_X1 U17050 ( .A(n13858), .ZN(n13859) );
  NAND2_X1 U17051 ( .A1(n13859), .A2(n9839), .ZN(n13860) );
  INV_X1 U17052 ( .A(n13862), .ZN(n13876) );
  NAND2_X1 U17053 ( .A1(n13863), .A2(n13876), .ZN(n13864) );
  NOR2_X1 U17054 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  OR2_X1 U17055 ( .A1(n13926), .A2(n13867), .ZN(n19286) );
  XNOR2_X1 U17056 ( .A(n13923), .B(n13890), .ZN(n13921) );
  XNOR2_X1 U17057 ( .A(n13922), .B(n13921), .ZN(n13901) );
  INV_X1 U17058 ( .A(n13868), .ZN(n13913) );
  NAND2_X1 U17059 ( .A1(n13913), .A2(n16444), .ZN(n13880) );
  NAND2_X1 U17060 ( .A1(n13872), .A2(n16480), .ZN(n13870) );
  NAND2_X1 U17061 ( .A1(n13871), .A2(n13870), .ZN(n13875) );
  INV_X1 U17062 ( .A(n13872), .ZN(n13873) );
  NAND2_X1 U17063 ( .A1(n13873), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13874) );
  NAND2_X1 U17064 ( .A1(n13869), .A2(n16497), .ZN(n16443) );
  INV_X1 U17065 ( .A(n16444), .ZN(n13877) );
  NAND2_X1 U17066 ( .A1(n13877), .A2(n13876), .ZN(n13879) );
  OAI21_X1 U17067 ( .B1(n13881), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13916), .ZN(n13882) );
  INV_X1 U17068 ( .A(n13882), .ZN(n13899) );
  OAI22_X1 U17069 ( .A1(n12535), .A2(n19294), .B1(n19503), .B2(n19283), .ZN(
        n13885) );
  INV_X1 U17070 ( .A(n19289), .ZN(n13896) );
  INV_X1 U17071 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13883) );
  OAI22_X1 U17072 ( .A1(n16438), .A2(n13896), .B1(n19514), .B2(n13883), .ZN(
        n13884) );
  AOI211_X1 U17073 ( .C1(n13899), .C2(n16449), .A(n13885), .B(n13884), .ZN(
        n13886) );
  OAI21_X1 U17074 ( .B1(n19493), .B2(n13901), .A(n13886), .ZN(P2_U3008) );
  NOR3_X1 U17075 ( .A1(n16480), .A2(n13547), .A3(n16497), .ZN(n13887) );
  NAND2_X1 U17076 ( .A1(n13887), .A2(n14274), .ZN(n13891) );
  NAND2_X1 U17077 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13887), .ZN(
        n14262) );
  AOI21_X1 U17078 ( .B1(n14262), .B2(n15517), .A(n13888), .ZN(n16471) );
  NAND2_X1 U17079 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19310), .ZN(n13889) );
  OAI221_X1 U17080 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n13891), .C1(
        n13890), .C2(n16471), .A(n13889), .ZN(n13898) );
  NOR2_X1 U17081 ( .A1(n13893), .A2(n13892), .ZN(n13894) );
  OR2_X1 U17082 ( .A1(n13895), .A2(n13894), .ZN(n19288) );
  OAI22_X1 U17083 ( .A1(n16469), .A2(n19288), .B1(n15640), .B2(n13896), .ZN(
        n13897) );
  AOI211_X1 U17084 ( .C1(n13899), .C2(n16493), .A(n13898), .B(n13897), .ZN(
        n13900) );
  OAI21_X1 U17085 ( .B1(n16477), .B2(n13901), .A(n13900), .ZN(P2_U3040) );
  OR2_X1 U17086 ( .A1(n13904), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13902) );
  NAND2_X1 U17087 ( .A1(n13904), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13905) );
  INV_X4 U17088 ( .A(n14334), .ZN(n16081) );
  XNOR2_X1 U17089 ( .A(n16081), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13906) );
  XNOR2_X1 U17090 ( .A(n14322), .B(n13906), .ZN(n16208) );
  AOI22_X1 U17091 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13907) );
  OAI21_X1 U17092 ( .B1(n20374), .B2(n13908), .A(n13907), .ZN(n13909) );
  AOI21_X1 U17093 ( .B1(n20265), .B2(n14411), .A(n13909), .ZN(n13910) );
  OAI21_X1 U17094 ( .B1(n16208), .B2(n20242), .A(n13910), .ZN(P1_U2990) );
  INV_X1 U17095 ( .A(n13911), .ZN(n13912) );
  NAND2_X1 U17096 ( .A1(n13912), .A2(n16444), .ZN(n13914) );
  NAND2_X1 U17097 ( .A1(n13914), .A2(n13913), .ZN(n13915) );
  XNOR2_X1 U17098 ( .A(n13917), .B(n14183), .ZN(n13919) );
  INV_X1 U17099 ( .A(n13919), .ZN(n13918) );
  NAND2_X1 U17100 ( .A1(n13918), .A2(n13927), .ZN(n14217) );
  OR2_X1 U17101 ( .A1(n10184), .A2(n14218), .ZN(n13920) );
  XNOR2_X1 U17102 ( .A(n14219), .B(n13920), .ZN(n16434) );
  INV_X1 U17103 ( .A(n16434), .ZN(n13939) );
  NAND2_X1 U17104 ( .A1(n13922), .A2(n13921), .ZN(n14100) );
  NAND2_X1 U17105 ( .A1(n13923), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14098) );
  NAND2_X1 U17106 ( .A1(n14100), .A2(n14098), .ZN(n16425) );
  INV_X1 U17107 ( .A(n13924), .ZN(n13925) );
  XNOR2_X1 U17108 ( .A(n13926), .B(n13925), .ZN(n19271) );
  NAND2_X1 U17109 ( .A1(n19271), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16422) );
  INV_X1 U17110 ( .A(n19271), .ZN(n13928) );
  NAND2_X1 U17111 ( .A1(n13928), .A2(n13927), .ZN(n16424) );
  NAND2_X1 U17112 ( .A1(n16422), .A2(n16424), .ZN(n13929) );
  XNOR2_X1 U17113 ( .A(n16425), .B(n13929), .ZN(n16435) );
  INV_X1 U17114 ( .A(n14262), .ZN(n13930) );
  NAND2_X1 U17115 ( .A1(n13930), .A2(n14274), .ZN(n16466) );
  NAND2_X1 U17116 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19310), .ZN(n13931) );
  OAI221_X1 U17117 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16466), .C1(
        n13927), .C2(n16471), .A(n13931), .ZN(n13937) );
  AOI21_X1 U17118 ( .B1(n13934), .B2(n13933), .A(n13932), .ZN(n19392) );
  INV_X1 U17119 ( .A(n19392), .ZN(n13935) );
  OAI22_X1 U17120 ( .A1(n16469), .A2(n13935), .B1(n15640), .B2(n19281), .ZN(
        n13936) );
  AOI211_X1 U17121 ( .C1(n16435), .C2(n16490), .A(n13937), .B(n13936), .ZN(
        n13938) );
  OAI21_X1 U17122 ( .B1(n13939), .B2(n16457), .A(n13938), .ZN(P2_U3039) );
  INV_X1 U17123 ( .A(n13940), .ZN(n13942) );
  OAI21_X1 U17124 ( .B1(n10404), .B2(n13942), .A(n15108), .ZN(n13987) );
  NOR2_X1 U17125 ( .A1(n13943), .A2(n20217), .ZN(n13944) );
  NAND2_X1 U17126 ( .A1(n13945), .A2(n13944), .ZN(n13946) );
  NAND2_X1 U17127 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  NAND2_X1 U17128 ( .A1(n14399), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17129 ( .A1(n14398), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13950) );
  INV_X1 U17130 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13956) );
  AOI22_X1 U17131 ( .A1(n14398), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13955) );
  INV_X1 U17132 ( .A(n13952), .ZN(n13953) );
  NAND2_X1 U17133 ( .A1(n13966), .A2(n13953), .ZN(n13954) );
  OAI211_X1 U17134 ( .C1(n12473), .C2(n13956), .A(n13955), .B(n13954), .ZN(
        n15606) );
  NOR2_X1 U17135 ( .A1(n12517), .A2(n15590), .ZN(n13961) );
  INV_X1 U17136 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13957) );
  OAI22_X1 U17137 ( .A1(n13959), .A2(n13958), .B1(n13957), .B2(n12473), .ZN(
        n13960) );
  AOI211_X1 U17138 ( .C1(P2_EAX_REG_13__SCAN_IN), .C2(n14398), .A(n13961), .B(
        n13960), .ZN(n15587) );
  NOR2_X4 U17139 ( .A1(n15607), .A2(n15587), .ZN(n15586) );
  INV_X1 U17140 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U17141 ( .A1(n12470), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13964) );
  NAND2_X1 U17142 ( .A1(n13966), .A2(n13962), .ZN(n13963) );
  OAI211_X1 U17143 ( .C1(n12473), .C2(n13965), .A(n13964), .B(n13963), .ZN(
        n15564) );
  NAND2_X2 U17144 ( .A1(n15586), .A2(n15564), .ZN(n15565) );
  AOI22_X1 U17145 ( .A1(n14399), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n13966), 
        .B2(n15082), .ZN(n13968) );
  AOI22_X1 U17146 ( .A1(n14398), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13967) );
  INV_X1 U17147 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20119) );
  AOI22_X1 U17148 ( .A1(n14398), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U17149 ( .B1(n12473), .B2(n20119), .A(n13969), .ZN(n14000) );
  XNOR2_X1 U17150 ( .A(n14018), .B(n14019), .ZN(n19184) );
  NOR2_X1 U17151 ( .A1(n19554), .A2(n19565), .ZN(n13970) );
  AOI22_X1 U17152 ( .A1(n19360), .A2(BUF2_REG_17__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17153 ( .A1(n19367), .A2(n13972), .B1(n19427), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13973) );
  OAI211_X1 U17154 ( .C1(n19365), .C2(n19184), .A(n13974), .B(n13973), .ZN(
        n13975) );
  INV_X1 U17155 ( .A(n13975), .ZN(n13976) );
  OAI21_X1 U17156 ( .B1(n13987), .B2(n19366), .A(n13976), .ZN(P2_U2902) );
  OR2_X1 U17157 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  NAND2_X1 U17158 ( .A1(n13977), .A2(n13980), .ZN(n14037) );
  XNOR2_X1 U17159 ( .A(n14037), .B(n14035), .ZN(n16100) );
  INV_X1 U17160 ( .A(n16100), .ZN(n14016) );
  INV_X1 U17161 ( .A(DATAI_11_), .ZN(n21195) );
  MUX2_X1 U17162 ( .A(n21195), .B(n16662), .S(n20415), .Z(n14622) );
  INV_X1 U17163 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13981) );
  OAI222_X1 U17164 ( .A1(n14016), .A2(n14672), .B1(n14622), .B2(n14676), .C1(
        n13981), .C2(n14674), .ZN(P1_U2893) );
  NAND2_X1 U17165 ( .A1(n9831), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13986) );
  NOR2_X1 U17166 ( .A1(n9929), .A2(n13983), .ZN(n13984) );
  NOR2_X1 U17167 ( .A1(n13982), .A2(n13984), .ZN(n19177) );
  NAND2_X1 U17168 ( .A1(n19177), .A2(n15104), .ZN(n13985) );
  OAI211_X1 U17169 ( .C1(n13987), .C2(n15106), .A(n13986), .B(n13985), .ZN(
        P2_U2870) );
  NOR2_X1 U17170 ( .A1(n13997), .A2(n13988), .ZN(n15107) );
  NOR2_X1 U17171 ( .A1(n13997), .A2(n13989), .ZN(n15098) );
  INV_X1 U17172 ( .A(n15098), .ZN(n13990) );
  OAI21_X1 U17173 ( .B1(n15107), .B2(n13991), .A(n13990), .ZN(n14034) );
  NAND2_X1 U17174 ( .A1(n9831), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13996) );
  NOR2_X1 U17175 ( .A1(n15112), .A2(n13993), .ZN(n13994) );
  NOR2_X1 U17176 ( .A1(n13992), .A2(n13994), .ZN(n19159) );
  NAND2_X1 U17177 ( .A1(n19159), .A2(n15104), .ZN(n13995) );
  OAI211_X1 U17178 ( .C1(n14034), .C2(n15106), .A(n13996), .B(n13995), .ZN(
        P2_U2868) );
  AOI21_X1 U17179 ( .B1(n13998), .B2(n13997), .A(n10404), .ZN(n14007) );
  OR2_X1 U17180 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  NAND2_X1 U17181 ( .A1(n14001), .A2(n14019), .ZN(n19196) );
  AOI22_X1 U17182 ( .A1(n19360), .A2(BUF2_REG_16__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U17183 ( .A1(n19367), .A2(n14002), .B1(n19427), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14003) );
  OAI211_X1 U17184 ( .C1(n19365), .C2(n19196), .A(n14004), .B(n14003), .ZN(
        n14005) );
  AOI21_X1 U17185 ( .B1(n14007), .B2(n19429), .A(n14005), .ZN(n14006) );
  INV_X1 U17186 ( .A(n14006), .ZN(P2_U2903) );
  NAND2_X1 U17187 ( .A1(n14007), .A2(n15110), .ZN(n14012) );
  NOR2_X1 U17188 ( .A1(n14009), .A2(n14008), .ZN(n14010) );
  NOR2_X1 U17189 ( .A1(n9929), .A2(n14010), .ZN(n19193) );
  NAND2_X1 U17190 ( .A1(n19193), .A2(n15104), .ZN(n14011) );
  OAI211_X1 U17191 ( .C1(n15104), .C2(n14145), .A(n14012), .B(n14011), .ZN(
        P2_U2871) );
  OR2_X1 U17192 ( .A1(n14014), .A2(n14013), .ZN(n14015) );
  NAND2_X1 U17193 ( .A1(n9935), .A2(n14015), .ZN(n16188) );
  INV_X1 U17194 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14017) );
  OAI222_X1 U17195 ( .A1(n16188), .A2(n14613), .B1(n14612), .B2(n14017), .C1(
        n14016), .C2(n14610), .ZN(P1_U2861) );
  INV_X1 U17196 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U17197 ( .A1(n12470), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14020) );
  OAI21_X1 U17198 ( .B1(n12473), .B2(n20123), .A(n14020), .ZN(n15208) );
  INV_X1 U17199 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17200 ( .A1(n12470), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14021) );
  OAI21_X1 U17201 ( .B1(n12473), .B2(n14022), .A(n14021), .ZN(n14024) );
  NOR2_X1 U17202 ( .A1(n14023), .A2(n14024), .ZN(n14025) );
  NOR2_X1 U17203 ( .A1(n15199), .A2(n14025), .ZN(n19158) );
  NAND2_X1 U17204 ( .A1(n19367), .A2(n14026), .ZN(n14027) );
  OAI21_X1 U17205 ( .B1(n19391), .B2(n14028), .A(n14027), .ZN(n14032) );
  INV_X1 U17206 ( .A(n19360), .ZN(n15193) );
  INV_X1 U17207 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14030) );
  INV_X1 U17208 ( .A(n19362), .ZN(n15191) );
  INV_X1 U17209 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14029) );
  OAI22_X1 U17210 ( .A1(n15193), .A2(n14030), .B1(n15191), .B2(n14029), .ZN(
        n14031) );
  AOI211_X1 U17211 ( .C1(n19428), .C2(n19158), .A(n14032), .B(n14031), .ZN(
        n14033) );
  OAI21_X1 U17212 ( .B1(n14034), .B2(n19366), .A(n14033), .ZN(P2_U2900) );
  INV_X1 U17213 ( .A(n14035), .ZN(n14036) );
  OAI21_X1 U17214 ( .B1(n14037), .B2(n14036), .A(n13977), .ZN(n14050) );
  AND2_X1 U17215 ( .A1(n14050), .A2(n14049), .ZN(n14052) );
  OAI21_X1 U17216 ( .B1(n14052), .B2(n14039), .A(n14038), .ZN(n14829) );
  AND2_X1 U17217 ( .A1(n9936), .A2(n14040), .ZN(n14041) );
  NOR2_X1 U17218 ( .A1(n14060), .A2(n14041), .ZN(n16169) );
  AOI22_X1 U17219 ( .A1(n14601), .A2(n16169), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14600), .ZN(n14042) );
  OAI21_X1 U17220 ( .B1(n14829), .B2(n14610), .A(n14042), .ZN(P1_U2859) );
  INV_X1 U17221 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21290) );
  INV_X1 U17222 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21453) );
  NOR2_X1 U17223 ( .A1(n21290), .A2(n21453), .ZN(n14057) );
  OAI21_X1 U17224 ( .B1(n14057), .B2(n20318), .A(n16055), .ZN(n16048) );
  INV_X1 U17225 ( .A(n16169), .ZN(n14044) );
  AOI21_X1 U17226 ( .B1(n20264), .B2(n14826), .A(n20306), .ZN(n14043) );
  OAI21_X1 U17227 ( .B1(n20313), .B2(n14044), .A(n14043), .ZN(n14047) );
  NAND3_X1 U17228 ( .A1(n20270), .A2(n16044), .A3(n14057), .ZN(n14056) );
  AOI22_X1 U17229 ( .A1(n20315), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20307), .ZN(n14045) );
  OAI21_X1 U17230 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n14056), .A(n14045), 
        .ZN(n14046) );
  AOI211_X1 U17231 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n16048), .A(n14047), 
        .B(n14046), .ZN(n14048) );
  OAI21_X1 U17232 ( .B1(n14829), .B2(n16051), .A(n14048), .ZN(P1_U2827) );
  NOR2_X1 U17233 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  INV_X1 U17234 ( .A(DATAI_12_), .ZN(n21208) );
  INV_X1 U17235 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16660) );
  MUX2_X1 U17236 ( .A(n21208), .B(n16660), .S(n20415), .Z(n14618) );
  INV_X1 U17237 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14053) );
  OAI222_X1 U17238 ( .A1(n16091), .A2(n14672), .B1(n14618), .B2(n14676), .C1(
        n14053), .C2(n14647), .ZN(P1_U2892) );
  OR2_X1 U17239 ( .A1(n14038), .A2(n14055), .ZN(n14077) );
  INV_X1 U17240 ( .A(n14077), .ZN(n14054) );
  AOI21_X1 U17241 ( .B1(n14055), .B2(n14038), .A(n14054), .ZN(n14811) );
  INV_X1 U17242 ( .A(n14811), .ZN(n14073) );
  INV_X1 U17243 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21289) );
  INV_X1 U17244 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21350) );
  OAI21_X1 U17245 ( .B1(n21289), .B2(n14056), .A(n21350), .ZN(n14066) );
  NAND4_X1 U17246 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(n16044), .A4(n14057), .ZN(n14555) );
  INV_X1 U17247 ( .A(n14555), .ZN(n14058) );
  OAI21_X1 U17248 ( .B1(n20318), .B2(n14058), .A(n20277), .ZN(n16036) );
  NOR2_X1 U17249 ( .A1(n14060), .A2(n14059), .ZN(n14061) );
  OR2_X1 U17250 ( .A1(n14607), .A2(n14061), .ZN(n14962) );
  AOI21_X1 U17251 ( .B1(n20307), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20306), .ZN(n14062) );
  OAI21_X1 U17252 ( .B1(n20324), .B2(n14809), .A(n14062), .ZN(n14063) );
  AOI21_X1 U17253 ( .B1(n20315), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14063), .ZN(
        n14064) );
  OAI21_X1 U17254 ( .B1(n20313), .B2(n14962), .A(n14064), .ZN(n14065) );
  AOI21_X1 U17255 ( .B1(n14066), .B2(n16036), .A(n14065), .ZN(n14067) );
  OAI21_X1 U17256 ( .B1(n14073), .B2(n16051), .A(n14067), .ZN(P1_U2826) );
  INV_X1 U17257 ( .A(n14962), .ZN(n14068) );
  AOI22_X1 U17258 ( .A1(n14068), .A2(n14601), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14600), .ZN(n14069) );
  OAI21_X1 U17259 ( .B1(n14073), .B2(n14610), .A(n14069), .ZN(P1_U2858) );
  NAND2_X1 U17260 ( .A1(n9935), .A2(n14070), .ZN(n14071) );
  NAND2_X1 U17261 ( .A1(n9936), .A2(n14071), .ZN(n16182) );
  INV_X1 U17262 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21482) );
  OAI222_X1 U17263 ( .A1(n16182), .A2(n14613), .B1(n14612), .B2(n21482), .C1(
        n16091), .C2(n14610), .ZN(P1_U2860) );
  INV_X1 U17264 ( .A(DATAI_14_), .ZN(n21253) );
  INV_X1 U17265 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16656) );
  MUX2_X1 U17266 ( .A(n21253), .B(n16656), .S(n20415), .Z(n14387) );
  INV_X1 U17267 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14072) );
  OAI222_X1 U17268 ( .A1(n14073), .A2(n14672), .B1(n14387), .B2(n14676), .C1(
        n14072), .C2(n14674), .ZN(P1_U2890) );
  INV_X1 U17269 ( .A(n14074), .ZN(n14075) );
  INV_X1 U17270 ( .A(n14075), .ZN(n14076) );
  AOI21_X1 U17271 ( .B1(n14078), .B2(n14077), .A(n14076), .ZN(n16085) );
  INV_X1 U17272 ( .A(n16085), .ZN(n14611) );
  OAI222_X1 U17273 ( .A1(n14672), .A2(n14611), .B1(n14676), .B2(n14080), .C1(
        n14647), .C2(n14079), .ZN(P1_U2889) );
  XOR2_X1 U17274 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14093), .Z(n14086)
         );
  OAI21_X1 U17275 ( .B1(n14083), .B2(n14082), .A(n14081), .ZN(n19306) );
  MUX2_X1 U17276 ( .A(n14084), .B(n19306), .S(n15104), .Z(n14085) );
  OAI21_X1 U17277 ( .B1(n14086), .B2(n15106), .A(n14085), .ZN(P2_U2882) );
  INV_X1 U17278 ( .A(n14087), .ZN(n14088) );
  NAND2_X1 U17279 ( .A1(n14089), .A2(n14088), .ZN(n14090) );
  OR2_X1 U17280 ( .A1(n14091), .A2(n14090), .ZN(n14092) );
  NAND2_X1 U17281 ( .A1(n14093), .A2(n14092), .ZN(n19405) );
  MUX2_X1 U17282 ( .A(n14094), .B(n19311), .S(n15104), .Z(n14095) );
  OAI21_X1 U17283 ( .B1(n19405), .B2(n15106), .A(n14095), .ZN(P2_U2883) );
  XNOR2_X1 U17284 ( .A(n14096), .B(n9952), .ZN(n19261) );
  AND2_X1 U17285 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14221) );
  NAND2_X1 U17286 ( .A1(n19261), .A2(n14221), .ZN(n16426) );
  AND2_X1 U17287 ( .A1(n16426), .A2(n16422), .ZN(n14097) );
  AND2_X1 U17288 ( .A1(n14098), .A2(n14097), .ZN(n14099) );
  NAND2_X1 U17289 ( .A1(n14100), .A2(n14099), .ZN(n14103) );
  NAND2_X1 U17290 ( .A1(n19261), .A2(n14183), .ZN(n14101) );
  NAND2_X1 U17291 ( .A1(n14101), .A2(n16470), .ZN(n16427) );
  AND2_X1 U17292 ( .A1(n16427), .A2(n16424), .ZN(n14102) );
  NAND2_X1 U17293 ( .A1(n19547), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14104) );
  XNOR2_X1 U17294 ( .A(n14105), .B(n14104), .ZN(n19250) );
  NAND2_X1 U17295 ( .A1(n19250), .A2(n14183), .ZN(n14116) );
  NAND2_X1 U17296 ( .A1(n19547), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14106) );
  OAI21_X1 U17297 ( .B1(n14107), .B2(n14106), .A(n14194), .ZN(n14108) );
  OR2_X1 U17298 ( .A1(n14109), .A2(n14108), .ZN(n19241) );
  OAI21_X1 U17299 ( .B1(n19241), .B2(n14110), .A(n15622), .ZN(n15617) );
  AOI21_X1 U17300 ( .B1(n14118), .B2(n14183), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16398) );
  NAND2_X1 U17301 ( .A1(n19547), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14111) );
  NAND3_X1 U17302 ( .A1(n14204), .A2(n9879), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n14113) );
  NAND2_X1 U17303 ( .A1(n14124), .A2(n14113), .ZN(n19231) );
  OAI21_X1 U17304 ( .B1(n19231), .B2(n14110), .A(n15589), .ZN(n15599) );
  NOR3_X1 U17305 ( .A1(n19231), .A2(n14110), .A3(n15589), .ZN(n15598) );
  INV_X1 U17306 ( .A(n19241), .ZN(n14115) );
  AND2_X1 U17307 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14114) );
  NAND2_X1 U17308 ( .A1(n14115), .A2(n14114), .ZN(n15616) );
  INV_X1 U17309 ( .A(n14116), .ZN(n14117) );
  NAND2_X1 U17310 ( .A1(n14117), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15615) );
  NAND2_X1 U17311 ( .A1(n15616), .A2(n15615), .ZN(n16394) );
  INV_X1 U17312 ( .A(n14118), .ZN(n14120) );
  NAND2_X1 U17313 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14119) );
  NOR2_X1 U17314 ( .A1(n14120), .A2(n14119), .ZN(n16397) );
  NOR2_X1 U17315 ( .A1(n14208), .A2(n14121), .ZN(n14123) );
  INV_X1 U17316 ( .A(n14123), .ZN(n14122) );
  XNOR2_X1 U17317 ( .A(n14124), .B(n14122), .ZN(n19219) );
  NOR2_X1 U17318 ( .A1(n14172), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15583) );
  NAND2_X1 U17319 ( .A1(n19547), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U17320 ( .A1(n14161), .A2(n14162), .ZN(n14151) );
  NOR2_X1 U17321 ( .A1(n14208), .A2(n14125), .ZN(n14150) );
  OR2_X2 U17322 ( .A1(n14151), .A2(n14150), .ZN(n14153) );
  NOR2_X1 U17323 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n14126) );
  AND2_X1 U17324 ( .A1(n11175), .A2(n14138), .ZN(n14127) );
  NOR2_X1 U17325 ( .A1(n14208), .A2(n14127), .ZN(n14128) );
  NOR2_X1 U17326 ( .A1(n14208), .A2(n14130), .ZN(n14131) );
  INV_X1 U17327 ( .A(n14194), .ZN(n14146) );
  AOI21_X1 U17328 ( .B1(n14132), .B2(n14131), .A(n14146), .ZN(n14133) );
  AND2_X1 U17329 ( .A1(n14133), .A2(n14181), .ZN(n19128) );
  AND2_X1 U17330 ( .A1(n19128), .A2(n14183), .ZN(n14166) );
  NOR2_X1 U17331 ( .A1(n14166), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15306) );
  NAND2_X1 U17332 ( .A1(n14204), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14134) );
  INV_X1 U17333 ( .A(n14158), .ZN(n14135) );
  MUX2_X1 U17334 ( .A(n14134), .B(n14204), .S(n14135), .Z(n14136) );
  NAND2_X1 U17335 ( .A1(n14135), .A2(n11175), .ZN(n14140) );
  NAND2_X1 U17336 ( .A1(n14136), .A2(n14140), .ZN(n19163) );
  OAI21_X1 U17337 ( .B1(n19163), .B2(n14110), .A(n14137), .ZN(n15337) );
  NOR2_X1 U17338 ( .A1(n14208), .A2(n14138), .ZN(n14139) );
  NAND2_X1 U17339 ( .A1(n14140), .A2(n14139), .ZN(n14142) );
  INV_X1 U17340 ( .A(n14141), .ZN(n14144) );
  NAND2_X1 U17341 ( .A1(n14142), .A2(n14144), .ZN(n19156) );
  NAND2_X1 U17342 ( .A1(n14174), .A2(n15478), .ZN(n15326) );
  NAND2_X1 U17343 ( .A1(n15337), .A2(n15326), .ZN(n15299) );
  NAND2_X1 U17344 ( .A1(n19547), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14143) );
  XNOR2_X1 U17345 ( .A(n14144), .B(n14143), .ZN(n19139) );
  AOI21_X1 U17346 ( .B1(n19139), .B2(n14183), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15302) );
  OR2_X1 U17347 ( .A1(n14153), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14157) );
  NOR2_X1 U17348 ( .A1(n14208), .A2(n14145), .ZN(n14147) );
  AOI21_X1 U17349 ( .B1(n14153), .B2(n14147), .A(n14146), .ZN(n14148) );
  NAND2_X1 U17350 ( .A1(n19185), .A2(n14183), .ZN(n14149) );
  XNOR2_X1 U17351 ( .A(n14149), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15358) );
  NAND2_X1 U17352 ( .A1(n14151), .A2(n14150), .ZN(n14152) );
  NAND2_X1 U17353 ( .A1(n14153), .A2(n14152), .ZN(n19200) );
  OR2_X1 U17354 ( .A1(n19200), .A2(n14110), .ZN(n14154) );
  NAND2_X1 U17355 ( .A1(n14154), .A2(n15549), .ZN(n15539) );
  NOR2_X1 U17356 ( .A1(n14208), .A2(n14155), .ZN(n14156) );
  NAND2_X1 U17357 ( .A1(n14157), .A2(n14156), .ZN(n14159) );
  NAND2_X1 U17358 ( .A1(n14159), .A2(n14158), .ZN(n19174) );
  OAI21_X1 U17359 ( .B1(n19174), .B2(n14110), .A(n14160), .ZN(n15298) );
  INV_X1 U17360 ( .A(n14161), .ZN(n14163) );
  XNOR2_X1 U17361 ( .A(n14163), .B(n14162), .ZN(n19208) );
  NAND2_X1 U17362 ( .A1(n19208), .A2(n14183), .ZN(n14164) );
  NAND2_X1 U17363 ( .A1(n14164), .A2(n15563), .ZN(n15557) );
  NAND4_X1 U17364 ( .A1(n15358), .A2(n15539), .A3(n15298), .A4(n15557), .ZN(
        n14165) );
  NOR4_X1 U17365 ( .A1(n15306), .A2(n15299), .A3(n15302), .A4(n14165), .ZN(
        n14179) );
  NAND2_X1 U17366 ( .A1(n14166), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15304) );
  INV_X1 U17367 ( .A(n19174), .ZN(n14168) );
  AND2_X1 U17368 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14167) );
  NAND2_X1 U17369 ( .A1(n14168), .A2(n14167), .ZN(n15297) );
  NAND2_X1 U17370 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14169) );
  OR2_X1 U17371 ( .A1(n19200), .A2(n14169), .ZN(n15538) );
  AND2_X1 U17372 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14170) );
  NAND2_X1 U17373 ( .A1(n19208), .A2(n14170), .ZN(n15556) );
  AND2_X1 U17374 ( .A1(n15538), .A2(n15556), .ZN(n15295) );
  AND2_X1 U17375 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14171) );
  NAND2_X1 U17376 ( .A1(n19185), .A2(n14171), .ZN(n15296) );
  INV_X1 U17377 ( .A(n14172), .ZN(n14173) );
  AND4_X1 U17378 ( .A1(n15297), .A2(n15295), .A3(n15296), .A4(n15581), .ZN(
        n14177) );
  OR2_X1 U17379 ( .A1(n14174), .A2(n15478), .ZN(n15327) );
  NAND2_X1 U17380 ( .A1(n14183), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14175) );
  OR2_X1 U17381 ( .A1(n19163), .A2(n14175), .ZN(n15336) );
  AND2_X1 U17382 ( .A1(n15327), .A2(n15336), .ZN(n15300) );
  INV_X1 U17383 ( .A(n19139), .ZN(n14176) );
  NAND4_X1 U17384 ( .A1(n15304), .A2(n14177), .A3(n15300), .A4(n15303), .ZN(
        n14178) );
  NOR2_X1 U17385 ( .A1(n14208), .A2(n14180), .ZN(n14182) );
  AOI21_X1 U17386 ( .B1(n14182), .B2(n14181), .A(n14185), .ZN(n15930) );
  AOI21_X1 U17387 ( .B1(n15930), .B2(n14183), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15448) );
  NAND3_X1 U17388 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14183), .ZN(n15449) );
  NAND2_X1 U17389 ( .A1(n19547), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14184) );
  XOR2_X1 U17390 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n14186), .Z(
        n15286) );
  NAND3_X1 U17391 ( .A1(n14187), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n19547), 
        .ZN(n14188) );
  NAND3_X1 U17392 ( .A1(n14189), .A2(n14194), .A3(n14188), .ZN(n16333) );
  NOR2_X1 U17393 ( .A1(n16333), .A2(n14110), .ZN(n15272) );
  NAND3_X1 U17394 ( .A1(n14189), .A2(P2_EBX_REG_25__SCAN_IN), .A3(n19547), 
        .ZN(n14190) );
  NAND2_X1 U17395 ( .A1(n14190), .A2(n14194), .ZN(n14191) );
  NOR2_X1 U17396 ( .A1(n14193), .A2(n14191), .ZN(n16322) );
  NAND2_X1 U17397 ( .A1(n16322), .A2(n12457), .ZN(n14200) );
  NAND2_X1 U17398 ( .A1(n19547), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14192) );
  OR2_X1 U17399 ( .A1(n14193), .A2(n14192), .ZN(n14195) );
  NAND2_X1 U17400 ( .A1(n16310), .A2(n14193), .ZN(n14243) );
  AND2_X1 U17401 ( .A1(n14195), .A2(n14213), .ZN(n14196) );
  INV_X1 U17402 ( .A(n14196), .ZN(n16311) );
  NOR2_X1 U17403 ( .A1(n16311), .A2(n14110), .ZN(n14197) );
  OAI21_X1 U17404 ( .B1(n14197), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14201), .ZN(n15243) );
  INV_X1 U17405 ( .A(n14213), .ZN(n14198) );
  NAND2_X1 U17406 ( .A1(n19547), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U17407 ( .A1(n14204), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14202) );
  XNOR2_X1 U17408 ( .A(n14246), .B(n14202), .ZN(n16289) );
  NAND2_X1 U17409 ( .A1(n16289), .A2(n12457), .ZN(n14250) );
  NOR2_X1 U17410 ( .A1(n14200), .A2(n14199), .ZN(n15264) );
  INV_X1 U17411 ( .A(n14202), .ZN(n14203) );
  NAND2_X1 U17412 ( .A1(n14204), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14205) );
  XNOR2_X1 U17413 ( .A(n14206), .B(n14205), .ZN(n16279) );
  OAI21_X1 U17414 ( .B1(n16279), .B2(n14110), .A(n15382), .ZN(n15225) );
  NOR3_X1 U17415 ( .A1(n16279), .A2(n14110), .A3(n15382), .ZN(n15224) );
  INV_X1 U17416 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n16278) );
  OAI21_X1 U17417 ( .B1(n16278), .B2(n14208), .A(n14206), .ZN(n14211) );
  NOR2_X1 U17418 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  XNOR2_X1 U17419 ( .A(n14211), .B(n14209), .ZN(n16266) );
  NOR2_X1 U17420 ( .A1(n16266), .A2(n14110), .ZN(n14210) );
  NAND2_X1 U17421 ( .A1(n14210), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15216) );
  NOR2_X1 U17422 ( .A1(n14211), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14212) );
  MUX2_X1 U17423 ( .A(n14213), .B(n14212), .S(n19547), .Z(n16258) );
  NAND2_X1 U17424 ( .A1(n16258), .A2(n12457), .ZN(n14214) );
  XNOR2_X1 U17425 ( .A(n14214), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14215) );
  XNOR2_X1 U17426 ( .A(n14216), .B(n14215), .ZN(n14406) );
  XNOR2_X1 U17427 ( .A(n14220), .B(n16470), .ZN(n16421) );
  INV_X1 U17428 ( .A(n14221), .ZN(n14222) );
  NAND3_X1 U17429 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U17430 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16460) );
  NOR2_X1 U17431 ( .A1(n15643), .A2(n16460), .ZN(n15562) );
  NAND3_X1 U17432 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n15562), .ZN(n15569) );
  NOR2_X1 U17433 ( .A1(n15563), .A2(n15569), .ZN(n15499) );
  NAND2_X1 U17434 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15499), .ZN(
        n14224) );
  NOR2_X1 U17435 ( .A1(n15500), .A2(n14224), .ZN(n14275) );
  AND2_X2 U17436 ( .A1(n15452), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15454) );
  NAND2_X1 U17437 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15401) );
  XOR2_X1 U17438 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14225), .Z(
        n14404) );
  AOI22_X1 U17439 ( .A1(n14227), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14230) );
  NAND2_X1 U17440 ( .A1(n14228), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14229) );
  OAI211_X1 U17441 ( .C1(n14232), .C2(n14231), .A(n14230), .B(n14229), .ZN(
        n14233) );
  NAND2_X1 U17442 ( .A1(n16263), .A2(n19510), .ZN(n14236) );
  INV_X1 U17443 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20150) );
  NOR2_X1 U17444 ( .A1(n19294), .A2(n20150), .ZN(n14402) );
  AOI21_X1 U17445 ( .B1(n19490), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14402), .ZN(n14235) );
  OAI211_X1 U17446 ( .C1(n19503), .C2(n14237), .A(n14236), .B(n14235), .ZN(
        n14238) );
  AOI21_X1 U17447 ( .B1(n14404), .B2(n16449), .A(n14238), .ZN(n14239) );
  OAI21_X1 U17448 ( .B1(n14406), .B2(n19493), .A(n14239), .ZN(P2_U2983) );
  INV_X1 U17449 ( .A(n14242), .ZN(n14244) );
  NAND2_X1 U17450 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  NAND2_X1 U17451 ( .A1(n14246), .A2(n14245), .ZN(n16300) );
  NOR2_X1 U17452 ( .A1(n16300), .A2(n14110), .ZN(n14248) );
  XOR2_X1 U17453 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14250), .Z(
        n14251) );
  XNOR2_X1 U17454 ( .A(n14252), .B(n14251), .ZN(n14300) );
  AOI21_X1 U17455 ( .B1(n15381), .B2(n15238), .A(n9880), .ZN(n14297) );
  AND2_X1 U17456 ( .A1(n15236), .A2(n14253), .ZN(n14254) );
  OR2_X1 U17457 ( .A1(n14254), .A2(n15228), .ZN(n16294) );
  NOR2_X1 U17458 ( .A1(n14255), .A2(n14256), .ZN(n14257) );
  INV_X1 U17459 ( .A(n15031), .ZN(n16291) );
  NAND2_X1 U17460 ( .A1(n16291), .A2(n19510), .ZN(n14259) );
  INV_X1 U17461 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20141) );
  NOR2_X1 U17462 ( .A1(n19294), .A2(n20141), .ZN(n14293) );
  AOI21_X1 U17463 ( .B1(n19490), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14293), .ZN(n14258) );
  OAI211_X1 U17464 ( .C1(n19503), .C2(n16294), .A(n14259), .B(n14258), .ZN(
        n14260) );
  AOI21_X1 U17465 ( .B1(n14297), .B2(n16449), .A(n14260), .ZN(n14261) );
  OAI21_X1 U17466 ( .B1(n14300), .B2(n19493), .A(n14261), .ZN(P2_U2986) );
  NOR3_X1 U17467 ( .A1(n13927), .A2(n16470), .A3(n14262), .ZN(n14273) );
  OAI221_X1 U17468 ( .B1(n15620), .B2(n14273), .C1(n15620), .C2(n14264), .A(
        n14263), .ZN(n15561) );
  INV_X1 U17469 ( .A(n14275), .ZN(n14265) );
  AND2_X1 U17470 ( .A1(n15517), .A2(n14265), .ZN(n14266) );
  OR2_X1 U17471 ( .A1(n15561), .A2(n14266), .ZN(n15509) );
  NOR2_X1 U17472 ( .A1(n15478), .A2(n15479), .ZN(n15477) );
  INV_X1 U17473 ( .A(n15477), .ZN(n14276) );
  AND2_X1 U17474 ( .A1(n15517), .A2(n14276), .ZN(n14267) );
  NOR2_X1 U17475 ( .A1(n15509), .A2(n14267), .ZN(n15466) );
  NAND2_X1 U17476 ( .A1(n15517), .A2(n15465), .ZN(n14268) );
  AND2_X1 U17477 ( .A1(n15466), .A2(n14268), .ZN(n15455) );
  NOR2_X1 U17478 ( .A1(n15458), .A2(n15437), .ZN(n15436) );
  INV_X1 U17479 ( .A(n15436), .ZN(n14269) );
  NAND2_X1 U17480 ( .A1(n15517), .A2(n14269), .ZN(n14270) );
  NAND2_X1 U17481 ( .A1(n15455), .A2(n14270), .ZN(n15430) );
  AND2_X1 U17482 ( .A1(n15517), .A2(n15278), .ZN(n14271) );
  AND2_X1 U17483 ( .A1(n15517), .A2(n15401), .ZN(n14272) );
  NOR2_X1 U17484 ( .A1(n15419), .A2(n14272), .ZN(n15389) );
  NAND2_X1 U17485 ( .A1(n15568), .A2(n14275), .ZN(n15493) );
  NAND2_X1 U17486 ( .A1(n15436), .A2(n15459), .ZN(n15426) );
  INV_X1 U17487 ( .A(n15379), .ZN(n15369) );
  NAND2_X1 U17488 ( .A1(n15369), .A2(n14392), .ZN(n15393) );
  NAND2_X1 U17489 ( .A1(n15389), .A2(n15393), .ZN(n15385) );
  NOR3_X1 U17490 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n14392), .ZN(n14296) );
  INV_X1 U17491 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U17492 ( .A1(n12470), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14277) );
  OAI21_X1 U17493 ( .B1(n12473), .B2(n20126), .A(n14277), .ZN(n15198) );
  NAND2_X1 U17494 ( .A1(n14399), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14279) );
  AOI22_X1 U17495 ( .A1(n12470), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14278) );
  NOR2_X2 U17496 ( .A1(n15200), .A2(n15186), .ZN(n15176) );
  INV_X1 U17497 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U17498 ( .A1(n12470), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14280) );
  OAI21_X1 U17499 ( .B1(n12473), .B2(n20130), .A(n14280), .ZN(n15177) );
  NAND2_X1 U17500 ( .A1(n14399), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17501 ( .A1(n12470), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U17502 ( .A1(n14282), .A2(n14281), .ZN(n15438) );
  NAND2_X1 U17503 ( .A1(n14399), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U17504 ( .A1(n12470), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14283) );
  AND2_X1 U17505 ( .A1(n14284), .A2(n14283), .ZN(n15167) );
  NAND2_X1 U17506 ( .A1(n14399), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U17507 ( .A1(n12470), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14285) );
  AND2_X1 U17508 ( .A1(n14286), .A2(n14285), .ZN(n15160) );
  INV_X1 U17509 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U17510 ( .A1(n12470), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14287) );
  OAI21_X1 U17511 ( .B1(n12473), .B2(n20137), .A(n14287), .ZN(n15151) );
  NAND2_X1 U17512 ( .A1(n14399), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U17513 ( .A1(n12470), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U17514 ( .A1(n14289), .A2(n14288), .ZN(n15143) );
  AOI22_X1 U17515 ( .A1(n12470), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14290) );
  OAI21_X1 U17516 ( .B1(n12473), .B2(n20141), .A(n14290), .ZN(n14291) );
  OR2_X1 U17517 ( .A1(n15145), .A2(n14291), .ZN(n14292) );
  AOI21_X1 U17518 ( .B1(n16485), .B2(n16290), .A(n14293), .ZN(n14294) );
  OAI21_X1 U17519 ( .B1(n15031), .B2(n15640), .A(n14294), .ZN(n14295) );
  AOI211_X1 U17520 ( .C1(n15385), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14296), .B(n14295), .ZN(n14299) );
  NAND2_X1 U17521 ( .A1(n14297), .A2(n16493), .ZN(n14298) );
  OAI211_X1 U17522 ( .C1(n14300), .C2(n16477), .A(n14299), .B(n14298), .ZN(
        P2_U3018) );
  INV_X1 U17523 ( .A(n14635), .ZN(n14301) );
  NAND2_X1 U17524 ( .A1(n14316), .A2(n14301), .ZN(n14319) );
  NAND2_X1 U17525 ( .A1(n20361), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14302) );
  OAI211_X1 U17526 ( .C1(n13661), .C2(n14320), .A(n14319), .B(n14302), .ZN(
        P1_U2960) );
  INV_X1 U17527 ( .A(n14387), .ZN(n14303) );
  NAND2_X1 U17528 ( .A1(n14316), .A2(n14303), .ZN(n20363) );
  NAND2_X1 U17529 ( .A1(n20361), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14304) );
  OAI211_X1 U17530 ( .C1(n21475), .C2(n14320), .A(n20363), .B(n14304), .ZN(
        P1_U2951) );
  INV_X1 U17531 ( .A(DATAI_13_), .ZN(n21358) );
  INV_X1 U17532 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16658) );
  MUX2_X1 U17533 ( .A(n21358), .B(n16658), .S(n20415), .Z(n14677) );
  INV_X1 U17534 ( .A(n14677), .ZN(n14305) );
  NAND2_X1 U17535 ( .A1(n14316), .A2(n14305), .ZN(n20359) );
  NAND2_X1 U17536 ( .A1(n20361), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14306) );
  OAI211_X1 U17537 ( .C1(n14307), .C2(n14320), .A(n20359), .B(n14306), .ZN(
        P1_U2950) );
  INV_X1 U17538 ( .A(n14618), .ZN(n14308) );
  NAND2_X1 U17539 ( .A1(n14316), .A2(n14308), .ZN(n20357) );
  NAND2_X1 U17540 ( .A1(n20361), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14309) );
  OAI211_X1 U17541 ( .C1(n21459), .C2(n14320), .A(n20357), .B(n14309), .ZN(
        P1_U2949) );
  INV_X1 U17542 ( .A(n14622), .ZN(n14310) );
  NAND2_X1 U17543 ( .A1(n14316), .A2(n14310), .ZN(n20355) );
  NAND2_X1 U17544 ( .A1(n20361), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14311) );
  OAI211_X1 U17545 ( .C1(n21484), .C2(n14320), .A(n20355), .B(n14311), .ZN(
        P1_U2948) );
  INV_X1 U17546 ( .A(n14627), .ZN(n14312) );
  NAND2_X1 U17547 ( .A1(n14316), .A2(n14312), .ZN(n20353) );
  NAND2_X1 U17548 ( .A1(n20361), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14313) );
  OAI211_X1 U17549 ( .C1(n14314), .C2(n14320), .A(n20353), .B(n14313), .ZN(
        P1_U2947) );
  INV_X1 U17550 ( .A(n14631), .ZN(n14315) );
  NAND2_X1 U17551 ( .A1(n14316), .A2(n14315), .ZN(n20351) );
  NAND2_X1 U17552 ( .A1(n20361), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14317) );
  OAI211_X1 U17553 ( .C1(n21466), .C2(n14320), .A(n20351), .B(n14317), .ZN(
        P1_U2946) );
  NAND2_X1 U17554 ( .A1(n20361), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14318) );
  OAI211_X1 U17555 ( .C1(n21478), .C2(n14320), .A(n14319), .B(n14318), .ZN(
        P1_U2945) );
  NOR2_X1 U17556 ( .A1(n16081), .A2(n16217), .ZN(n14321) );
  INV_X1 U17557 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16173) );
  NAND2_X1 U17558 ( .A1(n14805), .A2(n16173), .ZN(n14323) );
  NAND2_X1 U17559 ( .A1(n14803), .A2(n14323), .ZN(n14821) );
  NAND2_X1 U17560 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14324) );
  AND2_X1 U17561 ( .A1(n14336), .A2(n14324), .ZN(n14814) );
  INV_X1 U17562 ( .A(n14804), .ZN(n14326) );
  NAND2_X1 U17563 ( .A1(n14805), .A2(n14331), .ZN(n14325) );
  NAND2_X1 U17564 ( .A1(n14326), .A2(n14325), .ZN(n16068) );
  XNOR2_X1 U17565 ( .A(n16081), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14795) );
  NAND2_X1 U17566 ( .A1(n14805), .A2(n16159), .ZN(n14328) );
  NAND2_X1 U17567 ( .A1(n14795), .A2(n14328), .ZN(n16070) );
  NOR2_X1 U17568 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14329) );
  NAND2_X1 U17569 ( .A1(n14805), .A2(n16141), .ZN(n14330) );
  OR2_X1 U17570 ( .A1(n14805), .A2(n14331), .ZN(n14332) );
  NAND2_X1 U17571 ( .A1(n14803), .A2(n14332), .ZN(n14790) );
  NOR2_X1 U17572 ( .A1(n16081), .A2(n16159), .ZN(n16080) );
  NOR2_X1 U17573 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U17574 ( .A1(n14815), .A2(n14818), .ZN(n14333) );
  AND2_X1 U17575 ( .A1(n14334), .A2(n14333), .ZN(n14802) );
  XNOR2_X1 U17576 ( .A(n16081), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14783) );
  NAND2_X1 U17577 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14354) );
  INV_X1 U17578 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14933) );
  INV_X1 U17579 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16128) );
  INV_X1 U17580 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14944) );
  NAND4_X1 U17581 ( .A1(n16128), .A2(n14944), .A3(n14933), .A4(n14950), .ZN(
        n14337) );
  NAND2_X2 U17582 ( .A1(n14712), .A2(n14759), .ZN(n14699) );
  NAND3_X1 U17583 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U17584 ( .A1(n14712), .A2(n16081), .ZN(n14733) );
  NOR2_X2 U17585 ( .A1(n14699), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14734) );
  NOR2_X1 U17586 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14338) );
  AOI21_X2 U17587 ( .B1(n14734), .B2(n14338), .A(n16081), .ZN(n14724) );
  AND2_X1 U17588 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U17589 ( .A1(n14866), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14348) );
  INV_X1 U17590 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14857) );
  NAND2_X1 U17591 ( .A1(n14334), .A2(n14857), .ZN(n14687) );
  NOR2_X1 U17592 ( .A1(n14687), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14339) );
  NOR2_X1 U17593 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14678) );
  AOI22_X1 U17594 ( .A1(n14341), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14340), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14345) );
  MUX2_X1 U17595 ( .A(n14343), .B(n14342), .S(n14431), .Z(n14344) );
  XOR2_X1 U17596 ( .A(n14345), .B(n14344), .Z(n14568) );
  NOR2_X1 U17597 ( .A1(n14568), .A2(n16211), .ZN(n14366) );
  INV_X1 U17598 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16225) );
  NOR3_X1 U17599 ( .A1(n16225), .A2(n16231), .A3(n12259), .ZN(n16198) );
  AND3_X1 U17600 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16198), .ZN(n16192) );
  NAND2_X1 U17601 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16192), .ZN(
        n16179) );
  NOR2_X1 U17602 ( .A1(n14818), .A2(n16179), .ZN(n14352) );
  AND2_X1 U17603 ( .A1(n14352), .A2(n16197), .ZN(n16127) );
  NOR2_X1 U17604 ( .A1(n16173), .A2(n14331), .ZN(n16129) );
  NAND2_X1 U17605 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16152) );
  NOR2_X1 U17606 ( .A1(n16141), .A2(n16152), .ZN(n16133) );
  AND3_X1 U17607 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16129), .A3(
        n16133), .ZN(n14938) );
  AND2_X1 U17608 ( .A1(n16127), .A2(n14938), .ZN(n14350) );
  NAND2_X1 U17609 ( .A1(n16234), .A2(n14350), .ZN(n16126) );
  NAND2_X1 U17610 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14349) );
  INV_X1 U17611 ( .A(n14349), .ZN(n14346) );
  NOR2_X1 U17612 ( .A1(n14722), .A2(n14888), .ZN(n14347) );
  NAND2_X1 U17613 ( .A1(n14919), .A2(n14347), .ZN(n14874) );
  OR2_X1 U17614 ( .A1(n14874), .A2(n14348), .ZN(n14845) );
  INV_X1 U17615 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14846) );
  NOR3_X1 U17616 ( .A1(n14845), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14846), .ZN(n14365) );
  INV_X1 U17617 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21197) );
  NOR2_X1 U17618 ( .A1(n16210), .A2(n21197), .ZN(n14407) );
  AND2_X1 U17619 ( .A1(n16219), .A2(n14349), .ZN(n14359) );
  INV_X1 U17620 ( .A(n14350), .ZN(n14353) );
  NOR3_X1 U17621 ( .A1(n20411), .A2(n20397), .A3(n14351), .ZN(n16176) );
  NAND2_X1 U17622 ( .A1(n16176), .A2(n14352), .ZN(n14957) );
  INV_X1 U17623 ( .A(n14957), .ZN(n16168) );
  NAND2_X1 U17624 ( .A1(n16168), .A2(n14938), .ZN(n14941) );
  OAI21_X1 U17625 ( .B1(n20396), .B2(n14353), .A(n14941), .ZN(n14356) );
  INV_X1 U17626 ( .A(n14354), .ZN(n14355) );
  NAND2_X1 U17627 ( .A1(n14356), .A2(n14355), .ZN(n14357) );
  NAND2_X1 U17628 ( .A1(n16219), .A2(n14357), .ZN(n14358) );
  NAND2_X1 U17629 ( .A1(n14358), .A2(n14939), .ZN(n14929) );
  OR2_X1 U17630 ( .A1(n14359), .A2(n14929), .ZN(n14913) );
  NOR2_X1 U17631 ( .A1(n20398), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14360) );
  NOR2_X1 U17632 ( .A1(n14913), .A2(n14360), .ZN(n14904) );
  NAND2_X1 U17633 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14885) );
  AOI22_X1 U17634 ( .A1(n20396), .A2(n14885), .B1(n16180), .B2(n14909), .ZN(
        n14361) );
  NAND2_X1 U17635 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14362) );
  NAND2_X1 U17636 ( .A1(n16219), .A2(n14362), .ZN(n14363) );
  OAI21_X1 U17637 ( .B1(n16134), .B2(n14866), .A(n14873), .ZN(n14856) );
  AOI211_X1 U17638 ( .C1(n16219), .C2(n14857), .A(n14846), .B(n14856), .ZN(
        n14844) );
  AOI211_X1 U17639 ( .C1(n14887), .C2(n16134), .A(n12902), .B(n14844), .ZN(
        n14364) );
  NOR4_X1 U17640 ( .A1(n14366), .A2(n14365), .A3(n14407), .A4(n14364), .ZN(
        n14367) );
  OAI21_X1 U17641 ( .B1(n14413), .B2(n20387), .A(n14367), .ZN(P1_U3000) );
  INV_X1 U17642 ( .A(n14368), .ZN(n14972) );
  AOI22_X1 U17643 ( .A1(n14370), .A2(n14369), .B1(n14972), .B2(n15948), .ZN(
        n15946) );
  OAI21_X1 U17644 ( .B1(n15946), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21025), 
        .ZN(n14372) );
  INV_X1 U17645 ( .A(n14371), .ZN(n14981) );
  AOI22_X1 U17646 ( .A1(n14372), .A2(n14981), .B1(n15948), .B2(n14976), .ZN(
        n14376) );
  AOI21_X1 U17647 ( .B1(n14373), .B2(n16242), .A(n14375), .ZN(n14374) );
  OAI22_X1 U17648 ( .A1(n14376), .A2(n14375), .B1(n14374), .B2(n15948), .ZN(
        P1_U3474) );
  NAND2_X1 U17649 ( .A1(n14382), .A2(n20415), .ZN(n14386) );
  INV_X1 U17650 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U17651 ( .A1(n12180), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14378), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14379) );
  INV_X1 U17652 ( .A(n14379), .ZN(n14380) );
  XNOR2_X2 U17653 ( .A(n9894), .B(n14380), .ZN(n14414) );
  NAND3_X1 U17654 ( .A1(n14414), .A2(n14381), .A3(n14674), .ZN(n14385) );
  AOI22_X1 U17655 ( .A1(n14669), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14383), .ZN(n14384) );
  OAI211_X1 U17656 ( .C1(n14386), .C2(n19563), .A(n14385), .B(n14384), .ZN(
        P1_U2873) );
  INV_X1 U17657 ( .A(n14685), .ZN(n14391) );
  OAI22_X1 U17658 ( .A1(n14666), .A2(n14387), .B1(n14647), .B2(n21475), .ZN(
        n14388) );
  AOI21_X1 U17659 ( .B1(n14668), .B2(BUF1_REG_30__SCAN_IN), .A(n14388), .ZN(
        n14390) );
  NAND2_X1 U17660 ( .A1(n14669), .A2(DATAI_30_), .ZN(n14389) );
  OAI211_X1 U17661 ( .C1(n14391), .C2(n14672), .A(n14390), .B(n14389), .ZN(
        P1_U2874) );
  NOR3_X1 U17662 ( .A1(n15382), .A2(n15381), .A3(n14392), .ZN(n15368) );
  NAND2_X1 U17663 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15368), .ZN(
        n14395) );
  INV_X1 U17664 ( .A(n14395), .ZN(n14393) );
  OAI21_X1 U17665 ( .B1(n15620), .B2(n14393), .A(n15389), .ZN(n14394) );
  NAND2_X1 U17666 ( .A1(n14399), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17667 ( .A1(n12470), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12504), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14396) );
  AND2_X1 U17668 ( .A1(n14397), .A2(n14396), .ZN(n15131) );
  OR2_X2 U17669 ( .A1(n15130), .A2(n15131), .ZN(n15128) );
  AOI222_X1 U17670 ( .A1(n14399), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n14398), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n12504), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15120) );
  AOI222_X1 U17671 ( .A1(n14399), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14398), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n9842), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14400) );
  XNOR2_X1 U17672 ( .A(n14401), .B(n14400), .ZN(n19361) );
  NAND2_X1 U17673 ( .A1(n14404), .A2(n16493), .ZN(n14405) );
  OAI211_X1 U17674 ( .C1(n14406), .C2(n16477), .A(n9903), .B(n14405), .ZN(
        P2_U3015) );
  AOI21_X1 U17675 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14407), .ZN(n14408) );
  OAI21_X1 U17676 ( .B1(n20374), .B2(n14409), .A(n14408), .ZN(n14410) );
  OAI21_X1 U17677 ( .B1(n14413), .B2(n20242), .A(n14412), .ZN(P1_U2968) );
  NAND2_X1 U17678 ( .A1(n14414), .A2(n20292), .ZN(n14422) );
  INV_X1 U17679 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21353) );
  INV_X1 U17680 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21086) );
  NOR2_X1 U17681 ( .A1(n21353), .A2(n21086), .ZN(n14417) );
  INV_X1 U17682 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21447) );
  INV_X1 U17683 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21232) );
  INV_X1 U17684 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21068) );
  INV_X1 U17685 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21225) );
  INV_X1 U17686 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21062) );
  INV_X1 U17687 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21308) );
  NOR4_X1 U17688 ( .A1(n21225), .A2(n21062), .A3(n21308), .A4(n14555), .ZN(
        n16019) );
  NAND3_X1 U17689 ( .A1(n16019), .A2(P1_REIP_REG_18__SCAN_IN), .A3(
        P1_REIP_REG_19__SCAN_IN), .ZN(n14534) );
  NOR2_X1 U17690 ( .A1(n21068), .A2(n14534), .ZN(n16006) );
  NAND2_X1 U17691 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16006), .ZN(n14527) );
  NOR2_X1 U17692 ( .A1(n21232), .A2(n14527), .ZN(n14512) );
  NAND2_X1 U17693 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14512), .ZN(n14481) );
  NOR2_X1 U17694 ( .A1(n21447), .A2(n14481), .ZN(n14483) );
  NAND3_X1 U17695 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(n14483), .ZN(n14457) );
  INV_X1 U17696 ( .A(n14457), .ZN(n14415) );
  AND2_X1 U17697 ( .A1(n20277), .A2(n14415), .ZN(n14456) );
  AND3_X1 U17698 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14456), .A3(
        P1_REIP_REG_27__SCAN_IN), .ZN(n14416) );
  OR2_X1 U17699 ( .A1(n20279), .A2(n14416), .ZN(n14444) );
  OAI21_X1 U17700 ( .B1(n14417), .B2(n20318), .A(n14444), .ZN(n14425) );
  INV_X1 U17701 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14567) );
  INV_X1 U17702 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14418) );
  INV_X1 U17703 ( .A(n20307), .ZN(n16028) );
  OAI22_X1 U17704 ( .A1(n20297), .A2(n14567), .B1(n14418), .B2(n16028), .ZN(
        n14420) );
  INV_X1 U17705 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21079) );
  NOR3_X1 U17706 ( .A1(n20318), .A2(n14457), .A3(n21079), .ZN(n14446) );
  NAND2_X1 U17707 ( .A1(n14446), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14434) );
  NOR4_X1 U17708 ( .A1(n14434), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21353), 
        .A4(n21086), .ZN(n14419) );
  AOI211_X1 U17709 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14425), .A(n14420), 
        .B(n14419), .ZN(n14421) );
  OAI211_X1 U17710 ( .C1(n14568), .C2(n20313), .A(n14422), .B(n14421), .ZN(
        P1_U2809) );
  NAND2_X1 U17711 ( .A1(n14685), .A2(n20292), .ZN(n14428) );
  OAI21_X1 U17712 ( .B1(n14434), .B2(n21353), .A(n21086), .ZN(n14426) );
  AOI22_X1 U17713 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14681), .ZN(n14423) );
  OAI21_X1 U17714 ( .B1(n20297), .B2(n21192), .A(n14423), .ZN(n14424) );
  AOI21_X1 U17715 ( .B1(n14426), .B2(n14425), .A(n14424), .ZN(n14427) );
  OAI211_X1 U17716 ( .C1(n20313), .C2(n14842), .A(n14428), .B(n14427), .ZN(
        P1_U2810) );
  AOI21_X1 U17717 ( .B1(n14430), .B2(n14440), .A(n14429), .ZN(n14694) );
  INV_X1 U17718 ( .A(n14694), .ZN(n14617) );
  AOI21_X1 U17719 ( .B1(n14432), .B2(n9850), .A(n14431), .ZN(n14852) );
  OAI22_X1 U17720 ( .A1(n14433), .A2(n16028), .B1(n20324), .B2(n14692), .ZN(
        n14436) );
  NOR2_X1 U17721 ( .A1(n14434), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14435) );
  AOI211_X1 U17722 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n20315), .A(n14436), .B(
        n14435), .ZN(n14437) );
  OAI21_X1 U17723 ( .B1(n21353), .B2(n14444), .A(n14437), .ZN(n14438) );
  AOI21_X1 U17724 ( .B1(n14852), .B2(n20288), .A(n14438), .ZN(n14439) );
  OAI21_X1 U17725 ( .B1(n14617), .B2(n16051), .A(n14439), .ZN(P1_U2811) );
  OAI21_X1 U17726 ( .B1(n14454), .B2(n14441), .A(n14440), .ZN(n14710) );
  OR2_X1 U17727 ( .A1(n14453), .A2(n14442), .ZN(n14443) );
  AND2_X1 U17728 ( .A1(n9850), .A2(n14443), .ZN(n14865) );
  INV_X1 U17729 ( .A(n14444), .ZN(n14445) );
  OAI21_X1 U17730 ( .B1(n14446), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14445), 
        .ZN(n14448) );
  AOI22_X1 U17731 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14698), .ZN(n14447) );
  OAI211_X1 U17732 ( .C1(n20297), .C2(n14571), .A(n14448), .B(n14447), .ZN(
        n14449) );
  AOI21_X1 U17733 ( .B1(n14865), .B2(n20288), .A(n14449), .ZN(n14450) );
  OAI21_X1 U17734 ( .B1(n14710), .B2(n16051), .A(n14450), .ZN(P1_U2812) );
  NOR2_X1 U17735 ( .A1(n14475), .A2(n14451), .ZN(n14452) );
  OR2_X1 U17736 ( .A1(n14453), .A2(n14452), .ZN(n14876) );
  AOI21_X1 U17737 ( .B1(n14455), .B2(n14465), .A(n14454), .ZN(n14720) );
  NAND2_X1 U17738 ( .A1(n14720), .A2(n20292), .ZN(n14463) );
  NOR2_X1 U17739 ( .A1(n20279), .A2(n14456), .ZN(n14472) );
  INV_X1 U17740 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21481) );
  OR3_X1 U17741 ( .A1(n20318), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14457), .ZN(
        n14460) );
  INV_X1 U17742 ( .A(n14718), .ZN(n14458) );
  AOI22_X1 U17743 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14458), .ZN(n14459) );
  OAI211_X1 U17744 ( .C1(n20297), .C2(n21481), .A(n14460), .B(n14459), .ZN(
        n14461) );
  AOI21_X1 U17745 ( .B1(n14472), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14461), 
        .ZN(n14462) );
  OAI211_X1 U17746 ( .C1(n20313), .C2(n14876), .A(n14463), .B(n14462), .ZN(
        P1_U2813) );
  INV_X1 U17747 ( .A(n14479), .ZN(n14467) );
  INV_X1 U17748 ( .A(n14464), .ZN(n14466) );
  OAI21_X1 U17749 ( .B1(n14467), .B2(n14466), .A(n14465), .ZN(n14732) );
  INV_X1 U17750 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14726) );
  NAND3_X1 U17751 ( .A1(n14726), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14483), 
        .ZN(n14470) );
  INV_X1 U17752 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21260) );
  OR2_X1 U17753 ( .A1(n20297), .A2(n21260), .ZN(n14469) );
  AOI22_X1 U17754 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14729), .ZN(n14468) );
  OAI211_X1 U17755 ( .C1(n20318), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        n14471) );
  AOI21_X1 U17756 ( .B1(n14472), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14471), 
        .ZN(n14477) );
  AND2_X1 U17757 ( .A1(n14488), .A2(n14473), .ZN(n14474) );
  NOR2_X1 U17758 ( .A1(n14475), .A2(n14474), .ZN(n14884) );
  NAND2_X1 U17759 ( .A1(n14884), .A2(n20288), .ZN(n14476) );
  OAI211_X1 U17760 ( .C1(n14732), .C2(n16051), .A(n14477), .B(n14476), .ZN(
        P1_U2814) );
  OAI21_X1 U17761 ( .B1(n14478), .B2(n14480), .A(n14479), .ZN(n14742) );
  INV_X1 U17762 ( .A(n14481), .ZN(n14496) );
  AOI21_X1 U17763 ( .B1(n20277), .B2(n14496), .A(n20279), .ZN(n14511) );
  INV_X1 U17764 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U17765 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14482) );
  OAI211_X1 U17766 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14483), .A(n20270), 
        .B(n14482), .ZN(n14486) );
  INV_X1 U17767 ( .A(n14738), .ZN(n14484) );
  AOI22_X1 U17768 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14484), .ZN(n14485) );
  OAI211_X1 U17769 ( .C1(n14573), .C2(n20297), .A(n14486), .B(n14485), .ZN(
        n14492) );
  INV_X1 U17770 ( .A(n14499), .ZN(n14490) );
  INV_X1 U17771 ( .A(n14487), .ZN(n14489) );
  OAI21_X1 U17772 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14897) );
  NOR2_X1 U17773 ( .A1(n14897), .A2(n20313), .ZN(n14491) );
  AOI211_X1 U17774 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14511), .A(n14492), 
        .B(n14491), .ZN(n14493) );
  OAI21_X1 U17775 ( .B1(n14742), .B2(n16051), .A(n14493), .ZN(P1_U2815) );
  NOR2_X1 U17776 ( .A1(n14508), .A2(n14494), .ZN(n14495) );
  OR2_X1 U17777 ( .A1(n14478), .A2(n14495), .ZN(n14750) );
  NAND3_X1 U17778 ( .A1(n20270), .A2(n21447), .A3(n14496), .ZN(n14498) );
  AOI22_X1 U17779 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14747), .ZN(n14497) );
  OAI211_X1 U17780 ( .C1(n21479), .C2(n20297), .A(n14498), .B(n14497), .ZN(
        n14502) );
  OAI21_X1 U17781 ( .B1(n14506), .B2(n14500), .A(n14499), .ZN(n14905) );
  NOR2_X1 U17782 ( .A1(n14905), .A2(n20313), .ZN(n14501) );
  AOI211_X1 U17783 ( .C1(n14511), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14502), 
        .B(n14501), .ZN(n14503) );
  OAI21_X1 U17784 ( .B1(n14750), .B2(n16051), .A(n14503), .ZN(P1_U2816) );
  INV_X1 U17785 ( .A(n14579), .ZN(n14505) );
  AOI21_X1 U17786 ( .B1(n14505), .B2(n14522), .A(n14504), .ZN(n14507) );
  OR2_X1 U17787 ( .A1(n14507), .A2(n14506), .ZN(n14916) );
  AOI21_X1 U17788 ( .B1(n14509), .B2(n14519), .A(n14508), .ZN(n14757) );
  NAND2_X1 U17789 ( .A1(n14757), .A2(n20292), .ZN(n14518) );
  OAI22_X1 U17790 ( .A1(n14510), .A2(n16028), .B1(n20324), .B2(n14755), .ZN(
        n14516) );
  INV_X1 U17791 ( .A(n14511), .ZN(n14514) );
  AOI21_X1 U17792 ( .B1(n20270), .B2(n14512), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14513) );
  NOR2_X1 U17793 ( .A1(n14514), .A2(n14513), .ZN(n14515) );
  AOI211_X1 U17794 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20315), .A(n14516), .B(
        n14515), .ZN(n14517) );
  OAI211_X1 U17795 ( .C1(n20313), .C2(n14916), .A(n14518), .B(n14517), .ZN(
        P1_U2817) );
  INV_X1 U17796 ( .A(n14519), .ZN(n14520) );
  AOI21_X1 U17797 ( .B1(n14521), .B2(n14574), .A(n14520), .ZN(n14762) );
  INV_X1 U17798 ( .A(n14762), .ZN(n14646) );
  INV_X1 U17799 ( .A(n14522), .ZN(n14523) );
  XNOR2_X1 U17800 ( .A(n14579), .B(n14523), .ZN(n14922) );
  INV_X1 U17801 ( .A(n14922), .ZN(n14530) );
  INV_X1 U17802 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21340) );
  OAI21_X1 U17803 ( .B1(n16006), .B2(n20318), .A(n20277), .ZN(n16012) );
  AOI21_X1 U17804 ( .B1(n20270), .B2(n21340), .A(n16012), .ZN(n14526) );
  AOI22_X1 U17805 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14765), .ZN(n14525) );
  NAND2_X1 U17806 ( .A1(n20315), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14524) );
  OAI211_X1 U17807 ( .C1(n14526), .C2(n21232), .A(n14525), .B(n14524), .ZN(
        n14529) );
  NOR3_X1 U17808 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20318), .A3(n14527), 
        .ZN(n14528) );
  AOI211_X1 U17809 ( .C1(n14530), .C2(n20288), .A(n14529), .B(n14528), .ZN(
        n14531) );
  OAI21_X1 U17810 ( .B1(n14646), .B2(n16051), .A(n14531), .ZN(P1_U2818) );
  XNOR2_X1 U17811 ( .A(n14584), .B(n14533), .ZN(n14782) );
  OAI21_X1 U17812 ( .B1(n20318), .B2(n14534), .A(n21068), .ZN(n14540) );
  INV_X1 U17813 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14582) );
  NAND2_X1 U17814 ( .A1(n14588), .A2(n14535), .ZN(n14536) );
  AND2_X1 U17815 ( .A1(n9878), .A2(n14536), .ZN(n14949) );
  NAND2_X1 U17816 ( .A1(n14949), .A2(n20288), .ZN(n14538) );
  AOI22_X1 U17817 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20307), .B1(
        n20264), .B2(n14779), .ZN(n14537) );
  OAI211_X1 U17818 ( .C1(n14582), .C2(n20297), .A(n14538), .B(n14537), .ZN(
        n14539) );
  AOI21_X1 U17819 ( .B1(n16012), .B2(n14540), .A(n14539), .ZN(n14541) );
  OAI21_X1 U17820 ( .B1(n14782), .B2(n16051), .A(n14541), .ZN(P1_U2820) );
  XOR2_X1 U17821 ( .A(n14583), .B(n14593), .Z(n14788) );
  NOR2_X1 U17822 ( .A1(n14599), .A2(n14543), .ZN(n14544) );
  OR2_X1 U17823 ( .A1(n14587), .A2(n14544), .ZN(n16135) );
  INV_X1 U17824 ( .A(n16135), .ZN(n14552) );
  INV_X1 U17825 ( .A(n14545), .ZN(n14786) );
  NAND2_X1 U17826 ( .A1(n20307), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14547) );
  INV_X1 U17827 ( .A(n20306), .ZN(n14546) );
  OAI211_X1 U17828 ( .C1(n20324), .C2(n14786), .A(n14547), .B(n14546), .ZN(
        n14551) );
  NAND2_X1 U17829 ( .A1(n20270), .A2(n16019), .ZN(n14549) );
  OAI21_X1 U17830 ( .B1(n20318), .B2(n16019), .A(n20277), .ZN(n16027) );
  AOI22_X1 U17831 ( .A1(n16027), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n20315), .ZN(n14548) );
  OAI21_X1 U17832 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n14549), .A(n14548), 
        .ZN(n14550) );
  AOI211_X1 U17833 ( .C1(n14552), .C2(n20288), .A(n14551), .B(n14550), .ZN(
        n14553) );
  OAI21_X1 U17834 ( .B1(n14662), .B2(n16051), .A(n14553), .ZN(P1_U2822) );
  XOR2_X1 U17835 ( .A(n14554), .B(n14075), .Z(n14800) );
  NOR3_X1 U17836 ( .A1(n20318), .A2(n21308), .A3(n14555), .ZN(n16026) );
  INV_X1 U17837 ( .A(n16026), .ZN(n14557) );
  NOR3_X1 U17838 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n20318), .A3(n14555), 
        .ZN(n16037) );
  NOR2_X1 U17839 ( .A1(n16037), .A2(n16036), .ZN(n14556) );
  MUX2_X1 U17840 ( .A(n14557), .B(n14556), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14566) );
  NAND2_X1 U17841 ( .A1(n14609), .A2(n14558), .ZN(n14559) );
  NAND2_X1 U17842 ( .A1(n14597), .A2(n14559), .ZN(n16149) );
  INV_X1 U17843 ( .A(n16149), .ZN(n14564) );
  INV_X1 U17844 ( .A(n14560), .ZN(n14798) );
  NOR2_X1 U17845 ( .A1(n20324), .A2(n14798), .ZN(n14561) );
  AOI211_X1 U17846 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20306), .B(n14561), .ZN(n14562) );
  OAI21_X1 U17847 ( .B1(n14603), .B2(n20297), .A(n14562), .ZN(n14563) );
  AOI21_X1 U17848 ( .B1(n20288), .B2(n14564), .A(n14563), .ZN(n14565) );
  OAI211_X1 U17849 ( .C1(n14673), .C2(n16051), .A(n14566), .B(n14565), .ZN(
        P1_U2824) );
  OAI22_X1 U17850 ( .A1(n14568), .A2(n14613), .B1(n14612), .B2(n14567), .ZN(
        P1_U2841) );
  AOI22_X1 U17851 ( .A1(n14852), .A2(n14601), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14600), .ZN(n14569) );
  OAI21_X1 U17852 ( .B1(n14617), .B2(n14610), .A(n14569), .ZN(P1_U2843) );
  INV_X1 U17853 ( .A(n14865), .ZN(n14570) );
  OAI222_X1 U17854 ( .A1(n14610), .A2(n14710), .B1(n14571), .B2(n14612), .C1(
        n14570), .C2(n14613), .ZN(P1_U2844) );
  INV_X1 U17855 ( .A(n14720), .ZN(n14626) );
  OAI222_X1 U17856 ( .A1(n14610), .A2(n14626), .B1(n21481), .B2(n14612), .C1(
        n14876), .C2(n14613), .ZN(P1_U2845) );
  INV_X1 U17857 ( .A(n14884), .ZN(n14572) );
  OAI222_X1 U17858 ( .A1(n14610), .A2(n14732), .B1(n21260), .B2(n14612), .C1(
        n14572), .C2(n14613), .ZN(P1_U2846) );
  OAI222_X1 U17859 ( .A1(n14610), .A2(n14742), .B1(n14573), .B2(n14612), .C1(
        n14897), .C2(n14613), .ZN(P1_U2847) );
  OAI222_X1 U17860 ( .A1(n14610), .A2(n14750), .B1(n21479), .B2(n14612), .C1(
        n14905), .C2(n14613), .ZN(P1_U2848) );
  INV_X1 U17861 ( .A(n14757), .ZN(n14642) );
  OAI222_X1 U17862 ( .A1(n14610), .A2(n14642), .B1(n21336), .B2(n14612), .C1(
        n14916), .C2(n14613), .ZN(P1_U2849) );
  INV_X1 U17863 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n21468) );
  OAI222_X1 U17864 ( .A1(n14646), .A2(n14610), .B1(n14612), .B2(n21468), .C1(
        n14613), .C2(n14922), .ZN(P1_U2850) );
  OAI21_X1 U17865 ( .B1(n14576), .B2(n14575), .A(n14574), .ZN(n14771) );
  INV_X1 U17866 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U17867 ( .A1(n9878), .A2(n14577), .ZN(n14578) );
  NAND2_X1 U17868 ( .A1(n14579), .A2(n14578), .ZN(n16013) );
  OAI222_X1 U17869 ( .A1(n14610), .A2(n14771), .B1(n14612), .B2(n14580), .C1(
        n16013), .C2(n14613), .ZN(P1_U2851) );
  INV_X1 U17870 ( .A(n14949), .ZN(n14581) );
  OAI222_X1 U17871 ( .A1(n14782), .A2(n14610), .B1(n14612), .B2(n14582), .C1(
        n14581), .C2(n14613), .ZN(P1_U2852) );
  OR2_X1 U17872 ( .A1(n14593), .A2(n14583), .ZN(n14585) );
  AOI21_X1 U17873 ( .B1(n14586), .B2(n14585), .A(n14584), .ZN(n16064) );
  INV_X1 U17874 ( .A(n16064), .ZN(n14658) );
  INV_X1 U17875 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14592) );
  INV_X1 U17876 ( .A(n14587), .ZN(n14589) );
  AOI21_X1 U17877 ( .B1(n14590), .B2(n14589), .A(n10334), .ZN(n16122) );
  INV_X1 U17878 ( .A(n16122), .ZN(n14591) );
  OAI222_X1 U17879 ( .A1(n14658), .A2(n14610), .B1(n14612), .B2(n14592), .C1(
        n14591), .C2(n14613), .ZN(P1_U2853) );
  INV_X1 U17880 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21286) );
  OAI222_X1 U17881 ( .A1(n14662), .A2(n14610), .B1(n14612), .B2(n21286), .C1(
        n16135), .C2(n14613), .ZN(P1_U2854) );
  OAI21_X1 U17882 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n16031) );
  AND2_X1 U17883 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  NOR2_X1 U17884 ( .A1(n14599), .A2(n14598), .ZN(n16142) );
  AOI22_X1 U17885 ( .A1(n16142), .A2(n14601), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14600), .ZN(n14602) );
  OAI21_X1 U17886 ( .B1(n16031), .B2(n14610), .A(n14602), .ZN(P1_U2855) );
  OAI22_X1 U17887 ( .A1(n16149), .A2(n14613), .B1(n14603), .B2(n14612), .ZN(
        n14604) );
  INV_X1 U17888 ( .A(n14604), .ZN(n14605) );
  OAI21_X1 U17889 ( .B1(n14673), .B2(n14610), .A(n14605), .ZN(P1_U2856) );
  OR2_X1 U17890 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  NAND2_X1 U17891 ( .A1(n14609), .A2(n14608), .ZN(n16038) );
  INV_X1 U17892 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21313) );
  OAI222_X1 U17893 ( .A1(n16038), .A2(n14613), .B1(n14612), .B2(n21313), .C1(
        n14611), .C2(n14610), .ZN(P1_U2857) );
  OAI22_X1 U17894 ( .A1(n14666), .A2(n14677), .B1(n14647), .B2(n14307), .ZN(
        n14614) );
  AOI21_X1 U17895 ( .B1(n14668), .B2(BUF1_REG_29__SCAN_IN), .A(n14614), .ZN(
        n14616) );
  NAND2_X1 U17896 ( .A1(n14669), .A2(DATAI_29_), .ZN(n14615) );
  OAI211_X1 U17897 ( .C1(n14617), .C2(n14672), .A(n14616), .B(n14615), .ZN(
        P1_U2875) );
  OAI22_X1 U17898 ( .A1(n14666), .A2(n14618), .B1(n14647), .B2(n21459), .ZN(
        n14619) );
  AOI21_X1 U17899 ( .B1(n14668), .B2(BUF1_REG_28__SCAN_IN), .A(n14619), .ZN(
        n14621) );
  NAND2_X1 U17900 ( .A1(n14669), .A2(DATAI_28_), .ZN(n14620) );
  OAI211_X1 U17901 ( .C1(n14710), .C2(n14672), .A(n14621), .B(n14620), .ZN(
        P1_U2876) );
  OAI22_X1 U17902 ( .A1(n14666), .A2(n14622), .B1(n14647), .B2(n21484), .ZN(
        n14623) );
  AOI21_X1 U17903 ( .B1(n14668), .B2(BUF1_REG_27__SCAN_IN), .A(n14623), .ZN(
        n14625) );
  NAND2_X1 U17904 ( .A1(n14669), .A2(DATAI_27_), .ZN(n14624) );
  OAI211_X1 U17905 ( .C1(n14626), .C2(n14672), .A(n14625), .B(n14624), .ZN(
        P1_U2877) );
  OAI22_X1 U17906 ( .A1(n14666), .A2(n14627), .B1(n14647), .B2(n14314), .ZN(
        n14628) );
  AOI21_X1 U17907 ( .B1(n14668), .B2(BUF1_REG_26__SCAN_IN), .A(n14628), .ZN(
        n14630) );
  NAND2_X1 U17908 ( .A1(n14669), .A2(DATAI_26_), .ZN(n14629) );
  OAI211_X1 U17909 ( .C1(n14732), .C2(n14672), .A(n14630), .B(n14629), .ZN(
        P1_U2878) );
  OAI22_X1 U17910 ( .A1(n14666), .A2(n14631), .B1(n14674), .B2(n21466), .ZN(
        n14632) );
  AOI21_X1 U17911 ( .B1(n14668), .B2(BUF1_REG_25__SCAN_IN), .A(n14632), .ZN(
        n14634) );
  NAND2_X1 U17912 ( .A1(n14669), .A2(DATAI_25_), .ZN(n14633) );
  OAI211_X1 U17913 ( .C1(n14742), .C2(n14672), .A(n14634), .B(n14633), .ZN(
        P1_U2879) );
  OAI22_X1 U17914 ( .A1(n14666), .A2(n14635), .B1(n14647), .B2(n21478), .ZN(
        n14636) );
  AOI21_X1 U17915 ( .B1(n14668), .B2(BUF1_REG_24__SCAN_IN), .A(n14636), .ZN(
        n14638) );
  NAND2_X1 U17916 ( .A1(n14669), .A2(DATAI_24_), .ZN(n14637) );
  OAI211_X1 U17917 ( .C1(n14750), .C2(n14672), .A(n14638), .B(n14637), .ZN(
        P1_U2880) );
  OAI22_X1 U17918 ( .A1(n14666), .A2(n20482), .B1(n14647), .B2(n21238), .ZN(
        n14639) );
  AOI21_X1 U17919 ( .B1(n14668), .B2(BUF1_REG_23__SCAN_IN), .A(n14639), .ZN(
        n14641) );
  NAND2_X1 U17920 ( .A1(n14669), .A2(DATAI_23_), .ZN(n14640) );
  OAI211_X1 U17921 ( .C1(n14642), .C2(n14672), .A(n14641), .B(n14640), .ZN(
        P1_U2881) );
  OAI22_X1 U17922 ( .A1(n14666), .A2(n20473), .B1(n14647), .B2(n12815), .ZN(
        n14643) );
  AOI21_X1 U17923 ( .B1(n14668), .B2(BUF1_REG_22__SCAN_IN), .A(n14643), .ZN(
        n14645) );
  NAND2_X1 U17924 ( .A1(n14669), .A2(DATAI_22_), .ZN(n14644) );
  OAI211_X1 U17925 ( .C1(n14646), .C2(n14672), .A(n14645), .B(n14644), .ZN(
        P1_U2882) );
  OAI22_X1 U17926 ( .A1(n14666), .A2(n20465), .B1(n14647), .B2(n21226), .ZN(
        n14648) );
  AOI21_X1 U17927 ( .B1(n14668), .B2(BUF1_REG_21__SCAN_IN), .A(n14648), .ZN(
        n14650) );
  NAND2_X1 U17928 ( .A1(n14669), .A2(DATAI_21_), .ZN(n14649) );
  OAI211_X1 U17929 ( .C1(n14771), .C2(n14672), .A(n14650), .B(n14649), .ZN(
        P1_U2883) );
  OAI22_X1 U17930 ( .A1(n14666), .A2(n20459), .B1(n14674), .B2(n21323), .ZN(
        n14651) );
  AOI21_X1 U17931 ( .B1(n14668), .B2(BUF1_REG_20__SCAN_IN), .A(n14651), .ZN(
        n14653) );
  NAND2_X1 U17932 ( .A1(n14669), .A2(DATAI_20_), .ZN(n14652) );
  OAI211_X1 U17933 ( .C1(n14782), .C2(n14672), .A(n14653), .B(n14652), .ZN(
        P1_U2884) );
  OAI22_X1 U17934 ( .A1(n14666), .A2(n20454), .B1(n14674), .B2(n14654), .ZN(
        n14655) );
  AOI21_X1 U17935 ( .B1(n14668), .B2(BUF1_REG_19__SCAN_IN), .A(n14655), .ZN(
        n14657) );
  NAND2_X1 U17936 ( .A1(n14669), .A2(DATAI_19_), .ZN(n14656) );
  OAI211_X1 U17937 ( .C1(n14658), .C2(n14672), .A(n14657), .B(n14656), .ZN(
        P1_U2885) );
  OAI22_X1 U17938 ( .A1(n14666), .A2(n20448), .B1(n14674), .B2(n12823), .ZN(
        n14659) );
  AOI21_X1 U17939 ( .B1(n14668), .B2(BUF1_REG_18__SCAN_IN), .A(n14659), .ZN(
        n14661) );
  NAND2_X1 U17940 ( .A1(n14669), .A2(DATAI_18_), .ZN(n14660) );
  OAI211_X1 U17941 ( .C1(n14662), .C2(n14672), .A(n14661), .B(n14660), .ZN(
        P1_U2886) );
  OAI22_X1 U17942 ( .A1(n14666), .A2(n20442), .B1(n14674), .B2(n12821), .ZN(
        n14663) );
  AOI21_X1 U17943 ( .B1(n14668), .B2(BUF1_REG_17__SCAN_IN), .A(n14663), .ZN(
        n14665) );
  NAND2_X1 U17944 ( .A1(n14669), .A2(DATAI_17_), .ZN(n14664) );
  OAI211_X1 U17945 ( .C1(n16031), .C2(n14672), .A(n14665), .B(n14664), .ZN(
        P1_U2887) );
  OAI22_X1 U17946 ( .A1(n14666), .A2(n20431), .B1(n14674), .B2(n12812), .ZN(
        n14667) );
  AOI21_X1 U17947 ( .B1(n14668), .B2(BUF1_REG_16__SCAN_IN), .A(n14667), .ZN(
        n14671) );
  NAND2_X1 U17948 ( .A1(n14669), .A2(DATAI_16_), .ZN(n14670) );
  OAI211_X1 U17949 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        P1_U2888) );
  INV_X1 U17950 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14675) );
  OAI222_X1 U17951 ( .A1(n14829), .A2(n14672), .B1(n14677), .B2(n14676), .C1(
        n14675), .C2(n14674), .ZN(P1_U2891) );
  INV_X1 U17952 ( .A(n14678), .ZN(n14868) );
  NOR2_X1 U17953 ( .A1(n14687), .A2(n14868), .ZN(n14680) );
  NAND2_X1 U17954 ( .A1(n16094), .A2(n14681), .ZN(n14682) );
  NAND2_X1 U17955 ( .A1(n20380), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14843) );
  OAI211_X1 U17956 ( .C1(n14683), .C2(n14824), .A(n14682), .B(n14843), .ZN(
        n14684) );
  AOI21_X1 U17957 ( .B1(n14685), .B2(n14411), .A(n14684), .ZN(n14686) );
  OAI21_X1 U17958 ( .B1(n14851), .B2(n20242), .A(n14686), .ZN(P1_U2969) );
  INV_X1 U17959 ( .A(n14687), .ZN(n14688) );
  AOI21_X1 U17960 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16081), .A(
        n14688), .ZN(n14689) );
  XNOR2_X1 U17961 ( .A(n14690), .B(n14689), .ZN(n14860) );
  NOR2_X1 U17962 ( .A1(n16210), .A2(n21353), .ZN(n14855) );
  AOI21_X1 U17963 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14855), .ZN(n14691) );
  OAI21_X1 U17964 ( .B1(n20374), .B2(n14692), .A(n14691), .ZN(n14693) );
  AOI21_X1 U17965 ( .B1(n14694), .B2(n14411), .A(n14693), .ZN(n14695) );
  OAI21_X1 U17966 ( .B1(n14860), .B2(n20242), .A(n14695), .ZN(P1_U2970) );
  INV_X1 U17967 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21081) );
  NOR2_X1 U17968 ( .A1(n16210), .A2(n21081), .ZN(n14864) );
  NOR2_X1 U17969 ( .A1(n14824), .A2(n14696), .ZN(n14697) );
  AOI211_X1 U17970 ( .C1(n14698), .C2(n16094), .A(n14864), .B(n14697), .ZN(
        n14709) );
  NAND2_X1 U17971 ( .A1(n16081), .A2(n14722), .ZN(n14700) );
  NAND2_X1 U17972 ( .A1(n14699), .A2(n14700), .ZN(n14704) );
  NOR2_X1 U17973 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14701) );
  AND4_X1 U17974 ( .A1(n14701), .A2(n14909), .A3(n14918), .A4(n14888), .ZN(
        n14702) );
  AND2_X1 U17975 ( .A1(n14704), .A2(n14702), .ZN(n14706) );
  NAND2_X1 U17976 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14703) );
  NOR2_X1 U17977 ( .A1(n14704), .A2(n14703), .ZN(n14705) );
  MUX2_X1 U17978 ( .A(n14706), .B(n14705), .S(n14805), .Z(n14707) );
  XNOR2_X1 U17979 ( .A(n14707), .B(n14862), .ZN(n14861) );
  NAND2_X1 U17980 ( .A1(n14861), .A2(n20370), .ZN(n14708) );
  OAI211_X1 U17981 ( .C1(n14710), .C2(n20417), .A(n14709), .B(n14708), .ZN(
        P1_U2971) );
  INV_X1 U17982 ( .A(n14711), .ZN(n14713) );
  NOR2_X1 U17983 ( .A1(n14713), .A2(n14712), .ZN(n14715) );
  MUX2_X1 U17984 ( .A(n14715), .B(n14714), .S(n14334), .Z(n14716) );
  XNOR2_X1 U17985 ( .A(n14716), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14881) );
  OR2_X1 U17986 ( .A1(n16210), .A2(n21079), .ZN(n14875) );
  NAND2_X1 U17987 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14717) );
  OAI211_X1 U17988 ( .C1(n20374), .C2(n14718), .A(n14875), .B(n14717), .ZN(
        n14719) );
  AOI21_X1 U17989 ( .B1(n14720), .B2(n14411), .A(n14719), .ZN(n14721) );
  OAI21_X1 U17990 ( .B1(n14881), .B2(n20242), .A(n14721), .ZN(P1_U2972) );
  INV_X1 U17991 ( .A(n14722), .ZN(n14889) );
  AOI21_X1 U17992 ( .B1(n14699), .B2(n14889), .A(n14334), .ZN(n14723) );
  NOR2_X1 U17993 ( .A1(n14724), .A2(n14723), .ZN(n14725) );
  XNOR2_X1 U17994 ( .A(n14725), .B(n14888), .ZN(n14882) );
  NAND2_X1 U17995 ( .A1(n14882), .A2(n20370), .ZN(n14731) );
  NOR2_X1 U17996 ( .A1(n16210), .A2(n14726), .ZN(n14883) );
  INV_X1 U17997 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14727) );
  NOR2_X1 U17998 ( .A1(n14824), .A2(n14727), .ZN(n14728) );
  AOI211_X1 U17999 ( .C1(n16094), .C2(n14729), .A(n14883), .B(n14728), .ZN(
        n14730) );
  OAI211_X1 U18000 ( .C1(n20417), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        P1_U2973) );
  NAND2_X1 U18001 ( .A1(n14733), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14744) );
  INV_X1 U18002 ( .A(n14744), .ZN(n14736) );
  MUX2_X1 U18003 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14734), .S(
        n14334), .Z(n14735) );
  OAI21_X1 U18004 ( .B1(n14736), .B2(n14909), .A(n14735), .ZN(n14737) );
  XNOR2_X1 U18005 ( .A(n14737), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14894) );
  NAND2_X1 U18006 ( .A1(n14894), .A2(n20370), .ZN(n14741) );
  INV_X1 U18007 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21075) );
  NOR2_X1 U18008 ( .A1(n16210), .A2(n21075), .ZN(n14895) );
  NOR2_X1 U18009 ( .A1(n20374), .A2(n14738), .ZN(n14739) );
  AOI211_X1 U18010 ( .C1(n20365), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14895), .B(n14739), .ZN(n14740) );
  OAI211_X1 U18011 ( .C1(n20417), .C2(n14742), .A(n14741), .B(n14740), .ZN(
        P1_U2974) );
  INV_X1 U18012 ( .A(n14699), .ZN(n14743) );
  NAND2_X1 U18013 ( .A1(n14743), .A2(n14744), .ZN(n14745) );
  MUX2_X1 U18014 ( .A(n14745), .B(n14744), .S(n14805), .Z(n14746) );
  XNOR2_X1 U18015 ( .A(n14746), .B(n14909), .ZN(n14912) );
  NOR2_X1 U18016 ( .A1(n16210), .A2(n21447), .ZN(n14907) );
  AOI21_X1 U18017 ( .B1(n20365), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14907), .ZN(n14749) );
  NAND2_X1 U18018 ( .A1(n16094), .A2(n14747), .ZN(n14748) );
  OAI211_X1 U18019 ( .C1(n14750), .C2(n20417), .A(n14749), .B(n14748), .ZN(
        n14751) );
  INV_X1 U18020 ( .A(n14751), .ZN(n14752) );
  OAI21_X1 U18021 ( .B1(n14912), .B2(n20242), .A(n14752), .ZN(P1_U2975) );
  XNOR2_X1 U18022 ( .A(n16081), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14753) );
  XNOR2_X1 U18023 ( .A(n14699), .B(n14753), .ZN(n14921) );
  NAND2_X1 U18024 ( .A1(n20380), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U18025 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14754) );
  OAI211_X1 U18026 ( .C1(n20374), .C2(n14755), .A(n14915), .B(n14754), .ZN(
        n14756) );
  AOI21_X1 U18027 ( .B1(n14757), .B2(n14411), .A(n14756), .ZN(n14758) );
  OAI21_X1 U18028 ( .B1(n14921), .B2(n20242), .A(n14758), .ZN(P1_U2976) );
  NAND2_X1 U18029 ( .A1(n14760), .A2(n14759), .ZN(n14761) );
  XOR2_X1 U18030 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14761), .Z(
        n14928) );
  NAND2_X1 U18031 ( .A1(n14762), .A2(n14411), .ZN(n14767) );
  NOR2_X1 U18032 ( .A1(n16210), .A2(n21232), .ZN(n14924) );
  NOR2_X1 U18033 ( .A1(n14824), .A2(n14763), .ZN(n14764) );
  AOI211_X1 U18034 ( .C1(n16094), .C2(n14765), .A(n14924), .B(n14764), .ZN(
        n14766) );
  OAI211_X1 U18035 ( .C1(n14928), .C2(n20242), .A(n14767), .B(n14766), .ZN(
        P1_U2977) );
  OAI21_X1 U18036 ( .B1(n14805), .B2(n16128), .A(n14768), .ZN(n16063) );
  OR2_X1 U18037 ( .A1(n14805), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16059) );
  NOR2_X1 U18038 ( .A1(n14334), .A2(n14944), .ZN(n16061) );
  NAND3_X1 U18039 ( .A1(n14784), .A2(n14783), .A3(n16061), .ZN(n14769) );
  OAI21_X1 U18040 ( .B1(n16063), .B2(n16059), .A(n14769), .ZN(n14776) );
  NAND2_X1 U18041 ( .A1(n14776), .A2(n14950), .ZN(n14775) );
  OAI22_X1 U18042 ( .A1(n14775), .A2(n16081), .B1(n14950), .B2(n14769), .ZN(
        n14770) );
  XNOR2_X1 U18043 ( .A(n14770), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14936) );
  INV_X1 U18044 ( .A(n14771), .ZN(n16015) );
  NAND2_X1 U18045 ( .A1(n20380), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14931) );
  NAND2_X1 U18046 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14772) );
  OAI211_X1 U18047 ( .C1(n20374), .C2(n16018), .A(n14931), .B(n14772), .ZN(
        n14773) );
  AOI21_X1 U18048 ( .B1(n16015), .B2(n14411), .A(n14773), .ZN(n14774) );
  OAI21_X1 U18049 ( .B1(n14936), .B2(n20242), .A(n14774), .ZN(P1_U2978) );
  OAI21_X1 U18050 ( .B1(n14776), .B2(n14950), .A(n14775), .ZN(n14937) );
  NAND2_X1 U18051 ( .A1(n14937), .A2(n20370), .ZN(n14781) );
  NOR2_X1 U18052 ( .A1(n16210), .A2(n21068), .ZN(n14948) );
  INV_X1 U18053 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14777) );
  NOR2_X1 U18054 ( .A1(n14824), .A2(n14777), .ZN(n14778) );
  AOI211_X1 U18055 ( .C1(n16094), .C2(n14779), .A(n14948), .B(n14778), .ZN(
        n14780) );
  OAI211_X1 U18056 ( .C1(n20417), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        P1_U2979) );
  XNOR2_X1 U18057 ( .A(n14784), .B(n14783), .ZN(n16136) );
  AOI22_X1 U18058 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U18059 ( .B1(n20374), .B2(n14786), .A(n14785), .ZN(n14787) );
  AOI21_X1 U18060 ( .B1(n14788), .B2(n14411), .A(n14787), .ZN(n14789) );
  OAI21_X1 U18061 ( .B1(n16136), .B2(n20242), .A(n14789), .ZN(P1_U2981) );
  INV_X1 U18062 ( .A(n14790), .ZN(n14792) );
  INV_X1 U18063 ( .A(n14802), .ZN(n14791) );
  NAND3_X1 U18064 ( .A1(n14793), .A2(n14792), .A3(n14791), .ZN(n16083) );
  NOR2_X1 U18065 ( .A1(n16083), .A2(n16080), .ZN(n14794) );
  NOR2_X1 U18066 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16148) );
  NOR2_X1 U18067 ( .A1(n14794), .A2(n16148), .ZN(n14796) );
  OAI22_X1 U18068 ( .A1(n14796), .A2(n14795), .B1(n14794), .B2(n16070), .ZN(
        n16150) );
  AOI22_X1 U18069 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14797) );
  OAI21_X1 U18070 ( .B1(n20374), .B2(n14798), .A(n14797), .ZN(n14799) );
  AOI21_X1 U18071 ( .B1(n14800), .B2(n14411), .A(n14799), .ZN(n14801) );
  OAI21_X1 U18072 ( .B1(n16150), .B2(n20242), .A(n14801), .ZN(P1_U2983) );
  NOR2_X1 U18073 ( .A1(n9893), .A2(n14802), .ZN(n16069) );
  OAI21_X1 U18074 ( .B1(n16069), .B2(n14804), .A(n14803), .ZN(n14807) );
  MUX2_X1 U18075 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n14331), .S(
        n14805), .Z(n14806) );
  XNOR2_X1 U18076 ( .A(n14807), .B(n14806), .ZN(n14955) );
  INV_X1 U18077 ( .A(n14955), .ZN(n14813) );
  AOI22_X1 U18078 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14808) );
  OAI21_X1 U18079 ( .B1(n20374), .B2(n14809), .A(n14808), .ZN(n14810) );
  AOI21_X1 U18080 ( .B1(n14811), .B2(n14411), .A(n14810), .ZN(n14812) );
  OAI21_X1 U18081 ( .B1(n14813), .B2(n20242), .A(n14812), .ZN(P1_U2985) );
  OR2_X1 U18082 ( .A1(n10132), .A2(n14814), .ZN(n14817) );
  OR2_X1 U18083 ( .A1(n14805), .A2(n14815), .ZN(n14816) );
  NAND2_X1 U18084 ( .A1(n14817), .A2(n14816), .ZN(n16090) );
  NOR2_X1 U18085 ( .A1(n16081), .A2(n14818), .ZN(n14819) );
  OR2_X1 U18086 ( .A1(n14820), .A2(n14819), .ZN(n16089) );
  NOR2_X1 U18087 ( .A1(n16090), .A2(n16089), .ZN(n16088) );
  NOR2_X1 U18088 ( .A1(n16088), .A2(n14820), .ZN(n14822) );
  XNOR2_X1 U18089 ( .A(n14822), .B(n14821), .ZN(n16170) );
  NAND2_X1 U18090 ( .A1(n16170), .A2(n20370), .ZN(n14828) );
  INV_X1 U18091 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14823) );
  OAI22_X1 U18092 ( .A1(n14824), .A2(n14823), .B1(n16210), .B2(n21289), .ZN(
        n14825) );
  AOI21_X1 U18093 ( .B1(n16094), .B2(n14826), .A(n14825), .ZN(n14827) );
  OAI211_X1 U18094 ( .C1(n20417), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        P1_U2986) );
  XNOR2_X1 U18095 ( .A(n10132), .B(n16207), .ZN(n14831) );
  NAND2_X1 U18096 ( .A1(n14832), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14830) );
  MUX2_X1 U18097 ( .A(n14831), .B(n14830), .S(n14334), .Z(n14835) );
  INV_X1 U18098 ( .A(n14832), .ZN(n14834) );
  NAND3_X1 U18099 ( .A1(n14834), .A2(n14833), .A3(n16207), .ZN(n16097) );
  NAND2_X1 U18100 ( .A1(n14835), .A2(n16097), .ZN(n16205) );
  INV_X1 U18101 ( .A(n16205), .ZN(n14841) );
  AOI22_X1 U18102 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14836) );
  OAI21_X1 U18103 ( .B1(n20374), .B2(n14837), .A(n14836), .ZN(n14838) );
  AOI21_X1 U18104 ( .B1(n14839), .B2(n14411), .A(n14838), .ZN(n14840) );
  OAI21_X1 U18105 ( .B1(n14841), .B2(n20242), .A(n14840), .ZN(P1_U2989) );
  INV_X1 U18106 ( .A(n14842), .ZN(n14849) );
  INV_X1 U18107 ( .A(n14843), .ZN(n14848) );
  AOI21_X1 U18108 ( .B1(n14846), .B2(n14845), .A(n14844), .ZN(n14847) );
  AOI211_X1 U18109 ( .C1(n14849), .C2(n20404), .A(n14848), .B(n14847), .ZN(
        n14850) );
  OAI21_X1 U18110 ( .B1(n14851), .B2(n20387), .A(n14850), .ZN(P1_U3001) );
  INV_X1 U18111 ( .A(n14852), .ZN(n14853) );
  NOR2_X1 U18112 ( .A1(n14853), .A2(n16211), .ZN(n14854) );
  AOI211_X1 U18113 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14856), .A(
        n14855), .B(n14854), .ZN(n14859) );
  INV_X1 U18114 ( .A(n14874), .ZN(n14869) );
  NAND3_X1 U18115 ( .A1(n14869), .A2(n14866), .A3(n14857), .ZN(n14858) );
  OAI211_X1 U18116 ( .C1(n14860), .C2(n20387), .A(n14859), .B(n14858), .ZN(
        P1_U3002) );
  INV_X1 U18117 ( .A(n14861), .ZN(n14872) );
  NOR2_X1 U18118 ( .A1(n14873), .A2(n14862), .ZN(n14863) );
  AOI211_X1 U18119 ( .C1(n14865), .C2(n20404), .A(n14864), .B(n14863), .ZN(
        n14871) );
  INV_X1 U18120 ( .A(n14866), .ZN(n14867) );
  NAND3_X1 U18121 ( .A1(n14869), .A2(n14868), .A3(n14867), .ZN(n14870) );
  OAI211_X1 U18122 ( .C1(n14872), .C2(n20387), .A(n14871), .B(n14870), .ZN(
        P1_U3003) );
  INV_X1 U18123 ( .A(n14873), .ZN(n14879) );
  NOR2_X1 U18124 ( .A1(n14874), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14878) );
  OAI21_X1 U18125 ( .B1(n14876), .B2(n16211), .A(n14875), .ZN(n14877) );
  AOI211_X1 U18126 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14879), .A(
        n14878), .B(n14877), .ZN(n14880) );
  OAI21_X1 U18127 ( .B1(n14881), .B2(n20387), .A(n14880), .ZN(P1_U3004) );
  NAND2_X1 U18128 ( .A1(n14882), .A2(n20405), .ZN(n14893) );
  AOI21_X1 U18129 ( .B1(n14884), .B2(n20404), .A(n14883), .ZN(n14892) );
  INV_X1 U18130 ( .A(n14919), .ZN(n14886) );
  NOR3_X1 U18131 ( .A1(n14886), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14885), .ZN(n14898) );
  INV_X1 U18132 ( .A(n14887), .ZN(n14900) );
  OAI21_X1 U18133 ( .B1(n14898), .B2(n14900), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14891) );
  NAND3_X1 U18134 ( .A1(n14919), .A2(n14889), .A3(n14888), .ZN(n14890) );
  NAND4_X1 U18135 ( .A1(n14893), .A2(n14892), .A3(n14891), .A4(n14890), .ZN(
        P1_U3005) );
  INV_X1 U18136 ( .A(n14894), .ZN(n14902) );
  INV_X1 U18137 ( .A(n14895), .ZN(n14896) );
  OAI21_X1 U18138 ( .B1(n14897), .B2(n16211), .A(n14896), .ZN(n14899) );
  AOI211_X1 U18139 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n14900), .A(
        n14899), .B(n14898), .ZN(n14901) );
  OAI21_X1 U18140 ( .B1(n14902), .B2(n20387), .A(n14901), .ZN(P1_U3006) );
  INV_X1 U18141 ( .A(n14903), .ZN(n16181) );
  OAI21_X1 U18142 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16181), .A(
        n14904), .ZN(n14908) );
  NOR2_X1 U18143 ( .A1(n14905), .A2(n16211), .ZN(n14906) );
  AOI211_X1 U18144 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14908), .A(
        n14907), .B(n14906), .ZN(n14911) );
  NAND3_X1 U18145 ( .A1(n14919), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14909), .ZN(n14910) );
  OAI211_X1 U18146 ( .C1(n14912), .C2(n20387), .A(n14911), .B(n14910), .ZN(
        P1_U3007) );
  NAND2_X1 U18147 ( .A1(n14913), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14914) );
  OAI211_X1 U18148 ( .C1(n14916), .C2(n16211), .A(n14915), .B(n14914), .ZN(
        n14917) );
  AOI21_X1 U18149 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  OAI21_X1 U18150 ( .B1(n14921), .B2(n20387), .A(n14920), .ZN(P1_U3008) );
  NOR2_X1 U18151 ( .A1(n14922), .A2(n16211), .ZN(n14923) );
  AOI211_X1 U18152 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n14929), .A(
        n14924), .B(n14923), .ZN(n14927) );
  XNOR2_X1 U18153 ( .A(n14933), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14925) );
  NAND2_X1 U18154 ( .A1(n14934), .A2(n14925), .ZN(n14926) );
  OAI211_X1 U18155 ( .C1(n14928), .C2(n20387), .A(n14927), .B(n14926), .ZN(
        P1_U3009) );
  NAND2_X1 U18156 ( .A1(n14929), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14930) );
  OAI211_X1 U18157 ( .C1(n16013), .C2(n16211), .A(n14931), .B(n14930), .ZN(
        n14932) );
  AOI21_X1 U18158 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(n14935) );
  OAI21_X1 U18159 ( .B1(n14936), .B2(n20387), .A(n14935), .ZN(P1_U3010) );
  INV_X1 U18160 ( .A(n14937), .ZN(n14954) );
  NOR2_X1 U18161 ( .A1(n20398), .A2(n14938), .ZN(n14940) );
  OAI21_X1 U18162 ( .B1(n16127), .B2(n20398), .A(n14939), .ZN(n16130) );
  AOI211_X1 U18163 ( .C1(n14941), .C2(n20396), .A(n14940), .B(n16130), .ZN(
        n16120) );
  INV_X1 U18164 ( .A(n14942), .ZN(n14943) );
  AOI22_X1 U18165 ( .A1(n14943), .A2(n16168), .B1(n16127), .B2(n16180), .ZN(
        n14959) );
  INV_X1 U18166 ( .A(n14959), .ZN(n14945) );
  OAI21_X1 U18167 ( .B1(n14945), .B2(n14956), .A(n14944), .ZN(n14946) );
  AOI21_X1 U18168 ( .B1(n16120), .B2(n14946), .A(n14950), .ZN(n14947) );
  AOI211_X1 U18169 ( .C1(n20404), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        n14953) );
  INV_X1 U18170 ( .A(n16126), .ZN(n14951) );
  NAND3_X1 U18171 ( .A1(n14951), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14950), .ZN(n14952) );
  OAI211_X1 U18172 ( .C1(n14954), .C2(n20387), .A(n14953), .B(n14952), .ZN(
        P1_U3011) );
  INV_X1 U18173 ( .A(n16234), .ZN(n16201) );
  NAND3_X1 U18174 ( .A1(n16127), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n14331), .ZN(n14967) );
  NAND2_X1 U18175 ( .A1(n14955), .A2(n20405), .ZN(n14966) );
  NAND2_X1 U18176 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16168), .ZN(
        n16132) );
  AND2_X1 U18177 ( .A1(n14956), .A2(n16132), .ZN(n16167) );
  AOI211_X1 U18178 ( .C1(n14958), .C2(n14957), .A(n16167), .B(n16130), .ZN(
        n16174) );
  NOR2_X1 U18179 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14959), .ZN(
        n16165) );
  INV_X1 U18180 ( .A(n16165), .ZN(n14960) );
  AOI21_X1 U18181 ( .B1(n16174), .B2(n14960), .A(n14331), .ZN(n14964) );
  OR2_X1 U18182 ( .A1(n16210), .A2(n21350), .ZN(n14961) );
  OAI21_X1 U18183 ( .B1(n16211), .B2(n14962), .A(n14961), .ZN(n14963) );
  NOR2_X1 U18184 ( .A1(n14964), .A2(n14963), .ZN(n14965) );
  OAI211_X1 U18185 ( .C1(n16201), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        P1_U3017) );
  NOR2_X1 U18186 ( .A1(n13316), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14969) );
  OAI22_X1 U18187 ( .A1(n20808), .A2(n14969), .B1(n20932), .B2(n14968), .ZN(
        n14970) );
  MUX2_X1 U18188 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14970), .S(
        n20413), .Z(P1_U3477) );
  INV_X1 U18189 ( .A(n14971), .ZN(n14977) );
  NAND3_X1 U18190 ( .A1(n14972), .A2(n14978), .A3(n14977), .ZN(n14973) );
  OAI211_X1 U18191 ( .C1(n20932), .C2(n14975), .A(n14974), .B(n14973), .ZN(
        n15951) );
  NAND2_X1 U18192 ( .A1(n15951), .A2(n16242), .ZN(n14980) );
  NAND3_X1 U18193 ( .A1(n14978), .A2(n14977), .A3(n14976), .ZN(n14979) );
  OAI211_X1 U18194 ( .C1(n14982), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n14983) );
  MUX2_X1 U18195 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14983), .S(
        n16245), .Z(P1_U3473) );
  INV_X1 U18196 ( .A(n14984), .ZN(n14988) );
  OAI22_X1 U18197 ( .A1(n14988), .A2(n14987), .B1(n14986), .B2(n14985), .ZN(
        n14989) );
  MUX2_X1 U18198 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14989), .S(
        n16245), .Z(P1_U3469) );
  INV_X1 U18199 ( .A(n19356), .ZN(n19312) );
  NAND2_X1 U18200 ( .A1(n15010), .A2(n14990), .ZN(n14991) );
  XNOR2_X1 U18201 ( .A(n14992), .B(n14991), .ZN(n14993) );
  NAND2_X1 U18202 ( .A1(n14993), .A2(n19303), .ZN(n15003) );
  OAI22_X1 U18203 ( .A1(n19343), .A2(n14996), .B1(n14995), .B2(n19353), .ZN(
        n14998) );
  NOR2_X1 U18204 ( .A1(n19342), .A2(n13568), .ZN(n14997) );
  AOI211_X1 U18205 ( .C1(n19333), .C2(n20166), .A(n14998), .B(n14997), .ZN(
        n14999) );
  OAI21_X1 U18206 ( .B1(n15000), .B2(n19328), .A(n14999), .ZN(n15001) );
  AOI21_X1 U18207 ( .B1(n14994), .B2(n19290), .A(n15001), .ZN(n15002) );
  OAI211_X1 U18208 ( .C1(n19583), .C2(n19312), .A(n15003), .B(n15002), .ZN(
        P2_U2852) );
  INV_X1 U18209 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n15007) );
  NAND2_X1 U18210 ( .A1(n19346), .A2(n15004), .ZN(n15006) );
  AOI22_X1 U18211 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19324), .ZN(n15005) );
  OAI211_X1 U18212 ( .C1(n15007), .C2(n19342), .A(n15006), .B(n15005), .ZN(
        n15008) );
  AOI21_X1 U18213 ( .B1(n20179), .B2(n19333), .A(n15008), .ZN(n15009) );
  OAI21_X1 U18214 ( .B1(n13468), .B2(n19349), .A(n15009), .ZN(n15015) );
  INV_X1 U18215 ( .A(n19502), .ZN(n15013) );
  NOR2_X1 U18216 ( .A1(n19315), .A2(n15011), .ZN(n15658) );
  INV_X1 U18217 ( .A(n15658), .ZN(n15012) );
  AOI221_X1 U18218 ( .B1(n15013), .B2(n15658), .C1(n19502), .C2(n15012), .A(
        n19339), .ZN(n15014) );
  AOI211_X1 U18219 ( .C1(n20174), .C2(n19356), .A(n15015), .B(n15014), .ZN(
        n15016) );
  INV_X1 U18220 ( .A(n15016), .ZN(P2_U2853) );
  MUX2_X1 U18221 ( .A(n16263), .B(P2_EBX_REG_31__SCAN_IN), .S(n9831), .Z(
        P2_U2856) );
  OR2_X1 U18222 ( .A1(n15021), .A2(n15020), .ZN(n15124) );
  NAND3_X1 U18223 ( .A1(n15124), .A2(n15022), .A3(n15110), .ZN(n15024) );
  NAND2_X1 U18224 ( .A1(n9831), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15023) );
  OAI211_X1 U18225 ( .C1(n9831), .C2(n16288), .A(n15024), .B(n15023), .ZN(
        P2_U2858) );
  NOR2_X1 U18226 ( .A1(n15026), .A2(n15025), .ZN(n15028) );
  XNOR2_X1 U18227 ( .A(n15028), .B(n15027), .ZN(n15136) );
  NAND2_X1 U18228 ( .A1(n15136), .A2(n15110), .ZN(n15030) );
  NAND2_X1 U18229 ( .A1(n9831), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15029) );
  OAI211_X1 U18230 ( .C1(n9831), .C2(n15031), .A(n15030), .B(n15029), .ZN(
        P2_U2859) );
  OAI21_X1 U18231 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15150) );
  INV_X1 U18232 ( .A(n14255), .ZN(n15035) );
  OAI21_X1 U18233 ( .B1(n15041), .B2(n15036), .A(n15035), .ZN(n16309) );
  NOR2_X1 U18234 ( .A1(n16309), .A2(n9831), .ZN(n15037) );
  AOI21_X1 U18235 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9831), .A(n15037), .ZN(
        n15038) );
  OAI21_X1 U18236 ( .B1(n15150), .B2(n15106), .A(n15038), .ZN(P2_U2860) );
  NOR2_X1 U18237 ( .A1(n15052), .A2(n15039), .ZN(n15040) );
  OR2_X1 U18238 ( .A1(n15041), .A2(n15040), .ZN(n15247) );
  AOI21_X1 U18239 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15157) );
  NAND2_X1 U18240 ( .A1(n15157), .A2(n15110), .ZN(n15046) );
  NAND2_X1 U18241 ( .A1(n9831), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15045) );
  OAI211_X1 U18242 ( .C1(n9831), .C2(n15247), .A(n15046), .B(n15045), .ZN(
        P2_U2861) );
  OAI21_X1 U18243 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15159) );
  NOR2_X1 U18244 ( .A1(n15061), .A2(n15050), .ZN(n15051) );
  OR2_X1 U18245 ( .A1(n15052), .A2(n15051), .ZN(n16332) );
  NOR2_X1 U18246 ( .A1(n16332), .A2(n9831), .ZN(n15053) );
  AOI21_X1 U18247 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n9831), .A(n15053), .ZN(
        n15054) );
  OAI21_X1 U18248 ( .B1(n15159), .B2(n15106), .A(n15054), .ZN(P2_U2862) );
  AOI21_X1 U18249 ( .B1(n15056), .B2(n15055), .A(n9905), .ZN(n15057) );
  XOR2_X1 U18250 ( .A(n15058), .B(n15057), .Z(n15175) );
  NOR2_X1 U18251 ( .A1(n15070), .A2(n15059), .ZN(n15060) );
  OR2_X1 U18252 ( .A1(n15061), .A2(n15060), .ZN(n15275) );
  NOR2_X1 U18253 ( .A1(n15275), .A2(n9831), .ZN(n15062) );
  AOI21_X1 U18254 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n9831), .A(n15062), .ZN(
        n15063) );
  OAI21_X1 U18255 ( .B1(n15175), .B2(n15106), .A(n15063), .ZN(P2_U2863) );
  NOR2_X1 U18256 ( .A1(n15065), .A2(n15064), .ZN(n15066) );
  NOR2_X1 U18257 ( .A1(n15066), .A2(n9891), .ZN(n16357) );
  NAND2_X1 U18258 ( .A1(n16357), .A2(n15110), .ZN(n15073) );
  NOR2_X1 U18259 ( .A1(n15067), .A2(n15068), .ZN(n15069) );
  OR2_X1 U18260 ( .A1(n15070), .A2(n15069), .ZN(n16354) );
  INV_X1 U18261 ( .A(n16354), .ZN(n15071) );
  NAND2_X1 U18262 ( .A1(n15071), .A2(n15104), .ZN(n15072) );
  OAI211_X1 U18263 ( .C1(n15104), .C2(n15074), .A(n15073), .B(n15072), .ZN(
        P2_U2864) );
  NAND2_X1 U18264 ( .A1(n15083), .A2(n15075), .ZN(n15086) );
  AOI21_X1 U18265 ( .B1(n15077), .B2(n15086), .A(n15076), .ZN(n15183) );
  NAND2_X1 U18266 ( .A1(n15183), .A2(n15110), .ZN(n15081) );
  NOR2_X1 U18267 ( .A1(n15088), .A2(n15078), .ZN(n15079) );
  NOR2_X1 U18268 ( .A1(n15067), .A2(n15079), .ZN(n16364) );
  NAND2_X1 U18269 ( .A1(n16364), .A2(n15104), .ZN(n15080) );
  OAI211_X1 U18270 ( .C1(n15104), .C2(n14180), .A(n15081), .B(n15080), .ZN(
        P2_U2865) );
  AND2_X1 U18271 ( .A1(n15083), .A2(n15082), .ZN(n15085) );
  AND2_X1 U18272 ( .A1(n15085), .A2(n15084), .ZN(n15095) );
  OAI21_X1 U18273 ( .B1(n15095), .B2(n15087), .A(n15086), .ZN(n15197) );
  INV_X1 U18274 ( .A(n15088), .ZN(n15093) );
  INV_X1 U18275 ( .A(n15100), .ZN(n15091) );
  INV_X1 U18276 ( .A(n15089), .ZN(n15090) );
  NAND2_X1 U18277 ( .A1(n15091), .A2(n15090), .ZN(n15092) );
  NAND2_X1 U18278 ( .A1(n15093), .A2(n15092), .ZN(n19138) );
  MUX2_X1 U18279 ( .A(n14130), .B(n19138), .S(n15104), .Z(n15094) );
  OAI21_X1 U18280 ( .B1(n15197), .B2(n15106), .A(n15094), .ZN(P2_U2866) );
  INV_X1 U18281 ( .A(n15095), .ZN(n15096) );
  OAI21_X1 U18282 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15207) );
  INV_X1 U18283 ( .A(n15099), .ZN(n15102) );
  INV_X1 U18284 ( .A(n13992), .ZN(n15101) );
  AOI21_X1 U18285 ( .B1(n15102), .B2(n15101), .A(n15100), .ZN(n19148) );
  NOR2_X1 U18286 ( .A1(n15104), .A2(n14129), .ZN(n15103) );
  AOI21_X1 U18287 ( .B1(n19148), .B2(n15104), .A(n15103), .ZN(n15105) );
  OAI21_X1 U18288 ( .B1(n15207), .B2(n15106), .A(n15105), .ZN(P2_U2867) );
  AOI21_X1 U18289 ( .B1(n15109), .B2(n15108), .A(n15107), .ZN(n15214) );
  NAND2_X1 U18290 ( .A1(n15214), .A2(n15110), .ZN(n15116) );
  INV_X1 U18291 ( .A(n15111), .ZN(n15114) );
  INV_X1 U18292 ( .A(n13982), .ZN(n15113) );
  AOI21_X1 U18293 ( .B1(n15114), .B2(n15113), .A(n15112), .ZN(n19169) );
  NAND2_X1 U18294 ( .A1(n19169), .A2(n15104), .ZN(n15115) );
  OAI211_X1 U18295 ( .C1(n15104), .C2(n11175), .A(n15116), .B(n15115), .ZN(
        P2_U2869) );
  NAND2_X1 U18296 ( .A1(n15125), .A2(BUF2_REG_14__SCAN_IN), .ZN(n15119) );
  OR2_X1 U18297 ( .A1(n15125), .A2(n16656), .ZN(n15118) );
  NAND2_X1 U18298 ( .A1(n15119), .A2(n15118), .ZN(n19480) );
  AOI22_X1 U18299 ( .A1(n19367), .A2(n19480), .B1(n19427), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U18300 ( .A1(n19360), .A2(BUF2_REG_30__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U18301 ( .A1(n16268), .A2(n19428), .ZN(n15121) );
  NAND3_X1 U18302 ( .A1(n15124), .A2(n15022), .A3(n19429), .ZN(n15135) );
  NAND2_X1 U18303 ( .A1(n15125), .A2(BUF2_REG_13__SCAN_IN), .ZN(n15127) );
  OR2_X1 U18304 ( .A1(n15125), .A2(n16658), .ZN(n15126) );
  NAND2_X1 U18305 ( .A1(n15127), .A2(n15126), .ZN(n19478) );
  AOI22_X1 U18306 ( .A1(n19367), .A2(n19478), .B1(n19427), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15134) );
  AOI22_X1 U18307 ( .A1(n19360), .A2(BUF2_REG_29__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15133) );
  INV_X1 U18308 ( .A(n15128), .ZN(n15129) );
  AOI21_X1 U18309 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n16282) );
  NAND2_X1 U18310 ( .A1(n16282), .A2(n19428), .ZN(n15132) );
  NAND4_X1 U18311 ( .A1(n15135), .A2(n15134), .A3(n15133), .A4(n15132), .ZN(
        P2_U2890) );
  NAND2_X1 U18312 ( .A1(n15136), .A2(n19429), .ZN(n15141) );
  AOI22_X1 U18313 ( .A1(n19367), .A2(n15137), .B1(n19427), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15140) );
  AOI22_X1 U18314 ( .A1(n19360), .A2(BUF2_REG_28__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15139) );
  NAND2_X1 U18315 ( .A1(n19428), .A2(n16290), .ZN(n15138) );
  NAND4_X1 U18316 ( .A1(n15141), .A2(n15140), .A3(n15139), .A4(n15138), .ZN(
        P2_U2891) );
  NOR2_X1 U18317 ( .A1(n15142), .A2(n15143), .ZN(n15144) );
  OR2_X1 U18318 ( .A1(n15145), .A2(n15144), .ZN(n15390) );
  AOI22_X1 U18319 ( .A1(n19360), .A2(BUF2_REG_27__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15147) );
  AOI22_X1 U18320 ( .A1(n19367), .A2(n19379), .B1(n19427), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15146) );
  OAI211_X1 U18321 ( .C1(n19365), .C2(n15390), .A(n15147), .B(n15146), .ZN(
        n15148) );
  INV_X1 U18322 ( .A(n15148), .ZN(n15149) );
  OAI21_X1 U18323 ( .B1(n15150), .B2(n19366), .A(n15149), .ZN(P2_U2892) );
  NOR2_X1 U18324 ( .A1(n15162), .A2(n15151), .ZN(n15152) );
  OR2_X1 U18325 ( .A1(n15142), .A2(n15152), .ZN(n16320) );
  AOI22_X1 U18326 ( .A1(n19360), .A2(BUF2_REG_26__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15155) );
  AOI22_X1 U18327 ( .A1(n19367), .A2(n15153), .B1(n19427), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15154) );
  OAI211_X1 U18328 ( .C1(n19365), .C2(n16320), .A(n15155), .B(n15154), .ZN(
        n15156) );
  AOI21_X1 U18329 ( .B1(n15157), .B2(n19429), .A(n15156), .ZN(n15158) );
  INV_X1 U18330 ( .A(n15158), .ZN(P2_U2893) );
  OR2_X1 U18331 ( .A1(n15159), .A2(n19366), .ZN(n15166) );
  AOI22_X1 U18332 ( .A1(n19367), .A2(n19385), .B1(n19427), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U18333 ( .A1(n19360), .A2(BUF2_REG_25__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15164) );
  AND2_X1 U18334 ( .A1(n15169), .A2(n15160), .ZN(n15161) );
  NOR2_X1 U18335 ( .A1(n15162), .A2(n15161), .ZN(n16326) );
  NAND2_X1 U18336 ( .A1(n19428), .A2(n16326), .ZN(n15163) );
  NAND4_X1 U18337 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        P2_U2894) );
  NAND2_X1 U18338 ( .A1(n15441), .A2(n15167), .ZN(n15168) );
  NAND2_X1 U18339 ( .A1(n15169), .A2(n15168), .ZN(n16335) );
  AOI22_X1 U18340 ( .A1(n19360), .A2(BUF2_REG_24__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15172) );
  AOI22_X1 U18341 ( .A1(n19367), .A2(n15170), .B1(n19427), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15171) );
  OAI211_X1 U18342 ( .C1(n19365), .C2(n16335), .A(n15172), .B(n15171), .ZN(
        n15173) );
  INV_X1 U18343 ( .A(n15173), .ZN(n15174) );
  OAI21_X1 U18344 ( .B1(n15175), .B2(n19366), .A(n15174), .ZN(P2_U2895) );
  NOR2_X1 U18345 ( .A1(n15177), .A2(n15176), .ZN(n15178) );
  OR2_X1 U18346 ( .A1(n15439), .A2(n15178), .ZN(n15945) );
  AOI22_X1 U18347 ( .A1(n19360), .A2(BUF2_REG_22__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15181) );
  AOI22_X1 U18348 ( .A1(n19367), .A2(n15179), .B1(n19427), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15180) );
  OAI211_X1 U18349 ( .C1(n19365), .C2(n15945), .A(n15181), .B(n15180), .ZN(
        n15182) );
  AOI21_X1 U18350 ( .B1(n15183), .B2(n19429), .A(n15182), .ZN(n15184) );
  INV_X1 U18351 ( .A(n15184), .ZN(P2_U2897) );
  INV_X1 U18352 ( .A(n15200), .ZN(n15185) );
  XNOR2_X1 U18353 ( .A(n15186), .B(n15185), .ZN(n19132) );
  NAND2_X1 U18354 ( .A1(n19367), .A2(n15187), .ZN(n15188) );
  OAI21_X1 U18355 ( .B1(n19391), .B2(n15189), .A(n15188), .ZN(n15195) );
  INV_X1 U18356 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15192) );
  INV_X1 U18357 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15190) );
  OAI22_X1 U18358 ( .A1(n15193), .A2(n15192), .B1(n15191), .B2(n15190), .ZN(
        n15194) );
  AOI211_X1 U18359 ( .C1(n19428), .C2(n19132), .A(n15195), .B(n15194), .ZN(
        n15196) );
  OAI21_X1 U18360 ( .B1(n15197), .B2(n19366), .A(n15196), .ZN(P2_U2898) );
  OR2_X1 U18361 ( .A1(n15199), .A2(n15198), .ZN(n15201) );
  NAND2_X1 U18362 ( .A1(n15201), .A2(n15200), .ZN(n19151) );
  AOI22_X1 U18363 ( .A1(n19360), .A2(BUF2_REG_20__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U18364 ( .A1(n19367), .A2(n15202), .B1(n19427), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15203) );
  OAI211_X1 U18365 ( .C1(n19365), .C2(n19151), .A(n15204), .B(n15203), .ZN(
        n15205) );
  INV_X1 U18366 ( .A(n15205), .ZN(n15206) );
  OAI21_X1 U18367 ( .B1(n15207), .B2(n19366), .A(n15206), .ZN(P2_U2899) );
  NOR2_X1 U18368 ( .A1(n15208), .A2(n9939), .ZN(n15209) );
  OR2_X1 U18369 ( .A1(n14023), .A2(n15209), .ZN(n19172) );
  AOI22_X1 U18370 ( .A1(n19360), .A2(BUF2_REG_18__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15212) );
  AOI22_X1 U18371 ( .A1(n19367), .A2(n15210), .B1(n19427), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15211) );
  OAI211_X1 U18372 ( .C1(n19365), .C2(n19172), .A(n15212), .B(n15211), .ZN(
        n15213) );
  AOI21_X1 U18373 ( .B1(n15214), .B2(n19429), .A(n15213), .ZN(n15215) );
  INV_X1 U18374 ( .A(n15215), .ZN(P2_U2901) );
  NAND2_X1 U18375 ( .A1(n9897), .A2(n15216), .ZN(n15217) );
  XNOR2_X1 U18376 ( .A(n15218), .B(n15217), .ZN(n15375) );
  XNOR2_X1 U18377 ( .A(n15223), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15372) );
  XNOR2_X1 U18378 ( .A(n15229), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16272) );
  NAND2_X1 U18379 ( .A1(n16269), .A2(n19510), .ZN(n15220) );
  INV_X1 U18380 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20147) );
  NOR2_X1 U18381 ( .A1(n19294), .A2(n20147), .ZN(n15366) );
  AOI21_X1 U18382 ( .B1(n19490), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15366), .ZN(n15219) );
  OAI211_X1 U18383 ( .C1(n19503), .C2(n16272), .A(n15220), .B(n15219), .ZN(
        n15221) );
  AOI21_X1 U18384 ( .B1(n15372), .B2(n16449), .A(n15221), .ZN(n15222) );
  OAI21_X1 U18385 ( .B1(n15375), .B2(n19493), .A(n15222), .ZN(P2_U2984) );
  OAI21_X1 U18386 ( .B1(n9880), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15223), .ZN(n15388) );
  NAND2_X1 U18387 ( .A1(n10370), .A2(n15225), .ZN(n15226) );
  XNOR2_X1 U18388 ( .A(n15227), .B(n15226), .ZN(n15376) );
  NAND2_X1 U18389 ( .A1(n15376), .A2(n19504), .ZN(n15234) );
  INV_X1 U18390 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16277) );
  INV_X1 U18391 ( .A(n15228), .ZN(n15230) );
  AOI21_X1 U18392 ( .B1(n16277), .B2(n15230), .A(n15229), .ZN(n16254) );
  NAND2_X1 U18393 ( .A1(n19310), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15378) );
  OAI21_X1 U18394 ( .B1(n19514), .B2(n16277), .A(n15378), .ZN(n15232) );
  NOR2_X1 U18395 ( .A1(n16288), .A2(n16438), .ZN(n15231) );
  AOI211_X1 U18396 ( .C1(n16442), .C2(n16254), .A(n15232), .B(n15231), .ZN(
        n15233) );
  OAI211_X1 U18397 ( .C1(n19501), .C2(n15388), .A(n15234), .B(n15233), .ZN(
        P2_U2985) );
  XNOR2_X1 U18398 ( .A(n15235), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15399) );
  INV_X1 U18399 ( .A(n16309), .ZN(n15241) );
  OAI21_X1 U18400 ( .B1(n15248), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15236), .ZN(n16306) );
  AND2_X1 U18401 ( .A1(n19310), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15391) );
  AOI21_X1 U18402 ( .B1(n19490), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15391), .ZN(n15237) );
  OAI21_X1 U18403 ( .B1(n19503), .B2(n16306), .A(n15237), .ZN(n15240) );
  OAI21_X1 U18404 ( .B1(n15254), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15238), .ZN(n15394) );
  NOR2_X1 U18405 ( .A1(n15394), .A2(n19501), .ZN(n15239) );
  AOI211_X1 U18406 ( .C1(n19510), .C2(n15241), .A(n15240), .B(n15239), .ZN(
        n15242) );
  OAI21_X1 U18407 ( .B1(n15399), .B2(n19493), .A(n15242), .ZN(P2_U2987) );
  AOI21_X1 U18408 ( .B1(n15266), .B2(n10203), .A(n15263), .ZN(n15244) );
  MUX2_X1 U18409 ( .A(n10203), .B(n15244), .S(n15243), .Z(n15245) );
  NAND2_X1 U18410 ( .A1(n15246), .A2(n15245), .ZN(n15412) );
  INV_X1 U18411 ( .A(n15247), .ZN(n16314) );
  INV_X1 U18412 ( .A(n15248), .ZN(n15252) );
  INV_X1 U18413 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15250) );
  INV_X1 U18414 ( .A(n15267), .ZN(n15249) );
  NAND2_X1 U18415 ( .A1(n15250), .A2(n15249), .ZN(n15251) );
  NAND2_X1 U18416 ( .A1(n15252), .A2(n15251), .ZN(n16317) );
  NAND2_X1 U18417 ( .A1(n19310), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15402) );
  NAND2_X1 U18418 ( .A1(n19490), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15253) );
  OAI211_X1 U18419 ( .C1(n19503), .C2(n16317), .A(n15402), .B(n15253), .ZN(
        n15259) );
  INV_X1 U18420 ( .A(n15254), .ZN(n15257) );
  INV_X1 U18421 ( .A(n15280), .ZN(n15262) );
  NAND2_X1 U18422 ( .A1(n15262), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15261) );
  NAND2_X1 U18423 ( .A1(n15261), .A2(n15255), .ZN(n15256) );
  NAND2_X1 U18424 ( .A1(n15257), .A2(n15256), .ZN(n15409) );
  NOR2_X1 U18425 ( .A1(n15409), .A2(n19501), .ZN(n15258) );
  OAI21_X1 U18426 ( .B1(n15412), .B2(n19493), .A(n15260), .ZN(P2_U2988) );
  OAI21_X1 U18427 ( .B1(n15262), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15261), .ZN(n15422) );
  NOR2_X1 U18428 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  XNOR2_X1 U18429 ( .A(n15266), .B(n15265), .ZN(n15413) );
  NAND2_X1 U18430 ( .A1(n15413), .A2(n19504), .ZN(n15271) );
  AOI21_X1 U18431 ( .B1(n16321), .B2(n15276), .A(n15267), .ZN(n16255) );
  NAND2_X1 U18432 ( .A1(n19310), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15415) );
  OAI21_X1 U18433 ( .B1(n19514), .B2(n16321), .A(n15415), .ZN(n15269) );
  NOR2_X1 U18434 ( .A1(n16332), .A2(n16438), .ZN(n15268) );
  AOI211_X1 U18435 ( .C1(n16442), .C2(n16255), .A(n15269), .B(n15268), .ZN(
        n15270) );
  OAI211_X1 U18436 ( .C1(n19501), .C2(n15422), .A(n15271), .B(n15270), .ZN(
        P2_U2989) );
  XNOR2_X1 U18437 ( .A(n15272), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15273) );
  XNOR2_X1 U18438 ( .A(n15274), .B(n15273), .ZN(n15432) );
  INV_X1 U18439 ( .A(n15275), .ZN(n16337) );
  OAI21_X1 U18440 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n9947), .A(
        n15276), .ZN(n16340) );
  NAND2_X1 U18441 ( .A1(n19310), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U18442 ( .A1(n19490), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15277) );
  OAI211_X1 U18443 ( .C1(n19503), .C2(n16340), .A(n15423), .B(n15277), .ZN(
        n15282) );
  NAND2_X1 U18444 ( .A1(n15284), .A2(n15278), .ZN(n15279) );
  NAND2_X1 U18445 ( .A1(n15280), .A2(n15279), .ZN(n15427) );
  NOR2_X1 U18446 ( .A1(n15427), .A2(n19501), .ZN(n15281) );
  AOI211_X1 U18447 ( .C1(n16337), .C2(n19510), .A(n15282), .B(n15281), .ZN(
        n15283) );
  OAI21_X1 U18448 ( .B1(n15432), .B2(n19493), .A(n15283), .ZN(P2_U2990) );
  OAI21_X1 U18449 ( .B1(n15454), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15284), .ZN(n15434) );
  XOR2_X1 U18450 ( .A(n15286), .B(n15285), .Z(n15433) );
  NAND2_X1 U18451 ( .A1(n15433), .A2(n19504), .ZN(n15291) );
  AOI21_X1 U18452 ( .B1(n16345), .B2(n15934), .A(n9947), .ZN(n16256) );
  INV_X1 U18453 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n15287) );
  OAI22_X1 U18454 ( .A1(n19514), .A2(n16345), .B1(n15287), .B2(n19294), .ZN(
        n15289) );
  NOR2_X1 U18455 ( .A1(n16354), .A2(n16438), .ZN(n15288) );
  AOI211_X1 U18456 ( .C1(n16442), .C2(n16256), .A(n15289), .B(n15288), .ZN(
        n15290) );
  OAI211_X1 U18457 ( .C1(n19501), .C2(n15434), .A(n15291), .B(n15290), .ZN(
        P2_U2991) );
  INV_X1 U18458 ( .A(n15292), .ZN(n15293) );
  NAND2_X1 U18459 ( .A1(n15293), .A2(n15581), .ZN(n15558) );
  NAND2_X1 U18460 ( .A1(n15558), .A2(n15557), .ZN(n15540) );
  INV_X1 U18461 ( .A(n15539), .ZN(n15294) );
  AOI21_X1 U18462 ( .B1(n15540), .B2(n15295), .A(n15294), .ZN(n15359) );
  NAND2_X1 U18463 ( .A1(n15359), .A2(n15358), .ZN(n15357) );
  NAND2_X1 U18464 ( .A1(n15357), .A2(n15296), .ZN(n15347) );
  NAND2_X1 U18465 ( .A1(n15298), .A2(n15297), .ZN(n15348) );
  INV_X1 U18466 ( .A(n15303), .ZN(n15301) );
  NOR2_X1 U18467 ( .A1(n15302), .A2(n15301), .ZN(n15315) );
  NAND2_X1 U18468 ( .A1(n15316), .A2(n15315), .ZN(n15314) );
  NAND2_X1 U18469 ( .A1(n15314), .A2(n15303), .ZN(n15308) );
  INV_X1 U18470 ( .A(n15304), .ZN(n15305) );
  NOR2_X1 U18471 ( .A1(n15306), .A2(n15305), .ZN(n15307) );
  XNOR2_X1 U18472 ( .A(n15308), .B(n15307), .ZN(n15476) );
  INV_X1 U18473 ( .A(n15320), .ZN(n15309) );
  AOI21_X1 U18474 ( .B1(n15465), .B2(n15309), .A(n15452), .ZN(n15474) );
  AOI21_X1 U18475 ( .B1(n19127), .B2(n15317), .A(n15935), .ZN(n15936) );
  NAND2_X1 U18476 ( .A1(n19310), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15467) );
  OAI21_X1 U18477 ( .B1(n19514), .B2(n19127), .A(n15467), .ZN(n15310) );
  AOI21_X1 U18478 ( .B1(n16442), .B2(n15936), .A(n15310), .ZN(n15311) );
  OAI21_X1 U18479 ( .B1(n19138), .B2(n16438), .A(n15311), .ZN(n15312) );
  AOI21_X1 U18480 ( .B1(n15474), .B2(n16449), .A(n15312), .ZN(n15313) );
  OAI21_X1 U18481 ( .B1(n15476), .B2(n19493), .A(n15313), .ZN(P2_U2993) );
  OAI21_X1 U18482 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(n15487) );
  OAI21_X1 U18483 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15330), .A(
        n15317), .ZN(n19143) );
  NAND2_X1 U18484 ( .A1(n19310), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15480) );
  NAND2_X1 U18485 ( .A1(n19490), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15318) );
  OAI211_X1 U18486 ( .C1(n19503), .C2(n19143), .A(n15480), .B(n15318), .ZN(
        n15319) );
  AOI21_X1 U18487 ( .B1(n19148), .B2(n19510), .A(n15319), .ZN(n15322) );
  AOI21_X1 U18488 ( .B1(n15479), .B2(n15324), .A(n15320), .ZN(n15484) );
  NAND2_X1 U18489 ( .A1(n15484), .A2(n16449), .ZN(n15321) );
  OAI211_X1 U18490 ( .C1(n15487), .C2(n19493), .A(n15322), .B(n15321), .ZN(
        P2_U2994) );
  NAND2_X1 U18491 ( .A1(n15343), .A2(n15478), .ZN(n15323) );
  NAND2_X1 U18492 ( .A1(n15324), .A2(n15323), .ZN(n15497) );
  INV_X1 U18493 ( .A(n15337), .ZN(n15325) );
  AOI21_X1 U18494 ( .B1(n15339), .B2(n15336), .A(n15325), .ZN(n15329) );
  NAND2_X1 U18495 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  XNOR2_X1 U18496 ( .A(n15329), .B(n15328), .ZN(n15488) );
  NAND2_X1 U18497 ( .A1(n15488), .A2(n19504), .ZN(n15335) );
  AOI21_X1 U18498 ( .B1(n15340), .B2(n15332), .A(n15330), .ZN(n19154) );
  NAND2_X1 U18499 ( .A1(n19154), .A2(n16442), .ZN(n15331) );
  NAND2_X1 U18500 ( .A1(n19310), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15489) );
  OAI211_X1 U18501 ( .C1(n19514), .C2(n15332), .A(n15331), .B(n15489), .ZN(
        n15333) );
  AOI21_X1 U18502 ( .B1(n19159), .B2(n19510), .A(n15333), .ZN(n15334) );
  OAI211_X1 U18503 ( .C1(n19501), .C2(n15497), .A(n15335), .B(n15334), .ZN(
        P2_U2995) );
  NAND2_X1 U18504 ( .A1(n15337), .A2(n15336), .ZN(n15338) );
  XNOR2_X1 U18505 ( .A(n15339), .B(n15338), .ZN(n15511) );
  OAI21_X1 U18506 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15349), .A(
        n15340), .ZN(n19167) );
  NAND2_X1 U18507 ( .A1(n19310), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U18508 ( .A1(n19490), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15341) );
  OAI211_X1 U18509 ( .C1(n19167), .C2(n19503), .A(n15498), .B(n15341), .ZN(
        n15345) );
  INV_X1 U18510 ( .A(n15637), .ZN(n15342) );
  INV_X1 U18511 ( .A(n15499), .ZN(n15516) );
  NOR3_X1 U18512 ( .A1(n15342), .A2(n15516), .A3(n15500), .ZN(n15353) );
  OAI21_X1 U18513 ( .B1(n15353), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15343), .ZN(n15506) );
  NOR2_X1 U18514 ( .A1(n15506), .A2(n19501), .ZN(n15344) );
  AOI211_X1 U18515 ( .C1(n19510), .C2(n19169), .A(n15345), .B(n15344), .ZN(
        n15346) );
  OAI21_X1 U18516 ( .B1(n15511), .B2(n19493), .A(n15346), .ZN(P2_U2996) );
  XOR2_X1 U18517 ( .A(n15348), .B(n15347), .Z(n15527) );
  INV_X1 U18518 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20121) );
  NOR2_X1 U18519 ( .A1(n20121), .A2(n19294), .ZN(n15522) );
  AOI21_X1 U18520 ( .B1(n15350), .B2(n15360), .A(n15349), .ZN(n15941) );
  INV_X1 U18521 ( .A(n15941), .ZN(n19180) );
  OAI22_X1 U18522 ( .A1(n15350), .A2(n19514), .B1(n19503), .B2(n19180), .ZN(
        n15351) );
  AOI211_X1 U18523 ( .C1(n19510), .C2(n19177), .A(n15522), .B(n15351), .ZN(
        n15356) );
  INV_X1 U18524 ( .A(n15569), .ZN(n15352) );
  NAND2_X1 U18525 ( .A1(n15637), .A2(n15352), .ZN(n15578) );
  INV_X1 U18526 ( .A(n15353), .ZN(n15354) );
  OAI211_X1 U18527 ( .C1(n15515), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16449), .B(n15354), .ZN(n15355) );
  OAI211_X1 U18528 ( .C1(n15527), .C2(n19493), .A(n15356), .B(n15355), .ZN(
        P2_U2997) );
  OAI21_X1 U18529 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15537) );
  OAI21_X1 U18530 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9948), .A(
        n15360), .ZN(n19190) );
  AOI22_X1 U18531 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19310), .ZN(n15361) );
  OAI21_X1 U18532 ( .B1(n19503), .B2(n19190), .A(n15361), .ZN(n15362) );
  AOI21_X1 U18533 ( .B1(n19510), .B2(n19193), .A(n15362), .ZN(n15365) );
  INV_X1 U18534 ( .A(n15515), .ZN(n15363) );
  OAI211_X1 U18535 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15543), .A(
        n15363), .B(n16449), .ZN(n15364) );
  OAI211_X1 U18536 ( .C1(n15537), .C2(n19493), .A(n15365), .B(n15364), .ZN(
        P2_U2998) );
  OAI21_X1 U18537 ( .B1(n15620), .B2(n15368), .A(n15389), .ZN(n15371) );
  NAND2_X1 U18538 ( .A1(n15372), .A2(n16493), .ZN(n15373) );
  OAI211_X1 U18539 ( .C1(n15375), .C2(n16477), .A(n15374), .B(n15373), .ZN(
        P2_U3016) );
  NAND2_X1 U18540 ( .A1(n15376), .A2(n16490), .ZN(n15387) );
  NAND2_X1 U18541 ( .A1(n16282), .A2(n16485), .ZN(n15377) );
  OAI211_X1 U18542 ( .C1(n16288), .C2(n15640), .A(n15378), .B(n15377), .ZN(
        n15384) );
  AOI21_X1 U18543 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15382), .A(
        n15381), .ZN(n15380) );
  AOI211_X1 U18544 ( .C1(n15382), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        n15383) );
  AOI211_X1 U18545 ( .C1(n15385), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15384), .B(n15383), .ZN(n15386) );
  OAI211_X1 U18546 ( .C1(n15388), .C2(n16457), .A(n15387), .B(n15386), .ZN(
        P2_U3017) );
  INV_X1 U18547 ( .A(n15389), .ZN(n15397) );
  INV_X1 U18548 ( .A(n15390), .ZN(n16303) );
  AOI21_X1 U18549 ( .B1(n16485), .B2(n16303), .A(n15391), .ZN(n15392) );
  OAI211_X1 U18550 ( .C1(n16309), .C2(n15640), .A(n15393), .B(n15392), .ZN(
        n15396) );
  NOR2_X1 U18551 ( .A1(n15394), .A2(n16457), .ZN(n15395) );
  AOI211_X1 U18552 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15397), .A(
        n15396), .B(n15395), .ZN(n15398) );
  OAI21_X1 U18553 ( .B1(n15399), .B2(n16477), .A(n15398), .ZN(P2_U3019) );
  INV_X1 U18554 ( .A(n15426), .ZN(n15400) );
  NAND2_X1 U18555 ( .A1(n15400), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15416) );
  OAI21_X1 U18556 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15401), .ZN(n15407) );
  INV_X1 U18557 ( .A(n16320), .ZN(n15404) );
  INV_X1 U18558 ( .A(n15402), .ZN(n15403) );
  AOI21_X1 U18559 ( .B1(n16485), .B2(n15404), .A(n15403), .ZN(n15406) );
  NAND2_X1 U18560 ( .A1(n16314), .A2(n16492), .ZN(n15405) );
  OAI211_X1 U18561 ( .C1(n15416), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15408) );
  AOI21_X1 U18562 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15419), .A(
        n15408), .ZN(n15411) );
  OR2_X1 U18563 ( .A1(n15409), .A2(n16457), .ZN(n15410) );
  OAI211_X1 U18564 ( .C1(n15412), .C2(n16477), .A(n15411), .B(n15410), .ZN(
        P2_U3020) );
  NAND2_X1 U18565 ( .A1(n15413), .A2(n16490), .ZN(n15421) );
  NAND2_X1 U18566 ( .A1(n16485), .A2(n16326), .ZN(n15414) );
  OAI211_X1 U18567 ( .C1(n16332), .C2(n15640), .A(n15415), .B(n15414), .ZN(
        n15418) );
  NOR2_X1 U18568 ( .A1(n15416), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15417) );
  AOI211_X1 U18569 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15419), .A(
        n15418), .B(n15417), .ZN(n15420) );
  OAI211_X1 U18570 ( .C1(n15422), .C2(n16457), .A(n15421), .B(n15420), .ZN(
        P2_U3021) );
  OAI21_X1 U18571 ( .B1(n16469), .B2(n16335), .A(n15423), .ZN(n15424) );
  AOI21_X1 U18572 ( .B1(n16337), .B2(n16492), .A(n15424), .ZN(n15425) );
  OAI21_X1 U18573 ( .B1(n15426), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15425), .ZN(n15429) );
  NOR2_X1 U18574 ( .A1(n15427), .A2(n16457), .ZN(n15428) );
  AOI211_X1 U18575 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15430), .A(
        n15429), .B(n15428), .ZN(n15431) );
  OAI21_X1 U18576 ( .B1(n15432), .B2(n16477), .A(n15431), .ZN(P2_U3022) );
  INV_X1 U18577 ( .A(n15433), .ZN(n15447) );
  INV_X1 U18578 ( .A(n15434), .ZN(n15445) );
  OAI21_X1 U18579 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15459), .ZN(n15435) );
  OAI22_X1 U18580 ( .A1(n15455), .A2(n15437), .B1(n15436), .B2(n15435), .ZN(
        n15444) );
  OR2_X1 U18581 ( .A1(n15439), .A2(n15438), .ZN(n15440) );
  AND2_X1 U18582 ( .A1(n15441), .A2(n15440), .ZN(n16356) );
  AOI22_X1 U18583 ( .A1(n16485), .A2(n16356), .B1(n19310), .B2(
        P2_REIP_REG_23__SCAN_IN), .ZN(n15442) );
  OAI21_X1 U18584 ( .B1(n16354), .B2(n15640), .A(n15442), .ZN(n15443) );
  AOI211_X1 U18585 ( .C1(n15445), .C2(n16493), .A(n15444), .B(n15443), .ZN(
        n15446) );
  OAI21_X1 U18586 ( .B1(n15447), .B2(n16477), .A(n15446), .ZN(P2_U3023) );
  NAND2_X1 U18587 ( .A1(n10353), .A2(n15449), .ZN(n15450) );
  XNOR2_X1 U18588 ( .A(n15451), .B(n15450), .ZN(n16362) );
  NOR2_X1 U18589 ( .A1(n15452), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15453) );
  OR2_X1 U18590 ( .A1(n15454), .A2(n15453), .ZN(n16361) );
  INV_X1 U18591 ( .A(n15455), .ZN(n15457) );
  NOR2_X1 U18592 ( .A1(n20130), .A2(n19294), .ZN(n15456) );
  AOI221_X1 U18593 ( .B1(n15459), .B2(n15458), .C1(n15457), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15456), .ZN(n15462) );
  INV_X1 U18594 ( .A(n15945), .ZN(n15460) );
  AOI22_X1 U18595 ( .A1(n16364), .A2(n16492), .B1(n16485), .B2(n15460), .ZN(
        n15461) );
  OAI211_X1 U18596 ( .C1(n16361), .C2(n16457), .A(n15462), .B(n15461), .ZN(
        n15463) );
  INV_X1 U18597 ( .A(n15463), .ZN(n15464) );
  OAI21_X1 U18598 ( .B1(n16362), .B2(n16477), .A(n15464), .ZN(P2_U3024) );
  NOR2_X1 U18599 ( .A1(n15466), .A2(n15465), .ZN(n15473) );
  OR2_X1 U18600 ( .A1(n19138), .A2(n15640), .ZN(n15470) );
  INV_X1 U18601 ( .A(n15467), .ZN(n15468) );
  AOI21_X1 U18602 ( .B1(n16485), .B2(n19132), .A(n15468), .ZN(n15469) );
  OAI211_X1 U18603 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15471), .A(
        n15470), .B(n15469), .ZN(n15472) );
  AOI211_X1 U18604 ( .C1(n15474), .C2(n16493), .A(n15473), .B(n15472), .ZN(
        n15475) );
  OAI21_X1 U18605 ( .B1(n15476), .B2(n16477), .A(n15475), .ZN(P2_U3025) );
  AOI211_X1 U18606 ( .C1(n15479), .C2(n15478), .A(n15477), .B(n15493), .ZN(
        n15483) );
  NAND2_X1 U18607 ( .A1(n19148), .A2(n16492), .ZN(n15481) );
  OAI211_X1 U18608 ( .C1(n16469), .C2(n19151), .A(n15481), .B(n15480), .ZN(
        n15482) );
  AOI211_X1 U18609 ( .C1(n15509), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15483), .B(n15482), .ZN(n15486) );
  NAND2_X1 U18610 ( .A1(n15484), .A2(n16493), .ZN(n15485) );
  OAI211_X1 U18611 ( .C1(n15487), .C2(n16477), .A(n15486), .B(n15485), .ZN(
        P2_U3026) );
  NAND2_X1 U18612 ( .A1(n15488), .A2(n16490), .ZN(n15496) );
  INV_X1 U18613 ( .A(n15489), .ZN(n15490) );
  AOI21_X1 U18614 ( .B1(n16485), .B2(n19158), .A(n15490), .ZN(n15492) );
  NAND2_X1 U18615 ( .A1(n19159), .A2(n16492), .ZN(n15491) );
  OAI211_X1 U18616 ( .C1(n15493), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15492), .B(n15491), .ZN(n15494) );
  AOI21_X1 U18617 ( .B1(n15509), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15494), .ZN(n15495) );
  OAI211_X1 U18618 ( .C1(n15497), .C2(n16457), .A(n15496), .B(n15495), .ZN(
        P2_U3027) );
  INV_X1 U18619 ( .A(n19169), .ZN(n15505) );
  INV_X1 U18620 ( .A(n19172), .ZN(n15503) );
  INV_X1 U18621 ( .A(n15498), .ZN(n15502) );
  NAND2_X1 U18622 ( .A1(n15499), .A2(n15568), .ZN(n15524) );
  NOR3_X1 U18623 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15500), .A3(
        n15524), .ZN(n15501) );
  AOI211_X1 U18624 ( .C1(n16485), .C2(n15503), .A(n15502), .B(n15501), .ZN(
        n15504) );
  OAI21_X1 U18625 ( .B1(n15505), .B2(n15640), .A(n15504), .ZN(n15508) );
  NOR2_X1 U18626 ( .A1(n15506), .A2(n16457), .ZN(n15507) );
  AOI211_X1 U18627 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15509), .A(
        n15508), .B(n15507), .ZN(n15510) );
  OAI21_X1 U18628 ( .B1(n15511), .B2(n16477), .A(n15510), .ZN(P2_U3028) );
  INV_X1 U18629 ( .A(n15512), .ZN(n15513) );
  NOR2_X1 U18630 ( .A1(n15513), .A2(n16493), .ZN(n15514) );
  AND2_X1 U18631 ( .A1(n15517), .A2(n15516), .ZN(n15518) );
  OR2_X1 U18632 ( .A1(n15561), .A2(n15518), .ZN(n15544) );
  NOR2_X1 U18633 ( .A1(n15519), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15520) );
  NOR2_X1 U18634 ( .A1(n15544), .A2(n15520), .ZN(n15521) );
  OAI21_X1 U18635 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15620), .A(
        n15528), .ZN(n15523) );
  NAND2_X1 U18636 ( .A1(n15543), .A2(n16493), .ZN(n15526) );
  INV_X1 U18637 ( .A(n15524), .ZN(n15548) );
  NAND2_X1 U18638 ( .A1(n15548), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15525) );
  NAND2_X1 U18639 ( .A1(n15526), .A2(n15525), .ZN(n15530) );
  INV_X1 U18640 ( .A(n19193), .ZN(n15534) );
  NAND2_X1 U18641 ( .A1(n15530), .A2(n15529), .ZN(n15533) );
  INV_X1 U18642 ( .A(n19196), .ZN(n15531) );
  AOI22_X1 U18643 ( .A1(n16485), .A2(n15531), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19310), .ZN(n15532) );
  OAI211_X1 U18644 ( .C1(n15534), .C2(n15640), .A(n15533), .B(n15532), .ZN(
        n15535) );
  AOI21_X1 U18645 ( .B1(n10015), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15535), .ZN(n15536) );
  OAI21_X1 U18646 ( .B1(n15537), .B2(n16477), .A(n15536), .ZN(P2_U3030) );
  NAND2_X1 U18647 ( .A1(n15539), .A2(n15538), .ZN(n15542) );
  NAND2_X1 U18648 ( .A1(n15540), .A2(n15556), .ZN(n15541) );
  XOR2_X1 U18649 ( .A(n15542), .B(n15541), .Z(n16368) );
  AOI21_X1 U18650 ( .B1(n15549), .B2(n15555), .A(n15543), .ZN(n16369) );
  NAND2_X1 U18651 ( .A1(n15544), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15551) );
  INV_X1 U18652 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20117) );
  NOR2_X1 U18653 ( .A1(n20117), .A2(n19294), .ZN(n15547) );
  XNOR2_X1 U18654 ( .A(n15545), .B(n15565), .ZN(n19372) );
  NOR2_X1 U18655 ( .A1(n16469), .A2(n19372), .ZN(n15546) );
  AOI211_X1 U18656 ( .C1(n15549), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        n15550) );
  OAI211_X1 U18657 ( .C1(n19203), .C2(n15640), .A(n15551), .B(n15550), .ZN(
        n15552) );
  AOI21_X1 U18658 ( .B1(n16369), .B2(n16493), .A(n15552), .ZN(n15553) );
  OAI21_X1 U18659 ( .B1(n16368), .B2(n16477), .A(n15553), .ZN(P2_U3031) );
  NAND2_X1 U18660 ( .A1(n15578), .A2(n15563), .ZN(n15554) );
  NAND2_X1 U18661 ( .A1(n15555), .A2(n15554), .ZN(n16375) );
  NAND2_X1 U18662 ( .A1(n15557), .A2(n15556), .ZN(n15559) );
  XOR2_X1 U18663 ( .A(n15559), .B(n15558), .Z(n16376) );
  OR2_X1 U18664 ( .A1(n16376), .A2(n16477), .ZN(n15577) );
  NAND2_X1 U18665 ( .A1(n15562), .A2(n15568), .ZN(n15560) );
  NOR2_X1 U18666 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15560), .ZN(
        n15604) );
  INV_X1 U18667 ( .A(n15561), .ZN(n15642) );
  OAI21_X1 U18668 ( .B1(n15562), .B2(n15620), .A(n15642), .ZN(n15605) );
  NOR2_X1 U18669 ( .A1(n15604), .A2(n15605), .ZN(n15591) );
  NAND3_X1 U18670 ( .A1(n15562), .A2(n15568), .A3(n15590), .ZN(n15588) );
  AOI21_X1 U18671 ( .B1(n15591), .B2(n15588), .A(n15563), .ZN(n15575) );
  OR2_X1 U18672 ( .A1(n15564), .A2(n15586), .ZN(n15566) );
  NAND2_X1 U18673 ( .A1(n15566), .A2(n15565), .ZN(n19374) );
  INV_X1 U18674 ( .A(n19374), .ZN(n15567) );
  NAND2_X1 U18675 ( .A1(n16485), .A2(n15567), .ZN(n15572) );
  INV_X1 U18676 ( .A(n15568), .ZN(n15644) );
  NOR3_X1 U18677 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15569), .A3(
        n15644), .ZN(n15570) );
  AOI21_X1 U18678 ( .B1(n19310), .B2(P2_REIP_REG_14__SCAN_IN), .A(n15570), 
        .ZN(n15571) );
  OAI211_X1 U18679 ( .C1(n15640), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        n15574) );
  NOR2_X1 U18680 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  OAI211_X1 U18681 ( .C1(n16375), .C2(n16457), .A(n15577), .B(n15576), .ZN(
        P2_U3032) );
  NAND2_X1 U18682 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15636) );
  AOI21_X1 U18683 ( .B1(n16392), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15580) );
  INV_X1 U18684 ( .A(n15578), .ZN(n15579) );
  NOR2_X1 U18685 ( .A1(n15580), .A2(n15579), .ZN(n16380) );
  INV_X1 U18686 ( .A(n16380), .ZN(n15596) );
  INV_X1 U18687 ( .A(n15581), .ZN(n15582) );
  NOR2_X1 U18688 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  XNOR2_X1 U18689 ( .A(n15585), .B(n15584), .ZN(n16382) );
  NAND2_X1 U18690 ( .A1(n16382), .A2(n16490), .ZN(n15595) );
  AOI21_X1 U18691 ( .B1(n15587), .B2(n15607), .A(n15586), .ZN(n19375) );
  OAI22_X1 U18692 ( .A1(n15640), .A2(n19229), .B1(n13957), .B2(n19294), .ZN(
        n15593) );
  OAI22_X1 U18693 ( .A1(n15591), .A2(n15590), .B1(n15589), .B2(n15588), .ZN(
        n15592) );
  AOI211_X1 U18694 ( .C1(n16485), .C2(n19375), .A(n15593), .B(n15592), .ZN(
        n15594) );
  OAI211_X1 U18695 ( .C1(n15596), .C2(n16457), .A(n15595), .B(n15594), .ZN(
        P2_U3033) );
  XNOR2_X1 U18696 ( .A(n16392), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16386) );
  NOR2_X1 U18697 ( .A1(n9900), .A2(n15597), .ZN(n15602) );
  INV_X1 U18698 ( .A(n15598), .ZN(n15600) );
  NAND2_X1 U18699 ( .A1(n15600), .A2(n15599), .ZN(n15601) );
  XNOR2_X1 U18700 ( .A(n15602), .B(n15601), .ZN(n16387) );
  NOR2_X1 U18701 ( .A1(n13956), .A2(n19294), .ZN(n15603) );
  AOI211_X1 U18702 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15605), .A(
        n15604), .B(n15603), .ZN(n15611) );
  OR2_X1 U18703 ( .A1(n15606), .A2(n9933), .ZN(n15608) );
  NAND2_X1 U18704 ( .A1(n15608), .A2(n15607), .ZN(n19378) );
  INV_X1 U18705 ( .A(n19378), .ZN(n15609) );
  AOI22_X1 U18706 ( .A1(n19237), .A2(n16492), .B1(n16485), .B2(n15609), .ZN(
        n15610) );
  OAI211_X1 U18707 ( .C1(n16387), .C2(n16477), .A(n15611), .B(n15610), .ZN(
        n15612) );
  INV_X1 U18708 ( .A(n15612), .ZN(n15613) );
  OAI21_X1 U18709 ( .B1(n16457), .B2(n16386), .A(n15613), .ZN(P2_U3034) );
  XNOR2_X1 U18710 ( .A(n15636), .B(n15622), .ZN(n16409) );
  INV_X1 U18711 ( .A(n15615), .ZN(n15634) );
  OR2_X1 U18712 ( .A1(n15614), .A2(n15634), .ZN(n15619) );
  AND2_X1 U18713 ( .A1(n15617), .A2(n15616), .ZN(n15618) );
  XNOR2_X1 U18714 ( .A(n15619), .B(n15618), .ZN(n16408) );
  NOR2_X1 U18715 ( .A1(n15643), .A2(n15644), .ZN(n16461) );
  OAI21_X1 U18716 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15620), .A(
        n15642), .ZN(n16452) );
  NOR2_X1 U18717 ( .A1(n12543), .A2(n19294), .ZN(n15621) );
  AOI221_X1 U18718 ( .B1(n16461), .B2(n15622), .C1(n16452), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15621), .ZN(n15628) );
  OR2_X1 U18719 ( .A1(n15623), .A2(n15638), .ZN(n15625) );
  NAND2_X1 U18720 ( .A1(n15625), .A2(n15624), .ZN(n19383) );
  INV_X1 U18721 ( .A(n19383), .ZN(n15626) );
  AOI22_X1 U18722 ( .A1(n16492), .A2(n19247), .B1(n16485), .B2(n15626), .ZN(
        n15627) );
  OAI211_X1 U18723 ( .C1(n16408), .C2(n16477), .A(n15628), .B(n15627), .ZN(
        n15629) );
  INV_X1 U18724 ( .A(n15629), .ZN(n15630) );
  OAI21_X1 U18725 ( .B1(n16457), .B2(n16409), .A(n15630), .ZN(P2_U3036) );
  INV_X1 U18726 ( .A(n15614), .ZN(n15635) );
  OAI21_X1 U18727 ( .B1(n15632), .B2(n15634), .A(n15631), .ZN(n15633) );
  OAI21_X1 U18728 ( .B1(n15635), .B2(n15634), .A(n15633), .ZN(n16415) );
  INV_X1 U18729 ( .A(n15636), .ZN(n16413) );
  NOR2_X1 U18730 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16414) );
  OR3_X1 U18731 ( .A1(n16413), .A2(n16414), .A3(n16457), .ZN(n15648) );
  AOI21_X1 U18732 ( .B1(n15639), .B2(n16467), .A(n15638), .ZN(n19386) );
  NOR2_X1 U18733 ( .A1(n15640), .A2(n19260), .ZN(n15646) );
  NAND2_X1 U18734 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19310), .ZN(n15641) );
  OAI221_X1 U18735 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15644), .C1(
        n15643), .C2(n15642), .A(n15641), .ZN(n15645) );
  AOI211_X1 U18736 ( .C1(n16485), .C2(n19386), .A(n15646), .B(n15645), .ZN(
        n15647) );
  OAI211_X1 U18737 ( .C1(n16415), .C2(n16477), .A(n15648), .B(n15647), .ZN(
        P2_U3037) );
  INV_X1 U18738 ( .A(n20163), .ZN(n15744) );
  INV_X1 U18739 ( .A(n11108), .ZN(n15650) );
  NAND2_X1 U18740 ( .A1(n15650), .A2(n15649), .ZN(n15667) );
  MUX2_X1 U18741 ( .A(n15667), .B(n10646), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15651) );
  AOI21_X1 U18742 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n16506) );
  OAI22_X1 U18743 ( .A1(n15010), .A2(n15654), .B1(n19359), .B2(n19315), .ZN(
        n15661) );
  OAI222_X1 U18744 ( .A1(n15656), .A2(n15655), .B1(n15744), .B2(n16506), .C1(
        n20079), .C2(n15661), .ZN(n15657) );
  MUX2_X1 U18745 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15657), .S(
        n15749), .Z(P2_U3601) );
  OAI21_X1 U18746 ( .B1(n19359), .B2(n15659), .A(n15658), .ZN(n19338) );
  OAI21_X1 U18747 ( .B1(n9843), .B2(n15660), .A(n19338), .ZN(n15684) );
  INV_X1 U18748 ( .A(n15684), .ZN(n15669) );
  INV_X1 U18749 ( .A(n15661), .ZN(n15662) );
  NOR2_X1 U18750 ( .A1(n15662), .A2(n20079), .ZN(n15683) );
  NOR2_X1 U18751 ( .A1(n15663), .A2(n15664), .ZN(n15666) );
  AOI22_X1 U18752 ( .A1(n15667), .A2(n15666), .B1(n10646), .B2(n15665), .ZN(
        n15668) );
  OAI21_X1 U18753 ( .B1(n19330), .B2(n15682), .A(n15668), .ZN(n16508) );
  AOI222_X1 U18754 ( .A1(n20184), .A2(n16547), .B1(n15669), .B2(n15683), .C1(
        n16508), .C2(n20163), .ZN(n15671) );
  NAND2_X1 U18755 ( .A1(n15686), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15670) );
  OAI21_X1 U18756 ( .B1(n15671), .B2(n15686), .A(n15670), .ZN(P2_U3600) );
  NOR2_X1 U18757 ( .A1(n15673), .A2(n10894), .ZN(n15676) );
  OAI22_X1 U18758 ( .A1(n15677), .A2(n15676), .B1(n15675), .B2(n15674), .ZN(
        n15678) );
  AOI21_X1 U18759 ( .B1(n15680), .B2(n15679), .A(n15678), .ZN(n15681) );
  OAI21_X1 U18760 ( .B1(n13468), .B2(n15682), .A(n15681), .ZN(n16513) );
  AOI222_X1 U18761 ( .A1(n16513), .A2(n20163), .B1(n15684), .B2(n15683), .C1(
        n16547), .C2(n20174), .ZN(n15687) );
  NAND2_X1 U18762 ( .A1(n15686), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15685) );
  OAI21_X1 U18763 ( .B1(n15687), .B2(n15686), .A(n15685), .ZN(P2_U3599) );
  INV_X1 U18764 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16964) );
  INV_X1 U18765 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16986) );
  INV_X1 U18766 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17013) );
  NOR4_X1 U18767 ( .A1(n17013), .A2(n17437), .A3(n17436), .A4(n17392), .ZN(
        n17410) );
  NAND2_X1 U18768 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17410), .ZN(n17389) );
  NAND2_X1 U18769 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17375), .ZN(n15688) );
  NOR2_X1 U18770 ( .A1(n16964), .A2(n15688), .ZN(n17325) );
  INV_X1 U18771 ( .A(n15688), .ZN(n15689) );
  OAI21_X1 U18772 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15689), .A(n17451), .ZN(
        n15703) );
  AOI22_X1 U18773 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15690) );
  OAI21_X1 U18774 ( .B1(n13155), .B2(n15691), .A(n15690), .ZN(n15702) );
  AOI22_X1 U18775 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15699) );
  INV_X1 U18776 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18777 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U18778 ( .B1(n9846), .B2(n15693), .A(n15692), .ZN(n15697) );
  AOI22_X1 U18779 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15695) );
  AOI22_X1 U18780 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15694) );
  OAI211_X1 U18781 ( .C1(n15793), .C2(n17216), .A(n15695), .B(n15694), .ZN(
        n15696) );
  AOI211_X1 U18782 ( .C1(n9965), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15697), .B(n15696), .ZN(n15698) );
  OAI211_X1 U18783 ( .C1(n17344), .C2(n15700), .A(n15699), .B(n15698), .ZN(
        n15701) );
  AOI211_X1 U18784 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n15702), .B(n15701), .ZN(n17548) );
  OAI22_X1 U18785 ( .A1(n17325), .A2(n15703), .B1(n17548), .B2(n17451), .ZN(
        P3_U2690) );
  INV_X1 U18786 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19031) );
  NOR2_X1 U18787 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19031), .ZN(
        n18398) );
  NAND3_X1 U18788 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19029)
         );
  INV_X1 U18789 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17078) );
  OAI21_X1 U18790 ( .B1(n15704), .B2(n19055), .A(n17078), .ZN(n15742) );
  NOR2_X1 U18791 ( .A1(n9822), .A2(n15742), .ZN(n18397) );
  NOR2_X1 U18792 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19087) );
  AOI21_X1 U18793 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19087), .ZN(n18932) );
  NOR2_X1 U18794 ( .A1(n19056), .A2(n18932), .ZN(n18411) );
  INV_X1 U18795 ( .A(n18765), .ZN(n18565) );
  INV_X1 U18796 ( .A(n19029), .ZN(n15705) );
  NAND2_X1 U18797 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n15705), .ZN(n15741) );
  OAI211_X1 U18798 ( .C1(n19029), .C2(n18397), .A(n18565), .B(n15741), .ZN(
        n18404) );
  INV_X1 U18799 ( .A(n18404), .ZN(n18400) );
  NOR2_X1 U18800 ( .A1(n18398), .A2(n18400), .ZN(n15707) );
  INV_X1 U18801 ( .A(n18713), .ZN(n18762) );
  NOR2_X1 U18802 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19058) );
  INV_X1 U18803 ( .A(n19058), .ZN(n19095) );
  NAND2_X1 U18804 ( .A1(n18177), .A2(n19031), .ZN(n16727) );
  NAND2_X1 U18805 ( .A1(n19095), .A2(n16727), .ZN(n19077) );
  INV_X1 U18806 ( .A(n19077), .ZN(n16566) );
  NAND2_X1 U18807 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18044) );
  INV_X1 U18808 ( .A(n18044), .ZN(n17982) );
  OAI22_X1 U18809 ( .A1(n16566), .A2(n17982), .B1(n18897), .B2(n19031), .ZN(
        n15710) );
  NAND3_X1 U18810 ( .A1(n18898), .A2(n18404), .A3(n15710), .ZN(n15706) );
  OAI221_X1 U18811 ( .B1(n18898), .B2(n15707), .C1(n18898), .C2(n18762), .A(
        n15706), .ZN(P3_U2864) );
  NAND2_X1 U18812 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18406) );
  NOR2_X1 U18813 ( .A1(n16566), .A2(n17982), .ZN(n15709) );
  INV_X1 U18814 ( .A(n15707), .ZN(n15708) );
  AOI221_X1 U18815 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18406), .C1(n15709), 
        .C2(n18406), .A(n15708), .ZN(n18403) );
  OAI221_X1 U18816 ( .B1(n18713), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18713), .C2(n15710), .A(n18404), .ZN(n18401) );
  AOI22_X1 U18817 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18403), .B1(
        n18401), .B2(n18903), .ZN(P3_U2865) );
  NAND2_X1 U18818 ( .A1(n15714), .A2(n15713), .ZN(n15711) );
  OAI211_X1 U18819 ( .C1(n15714), .C2(n15713), .A(n15712), .B(n15711), .ZN(
        n15875) );
  NAND2_X1 U18820 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19085) );
  NOR2_X1 U18821 ( .A1(n16731), .A2(n18938), .ZN(n15740) );
  NAND3_X1 U18822 ( .A1(n15728), .A2(n17463), .A3(n15872), .ZN(n15731) );
  NOR2_X1 U18823 ( .A1(n15715), .A2(n17463), .ZN(n15720) );
  NAND2_X1 U18824 ( .A1(n19084), .A2(n9877), .ZN(n17647) );
  INV_X2 U18825 ( .A(n19093), .ZN(n19092) );
  NAND2_X2 U18826 ( .A1(n19092), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19015) );
  OAI211_X1 U18827 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18950), .B(n19015), .ZN(n19082) );
  NAND2_X1 U18828 ( .A1(n17463), .A2(n18437), .ZN(n16003) );
  NAND2_X1 U18829 ( .A1(n19084), .A2(n18412), .ZN(n15886) );
  AOI21_X1 U18830 ( .B1(n18449), .B2(n16003), .A(n15886), .ZN(n15730) );
  NAND2_X1 U18831 ( .A1(n15728), .A2(n15887), .ZN(n15724) );
  AOI211_X1 U18832 ( .C1(n18432), .C2(n16003), .A(n15717), .B(n15729), .ZN(
        n15718) );
  INV_X1 U18833 ( .A(n15718), .ZN(n15719) );
  INV_X1 U18834 ( .A(n15720), .ZN(n15725) );
  NAND2_X1 U18835 ( .A1(n15728), .A2(n15720), .ZN(n15871) );
  AOI21_X1 U18836 ( .B1(n15731), .B2(n15871), .A(n18412), .ZN(n15723) );
  NAND2_X1 U18837 ( .A1(n18449), .A2(n15725), .ZN(n15722) );
  AOI21_X1 U18838 ( .B1(n15869), .B2(n15732), .A(n15726), .ZN(n15727) );
  NOR2_X1 U18839 ( .A1(n15730), .A2(n15727), .ZN(n15881) );
  NAND2_X1 U18840 ( .A1(n15734), .A2(n15728), .ZN(n15890) );
  AOI21_X1 U18841 ( .B1(n15879), .B2(n15731), .A(n15730), .ZN(n15733) );
  OAI211_X1 U18842 ( .C1(n15888), .C2(n18869), .A(n15881), .B(n16002), .ZN(
        n15739) );
  NAND2_X1 U18843 ( .A1(n18923), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18410) );
  AND2_X1 U18844 ( .A1(n15742), .A2(n18881), .ZN(n18871) );
  NAND3_X1 U18845 ( .A1(n19060), .A2(n19058), .A3(n18871), .ZN(n15743) );
  OAI21_X1 U18846 ( .B1(n19060), .B2(n17078), .A(n15743), .ZN(P3_U3284) );
  NOR4_X1 U18847 ( .A1(n15745), .A2(n16522), .A3(n9833), .A4(n15744), .ZN(
        n15746) );
  NAND2_X1 U18848 ( .A1(n15749), .A2(n15746), .ZN(n15747) );
  OAI21_X1 U18849 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(P2_U3595) );
  INV_X1 U18850 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U18851 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15750) );
  OAI21_X1 U18852 ( .B1(n17396), .B2(n18827), .A(n15750), .ZN(n15757) );
  AOI22_X1 U18853 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U18854 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15751) );
  OAI21_X1 U18855 ( .B1(n9846), .B2(n15752), .A(n15751), .ZN(n15754) );
  AOI22_X1 U18856 ( .A1(n13142), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15753) );
  AOI211_X2 U18857 ( .C1(n17281), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n15757), .B(n15756), .ZN(n17591) );
  AOI22_X1 U18858 ( .A1(n13142), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15759) );
  AOI22_X1 U18859 ( .A1(n17359), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15758) );
  OAI211_X1 U18860 ( .C1(n9828), .C2(n18419), .A(n15759), .B(n15758), .ZN(
        n15760) );
  AOI22_X1 U18861 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15763) );
  NAND3_X1 U18862 ( .A1(n15764), .A2(n15763), .A3(n15762), .ZN(n15770) );
  AOI22_X1 U18863 ( .A1(n17360), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U18864 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15767) );
  AOI22_X1 U18865 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17311), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15766) );
  NAND2_X1 U18866 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n15765) );
  NAND4_X1 U18867 ( .A1(n15768), .A2(n15767), .A3(n15766), .A4(n15765), .ZN(
        n15769) );
  OR2_X2 U18868 ( .A1(n15770), .A2(n15769), .ZN(n15802) );
  INV_X1 U18869 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18424) );
  AOI22_X1 U18870 ( .A1(n13142), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15771) );
  AOI22_X1 U18871 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15775) );
  AOI22_X1 U18872 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17360), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U18873 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15773) );
  AOI22_X1 U18874 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15776) );
  NAND2_X1 U18875 ( .A1(n15802), .A2(n17597), .ZN(n15903) );
  INV_X1 U18876 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U18877 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U18878 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18879 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15777) );
  OAI211_X1 U18880 ( .C1(n9828), .C2(n18435), .A(n15778), .B(n15777), .ZN(
        n15784) );
  AOI22_X1 U18881 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18882 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15781) );
  AOI22_X1 U18883 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15780) );
  NAND2_X1 U18884 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n15779) );
  NAND4_X1 U18885 ( .A1(n15782), .A2(n15781), .A3(n15780), .A4(n15779), .ZN(
        n15783) );
  AOI211_X1 U18886 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15784), .B(n15783), .ZN(n15785) );
  NAND2_X1 U18887 ( .A1(n15801), .A2(n15898), .ZN(n15823) );
  AOI22_X1 U18888 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15788) );
  OAI21_X1 U18889 ( .B1(n17415), .B2(n17221), .A(n15788), .ZN(n15800) );
  AOI22_X1 U18890 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15797) );
  AOI22_X1 U18891 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15789) );
  OAI21_X1 U18892 ( .B1(n9828), .B2(n18441), .A(n15789), .ZN(n15795) );
  AOI22_X1 U18893 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15791) );
  AOI22_X1 U18894 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15790) );
  OAI211_X1 U18895 ( .C1(n15793), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15794) );
  AOI211_X1 U18896 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15795), .B(n15794), .ZN(n15796) );
  OAI211_X1 U18897 ( .C1(n17344), .C2(n15798), .A(n15797), .B(n15796), .ZN(
        n15799) );
  XNOR2_X1 U18898 ( .A(n15823), .B(n17584), .ZN(n15820) );
  XNOR2_X1 U18899 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n15802), .ZN(
        n18073) );
  INV_X1 U18900 ( .A(n18073), .ZN(n18075) );
  INV_X1 U18901 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U18902 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U18903 ( .A1(n17360), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15804) );
  AOI22_X1 U18904 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15803) );
  OAI211_X1 U18905 ( .C1(n9828), .C2(n18415), .A(n15804), .B(n15803), .ZN(
        n15811) );
  AOI22_X1 U18906 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15805) );
  INV_X1 U18907 ( .A(n15805), .ZN(n15810) );
  AOI22_X1 U18908 ( .A1(n17418), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15808) );
  AOI22_X1 U18909 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15807) );
  NAND3_X1 U18910 ( .A1(n15808), .A2(n15807), .A3(n15806), .ZN(n15809) );
  OAI211_X1 U18911 ( .C1(n13155), .C2(n17413), .A(n15813), .B(n15812), .ZN(
        n16004) );
  NAND2_X1 U18912 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16004), .ZN(
        n18082) );
  AOI21_X1 U18913 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17608), .A(
        n18074), .ZN(n18063) );
  INV_X1 U18914 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18372) );
  XNOR2_X1 U18915 ( .A(n18372), .B(n15814), .ZN(n18062) );
  NOR2_X1 U18916 ( .A1(n18063), .A2(n18062), .ZN(n18061) );
  NOR2_X1 U18917 ( .A1(n18372), .A2(n15814), .ZN(n15815) );
  NOR2_X1 U18918 ( .A1(n18061), .A2(n15815), .ZN(n15817) );
  XNOR2_X1 U18919 ( .A(n15903), .B(n17591), .ZN(n15816) );
  NOR2_X1 U18920 ( .A1(n15817), .A2(n15816), .ZN(n15818) );
  INV_X1 U18921 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18358) );
  XNOR2_X1 U18922 ( .A(n15817), .B(n15816), .ZN(n18053) );
  XNOR2_X1 U18923 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15819), .ZN(
        n18040) );
  AOI22_X1 U18924 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15833) );
  INV_X1 U18925 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U18926 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U18927 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15824) );
  OAI211_X1 U18928 ( .C1(n17298), .C2(n17327), .A(n15825), .B(n15824), .ZN(
        n15831) );
  AOI22_X1 U18929 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U18930 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15828) );
  AOI22_X1 U18931 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15827) );
  NAND2_X1 U18932 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n15826) );
  NAND4_X1 U18933 ( .A1(n15829), .A2(n15828), .A3(n15827), .A4(n15826), .ZN(
        n15830) );
  AOI211_X1 U18934 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n15831), .B(n15830), .ZN(n15832) );
  XOR2_X1 U18935 ( .A(n15836), .B(n18008), .Z(n15834) );
  XNOR2_X1 U18936 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15834), .ZN(
        n18017) );
  NAND2_X1 U18937 ( .A1(n15836), .A2(n18008), .ZN(n16621) );
  INV_X1 U18938 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U18939 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15837), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15847) );
  AOI22_X1 U18940 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15839) );
  AOI22_X1 U18941 ( .A1(n17359), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15838) );
  OAI211_X1 U18942 ( .C1(n9828), .C2(n18454), .A(n15839), .B(n15838), .ZN(
        n15845) );
  AOI22_X1 U18943 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17412), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15843) );
  AOI22_X1 U18944 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15842) );
  AOI22_X1 U18945 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15841) );
  NAND2_X1 U18946 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n15840) );
  NAND4_X1 U18947 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        n15844) );
  AOI211_X1 U18948 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n15845), .B(n15844), .ZN(n15846) );
  AOI21_X1 U18949 ( .B1(n16621), .B2(n17578), .A(n15851), .ZN(n15848) );
  INV_X1 U18950 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18301) );
  NOR2_X1 U18951 ( .A1(n15849), .A2(n10072), .ZN(n15852) );
  INV_X1 U18952 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15850) );
  INV_X1 U18953 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17903) );
  INV_X1 U18954 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18231) );
  INV_X1 U18955 ( .A(n15851), .ZN(n17951) );
  NAND2_X1 U18956 ( .A1(n17870), .A2(n17951), .ZN(n15857) );
  INV_X1 U18957 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18319) );
  INV_X1 U18958 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U18959 ( .A1(n18290), .A2(n17950), .ZN(n18276) );
  NAND2_X1 U18960 ( .A1(n18276), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18260) );
  NOR2_X1 U18961 ( .A1(n18260), .A2(n18267), .ZN(n17910) );
  NAND2_X1 U18962 ( .A1(n17910), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18237) );
  NOR2_X1 U18963 ( .A1(n18237), .A2(n17903), .ZN(n17900) );
  NAND2_X1 U18964 ( .A1(n17900), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18148) );
  NAND2_X1 U18965 ( .A1(n17799), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15856) );
  INV_X1 U18966 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18216) );
  NAND2_X1 U18967 ( .A1(n15863), .A2(n18216), .ZN(n15855) );
  INV_X1 U18968 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18203) );
  INV_X1 U18969 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18133) );
  NAND2_X1 U18970 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18197) );
  INV_X1 U18971 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18147) );
  NOR2_X1 U18972 ( .A1(n18197), .A2(n18147), .ZN(n18149) );
  INV_X1 U18973 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17830) );
  INV_X1 U18974 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17822) );
  NOR2_X1 U18975 ( .A1(n17830), .A2(n17822), .ZN(n18156) );
  NAND2_X1 U18976 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18156), .ZN(
        n17796) );
  INV_X1 U18977 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18159) );
  NOR2_X1 U18978 ( .A1(n17796), .A2(n18159), .ZN(n15862) );
  NAND2_X1 U18979 ( .A1(n18149), .A2(n15862), .ZN(n18140) );
  NOR2_X1 U18980 ( .A1(n18133), .A2(n18140), .ZN(n15921) );
  NAND2_X1 U18981 ( .A1(n17853), .A2(n17830), .ZN(n15858) );
  NOR2_X1 U18982 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15858), .ZN(
        n17817) );
  INV_X1 U18983 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17809) );
  NAND2_X1 U18984 ( .A1(n17817), .A2(n17809), .ZN(n17798) );
  NAND2_X1 U18985 ( .A1(n15859), .A2(n10420), .ZN(n15860) );
  INV_X1 U18986 ( .A(n18197), .ZN(n17852) );
  NAND2_X1 U18987 ( .A1(n17852), .A2(n15861), .ZN(n17816) );
  INV_X1 U18988 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18119) );
  NAND2_X1 U18989 ( .A1(n15863), .A2(n18119), .ZN(n15864) );
  NAND2_X1 U18990 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18091) );
  NOR2_X1 U18991 ( .A1(n17744), .A2(n15866), .ZN(n15867) );
  NAND2_X1 U18992 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15867), .ZN(
        n17732) );
  NAND2_X1 U18993 ( .A1(n15863), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16615) );
  NOR2_X2 U18994 ( .A1(n15867), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17731) );
  INV_X1 U18995 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17719) );
  NAND3_X1 U18996 ( .A1(n17731), .A2(n17951), .A3(n17719), .ZN(n15985) );
  OAI21_X1 U18997 ( .B1(n17732), .B2(n16615), .A(n15985), .ZN(n15868) );
  NOR2_X1 U18998 ( .A1(n19084), .A2(n18421), .ZN(n15877) );
  NAND2_X1 U18999 ( .A1(n15877), .A2(n18443), .ZN(n15882) );
  INV_X1 U19000 ( .A(n15869), .ZN(n15870) );
  AOI21_X1 U19001 ( .B1(n15872), .B2(n15871), .A(n18869), .ZN(n15884) );
  INV_X1 U19002 ( .A(n15873), .ZN(n15876) );
  OAI21_X1 U19003 ( .B1(n15876), .B2(n15875), .A(n15874), .ZN(n18864) );
  AOI21_X1 U19004 ( .B1(n19084), .B2(n18421), .A(n15877), .ZN(n15878) );
  AOI21_X1 U19005 ( .B1(n15878), .B2(n19082), .A(n18938), .ZN(n16730) );
  NAND3_X1 U19006 ( .A1(n16730), .A2(n15879), .A3(n18865), .ZN(n15880) );
  INV_X1 U19007 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18097) );
  NAND2_X1 U19008 ( .A1(n15887), .A2(n15886), .ZN(n19081) );
  NAND2_X1 U19009 ( .A1(n9820), .A2(n10174), .ZN(n18283) );
  INV_X1 U19010 ( .A(n18892), .ZN(n18882) );
  NOR2_X1 U19011 ( .A1(n18882), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18192) );
  INV_X1 U19012 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18105) );
  INV_X1 U19013 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15920) );
  NOR2_X1 U19014 ( .A1(n18133), .A2(n15920), .ZN(n18112) );
  NAND2_X1 U19015 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18112), .ZN(
        n18104) );
  NOR2_X1 U19016 ( .A1(n18105), .A2(n18104), .ZN(n16586) );
  AOI21_X1 U19017 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18304) );
  INV_X1 U19018 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18007) );
  NAND3_X1 U19019 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18329) );
  NOR2_X1 U19020 ( .A1(n18007), .A2(n18329), .ZN(n18188) );
  NOR2_X1 U19021 ( .A1(n18319), .A2(n18301), .ZN(n18189) );
  NAND2_X1 U19022 ( .A1(n18188), .A2(n18189), .ZN(n15891) );
  NOR2_X1 U19023 ( .A1(n18304), .A2(n15891), .ZN(n18270) );
  NAND2_X1 U19024 ( .A1(n18190), .A2(n18270), .ZN(n18193) );
  NOR2_X1 U19025 ( .A1(n18140), .A2(n18193), .ZN(n18132) );
  AOI21_X1 U19026 ( .B1(n16586), .B2(n18132), .A(n10174), .ZN(n18089) );
  NAND2_X1 U19027 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18366) );
  NOR2_X1 U19028 ( .A1(n18366), .A2(n15891), .ZN(n18209) );
  NAND2_X1 U19029 ( .A1(n18190), .A2(n18209), .ZN(n18191) );
  NOR2_X1 U19030 ( .A1(n18140), .A2(n18191), .ZN(n18127) );
  INV_X1 U19031 ( .A(n16586), .ZN(n17740) );
  NOR2_X1 U19032 ( .A1(n18097), .A2(n17740), .ZN(n16618) );
  AOI21_X1 U19033 ( .B1(n18127), .B2(n16618), .A(n18882), .ZN(n15893) );
  AOI21_X1 U19034 ( .B1(n16586), .B2(n18127), .A(n9820), .ZN(n15892) );
  NOR4_X1 U19035 ( .A1(n18192), .A2(n18089), .A3(n15893), .A4(n15892), .ZN(
        n15988) );
  INV_X1 U19036 ( .A(n15988), .ZN(n15894) );
  AOI21_X1 U19037 ( .B1(n18097), .B2(n18283), .A(n15894), .ZN(n16622) );
  AOI21_X1 U19038 ( .B1(n18309), .B2(n17719), .A(n18392), .ZN(n15924) );
  NOR2_X1 U19039 ( .A1(n18097), .A2(n17719), .ZN(n16587) );
  NAND2_X1 U19040 ( .A1(n16587), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15990) );
  INV_X1 U19041 ( .A(n15898), .ZN(n17588) );
  INV_X1 U19042 ( .A(n16004), .ZN(n15904) );
  NOR2_X1 U19043 ( .A1(n17608), .A2(n15904), .ZN(n15905) );
  NOR2_X1 U19044 ( .A1(n17597), .A2(n15905), .ZN(n15901) );
  OR2_X1 U19045 ( .A1(n17591), .A2(n15901), .ZN(n15897) );
  NAND2_X1 U19046 ( .A1(n18008), .A2(n18012), .ZN(n15913) );
  NOR2_X1 U19047 ( .A1(n15913), .A2(n17578), .ZN(n15918) );
  INV_X1 U19048 ( .A(n15918), .ZN(n15914) );
  INV_X1 U19049 ( .A(n18012), .ZN(n18010) );
  XNOR2_X1 U19050 ( .A(n18008), .B(n18010), .ZN(n15912) );
  XOR2_X1 U19051 ( .A(n17584), .B(n15895), .Z(n15896) );
  NAND2_X1 U19052 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15896), .ZN(
        n15911) );
  XNOR2_X1 U19053 ( .A(n18028), .B(n15896), .ZN(n18031) );
  XNOR2_X1 U19054 ( .A(n15898), .B(n15897), .ZN(n15899) );
  NAND2_X1 U19055 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15899), .ZN(
        n15910) );
  INV_X1 U19056 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18348) );
  XNOR2_X1 U19057 ( .A(n18348), .B(n15899), .ZN(n18039) );
  XOR2_X1 U19058 ( .A(n15901), .B(n17591), .Z(n15900) );
  NAND2_X1 U19059 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15900), .ZN(
        n15909) );
  XNOR2_X1 U19060 ( .A(n18358), .B(n15900), .ZN(n18051) );
  INV_X1 U19061 ( .A(n15901), .ZN(n15902) );
  OAI21_X1 U19062 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(n15907) );
  NAND2_X1 U19063 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15907), .ZN(
        n15908) );
  NOR2_X1 U19064 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15802), .ZN(
        n15906) );
  INV_X1 U19065 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19059) );
  NAND2_X1 U19066 ( .A1(n15904), .A2(n19059), .ZN(n18081) );
  NOR2_X1 U19067 ( .A1(n18073), .A2(n18081), .ZN(n18072) );
  NOR3_X1 U19068 ( .A1(n15906), .A2(n15905), .A3(n18072), .ZN(n18066) );
  XNOR2_X1 U19069 ( .A(n18372), .B(n15907), .ZN(n18065) );
  NAND2_X1 U19070 ( .A1(n18066), .A2(n18065), .ZN(n18064) );
  NAND2_X1 U19071 ( .A1(n15908), .A2(n18064), .ZN(n18050) );
  NAND2_X1 U19072 ( .A1(n18051), .A2(n18050), .ZN(n18049) );
  NAND2_X1 U19073 ( .A1(n15909), .A2(n18049), .ZN(n18038) );
  NAND2_X1 U19074 ( .A1(n18039), .A2(n18038), .ZN(n18037) );
  NAND2_X1 U19075 ( .A1(n15910), .A2(n18037), .ZN(n18030) );
  NAND2_X1 U19076 ( .A1(n18031), .A2(n18030), .ZN(n18029) );
  NAND2_X1 U19077 ( .A1(n15911), .A2(n18029), .ZN(n18011) );
  AOI222_X1 U19078 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15912), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18011), .C1(n15912), .C2(
        n18011), .ZN(n17996) );
  XOR2_X1 U19079 ( .A(n16619), .B(n15913), .Z(n17997) );
  NAND2_X1 U19080 ( .A1(n17996), .A2(n17997), .ZN(n17995) );
  NAND2_X1 U19081 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17995), .ZN(
        n15917) );
  NOR2_X1 U19082 ( .A1(n15914), .A2(n15917), .ZN(n15919) );
  NOR2_X1 U19083 ( .A1(n17996), .A2(n17997), .ZN(n15916) );
  NOR2_X1 U19084 ( .A1(n15918), .A2(n15917), .ZN(n15915) );
  AOI211_X1 U19085 ( .C1(n15918), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        n17980) );
  NOR2_X1 U19086 ( .A1(n17980), .A2(n18319), .ZN(n17979) );
  NOR2_X1 U19087 ( .A1(n18273), .A2(n18148), .ZN(n18157) );
  NAND2_X1 U19088 ( .A1(n15921), .A2(n18157), .ZN(n18129) );
  NOR2_X1 U19089 ( .A1(n15920), .A2(n18129), .ZN(n17767) );
  NAND3_X1 U19090 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n17767), .ZN(n18095) );
  NOR2_X1 U19091 ( .A1(n15990), .A2(n18095), .ZN(n16573) );
  INV_X1 U19092 ( .A(n16573), .ZN(n16578) );
  NAND2_X1 U19093 ( .A1(n18271), .A2(n18190), .ZN(n18218) );
  INV_X1 U19094 ( .A(n15921), .ZN(n15922) );
  NAND2_X1 U19095 ( .A1(n18131), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17766) );
  NOR2_X1 U19096 ( .A1(n18119), .A2(n17766), .ZN(n17765) );
  NAND2_X1 U19097 ( .A1(n17765), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17717) );
  NOR2_X1 U19098 ( .A1(n17717), .A2(n15990), .ZN(n16577) );
  NOR2_X1 U19099 ( .A1(n16619), .A2(n18863), .ZN(n18248) );
  INV_X1 U19100 ( .A(n18248), .ZN(n18313) );
  NOR3_X1 U19101 ( .A1(n16577), .A2(n18392), .A3(n18313), .ZN(n15923) );
  AOI21_X1 U19102 ( .B1(n18322), .B2(n16578), .A(n15923), .ZN(n15991) );
  OAI221_X1 U19103 ( .B1(n9832), .B2(n16622), .C1(n9832), .C2(n15924), .A(
        n15991), .ZN(n15928) );
  INV_X1 U19104 ( .A(n16587), .ZN(n15925) );
  NOR2_X1 U19105 ( .A1(n15925), .A2(n18095), .ZN(n16624) );
  NOR2_X1 U19106 ( .A1(n17717), .A2(n15925), .ZN(n16625) );
  AOI22_X1 U19107 ( .A1(n18868), .A2(n16624), .B1(n18248), .B2(n16625), .ZN(
        n15927) );
  INV_X1 U19108 ( .A(n9820), .ZN(n18874) );
  AOI21_X1 U19109 ( .B1(n18892), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18874), .ZN(n18187) );
  OAI22_X1 U19110 ( .A1(n10174), .A2(n18193), .B1(n18187), .B2(n18191), .ZN(
        n15926) );
  INV_X1 U19111 ( .A(n15926), .ZN(n16617) );
  NOR2_X1 U19112 ( .A1(n16617), .A2(n18140), .ZN(n18111) );
  NAND3_X1 U19113 ( .A1(n16587), .A2(n18111), .A3(n16586), .ZN(n16607) );
  AOI21_X1 U19114 ( .B1(n15927), .B2(n16607), .A(n18392), .ZN(n15993) );
  INV_X1 U19115 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16609) );
  AOI22_X1 U19116 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15928), .B1(
        n15993), .B2(n16609), .ZN(n15929) );
  NAND2_X1 U19117 ( .A1(n9832), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16602) );
  OAI211_X1 U19118 ( .C1(n16593), .C2(n18299), .A(n15929), .B(n16602), .ZN(
        P3_U2833) );
  OAI22_X1 U19119 ( .A1(n10228), .A2(n19353), .B1(n20130), .B2(n19342), .ZN(
        n15933) );
  INV_X1 U19120 ( .A(n15930), .ZN(n15931) );
  OAI22_X1 U19121 ( .A1(n15931), .A2(n19328), .B1(n14180), .B2(n19343), .ZN(
        n15932) );
  AOI211_X1 U19122 ( .C1(n16364), .C2(n19290), .A(n15933), .B(n15932), .ZN(
        n15944) );
  OAI21_X1 U19123 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15935), .A(
        n15934), .ZN(n16367) );
  INV_X1 U19124 ( .A(n15936), .ZN(n19135) );
  AOI21_X1 U19125 ( .B1(n16374), .B2(n15939), .A(n9948), .ZN(n19198) );
  AOI21_X1 U19126 ( .B1(n16385), .B2(n15937), .A(n15940), .ZN(n19226) );
  OAI21_X1 U19127 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15938), .A(
        n15937), .ZN(n19234) );
  NAND2_X1 U19128 ( .A1(n19233), .A2(n19234), .ZN(n19218) );
  NOR2_X1 U19129 ( .A1(n19226), .A2(n19218), .ZN(n19211) );
  OAI21_X1 U19130 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15940), .A(
        n15939), .ZN(n19212) );
  NAND2_X1 U19131 ( .A1(n19211), .A2(n19212), .ZN(n19197) );
  NOR2_X1 U19132 ( .A1(n19198), .A2(n19197), .ZN(n19189) );
  NAND2_X1 U19133 ( .A1(n19189), .A2(n19190), .ZN(n19178) );
  NOR2_X1 U19134 ( .A1(n15941), .A2(n19178), .ZN(n19166) );
  NAND2_X1 U19135 ( .A1(n19166), .A2(n19167), .ZN(n19152) );
  NOR2_X1 U19136 ( .A1(n19154), .A2(n19152), .ZN(n19144) );
  NAND2_X1 U19137 ( .A1(n19144), .A2(n19143), .ZN(n19142) );
  NAND2_X1 U19138 ( .A1(n15010), .A2(n19142), .ZN(n19134) );
  NAND2_X1 U19139 ( .A1(n19135), .A2(n19134), .ZN(n19133) );
  NAND2_X1 U19140 ( .A1(n9843), .A2(n19133), .ZN(n15942) );
  NAND2_X1 U19141 ( .A1(n16367), .A2(n15942), .ZN(n16257) );
  OAI211_X1 U19142 ( .C1(n16367), .C2(n15942), .A(n19303), .B(n16257), .ZN(
        n15943) );
  OAI211_X1 U19143 ( .C1(n19340), .C2(n15945), .A(n15944), .B(n15943), .ZN(
        P2_U2833) );
  OAI211_X1 U19144 ( .C1(n15948), .C2(n15947), .A(n15946), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15950) );
  INV_X1 U19145 ( .A(n15950), .ZN(n15954) );
  INV_X1 U19146 ( .A(n15949), .ZN(n15952) );
  AOI22_X1 U19147 ( .A1(n15952), .A2(n15951), .B1(n20839), .B2(n15950), .ZN(
        n15953) );
  AOI21_X1 U19148 ( .B1(n15954), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15953), .ZN(n15956) );
  INV_X1 U19149 ( .A(n15956), .ZN(n15958) );
  OAI21_X1 U19150 ( .B1(n15956), .B2(n20764), .A(n15955), .ZN(n15957) );
  OAI21_X1 U19151 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15958), .A(
        n15957), .ZN(n15960) );
  AOI222_X1 U19152 ( .A1(n15960), .A2(n15959), .B1(n15960), .B2(n20804), .C1(
        n15959), .C2(n20804), .ZN(n15969) );
  INV_X1 U19153 ( .A(n15961), .ZN(n15966) );
  AOI21_X1 U19154 ( .B1(n21311), .B2(n21252), .A(n15962), .ZN(n15964) );
  NOR4_X1 U19155 ( .A1(n15966), .A2(n15965), .A3(n15964), .A4(n15963), .ZN(
        n15967) );
  OAI211_X1 U19156 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15969), .A(
        n15968), .B(n15967), .ZN(n15975) );
  NOR3_X1 U19157 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21028), .A3(n21110), 
        .ZN(n15974) );
  OR2_X1 U19158 ( .A1(n15971), .A2(n15970), .ZN(n15973) );
  OAI22_X1 U19159 ( .A1(n15976), .A2(n15974), .B1(n15973), .B2(n15972), .ZN(
        n16250) );
  AOI221_X1 U19160 ( .B1(n21026), .B2(n21025), .C1(n15975), .C2(n21025), .A(
        n16250), .ZN(n15977) );
  NOR2_X1 U19161 ( .A1(n15977), .A2(n21026), .ZN(n16253) );
  OAI211_X1 U19162 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21110), .A(n16253), 
        .B(n15979), .ZN(n16251) );
  AOI21_X1 U19163 ( .B1(n15976), .B2(n15975), .A(n16251), .ZN(n15983) );
  INV_X1 U19164 ( .A(n15977), .ZN(n15978) );
  OAI21_X1 U19165 ( .B1(n15980), .B2(n15979), .A(n15978), .ZN(n15981) );
  AOI22_X1 U19166 ( .A1(n15983), .A2(n15982), .B1(n21026), .B2(n15981), .ZN(
        P1_U3161) );
  NOR2_X1 U19167 ( .A1(n17732), .A2(n16615), .ZN(n15984) );
  NAND2_X1 U19168 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15984), .ZN(
        n16559) );
  INV_X1 U19169 ( .A(n16559), .ZN(n15986) );
  INV_X1 U19170 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16608) );
  XNOR2_X1 U19171 ( .A(n15987), .B(n16608), .ZN(n16590) );
  NOR2_X1 U19172 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16609), .ZN(
        n16585) );
  INV_X1 U19173 ( .A(n18309), .ZN(n18308) );
  NOR2_X1 U19174 ( .A1(n18308), .A2(n18392), .ZN(n18347) );
  NAND2_X1 U19175 ( .A1(n18388), .A2(n18392), .ZN(n18371) );
  OAI21_X1 U19176 ( .B1(n15988), .B2(n18392), .A(n18371), .ZN(n15989) );
  AOI21_X1 U19177 ( .B1(n18347), .B2(n15990), .A(n15989), .ZN(n16603) );
  AOI21_X1 U19178 ( .B1(n16603), .B2(n15991), .A(n16608), .ZN(n15992) );
  AOI21_X1 U19179 ( .B1(n15993), .B2(n16585), .A(n15992), .ZN(n15994) );
  NAND2_X1 U19180 ( .A1(n9832), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16580) );
  OAI211_X1 U19181 ( .C1(n16590), .C2(n18299), .A(n15994), .B(n16580), .ZN(
        P3_U2832) );
  NOR2_X1 U19182 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20232), .ZN(n21036) );
  INV_X1 U19183 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21038) );
  INV_X1 U19184 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21327) );
  AOI211_X1 U19185 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21038), .B(
        n21327), .ZN(n15995) );
  AOI211_X1 U19186 ( .C1(HOLD), .C2(n21036), .A(n15996), .B(n15995), .ZN(
        n15998) );
  NAND2_X1 U19187 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15997), .ZN(n21043) );
  NAND2_X1 U19188 ( .A1(n15998), .A2(n21043), .ZN(P1_U3195) );
  AND2_X1 U19189 ( .A1(n15999), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI221_X1 U19190 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n20216), .C1(n20218), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(
        n20072) );
  NOR3_X1 U19191 ( .A1(n16548), .A2(n16554), .A3(n20072), .ZN(P2_U3178) );
  AOI221_X1 U19192 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16554), .C1(n20205), .C2(
        n16554), .A(n19975), .ZN(n20197) );
  INV_X1 U19193 ( .A(n20197), .ZN(n20198) );
  NOR2_X1 U19194 ( .A1(n16517), .A2(n20198), .ZN(P2_U3047) );
  NAND3_X1 U19195 ( .A1(n17068), .A2(n19084), .A3(n16000), .ZN(n16001) );
  NAND2_X1 U19196 ( .A1(n17577), .A2(n17460), .ZN(n17502) );
  INV_X1 U19197 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17679) );
  INV_X1 U19198 ( .A(n16003), .ZN(n18893) );
  AOI22_X1 U19199 ( .A1(n17605), .A2(BUF2_REG_0__SCAN_IN), .B1(n17573), .B2(
        n16004), .ZN(n16005) );
  OAI221_X1 U19200 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17502), .C1(n17679), 
        .C2(n17460), .A(n16005), .ZN(P3_U2735) );
  INV_X1 U19201 ( .A(n16006), .ZN(n16007) );
  NOR3_X1 U19202 ( .A1(n20318), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n16007), 
        .ZN(n16008) );
  AOI21_X1 U19203 ( .B1(n20315), .B2(P1_EBX_REG_21__SCAN_IN), .A(n16008), .ZN(
        n16009) );
  OAI21_X1 U19204 ( .B1(n16010), .B2(n16028), .A(n16009), .ZN(n16011) );
  AOI21_X1 U19205 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n16012), .A(n16011), 
        .ZN(n16017) );
  INV_X1 U19206 ( .A(n16013), .ZN(n16014) );
  AOI22_X1 U19207 ( .A1(n16015), .A2(n20292), .B1(n16014), .B2(n20288), .ZN(
        n16016) );
  OAI211_X1 U19208 ( .C1(n16018), .C2(n20324), .A(n16017), .B(n16016), .ZN(
        P1_U2819) );
  INV_X1 U19209 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21236) );
  INV_X1 U19210 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21180) );
  NOR2_X1 U19211 ( .A1(n21236), .A2(n21180), .ZN(n16022) );
  OAI211_X1 U19212 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(P1_REIP_REG_19__SCAN_IN), .A(n16019), .B(n20270), .ZN(n16021) );
  AOI22_X1 U19213 ( .A1(n16027), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(n20315), .ZN(n16020) );
  OAI21_X1 U19214 ( .B1(n16022), .B2(n16021), .A(n16020), .ZN(n16023) );
  AOI211_X1 U19215 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20306), .B(n16023), .ZN(n16025) );
  AOI22_X1 U19216 ( .A1(n16064), .A2(n20292), .B1(n20288), .B2(n16122), .ZN(
        n16024) );
  OAI211_X1 U19217 ( .C1(n16067), .C2(n20324), .A(n16025), .B(n16024), .ZN(
        P1_U2821) );
  AOI21_X1 U19218 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n16026), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16035) );
  INV_X1 U19219 ( .A(n16027), .ZN(n16034) );
  OAI22_X1 U19220 ( .A1(n20297), .A2(n21485), .B1(n16029), .B2(n16028), .ZN(
        n16030) );
  AOI211_X1 U19221 ( .C1(n20264), .C2(n16076), .A(n20306), .B(n16030), .ZN(
        n16033) );
  INV_X1 U19222 ( .A(n16031), .ZN(n16077) );
  AOI22_X1 U19223 ( .A1(n16077), .A2(n20292), .B1(n20288), .B2(n16142), .ZN(
        n16032) );
  OAI211_X1 U19224 ( .C1(n16035), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        P1_U2823) );
  AOI22_X1 U19225 ( .A1(n16036), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n20315), .ZN(n16042) );
  AOI211_X1 U19226 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20306), .B(n16037), .ZN(n16041) );
  AOI22_X1 U19227 ( .A1(n16085), .A2(n20292), .B1(n20264), .B2(n16084), .ZN(
        n16040) );
  INV_X1 U19228 ( .A(n16038), .ZN(n16162) );
  NAND2_X1 U19229 ( .A1(n20288), .A2(n16162), .ZN(n16039) );
  NAND4_X1 U19230 ( .A1(n16042), .A2(n16041), .A3(n16040), .A4(n16039), .ZN(
        P1_U2825) );
  OAI22_X1 U19231 ( .A1(n21482), .A2(n20297), .B1(n20313), .B2(n16182), .ZN(
        n16043) );
  AOI211_X1 U19232 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20306), .B(n16043), .ZN(n16050) );
  INV_X1 U19233 ( .A(n16044), .ZN(n16045) );
  NOR2_X1 U19234 ( .A1(n20318), .A2(n16045), .ZN(n16053) );
  AOI21_X1 U19235 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16053), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16046) );
  INV_X1 U19236 ( .A(n16046), .ZN(n16047) );
  AOI22_X1 U19237 ( .A1(n16093), .A2(n20264), .B1(n16048), .B2(n16047), .ZN(
        n16049) );
  OAI211_X1 U19238 ( .C1(n16051), .C2(n16091), .A(n16050), .B(n16049), .ZN(
        P1_U2828) );
  INV_X1 U19239 ( .A(n16188), .ZN(n16052) );
  AOI22_X1 U19240 ( .A1(n16053), .A2(n21290), .B1(n20288), .B2(n16052), .ZN(
        n16058) );
  AOI22_X1 U19241 ( .A1(n20315), .A2(P1_EBX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20307), .ZN(n16054) );
  OAI21_X1 U19242 ( .B1(n16055), .B2(n21290), .A(n16054), .ZN(n16056) );
  AOI211_X1 U19243 ( .C1(n16100), .C2(n20292), .A(n20306), .B(n16056), .ZN(
        n16057) );
  OAI211_X1 U19244 ( .C1(n16103), .C2(n20324), .A(n16058), .B(n16057), .ZN(
        P1_U2829) );
  AOI22_X1 U19245 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16066) );
  INV_X1 U19246 ( .A(n16059), .ZN(n16060) );
  NOR2_X1 U19247 ( .A1(n16061), .A2(n16060), .ZN(n16062) );
  XNOR2_X1 U19248 ( .A(n16063), .B(n16062), .ZN(n16123) );
  AOI22_X1 U19249 ( .A1(n16123), .A2(n20370), .B1(n16064), .B2(n14411), .ZN(
        n16065) );
  OAI211_X1 U19250 ( .C1(n20374), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        P1_U2980) );
  NOR2_X1 U19251 ( .A1(n16081), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16074) );
  NOR2_X1 U19252 ( .A1(n16069), .A2(n16068), .ZN(n16072) );
  OAI21_X1 U19253 ( .B1(n16072), .B2(n16071), .A(n10402), .ZN(n16073) );
  MUX2_X1 U19254 ( .A(n14336), .B(n16074), .S(n16073), .Z(n16075) );
  XNOR2_X1 U19255 ( .A(n16075), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16147) );
  AOI22_X1 U19256 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16079) );
  AOI22_X1 U19257 ( .A1(n16077), .A2(n14411), .B1(n16076), .B2(n16094), .ZN(
        n16078) );
  OAI211_X1 U19258 ( .C1(n20242), .C2(n16147), .A(n16079), .B(n16078), .ZN(
        P1_U2982) );
  AOI21_X1 U19259 ( .B1(n16159), .B2(n16081), .A(n16080), .ZN(n16082) );
  XNOR2_X1 U19260 ( .A(n16083), .B(n16082), .ZN(n16164) );
  AOI22_X1 U19261 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16087) );
  AOI22_X1 U19262 ( .A1(n16085), .A2(n14411), .B1(n16094), .B2(n16084), .ZN(
        n16086) );
  OAI211_X1 U19263 ( .C1(n16164), .C2(n20242), .A(n16087), .B(n16086), .ZN(
        P1_U2984) );
  AOI21_X1 U19264 ( .B1(n16090), .B2(n16089), .A(n16088), .ZN(n16187) );
  AOI22_X1 U19265 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16096) );
  INV_X1 U19266 ( .A(n16091), .ZN(n16092) );
  AOI22_X1 U19267 ( .A1(n16094), .A2(n16093), .B1(n14411), .B2(n16092), .ZN(
        n16095) );
  OAI211_X1 U19268 ( .C1(n16187), .C2(n20242), .A(n16096), .B(n16095), .ZN(
        P1_U2987) );
  AOI22_X1 U19269 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16102) );
  NAND3_X1 U19270 ( .A1(n9893), .A2(n14805), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U19271 ( .A1(n16098), .A2(n16097), .ZN(n16099) );
  INV_X1 U19272 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16195) );
  XNOR2_X1 U19273 ( .A(n16099), .B(n16195), .ZN(n16190) );
  AOI22_X1 U19274 ( .A1(n20370), .A2(n16190), .B1(n14411), .B2(n16100), .ZN(
        n16101) );
  OAI211_X1 U19275 ( .C1(n20374), .C2(n16103), .A(n16102), .B(n16101), .ZN(
        P1_U2988) );
  AOI22_X1 U19276 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16109) );
  NAND2_X1 U19277 ( .A1(n16105), .A2(n16104), .ZN(n16106) );
  XNOR2_X1 U19278 ( .A(n16107), .B(n16106), .ZN(n16227) );
  AOI22_X1 U19279 ( .A1(n16227), .A2(n20370), .B1(n14411), .B2(n20281), .ZN(
        n16108) );
  OAI211_X1 U19280 ( .C1(n20374), .C2(n20284), .A(n16109), .B(n16108), .ZN(
        P1_U2992) );
  AOI22_X1 U19281 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16113) );
  INV_X1 U19282 ( .A(n16110), .ZN(n16111) );
  AOI22_X1 U19283 ( .A1(n16111), .A2(n20370), .B1(n14411), .B2(n20291), .ZN(
        n16112) );
  OAI211_X1 U19284 ( .C1(n20374), .C2(n20296), .A(n16113), .B(n16112), .ZN(
        P1_U2993) );
  AOI22_X1 U19285 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16119) );
  INV_X1 U19286 ( .A(n16114), .ZN(n16115) );
  AOI21_X1 U19287 ( .B1(n16117), .B2(n16116), .A(n16115), .ZN(n16236) );
  AOI22_X1 U19288 ( .A1(n16236), .A2(n20370), .B1(n14411), .B2(n20302), .ZN(
        n16118) );
  OAI211_X1 U19289 ( .C1(n20374), .C2(n20305), .A(n16119), .B(n16118), .ZN(
        P1_U2994) );
  INV_X1 U19290 ( .A(n16120), .ZN(n16121) );
  AOI22_X1 U19291 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16121), .B1(
        n20380), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U19292 ( .A1(n16123), .A2(n20405), .B1(n20404), .B2(n16122), .ZN(
        n16124) );
  OAI211_X1 U19293 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16126), .A(
        n16125), .B(n16124), .ZN(P1_U3012) );
  NAND3_X1 U19294 ( .A1(n16127), .A2(n16129), .A3(n16234), .ZN(n16160) );
  NAND2_X1 U19295 ( .A1(n16133), .A2(n16128), .ZN(n16140) );
  NOR2_X1 U19296 ( .A1(n16134), .A2(n16129), .ZN(n16131) );
  AOI211_X1 U19297 ( .C1(n20396), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        n16158) );
  OAI21_X1 U19298 ( .B1(n16134), .B2(n16133), .A(n16158), .ZN(n16144) );
  NOR2_X1 U19299 ( .A1(n16210), .A2(n21236), .ZN(n16138) );
  OAI22_X1 U19300 ( .A1(n16136), .A2(n20387), .B1(n16211), .B2(n16135), .ZN(
        n16137) );
  AOI211_X1 U19301 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16144), .A(
        n16138), .B(n16137), .ZN(n16139) );
  OAI21_X1 U19302 ( .B1(n16160), .B2(n16140), .A(n16139), .ZN(P1_U3013) );
  OAI21_X1 U19303 ( .B1(n16152), .B2(n16160), .A(n16141), .ZN(n16143) );
  AOI22_X1 U19304 ( .A1(n16144), .A2(n16143), .B1(n20404), .B2(n16142), .ZN(
        n16146) );
  NAND2_X1 U19305 ( .A1(n20380), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16145) );
  OAI211_X1 U19306 ( .C1(n16147), .C2(n20387), .A(n16146), .B(n16145), .ZN(
        P1_U3014) );
  NOR2_X1 U19307 ( .A1(n16148), .A2(n16160), .ZN(n16153) );
  OAI22_X1 U19308 ( .A1(n16150), .A2(n20387), .B1(n16211), .B2(n16149), .ZN(
        n16151) );
  AOI21_X1 U19309 ( .B1(n16153), .B2(n16152), .A(n16151), .ZN(n16155) );
  NAND2_X1 U19310 ( .A1(n20380), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n16154) );
  OAI211_X1 U19311 ( .C1(n16158), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        P1_U3015) );
  NAND2_X1 U19312 ( .A1(n20380), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16157) );
  OAI221_X1 U19313 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16160), 
        .C1(n16159), .C2(n16158), .A(n16157), .ZN(n16161) );
  AOI21_X1 U19314 ( .B1(n16162), .B2(n20404), .A(n16161), .ZN(n16163) );
  OAI21_X1 U19315 ( .B1(n16164), .B2(n20387), .A(n16163), .ZN(P1_U3016) );
  NOR2_X1 U19316 ( .A1(n16210), .A2(n21289), .ZN(n16166) );
  AOI211_X1 U19317 ( .C1(n16168), .C2(n16167), .A(n16166), .B(n16165), .ZN(
        n16172) );
  AOI22_X1 U19318 ( .A1(n16170), .A2(n20405), .B1(n20404), .B2(n16169), .ZN(
        n16171) );
  OAI211_X1 U19319 ( .C1(n16174), .C2(n16173), .A(n16172), .B(n16171), .ZN(
        P1_U3018) );
  NOR2_X1 U19320 ( .A1(n16179), .A2(n16222), .ZN(n16185) );
  AOI21_X1 U19321 ( .B1(n16192), .B2(n16176), .A(n16175), .ZN(n16178) );
  AOI211_X1 U19322 ( .C1(n16180), .C2(n16179), .A(n16178), .B(n16177), .ZN(
        n16196) );
  OAI21_X1 U19323 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16181), .A(
        n16196), .ZN(n16184) );
  OAI22_X1 U19324 ( .A1(n16211), .A2(n16182), .B1(n21453), .B2(n16210), .ZN(
        n16183) );
  AOI221_X1 U19325 ( .B1(n16185), .B2(n14818), .C1(n16184), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16183), .ZN(n16186) );
  OAI21_X1 U19326 ( .B1(n16187), .B2(n20387), .A(n16186), .ZN(P1_U3019) );
  OAI22_X1 U19327 ( .A1(n16211), .A2(n16188), .B1(n16210), .B2(n21290), .ZN(
        n16189) );
  INV_X1 U19328 ( .A(n16189), .ZN(n16194) );
  NOR2_X1 U19329 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16222), .ZN(
        n16191) );
  AOI22_X1 U19330 ( .A1(n16192), .A2(n16191), .B1(n20405), .B2(n16190), .ZN(
        n16193) );
  OAI211_X1 U19331 ( .C1(n16196), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        P1_U3020) );
  INV_X1 U19332 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16207) );
  NAND2_X1 U19333 ( .A1(n16198), .A2(n16197), .ZN(n16200) );
  OAI22_X1 U19334 ( .A1(n16219), .A2(n20395), .B1(n16199), .B2(n16200), .ZN(
        n16216) );
  OR2_X1 U19335 ( .A1(n16201), .A2(n16200), .ZN(n16209) );
  AOI221_X1 U19336 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16207), .C2(n16217), .A(
        n16209), .ZN(n16204) );
  OAI22_X1 U19337 ( .A1(n16211), .A2(n16202), .B1(n21054), .B2(n16210), .ZN(
        n16203) );
  AOI211_X1 U19338 ( .C1(n16205), .C2(n20405), .A(n16204), .B(n16203), .ZN(
        n16206) );
  OAI21_X1 U19339 ( .B1(n16207), .B2(n16216), .A(n16206), .ZN(P1_U3021) );
  INV_X1 U19340 ( .A(n16208), .ZN(n16214) );
  NOR2_X1 U19341 ( .A1(n16209), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16213) );
  INV_X1 U19342 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21326) );
  OAI22_X1 U19343 ( .A1(n16211), .A2(n20258), .B1(n21326), .B2(n16210), .ZN(
        n16212) );
  AOI211_X1 U19344 ( .C1(n16214), .C2(n20405), .A(n16213), .B(n16212), .ZN(
        n16215) );
  OAI21_X1 U19345 ( .B1(n16217), .B2(n16216), .A(n16215), .ZN(P1_U3022) );
  OAI21_X1 U19346 ( .B1(n20395), .B2(n16219), .A(n16218), .ZN(n16230) );
  AOI222_X1 U19347 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20380), .B1(n20404), 
        .B2(n16221), .C1(n20405), .C2(n16220), .ZN(n16224) );
  NOR2_X1 U19348 ( .A1(n12259), .A2(n16222), .ZN(n16226) );
  OAI221_X1 U19349 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16225), .C2(n16231), .A(
        n16226), .ZN(n16223) );
  OAI211_X1 U19350 ( .C1(n16230), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        P1_U3023) );
  AOI22_X1 U19351 ( .A1(n20404), .A2(n20269), .B1(n20380), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U19352 ( .A1(n16227), .A2(n20405), .B1(n16226), .B2(n16231), .ZN(
        n16228) );
  OAI211_X1 U19353 ( .C1(n16231), .C2(n16230), .A(n16229), .B(n16228), .ZN(
        P1_U3024) );
  AOI22_X1 U19354 ( .A1(n20404), .A2(n16232), .B1(n20380), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16238) );
  INV_X1 U19355 ( .A(n16233), .ZN(n20400) );
  NAND2_X1 U19356 ( .A1(n16234), .A2(n20400), .ZN(n20389) );
  INV_X1 U19357 ( .A(n20389), .ZN(n20382) );
  AOI22_X1 U19358 ( .A1(n16236), .A2(n20405), .B1(n20382), .B2(n16235), .ZN(
        n16237) );
  OAI211_X1 U19359 ( .C1(n16240), .C2(n16239), .A(n16238), .B(n16237), .ZN(
        P1_U3026) );
  NAND3_X1 U19360 ( .A1(n16243), .A2(n16242), .A3(n16241), .ZN(n16244) );
  OAI21_X1 U19361 ( .B1(n16245), .B2(n11600), .A(n16244), .ZN(P1_U3468) );
  NAND4_X1 U19362 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21028), .A4(n21110), .ZN(n16246) );
  AND2_X1 U19363 ( .A1(n16247), .A2(n16246), .ZN(n21027) );
  NAND2_X1 U19364 ( .A1(n21027), .A2(n16248), .ZN(n16249) );
  AOI22_X1 U19365 ( .A1(n21025), .A2(n16251), .B1(n16250), .B2(n16249), .ZN(
        P1_U3162) );
  OAI21_X1 U19366 ( .B1(n16253), .B2(n20847), .A(n16252), .ZN(P1_U3466) );
  INV_X1 U19367 ( .A(n16254), .ZN(n16285) );
  INV_X1 U19368 ( .A(n16255), .ZN(n16329) );
  INV_X1 U19369 ( .A(n16256), .ZN(n16351) );
  NAND2_X1 U19370 ( .A1(n9843), .A2(n16257), .ZN(n16350) );
  NAND2_X1 U19371 ( .A1(n16351), .A2(n16350), .ZN(n16349) );
  NAND2_X1 U19372 ( .A1(n9843), .A2(n16349), .ZN(n16339) );
  NAND2_X1 U19373 ( .A1(n16340), .A2(n16339), .ZN(n16338) );
  NAND2_X1 U19374 ( .A1(n9843), .A2(n16338), .ZN(n16328) );
  NAND2_X1 U19375 ( .A1(n16329), .A2(n16328), .ZN(n16327) );
  NAND2_X1 U19376 ( .A1(n9843), .A2(n16327), .ZN(n16316) );
  NAND2_X1 U19377 ( .A1(n16317), .A2(n16316), .ZN(n16315) );
  NAND2_X1 U19378 ( .A1(n9843), .A2(n16315), .ZN(n16305) );
  NAND2_X1 U19379 ( .A1(n16306), .A2(n16305), .ZN(n16304) );
  NAND2_X1 U19380 ( .A1(n9843), .A2(n16304), .ZN(n16293) );
  NAND2_X1 U19381 ( .A1(n16294), .A2(n16293), .ZN(n16292) );
  NAND2_X1 U19382 ( .A1(n15010), .A2(n16292), .ZN(n16284) );
  NAND2_X1 U19383 ( .A1(n16285), .A2(n16284), .ZN(n16283) );
  NAND2_X1 U19384 ( .A1(n9843), .A2(n16283), .ZN(n16271) );
  NAND2_X1 U19385 ( .A1(n16272), .A2(n16271), .ZN(n16270) );
  AND2_X1 U19386 ( .A1(n16258), .A2(n19346), .ZN(n16262) );
  OAI22_X1 U19387 ( .A1(n16260), .A2(n16259), .B1(n20150), .B2(n19342), .ZN(
        n16261) );
  AOI211_X1 U19388 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19324), .A(
        n16262), .B(n16261), .ZN(n16265) );
  AOI22_X1 U19389 ( .A1(n19333), .A2(n19361), .B1(n19290), .B2(n16263), .ZN(
        n16264) );
  OAI211_X1 U19390 ( .C1(n19358), .C2(n16270), .A(n16265), .B(n16264), .ZN(
        P2_U2824) );
  AOI22_X1 U19391 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19324), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19323), .ZN(n16276) );
  INV_X1 U19392 ( .A(n16266), .ZN(n16267) );
  AOI22_X1 U19393 ( .A1(n16267), .A2(n19346), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19325), .ZN(n16275) );
  AOI22_X1 U19394 ( .A1(n16269), .A2(n19290), .B1(n16268), .B2(n19333), .ZN(
        n16274) );
  OAI211_X1 U19395 ( .C1(n16272), .C2(n16271), .A(n19303), .B(n16270), .ZN(
        n16273) );
  NAND4_X1 U19396 ( .A1(n16276), .A2(n16275), .A3(n16274), .A4(n16273), .ZN(
        P2_U2825) );
  INV_X1 U19397 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20143) );
  OAI22_X1 U19398 ( .A1(n16277), .A2(n19353), .B1(n20143), .B2(n19342), .ZN(
        n16281) );
  OAI22_X1 U19399 ( .A1(n16279), .A2(n19328), .B1(n16278), .B2(n19343), .ZN(
        n16280) );
  AOI211_X1 U19400 ( .C1(n16282), .C2(n19333), .A(n16281), .B(n16280), .ZN(
        n16287) );
  OAI211_X1 U19401 ( .C1(n16285), .C2(n16284), .A(n19303), .B(n16283), .ZN(
        n16286) );
  OAI211_X1 U19402 ( .C1(n19349), .C2(n16288), .A(n16287), .B(n16286), .ZN(
        P2_U2826) );
  AOI22_X1 U19403 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19324), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19323), .ZN(n16298) );
  AOI22_X1 U19404 ( .A1(n16289), .A2(n19346), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19325), .ZN(n16297) );
  AOI22_X1 U19405 ( .A1(n16291), .A2(n19290), .B1(n16290), .B2(n19333), .ZN(
        n16296) );
  OAI211_X1 U19406 ( .C1(n16294), .C2(n16293), .A(n19303), .B(n16292), .ZN(
        n16295) );
  NAND4_X1 U19407 ( .A1(n16298), .A2(n16297), .A3(n16296), .A4(n16295), .ZN(
        P2_U2827) );
  INV_X1 U19408 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16299) );
  INV_X1 U19409 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20140) );
  OAI22_X1 U19410 ( .A1(n16299), .A2(n19353), .B1(n20140), .B2(n19342), .ZN(
        n16302) );
  OAI22_X1 U19411 ( .A1(n16300), .A2(n19328), .B1(n19343), .B2(n11195), .ZN(
        n16301) );
  AOI211_X1 U19412 ( .C1(n16303), .C2(n19333), .A(n16302), .B(n16301), .ZN(
        n16308) );
  OAI211_X1 U19413 ( .C1(n16306), .C2(n16305), .A(n19303), .B(n16304), .ZN(
        n16307) );
  OAI211_X1 U19414 ( .C1(n19349), .C2(n16309), .A(n16308), .B(n16307), .ZN(
        P2_U2828) );
  OAI22_X1 U19415 ( .A1(n15250), .A2(n19353), .B1(n20137), .B2(n19342), .ZN(
        n16313) );
  OAI22_X1 U19416 ( .A1(n16311), .A2(n19328), .B1(n19343), .B2(n16310), .ZN(
        n16312) );
  AOI211_X1 U19417 ( .C1(n16314), .C2(n19290), .A(n16313), .B(n16312), .ZN(
        n16319) );
  OAI211_X1 U19418 ( .C1(n16317), .C2(n16316), .A(n19303), .B(n16315), .ZN(
        n16318) );
  OAI211_X1 U19419 ( .C1(n19340), .C2(n16320), .A(n16319), .B(n16318), .ZN(
        P2_U2829) );
  INV_X1 U19420 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20135) );
  OAI22_X1 U19421 ( .A1(n16321), .A2(n19353), .B1(n20135), .B2(n19342), .ZN(
        n16325) );
  INV_X1 U19422 ( .A(n16322), .ZN(n16323) );
  OAI22_X1 U19423 ( .A1(n16323), .A2(n19328), .B1(n19343), .B2(n11190), .ZN(
        n16324) );
  AOI211_X1 U19424 ( .C1(n16326), .C2(n19333), .A(n16325), .B(n16324), .ZN(
        n16331) );
  OAI211_X1 U19425 ( .C1(n16329), .C2(n16328), .A(n19303), .B(n16327), .ZN(
        n16330) );
  OAI211_X1 U19426 ( .C1(n19349), .C2(n16332), .A(n16331), .B(n16330), .ZN(
        P2_U2830) );
  AOI22_X1 U19427 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19324), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19323), .ZN(n16344) );
  OAI22_X1 U19428 ( .A1(n16333), .A2(n19328), .B1(n19343), .B2(n10208), .ZN(
        n16334) );
  INV_X1 U19429 ( .A(n16334), .ZN(n16343) );
  INV_X1 U19430 ( .A(n16335), .ZN(n16336) );
  AOI22_X1 U19431 ( .A1(n16337), .A2(n19290), .B1(n16336), .B2(n19333), .ZN(
        n16342) );
  OAI211_X1 U19432 ( .C1(n16340), .C2(n16339), .A(n19303), .B(n16338), .ZN(
        n16341) );
  NAND4_X1 U19433 ( .A1(n16344), .A2(n16343), .A3(n16342), .A4(n16341), .ZN(
        P2_U2831) );
  OAI22_X1 U19434 ( .A1(n16345), .A2(n19353), .B1(n15287), .B2(n19342), .ZN(
        n16348) );
  OAI22_X1 U19435 ( .A1(n16346), .A2(n19328), .B1(n19343), .B2(n15074), .ZN(
        n16347) );
  AOI211_X1 U19436 ( .C1(n16356), .C2(n19333), .A(n16348), .B(n16347), .ZN(
        n16353) );
  OAI211_X1 U19437 ( .C1(n16351), .C2(n16350), .A(n19303), .B(n16349), .ZN(
        n16352) );
  OAI211_X1 U19438 ( .C1(n19349), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        P2_U2832) );
  AOI22_X1 U19439 ( .A1(n19367), .A2(n16355), .B1(n19427), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16360) );
  AOI22_X1 U19440 ( .A1(n19360), .A2(BUF2_REG_23__SCAN_IN), .B1(n19362), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19441 ( .A1(n16357), .A2(n19429), .B1(n19428), .B2(n16356), .ZN(
        n16358) );
  NAND3_X1 U19442 ( .A1(n16360), .A2(n16359), .A3(n16358), .ZN(P2_U2896) );
  AOI22_X1 U19443 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19310), .ZN(n16366) );
  OAI22_X1 U19444 ( .A1(n16362), .A2(n19493), .B1(n19501), .B2(n16361), .ZN(
        n16363) );
  AOI21_X1 U19445 ( .B1(n19510), .B2(n16364), .A(n16363), .ZN(n16365) );
  OAI211_X1 U19446 ( .C1(n19503), .C2(n16367), .A(n16366), .B(n16365), .ZN(
        P2_U2992) );
  AOI22_X1 U19447 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n19198), .ZN(n16373) );
  INV_X1 U19448 ( .A(n16368), .ZN(n16371) );
  INV_X1 U19449 ( .A(n19203), .ZN(n16370) );
  AOI222_X1 U19450 ( .A1(n16371), .A2(n19504), .B1(n19510), .B2(n16370), .C1(
        n16449), .C2(n16369), .ZN(n16372) );
  OAI211_X1 U19451 ( .C1(n16374), .C2(n19514), .A(n16373), .B(n16372), .ZN(
        P2_U2999) );
  AOI22_X1 U19452 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19310), .ZN(n16379) );
  OAI22_X1 U19453 ( .A1(n16376), .A2(n19493), .B1(n19501), .B2(n16375), .ZN(
        n16377) );
  AOI21_X1 U19454 ( .B1(n19510), .B2(n19214), .A(n16377), .ZN(n16378) );
  OAI211_X1 U19455 ( .C1(n19503), .C2(n19212), .A(n16379), .B(n16378), .ZN(
        P2_U3000) );
  AOI22_X1 U19456 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n19226), .ZN(n16384) );
  INV_X1 U19457 ( .A(n19229), .ZN(n16381) );
  AOI222_X1 U19458 ( .A1(n16382), .A2(n19504), .B1(n19510), .B2(n16381), .C1(
        n16449), .C2(n16380), .ZN(n16383) );
  OAI211_X1 U19459 ( .C1(n16385), .C2(n19514), .A(n16384), .B(n16383), .ZN(
        P2_U3001) );
  AOI22_X1 U19460 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19310), .ZN(n16390) );
  OAI22_X1 U19461 ( .A1(n16387), .A2(n19493), .B1(n16386), .B2(n19501), .ZN(
        n16388) );
  AOI21_X1 U19462 ( .B1(n19510), .B2(n19237), .A(n16388), .ZN(n16389) );
  OAI211_X1 U19463 ( .C1(n19503), .C2(n19234), .A(n16390), .B(n16389), .ZN(
        P2_U3002) );
  AOI22_X1 U19464 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n16391), .ZN(n16406) );
  AOI21_X1 U19465 ( .B1(n16413), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16393) );
  OR2_X1 U19466 ( .A1(n16393), .A2(n16392), .ZN(n16458) );
  INV_X1 U19467 ( .A(n16394), .ZN(n16395) );
  NAND2_X1 U19468 ( .A1(n16396), .A2(n16395), .ZN(n16400) );
  OR2_X1 U19469 ( .A1(n16398), .A2(n16397), .ZN(n16399) );
  XNOR2_X1 U19470 ( .A(n16400), .B(n16399), .ZN(n16453) );
  NAND2_X1 U19471 ( .A1(n16453), .A2(n19504), .ZN(n16403) );
  INV_X1 U19472 ( .A(n16401), .ZN(n16454) );
  NAND2_X1 U19473 ( .A1(n19510), .A2(n16454), .ZN(n16402) );
  OAI211_X1 U19474 ( .C1(n16458), .C2(n19501), .A(n16403), .B(n16402), .ZN(
        n16404) );
  INV_X1 U19475 ( .A(n16404), .ZN(n16405) );
  OAI211_X1 U19476 ( .C1(n16407), .C2(n19514), .A(n16406), .B(n16405), .ZN(
        P2_U3003) );
  AOI22_X1 U19477 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19310), .ZN(n16412) );
  OAI22_X1 U19478 ( .A1(n16409), .A2(n19501), .B1(n16408), .B2(n19493), .ZN(
        n16410) );
  AOI21_X1 U19479 ( .B1(n19510), .B2(n19247), .A(n16410), .ZN(n16411) );
  OAI211_X1 U19480 ( .C1(n19503), .C2(n19244), .A(n16412), .B(n16411), .ZN(
        P2_U3004) );
  AOI22_X1 U19481 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n19256), .ZN(n16419) );
  NOR3_X1 U19482 ( .A1(n16414), .A2(n16413), .A3(n19501), .ZN(n16417) );
  OAI22_X1 U19483 ( .A1(n16415), .A2(n19493), .B1(n16438), .B2(n19260), .ZN(
        n16416) );
  NOR2_X1 U19484 ( .A1(n16417), .A2(n16416), .ZN(n16418) );
  OAI211_X1 U19485 ( .C1(n19252), .C2(n19514), .A(n16419), .B(n16418), .ZN(
        P2_U3005) );
  AOI22_X1 U19486 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19310), .ZN(n16433) );
  XOR2_X1 U19487 ( .A(n16421), .B(n16420), .Z(n16474) );
  INV_X1 U19488 ( .A(n16474), .ZN(n16430) );
  INV_X1 U19489 ( .A(n16422), .ZN(n16423) );
  AOI21_X1 U19490 ( .B1(n16425), .B2(n16424), .A(n16423), .ZN(n16429) );
  NAND2_X1 U19491 ( .A1(n16427), .A2(n16426), .ZN(n16428) );
  XNOR2_X1 U19492 ( .A(n16429), .B(n16428), .ZN(n16478) );
  OAI22_X1 U19493 ( .A1(n16430), .A2(n19501), .B1(n16478), .B2(n19493), .ZN(
        n16431) );
  AOI21_X1 U19494 ( .B1(n19510), .B2(n19267), .A(n16431), .ZN(n16432) );
  OAI211_X1 U19495 ( .C1(n19503), .C2(n19265), .A(n16433), .B(n16432), .ZN(
        P2_U3006) );
  AOI22_X1 U19496 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n19277), .ZN(n16441) );
  NAND2_X1 U19497 ( .A1(n16434), .A2(n16449), .ZN(n16437) );
  NAND2_X1 U19498 ( .A1(n16435), .A2(n19504), .ZN(n16436) );
  OAI211_X1 U19499 ( .C1(n16438), .C2(n19281), .A(n16437), .B(n16436), .ZN(
        n16439) );
  INV_X1 U19500 ( .A(n16439), .ZN(n16440) );
  OAI211_X1 U19501 ( .C1(n19273), .C2(n19514), .A(n16441), .B(n16440), .ZN(
        P2_U3007) );
  AOI22_X1 U19502 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19310), .B1(n16442), 
        .B2(n19301), .ZN(n16451) );
  NAND2_X1 U19503 ( .A1(n16444), .A2(n16443), .ZN(n16446) );
  XNOR2_X1 U19504 ( .A(n16446), .B(n16445), .ZN(n16494) );
  INV_X1 U19505 ( .A(n19306), .ZN(n16491) );
  XOR2_X1 U19506 ( .A(n16448), .B(n16447), .Z(n16489) );
  AOI222_X1 U19507 ( .A1(n16494), .A2(n16449), .B1(n19510), .B2(n16491), .C1(
        n19504), .C2(n16489), .ZN(n16450) );
  OAI211_X1 U19508 ( .C1(n19295), .C2(n19514), .A(n16451), .B(n16450), .ZN(
        P2_U3009) );
  AOI22_X1 U19509 ( .A1(n16452), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16485), .B2(n19380), .ZN(n16465) );
  NAND2_X1 U19510 ( .A1(n16453), .A2(n16490), .ZN(n16456) );
  NAND2_X1 U19511 ( .A1(n16492), .A2(n16454), .ZN(n16455) );
  OAI211_X1 U19512 ( .C1(n16458), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        n16459) );
  INV_X1 U19513 ( .A(n16459), .ZN(n16464) );
  NAND2_X1 U19514 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19310), .ZN(n16463) );
  OAI211_X1 U19515 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16461), .B(n16460), .ZN(
        n16462) );
  NAND4_X1 U19516 ( .A1(n16465), .A2(n16464), .A3(n16463), .A4(n16462), .ZN(
        P2_U3035) );
  AOI221_X1 U19517 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n13927), .C2(n16470), .A(
        n16466), .ZN(n16473) );
  OAI21_X1 U19518 ( .B1(n16468), .B2(n13932), .A(n16467), .ZN(n19390) );
  OAI22_X1 U19519 ( .A1(n16471), .A2(n16470), .B1(n16469), .B2(n19390), .ZN(
        n16472) );
  AOI211_X1 U19520 ( .C1(n19310), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16473), .B(
        n16472), .ZN(n16476) );
  AOI22_X1 U19521 ( .A1(n16474), .A2(n16493), .B1(n16492), .B2(n19267), .ZN(
        n16475) );
  OAI211_X1 U19522 ( .C1(n16478), .C2(n16477), .A(n16476), .B(n16475), .ZN(
        P2_U3038) );
  AOI221_X1 U19523 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16480), .C2(n16497), .A(
        n16479), .ZN(n16488) );
  OR2_X1 U19524 ( .A1(n16482), .A2(n16481), .ZN(n16483) );
  AND2_X1 U19525 ( .A1(n16484), .A2(n16483), .ZN(n19397) );
  NAND2_X1 U19526 ( .A1(n16485), .A2(n19397), .ZN(n16486) );
  OAI21_X1 U19527 ( .B1(n12476), .B2(n19294), .A(n16486), .ZN(n16487) );
  NOR2_X1 U19528 ( .A1(n16488), .A2(n16487), .ZN(n16496) );
  AOI222_X1 U19529 ( .A1(n16494), .A2(n16493), .B1(n16492), .B2(n16491), .C1(
        n16490), .C2(n16489), .ZN(n16495) );
  OAI211_X1 U19530 ( .C1(n16498), .C2(n16497), .A(n16496), .B(n16495), .ZN(
        P2_U3041) );
  NOR2_X1 U19531 ( .A1(n16499), .A2(n20013), .ZN(n20210) );
  INV_X1 U19532 ( .A(n20210), .ZN(n16500) );
  NOR2_X1 U19533 ( .A1(n16501), .A2(n16500), .ZN(n16545) );
  INV_X1 U19534 ( .A(n16505), .ZN(n16537) );
  NAND2_X1 U19535 ( .A1(n16537), .A2(n16502), .ZN(n16503) );
  OAI21_X1 U19536 ( .B1(n16504), .B2(n16537), .A(n16503), .ZN(n16541) );
  MUX2_X1 U19537 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16513), .S(
        n16505), .Z(n16514) );
  INV_X1 U19538 ( .A(n16514), .ZN(n16540) );
  INV_X1 U19539 ( .A(n16508), .ZN(n16510) );
  INV_X1 U19540 ( .A(n16506), .ZN(n16507) );
  AOI211_X1 U19541 ( .C1(n16508), .C2(n20190), .A(n20199), .B(n16507), .ZN(
        n16509) );
  AOI211_X1 U19542 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16510), .A(
        n16537), .B(n16509), .ZN(n16512) );
  NAND2_X1 U19543 ( .A1(n16541), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16511) );
  OAI211_X1 U19544 ( .C1(n16513), .C2(n20181), .A(n16512), .B(n16511), .ZN(
        n16516) );
  NOR2_X1 U19545 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19573) );
  NAND2_X1 U19546 ( .A1(n16514), .A2(n19573), .ZN(n16515) );
  OAI211_X1 U19547 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n16541), .A(
        n16516), .B(n16515), .ZN(n16518) );
  NAND2_X1 U19548 ( .A1(n16518), .A2(n16517), .ZN(n16539) );
  INV_X1 U19549 ( .A(n16529), .ZN(n16520) );
  NOR4_X1 U19550 ( .A1(n16530), .A2(n16521), .A3(n16520), .A4(n16519), .ZN(
        n19107) );
  OAI21_X1 U19551 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19107), .ZN(n16526) );
  INV_X1 U19552 ( .A(n16522), .ZN(n16523) );
  NAND3_X1 U19553 ( .A1(n16524), .A2(n9838), .A3(n16523), .ZN(n16525) );
  OAI211_X1 U19554 ( .C1(n16528), .C2(n16527), .A(n16526), .B(n16525), .ZN(
        n16536) );
  OAI22_X1 U19555 ( .A1(n16534), .A2(n16531), .B1(n16530), .B2(n16529), .ZN(
        n16532) );
  AOI21_X1 U19556 ( .B1(n16534), .B2(n16533), .A(n16532), .ZN(n20207) );
  INV_X1 U19557 ( .A(n20207), .ZN(n16535) );
  AOI211_X1 U19558 ( .C1(n16537), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16536), .B(n16535), .ZN(n16538) );
  OAI211_X1 U19559 ( .C1(n16541), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        n16550) );
  OAI21_X1 U19560 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n16550), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n20073) );
  NAND2_X1 U19561 ( .A1(n16545), .A2(n20073), .ZN(n20076) );
  NOR3_X1 U19562 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20218), .A3(n20216), 
        .ZN(n16543) );
  AOI211_X1 U19563 ( .C1(n16544), .C2(n16554), .A(n16543), .B(n16542), .ZN(
        n16553) );
  INV_X1 U19564 ( .A(n16545), .ZN(n16546) );
  NOR2_X1 U19565 ( .A1(n20216), .A2(n16546), .ZN(n20074) );
  AOI211_X1 U19566 ( .C1(n16548), .C2(n16547), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n20074), .ZN(n16549) );
  AOI21_X1 U19567 ( .B1(n16551), .B2(n16550), .A(n16549), .ZN(n16552) );
  OAI211_X1 U19568 ( .C1(n20218), .C2(n20076), .A(n16553), .B(n16552), .ZN(
        P2_U3176) );
  AOI21_X1 U19569 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20218), .A(n16554), 
        .ZN(n16555) );
  OAI21_X1 U19570 ( .B1(n12466), .B2(n20076), .A(n16555), .ZN(P2_U3593) );
  OAI21_X1 U19571 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15863), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16558) );
  OAI221_X1 U19572 ( .B1(n16608), .B2(n16559), .C1(n15863), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16558), .ZN(n16564) );
  OAI21_X1 U19573 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16608), .A(
        n16559), .ZN(n16562) );
  NAND2_X1 U19574 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15863), .ZN(
        n16560) );
  OAI22_X1 U19575 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15863), .B1(
        n16560), .B2(n16608), .ZN(n16561) );
  OAI21_X1 U19576 ( .B1(n16565), .B2(n16562), .A(n16561), .ZN(n16563) );
  OAI21_X1 U19577 ( .B1(n16565), .B2(n16564), .A(n16563), .ZN(n16614) );
  INV_X1 U19578 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16597) );
  NAND2_X1 U19579 ( .A1(n18045), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18024) );
  NAND4_X1 U19580 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17940) );
  NOR2_X1 U19581 ( .A1(n17932), .A2(n17914), .ZN(n17916) );
  NAND2_X1 U19582 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17876) );
  NAND2_X1 U19583 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17836) );
  NAND2_X1 U19584 ( .A1(n17824), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17805) );
  NAND2_X1 U19585 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17806) );
  NAND2_X1 U19586 ( .A1(n16760), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17760) );
  NAND2_X1 U19587 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17761) );
  NAND2_X1 U19588 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17727) );
  NAND2_X1 U19589 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16595), .ZN(
        n16567) );
  INV_X1 U19590 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19012) );
  NOR2_X1 U19591 ( .A1(n19012), .A2(n18388), .ZN(n16605) );
  NAND2_X1 U19592 ( .A1(n9967), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16568) );
  INV_X1 U19593 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18077) );
  NAND2_X1 U19594 ( .A1(n18923), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18936) );
  OR2_X1 U19595 ( .A1(n16568), .A2(n17875), .ZN(n16582) );
  INV_X1 U19596 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16773) );
  XOR2_X1 U19597 ( .A(n16773), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16570) );
  NOR2_X1 U19598 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17823), .ZN(
        n16598) );
  INV_X1 U19599 ( .A(n16596), .ZN(n16753) );
  NAND2_X1 U19600 ( .A1(n18741), .A2(n16568), .ZN(n16569) );
  OAI211_X1 U19601 ( .C1(n16753), .C2(n18936), .A(n18083), .B(n16569), .ZN(
        n16599) );
  NOR2_X1 U19602 ( .A1(n16598), .A2(n16599), .ZN(n16581) );
  OAI22_X1 U19603 ( .A1(n16582), .A2(n16570), .B1(n16581), .B2(n16773), .ZN(
        n16571) );
  AOI211_X1 U19604 ( .C1(n17929), .C2(n17045), .A(n16605), .B(n16571), .ZN(
        n16576) );
  NOR2_X2 U19605 ( .A1(n16619), .A2(n18086), .ZN(n17911) );
  NAND2_X1 U19606 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16577), .ZN(
        n16572) );
  XNOR2_X1 U19607 ( .A(n16572), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16610) );
  NOR2_X2 U19608 ( .A1(n18416), .A2(n16733), .ZN(n17999) );
  NAND2_X1 U19609 ( .A1(n16573), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16574) );
  XNOR2_X1 U19610 ( .A(n16574), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16606) );
  AOI22_X1 U19611 ( .A1(n17911), .A2(n16610), .B1(n17999), .B2(n16606), .ZN(
        n16575) );
  OAI211_X1 U19612 ( .C1(n17978), .C2(n16614), .A(n16576), .B(n16575), .ZN(
        P3_U2799) );
  XOR2_X1 U19613 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16595), .Z(
        n16776) );
  NOR2_X1 U19614 ( .A1(n17992), .A2(n16577), .ZN(n16594) );
  INV_X1 U19615 ( .A(n16594), .ZN(n16579) );
  NAND2_X1 U19616 ( .A1(n17999), .A2(n16578), .ZN(n16591) );
  AOI21_X1 U19617 ( .B1(n16579), .B2(n16591), .A(n16608), .ZN(n16584) );
  INV_X1 U19618 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16777) );
  OAI221_X1 U19619 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16582), .C1(
        n16777), .C2(n16581), .A(n16580), .ZN(n16583) );
  AOI211_X1 U19620 ( .C1(n17929), .C2(n16776), .A(n16584), .B(n16583), .ZN(
        n16589) );
  INV_X2 U19621 ( .A(n17999), .ZN(n18088) );
  NAND4_X1 U19622 ( .A1(n16587), .A2(n16586), .A3(n17794), .A4(n16585), .ZN(
        n16588) );
  OAI211_X1 U19623 ( .C1(n16590), .C2(n17978), .A(n16589), .B(n16588), .ZN(
        P3_U2800) );
  NOR2_X1 U19624 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16624), .ZN(
        n16592) );
  AOI21_X1 U19625 ( .B1(n16597), .B2(n16596), .A(n16595), .ZN(n16785) );
  OAI21_X1 U19626 ( .B1(n16598), .B2(n17929), .A(n16785), .ZN(n16601) );
  OAI221_X1 U19627 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9967), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18741), .A(n16599), .ZN(
        n16600) );
  INV_X1 U19628 ( .A(n18347), .ZN(n18378) );
  INV_X1 U19629 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19040) );
  AOI221_X1 U19630 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16603), 
        .C1(n18378), .C2(n16603), .A(n19040), .ZN(n16604) );
  AOI211_X1 U19631 ( .C1(n16606), .C2(n18322), .A(n16605), .B(n16604), .ZN(
        n16613) );
  NOR4_X1 U19632 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16609), .A3(
        n16608), .A4(n16607), .ZN(n16611) );
  OAI221_X1 U19633 ( .B1(n16611), .B2(n16610), .C1(n16611), .C2(n18248), .A(
        n18328), .ZN(n16612) );
  OAI211_X1 U19634 ( .C1(n16614), .C2(n18299), .A(n16613), .B(n16612), .ZN(
        P3_U2831) );
  AOI21_X1 U19635 ( .B1(n15863), .B2(n17732), .A(n17731), .ZN(n17723) );
  OAI21_X1 U19636 ( .B1(n15863), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16615), .ZN(n17722) );
  NOR2_X1 U19637 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17951), .ZN(
        n16616) );
  AOI22_X1 U19638 ( .A1(n17731), .A2(n18315), .B1(n18391), .B2(n16616), .ZN(
        n16630) );
  INV_X1 U19639 ( .A(n18273), .ZN(n17947) );
  AOI22_X1 U19640 ( .A1(n18868), .A2(n17947), .B1(n18271), .B2(n18248), .ZN(
        n18262) );
  OAI21_X1 U19641 ( .B1(n18262), .B2(n18148), .A(n16617), .ZN(n18142) );
  NAND2_X1 U19642 ( .A1(n18328), .A2(n18142), .ZN(n18165) );
  NOR2_X1 U19643 ( .A1(n18140), .A2(n18165), .ZN(n18126) );
  AND2_X1 U19644 ( .A1(n16618), .A2(n17719), .ZN(n17725) );
  AOI22_X1 U19645 ( .A1(n9832), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18126), 
        .B2(n17725), .ZN(n16629) );
  OAI211_X1 U19646 ( .C1(n16621), .C2(n17732), .A(n16620), .B(n16619), .ZN(
        n16623) );
  OAI211_X1 U19647 ( .C1(n17721), .C2(n16623), .A(n16622), .B(n18371), .ZN(
        n16627) );
  OAI22_X1 U19648 ( .A1(n16625), .A2(n18313), .B1(n16624), .B2(n10170), .ZN(
        n16626) );
  OAI211_X1 U19649 ( .C1(n16627), .C2(n16626), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n9975), .ZN(n16628) );
  OAI211_X1 U19650 ( .C1(n17721), .C2(n16630), .A(n16629), .B(n16628), .ZN(
        P3_U2834) );
  NOR3_X1 U19651 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16632) );
  NOR4_X1 U19652 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16631) );
  INV_X2 U19653 ( .A(n16717), .ZN(U215) );
  NAND4_X1 U19654 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16632), .A3(n16631), .A4(
        U215), .ZN(U213) );
  INV_X1 U19655 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19436) );
  INV_X2 U19656 ( .A(U214), .ZN(n16682) );
  INV_X1 U19657 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16720) );
  OAI222_X1 U19658 ( .A1(U212), .A2(n19436), .B1(n16685), .B2(n19563), .C1(
        U214), .C2(n16720), .ZN(U216) );
  INV_X1 U19659 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16634) );
  INV_X1 U19660 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20470) );
  INV_X1 U19661 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19439) );
  OAI222_X1 U19662 ( .A1(U214), .A2(n16634), .B1(n16685), .B2(n20470), .C1(
        U212), .C2(n19439), .ZN(U217) );
  INV_X1 U19663 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n16635) );
  INV_X1 U19664 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20462) );
  INV_X1 U19665 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19442) );
  OAI222_X1 U19666 ( .A1(U214), .A2(n16635), .B1(n16685), .B2(n20462), .C1(
        U212), .C2(n19442), .ZN(U218) );
  INV_X1 U19667 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20457) );
  INV_X2 U19668 ( .A(U212), .ZN(n16683) );
  AOI22_X1 U19669 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16682), .ZN(n16636) );
  OAI21_X1 U19670 ( .B1(n20457), .B2(n16685), .A(n16636), .ZN(U219) );
  INV_X1 U19671 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20451) );
  AOI22_X1 U19672 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16682), .ZN(n16637) );
  OAI21_X1 U19673 ( .B1(n20451), .B2(n16685), .A(n16637), .ZN(U220) );
  INV_X1 U19674 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20445) );
  AOI22_X1 U19675 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16682), .ZN(n16638) );
  OAI21_X1 U19676 ( .B1(n20445), .B2(n16685), .A(n16638), .ZN(U221) );
  INV_X1 U19677 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U19678 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16682), .ZN(n16639) );
  OAI21_X1 U19679 ( .B1(n20439), .B2(n16685), .A(n16639), .ZN(U222) );
  AOI22_X1 U19680 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16682), .ZN(n16640) );
  OAI21_X1 U19681 ( .B1(n20421), .B2(n16685), .A(n16640), .ZN(U223) );
  INV_X1 U19682 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16642) );
  AOI22_X1 U19683 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16682), .ZN(n16641) );
  OAI21_X1 U19684 ( .B1(n16642), .B2(n16685), .A(n16641), .ZN(U224) );
  INV_X1 U19685 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16644) );
  AOI22_X1 U19686 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16682), .ZN(n16643) );
  OAI21_X1 U19687 ( .B1(n16644), .B2(n16685), .A(n16643), .ZN(U225) );
  AOI22_X1 U19688 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16682), .ZN(n16645) );
  OAI21_X1 U19689 ( .B1(n15190), .B2(n16685), .A(n16645), .ZN(U226) );
  INV_X1 U19690 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19540) );
  AOI22_X1 U19691 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16682), .ZN(n16646) );
  OAI21_X1 U19692 ( .B1(n19540), .B2(n16685), .A(n16646), .ZN(U227) );
  AOI22_X1 U19693 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16682), .ZN(n16647) );
  OAI21_X1 U19694 ( .B1(n14029), .B2(n16685), .A(n16647), .ZN(U228) );
  INV_X1 U19695 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U19696 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16682), .ZN(n16648) );
  OAI21_X1 U19697 ( .B1(n16649), .B2(n16685), .A(n16648), .ZN(U229) );
  INV_X1 U19698 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16651) );
  AOI22_X1 U19699 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16682), .ZN(n16650) );
  OAI21_X1 U19700 ( .B1(n16651), .B2(n16685), .A(n16650), .ZN(U230) );
  INV_X1 U19701 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16653) );
  AOI22_X1 U19702 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16682), .ZN(n16652) );
  OAI21_X1 U19703 ( .B1(n16653), .B2(n16685), .A(n16652), .ZN(U231) );
  AOI22_X1 U19704 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16682), .ZN(n16654) );
  OAI21_X1 U19705 ( .B1(n12869), .B2(n16685), .A(n16654), .ZN(U232) );
  AOI22_X1 U19706 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16682), .ZN(n16655) );
  OAI21_X1 U19707 ( .B1(n16656), .B2(n16685), .A(n16655), .ZN(U233) );
  AOI22_X1 U19708 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16682), .ZN(n16657) );
  OAI21_X1 U19709 ( .B1(n16658), .B2(n16685), .A(n16657), .ZN(U234) );
  AOI22_X1 U19710 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16682), .ZN(n16659) );
  OAI21_X1 U19711 ( .B1(n16660), .B2(n16685), .A(n16659), .ZN(U235) );
  AOI22_X1 U19712 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16682), .ZN(n16661) );
  OAI21_X1 U19713 ( .B1(n16662), .B2(n16685), .A(n16661), .ZN(U236) );
  AOI22_X1 U19714 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16682), .ZN(n16663) );
  OAI21_X1 U19715 ( .B1(n16664), .B2(n16685), .A(n16663), .ZN(U237) );
  AOI22_X1 U19716 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16682), .ZN(n16665) );
  OAI21_X1 U19717 ( .B1(n16666), .B2(n16685), .A(n16665), .ZN(U238) );
  AOI22_X1 U19718 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16682), .ZN(n16667) );
  OAI21_X1 U19719 ( .B1(n12674), .B2(n16685), .A(n16667), .ZN(U239) );
  AOI22_X1 U19720 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16682), .ZN(n16668) );
  OAI21_X1 U19721 ( .B1(n16669), .B2(n16685), .A(n16668), .ZN(U240) );
  AOI22_X1 U19722 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16682), .ZN(n16670) );
  OAI21_X1 U19723 ( .B1(n16671), .B2(n16685), .A(n16670), .ZN(U241) );
  AOI22_X1 U19724 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16682), .ZN(n16672) );
  OAI21_X1 U19725 ( .B1(n16673), .B2(n16685), .A(n16672), .ZN(U242) );
  AOI22_X1 U19726 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16682), .ZN(n16674) );
  OAI21_X1 U19727 ( .B1(n16675), .B2(n16685), .A(n16674), .ZN(U243) );
  AOI22_X1 U19728 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16682), .ZN(n16676) );
  OAI21_X1 U19729 ( .B1(n16677), .B2(n16685), .A(n16676), .ZN(U244) );
  INV_X1 U19730 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16679) );
  AOI22_X1 U19731 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16682), .ZN(n16678) );
  OAI21_X1 U19732 ( .B1(n16679), .B2(n16685), .A(n16678), .ZN(U245) );
  AOI22_X1 U19733 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16682), .ZN(n16680) );
  OAI21_X1 U19734 ( .B1(n16681), .B2(n16685), .A(n16680), .ZN(U246) );
  AOI22_X1 U19735 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16683), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16682), .ZN(n16684) );
  OAI21_X1 U19736 ( .B1(n16686), .B2(n16685), .A(n16684), .ZN(U247) );
  OAI22_X1 U19737 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16717), .ZN(n16687) );
  INV_X1 U19738 ( .A(n16687), .ZN(U251) );
  OAI22_X1 U19739 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16717), .ZN(n16688) );
  INV_X1 U19740 ( .A(n16688), .ZN(U252) );
  INV_X1 U19741 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16689) );
  INV_X1 U19742 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18420) );
  AOI22_X1 U19743 ( .A1(n16717), .A2(n16689), .B1(n18420), .B2(U215), .ZN(U253) );
  INV_X1 U19744 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16690) );
  INV_X1 U19745 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U19746 ( .A1(n16717), .A2(n16690), .B1(n18425), .B2(U215), .ZN(U254) );
  INV_X1 U19747 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16691) );
  INV_X1 U19748 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U19749 ( .A1(n16717), .A2(n16691), .B1(n18430), .B2(U215), .ZN(U255) );
  INV_X1 U19750 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16692) );
  INV_X1 U19751 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U19752 ( .A1(n16717), .A2(n16692), .B1(n18436), .B2(U215), .ZN(U256) );
  INV_X1 U19753 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16693) );
  INV_X1 U19754 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U19755 ( .A1(n16718), .A2(n16693), .B1(n18442), .B2(U215), .ZN(U257) );
  INV_X1 U19756 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16694) );
  INV_X1 U19757 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18447) );
  AOI22_X1 U19758 ( .A1(n16718), .A2(n16694), .B1(n18447), .B2(U215), .ZN(U258) );
  OAI22_X1 U19759 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16717), .ZN(n16695) );
  INV_X1 U19760 ( .A(n16695), .ZN(U259) );
  INV_X1 U19761 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16696) );
  INV_X1 U19762 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U19763 ( .A1(n16718), .A2(n16696), .B1(n17570), .B2(U215), .ZN(U260) );
  OAI22_X1 U19764 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16717), .ZN(n16697) );
  INV_X1 U19765 ( .A(n16697), .ZN(U261) );
  INV_X1 U19766 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16698) );
  INV_X1 U19767 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17560) );
  AOI22_X1 U19768 ( .A1(n16718), .A2(n16698), .B1(n17560), .B2(U215), .ZN(U262) );
  INV_X1 U19769 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16699) );
  INV_X1 U19770 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U19771 ( .A1(n16717), .A2(n16699), .B1(n17556), .B2(U215), .ZN(U263) );
  INV_X1 U19772 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16700) );
  INV_X1 U19773 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U19774 ( .A1(n16718), .A2(n16700), .B1(n17551), .B2(U215), .ZN(U264) );
  OAI22_X1 U19775 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16717), .ZN(n16701) );
  INV_X1 U19776 ( .A(n16701), .ZN(U265) );
  OAI22_X1 U19777 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16718), .ZN(n16702) );
  INV_X1 U19778 ( .A(n16702), .ZN(U266) );
  OAI22_X1 U19779 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16718), .ZN(n16703) );
  INV_X1 U19780 ( .A(n16703), .ZN(U267) );
  OAI22_X1 U19781 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16718), .ZN(n16704) );
  INV_X1 U19782 ( .A(n16704), .ZN(U268) );
  OAI22_X1 U19783 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16717), .ZN(n16705) );
  INV_X1 U19784 ( .A(n16705), .ZN(U269) );
  INV_X1 U19785 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16706) );
  AOI22_X1 U19786 ( .A1(n16717), .A2(n16706), .B1(n14030), .B2(U215), .ZN(U270) );
  INV_X1 U19787 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16707) );
  INV_X1 U19788 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19539) );
  AOI22_X1 U19789 ( .A1(n16717), .A2(n16707), .B1(n19539), .B2(U215), .ZN(U271) );
  INV_X1 U19790 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16708) );
  AOI22_X1 U19791 ( .A1(n16717), .A2(n16708), .B1(n15192), .B2(U215), .ZN(U272) );
  OAI22_X1 U19792 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16717), .ZN(n16709) );
  INV_X1 U19793 ( .A(n16709), .ZN(U273) );
  OAI22_X1 U19794 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16717), .ZN(n16710) );
  INV_X1 U19795 ( .A(n16710), .ZN(U274) );
  INV_X1 U19796 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16711) );
  AOI22_X1 U19797 ( .A1(n16717), .A2(n16711), .B1(n18409), .B2(U215), .ZN(U275) );
  INV_X1 U19798 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16712) );
  INV_X1 U19799 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19525) );
  AOI22_X1 U19800 ( .A1(n16718), .A2(n16712), .B1(n19525), .B2(U215), .ZN(U276) );
  INV_X1 U19801 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n16713) );
  INV_X1 U19802 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19530) );
  AOI22_X1 U19803 ( .A1(n16717), .A2(n16713), .B1(n19530), .B2(U215), .ZN(U277) );
  OAI22_X1 U19804 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16717), .ZN(n16715) );
  INV_X1 U19805 ( .A(n16715), .ZN(U278) );
  INV_X1 U19806 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16716) );
  INV_X1 U19807 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U19808 ( .A1(n16717), .A2(n16716), .B1(n18431), .B2(U215), .ZN(U279) );
  INV_X1 U19809 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19546) );
  AOI22_X1 U19810 ( .A1(n16717), .A2(n19442), .B1(n19546), .B2(U215), .ZN(U280) );
  INV_X1 U19811 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19553) );
  AOI22_X1 U19812 ( .A1(n16717), .A2(n19439), .B1(n19553), .B2(U215), .ZN(U281) );
  INV_X1 U19813 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19561) );
  AOI22_X1 U19814 ( .A1(n16718), .A2(n19436), .B1(n19561), .B2(U215), .ZN(U282) );
  INV_X1 U19815 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16719) );
  AOI222_X1 U19816 ( .A1(n19436), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16720), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16719), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16721) );
  INV_X2 U19817 ( .A(n16723), .ZN(n16722) );
  INV_X1 U19818 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18972) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U19820 ( .A1(n16722), .A2(n18972), .B1(n20111), .B2(n16723), .ZN(
        U347) );
  INV_X1 U19821 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18970) );
  INV_X1 U19822 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U19823 ( .A1(n16722), .A2(n18970), .B1(n20110), .B2(n16723), .ZN(
        U348) );
  INV_X1 U19824 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18967) );
  INV_X1 U19825 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U19826 ( .A1(n16722), .A2(n18967), .B1(n20109), .B2(n16723), .ZN(
        U349) );
  INV_X1 U19827 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18966) );
  INV_X1 U19828 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U19829 ( .A1(n16722), .A2(n18966), .B1(n20107), .B2(n16723), .ZN(
        U350) );
  INV_X1 U19830 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18964) );
  INV_X1 U19831 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20105) );
  AOI22_X1 U19832 ( .A1(n16722), .A2(n18964), .B1(n20105), .B2(n16723), .ZN(
        U351) );
  INV_X1 U19833 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18961) );
  INV_X1 U19834 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20104) );
  AOI22_X1 U19835 ( .A1(n16722), .A2(n18961), .B1(n20104), .B2(n16723), .ZN(
        U352) );
  INV_X1 U19836 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18960) );
  INV_X1 U19837 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U19838 ( .A1(n16722), .A2(n18960), .B1(n20103), .B2(n16723), .ZN(
        U353) );
  INV_X1 U19839 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18958) );
  AOI22_X1 U19840 ( .A1(n16722), .A2(n18958), .B1(n20102), .B2(n16723), .ZN(
        U354) );
  INV_X1 U19841 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19010) );
  INV_X1 U19842 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U19843 ( .A1(n16722), .A2(n19010), .B1(n20144), .B2(n16723), .ZN(
        U356) );
  INV_X1 U19844 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19007) );
  INV_X1 U19845 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U19846 ( .A1(n16722), .A2(n19007), .B1(n20142), .B2(n16723), .ZN(
        U357) );
  INV_X1 U19847 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19006) );
  INV_X1 U19848 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U19849 ( .A1(n16722), .A2(n19006), .B1(n20139), .B2(n16723), .ZN(
        U358) );
  INV_X1 U19850 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19004) );
  INV_X1 U19851 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20138) );
  AOI22_X1 U19852 ( .A1(n16722), .A2(n19004), .B1(n20138), .B2(n16723), .ZN(
        U359) );
  INV_X1 U19853 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19002) );
  INV_X1 U19854 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20136) );
  AOI22_X1 U19855 ( .A1(n16722), .A2(n19002), .B1(n20136), .B2(n16723), .ZN(
        U360) );
  INV_X1 U19856 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19000) );
  INV_X1 U19857 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U19858 ( .A1(n16722), .A2(n19000), .B1(n20134), .B2(n16723), .ZN(
        U361) );
  INV_X1 U19859 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18997) );
  INV_X1 U19860 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U19861 ( .A1(n16722), .A2(n18997), .B1(n20132), .B2(n16723), .ZN(
        U362) );
  INV_X1 U19862 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18996) );
  INV_X1 U19863 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U19864 ( .A1(n16722), .A2(n18996), .B1(n20131), .B2(n16723), .ZN(
        U363) );
  INV_X1 U19865 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18994) );
  INV_X1 U19866 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20129) );
  AOI22_X1 U19867 ( .A1(n16722), .A2(n18994), .B1(n20129), .B2(n16723), .ZN(
        U364) );
  INV_X1 U19868 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18956) );
  INV_X1 U19869 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20101) );
  AOI22_X1 U19870 ( .A1(n16722), .A2(n18956), .B1(n20101), .B2(n16723), .ZN(
        U365) );
  INV_X1 U19871 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18991) );
  INV_X1 U19872 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20127) );
  AOI22_X1 U19873 ( .A1(n16722), .A2(n18991), .B1(n20127), .B2(n16723), .ZN(
        U366) );
  INV_X1 U19874 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18990) );
  INV_X1 U19875 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20125) );
  AOI22_X1 U19876 ( .A1(n16722), .A2(n18990), .B1(n20125), .B2(n16723), .ZN(
        U367) );
  INV_X1 U19877 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18988) );
  INV_X1 U19878 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U19879 ( .A1(n16722), .A2(n18988), .B1(n20124), .B2(n16723), .ZN(
        U368) );
  INV_X1 U19880 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18985) );
  INV_X1 U19881 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U19882 ( .A1(n16722), .A2(n18985), .B1(n20122), .B2(n16723), .ZN(
        U369) );
  INV_X1 U19883 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18984) );
  INV_X1 U19884 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U19885 ( .A1(n16722), .A2(n18984), .B1(n20120), .B2(n16723), .ZN(
        U370) );
  INV_X1 U19886 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18982) );
  INV_X1 U19887 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U19888 ( .A1(n16722), .A2(n18982), .B1(n20118), .B2(n16723), .ZN(
        U371) );
  INV_X1 U19889 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18979) );
  INV_X1 U19890 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20116) );
  AOI22_X1 U19891 ( .A1(n16722), .A2(n18979), .B1(n20116), .B2(n16723), .ZN(
        U372) );
  INV_X1 U19892 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18978) );
  INV_X1 U19893 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U19894 ( .A1(n16722), .A2(n18978), .B1(n20115), .B2(n16723), .ZN(
        U373) );
  INV_X1 U19895 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18976) );
  INV_X1 U19896 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U19897 ( .A1(n16722), .A2(n18976), .B1(n20114), .B2(n16723), .ZN(
        U374) );
  INV_X1 U19898 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18974) );
  INV_X1 U19899 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20113) );
  AOI22_X1 U19900 ( .A1(n16722), .A2(n18974), .B1(n20113), .B2(n16723), .ZN(
        U375) );
  INV_X1 U19901 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18954) );
  INV_X1 U19902 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20100) );
  AOI22_X1 U19903 ( .A1(n16722), .A2(n18954), .B1(n20100), .B2(n16723), .ZN(
        U376) );
  INV_X1 U19904 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16725) );
  INV_X1 U19905 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18953) );
  AND3_X1 U19906 ( .A1(n18953), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n16724) );
  NOR2_X1 U19907 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18939) );
  NOR2_X1 U19908 ( .A1(n16724), .A2(n18939), .ZN(n19024) );
  OAI21_X1 U19909 ( .B1(n18950), .B2(n16725), .A(n19024), .ZN(P3_U2633) );
  OAI21_X1 U19910 ( .B1(n16732), .B2(n17609), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16726) );
  OAI21_X1 U19911 ( .B1(n16727), .B2(n18925), .A(n16726), .ZN(P3_U2634) );
  AOI22_X1 U19912 ( .A1(n18939), .A2(n18953), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n19093), .ZN(n16728) );
  OAI21_X1 U19913 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19093), .A(n16728), 
        .ZN(P3_U2635) );
  INV_X1 U19914 ( .A(n19024), .ZN(n19027) );
  NOR2_X1 U19915 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16729) );
  OAI21_X1 U19916 ( .B1(n16729), .B2(BS16), .A(n19027), .ZN(n19025) );
  OAI21_X1 U19917 ( .B1(n19027), .B2(n19083), .A(n19025), .ZN(P3_U2636) );
  NOR3_X1 U19918 ( .A1(n16732), .A2(n16731), .A3(n16730), .ZN(n18911) );
  NOR2_X1 U19919 ( .A1(n18911), .A2(n19078), .ZN(n19073) );
  INV_X1 U19920 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16734) );
  OAI21_X1 U19921 ( .B1(n19073), .B2(n16734), .A(n16733), .ZN(P3_U2637) );
  NOR4_X1 U19922 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16738) );
  NOR4_X1 U19923 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16737) );
  NOR4_X1 U19924 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16736) );
  NOR4_X1 U19925 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16735) );
  NAND4_X1 U19926 ( .A1(n16738), .A2(n16737), .A3(n16736), .A4(n16735), .ZN(
        n16744) );
  NOR4_X1 U19927 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16742) );
  AOI211_X1 U19928 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16741) );
  NOR4_X1 U19929 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16740) );
  NOR4_X1 U19930 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16739) );
  NAND4_X1 U19931 ( .A1(n16742), .A2(n16741), .A3(n16740), .A4(n16739), .ZN(
        n16743) );
  NOR2_X1 U19932 ( .A1(n16744), .A2(n16743), .ZN(n19067) );
  INV_X1 U19933 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19020) );
  NOR3_X1 U19934 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16746) );
  OAI21_X1 U19935 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16746), .A(n19067), .ZN(
        n16745) );
  OAI21_X1 U19936 ( .B1(n19067), .B2(n19020), .A(n16745), .ZN(P3_U2638) );
  INV_X1 U19937 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19063) );
  INV_X1 U19938 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19026) );
  AOI21_X1 U19939 ( .B1(n19063), .B2(n19026), .A(n16746), .ZN(n16747) );
  INV_X1 U19940 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19017) );
  INV_X1 U19941 ( .A(n19067), .ZN(n19070) );
  AOI22_X1 U19942 ( .A1(n19067), .A2(n16747), .B1(n19017), .B2(n19070), .ZN(
        P3_U2639) );
  NAND2_X1 U19943 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18177), .ZN(n18926) );
  NOR2_X1 U19944 ( .A1(n9832), .A2(n17076), .ZN(n17057) );
  AOI211_X1 U19945 ( .C1(n19084), .C2(n19082), .A(n18938), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18914) );
  NOR2_X1 U19946 ( .A1(n19097), .A2(n17068), .ZN(n16749) );
  INV_X1 U19947 ( .A(n16749), .ZN(n16752) );
  AOI211_X4 U19948 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18416), .A(n18914), .B(
        n16752), .ZN(n17081) );
  INV_X1 U19949 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19014) );
  INV_X1 U19950 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18999) );
  INV_X1 U19951 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18980) );
  INV_X1 U19952 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18977) );
  INV_X1 U19953 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18973) );
  INV_X1 U19954 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18962) );
  INV_X1 U19955 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18959) );
  NAND3_X1 U19956 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17065) );
  NOR3_X1 U19957 ( .A1(n18962), .A2(n18959), .A3(n17065), .ZN(n17027) );
  NAND4_X1 U19958 ( .A1(n17027), .A2(P3_REIP_REG_8__SCAN_IN), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n16999) );
  NAND2_X1 U19959 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16980) );
  NOR3_X1 U19960 ( .A1(n18973), .A2(n16999), .A3(n16980), .ZN(n16976) );
  NAND2_X1 U19961 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16976), .ZN(n16960) );
  NOR3_X1 U19962 ( .A1(n18980), .A2(n18977), .A3(n16960), .ZN(n16859) );
  NAND3_X1 U19963 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16890) );
  NAND3_X1 U19964 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16846) );
  NOR2_X1 U19965 ( .A1(n16890), .A2(n16846), .ZN(n16860) );
  INV_X1 U19966 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18995) );
  INV_X1 U19967 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18993) );
  NOR2_X1 U19968 ( .A1(n18995), .A2(n18993), .ZN(n16864) );
  NAND4_X1 U19969 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16859), .A3(n16860), 
        .A4(n16864), .ZN(n16835) );
  NOR2_X1 U19970 ( .A1(n18999), .A2(n16835), .ZN(n16826) );
  NAND2_X1 U19971 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16826), .ZN(n16766) );
  NOR2_X1 U19972 ( .A1(n17120), .A2(n16766), .ZN(n16814) );
  NAND2_X1 U19973 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16814), .ZN(n16813) );
  NAND2_X1 U19974 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16800) );
  NOR2_X1 U19975 ( .A1(n16813), .A2(n16800), .ZN(n16790) );
  NAND2_X1 U19976 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16790), .ZN(n16765) );
  NOR3_X1 U19977 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19014), .A3(n16765), 
        .ZN(n16750) );
  AOI21_X1 U19978 ( .B1(n17081), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16750), .ZN(
        n16772) );
  NAND2_X1 U19979 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18416), .ZN(n16751) );
  AOI211_X4 U19980 ( .C1(n19083), .C2(n19085), .A(n16752), .B(n16751), .ZN(
        n17115) );
  NOR3_X1 U19981 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17095) );
  INV_X1 U19982 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17441) );
  NAND2_X1 U19983 ( .A1(n17095), .A2(n17441), .ZN(n17092) );
  NOR2_X1 U19984 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17092), .ZN(n17066) );
  INV_X1 U19985 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U19986 ( .A1(n17066), .A2(n17064), .ZN(n17061) );
  INV_X1 U19987 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17037) );
  NAND2_X1 U19988 ( .A1(n17040), .A2(n17037), .ZN(n17036) );
  NOR2_X1 U19989 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17036), .ZN(n17010) );
  NAND2_X1 U19990 ( .A1(n17010), .A2(n17013), .ZN(n16996) );
  NAND2_X1 U19991 ( .A1(n16995), .A2(n16986), .ZN(n16985) );
  NAND2_X1 U19992 ( .A1(n16970), .A2(n16964), .ZN(n16963) );
  INV_X1 U19993 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17272) );
  NAND2_X1 U19994 ( .A1(n16949), .A2(n17272), .ZN(n16943) );
  NAND2_X1 U19995 ( .A1(n16925), .A2(n17278), .ZN(n16920) );
  INV_X1 U19996 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16898) );
  NAND2_X1 U19997 ( .A1(n16905), .A2(n16898), .ZN(n16897) );
  NAND2_X1 U19998 ( .A1(n16883), .A2(n16875), .ZN(n16874) );
  NOR2_X1 U19999 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16874), .ZN(n16857) );
  NAND2_X1 U20000 ( .A1(n16857), .A2(n16851), .ZN(n16849) );
  NOR2_X1 U20001 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16849), .ZN(n16840) );
  INV_X1 U20002 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17135) );
  NAND2_X1 U20003 ( .A1(n16840), .A2(n17135), .ZN(n16831) );
  NOR2_X1 U20004 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16831), .ZN(n16815) );
  INV_X1 U20005 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16810) );
  NAND2_X1 U20006 ( .A1(n16815), .A2(n16810), .ZN(n16809) );
  NOR2_X1 U20007 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16809), .ZN(n16797) );
  INV_X1 U20008 ( .A(n16797), .ZN(n16787) );
  NOR2_X1 U20009 ( .A1(n17126), .A2(n16774), .ZN(n16780) );
  INV_X1 U20010 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17140) );
  INV_X1 U20011 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16804) );
  NAND3_X1 U20012 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16760), .A3(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16758) );
  NOR2_X1 U20013 ( .A1(n17761), .A2(n16758), .ZN(n17714) );
  INV_X1 U20014 ( .A(n17714), .ZN(n16756) );
  NOR2_X1 U20015 ( .A1(n10091), .A2(n16756), .ZN(n16755) );
  NAND2_X1 U20016 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16755), .ZN(
        n16754) );
  AOI21_X1 U20017 ( .B1(n16804), .B2(n16754), .A(n16753), .ZN(n17716) );
  OAI21_X1 U20018 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16755), .A(
        n16754), .ZN(n17735) );
  INV_X1 U20019 ( .A(n17735), .ZN(n16806) );
  AOI21_X1 U20020 ( .B1(n10091), .B2(n16756), .A(n16755), .ZN(n17748) );
  INV_X1 U20021 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U20022 ( .A1(n17775), .A2(n16758), .ZN(n16757) );
  OAI21_X1 U20023 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16757), .A(
        n16756), .ZN(n17763) );
  INV_X1 U20024 ( .A(n17763), .ZN(n16825) );
  AOI21_X1 U20025 ( .B1(n17775), .B2(n16758), .A(n16757), .ZN(n17772) );
  INV_X1 U20026 ( .A(n16758), .ZN(n17759) );
  AOI21_X1 U20027 ( .B1(n16760), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16759) );
  NOR2_X1 U20028 ( .A1(n17759), .A2(n16759), .ZN(n17788) );
  INV_X1 U20029 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16869) );
  INV_X1 U20030 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17814) );
  AND2_X1 U20031 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17824), .ZN(
        n17802) );
  NAND2_X1 U20032 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17802), .ZN(
        n16762) );
  OR2_X1 U20033 ( .A1(n17814), .A2(n16762), .ZN(n16761) );
  INV_X1 U20034 ( .A(n16760), .ZN(n17790) );
  NOR2_X1 U20035 ( .A1(n18077), .A2(n17790), .ZN(n17784) );
  AOI21_X1 U20036 ( .B1(n16869), .B2(n16761), .A(n17784), .ZN(n17804) );
  XNOR2_X1 U20037 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16762), .ZN(
        n17810) );
  OAI21_X1 U20038 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17802), .A(
        n16762), .ZN(n16763) );
  INV_X1 U20039 ( .A(n16763), .ZN(n17828) );
  NOR2_X1 U20040 ( .A1(n18077), .A2(n17874), .ZN(n17872) );
  NAND2_X1 U20041 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17872), .ZN(
        n16936) );
  OAI21_X1 U20042 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16936), .A(
        n17045), .ZN(n16937) );
  OAI21_X1 U20043 ( .B1(n17802), .B2(n9840), .A(n16937), .ZN(n16881) );
  NOR2_X1 U20044 ( .A1(n17828), .A2(n16881), .ZN(n16880) );
  NOR2_X1 U20045 ( .A1(n16880), .A2(n9840), .ZN(n16871) );
  NOR2_X1 U20046 ( .A1(n17810), .A2(n16871), .ZN(n16870) );
  NOR2_X1 U20047 ( .A1(n16870), .A2(n9840), .ZN(n16862) );
  NOR2_X1 U20048 ( .A1(n17804), .A2(n16862), .ZN(n16861) );
  NOR2_X1 U20049 ( .A1(n16861), .A2(n9840), .ZN(n16848) );
  NOR2_X1 U20050 ( .A1(n17788), .A2(n16848), .ZN(n16847) );
  NOR2_X1 U20051 ( .A1(n16847), .A2(n9840), .ZN(n16839) );
  NOR2_X1 U20052 ( .A1(n17772), .A2(n16839), .ZN(n16838) );
  NOR2_X1 U20053 ( .A1(n16838), .A2(n9840), .ZN(n16824) );
  NOR2_X1 U20054 ( .A1(n16825), .A2(n16824), .ZN(n16823) );
  NOR2_X1 U20055 ( .A1(n16823), .A2(n9840), .ZN(n16817) );
  NOR2_X1 U20056 ( .A1(n17748), .A2(n16817), .ZN(n16816) );
  NOR2_X1 U20057 ( .A1(n16795), .A2(n9840), .ZN(n16784) );
  INV_X1 U20058 ( .A(n17076), .ZN(n18931) );
  NOR4_X1 U20059 ( .A1(n16776), .A2(n16775), .A3(n9840), .A4(n18931), .ZN(
        n16770) );
  NOR2_X1 U20060 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16765), .ZN(n16779) );
  INV_X1 U20061 ( .A(n16779), .ZN(n16768) );
  INV_X1 U20062 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19003) );
  INV_X1 U20063 ( .A(n17130), .ZN(n17114) );
  OR3_X1 U20064 ( .A1(n16766), .A2(n19003), .A3(n17114), .ZN(n16794) );
  NAND3_X1 U20065 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U20066 ( .A1(n17120), .A2(n17130), .ZN(n17128) );
  OAI21_X1 U20067 ( .B1(n16794), .B2(n16767), .A(n17128), .ZN(n16793) );
  AOI21_X1 U20068 ( .B1(n16768), .B2(n16793), .A(n19012), .ZN(n16769) );
  AOI211_X1 U20069 ( .C1(n16780), .C2(n17140), .A(n16770), .B(n16769), .ZN(
        n16771) );
  OAI211_X1 U20070 ( .C1(n16773), .C2(n17116), .A(n16772), .B(n16771), .ZN(
        P3_U2640) );
  NAND2_X1 U20071 ( .A1(n17115), .A2(n16774), .ZN(n16786) );
  OAI22_X1 U20072 ( .A1(n16777), .A2(n17116), .B1(n19014), .B2(n16793), .ZN(
        n16778) );
  OAI21_X1 U20073 ( .B1(n17081), .B2(n16780), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16781) );
  OAI211_X1 U20074 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16786), .A(n16782), .B(
        n16781), .ZN(P3_U2641) );
  INV_X1 U20075 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19009) );
  AOI22_X1 U20076 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17091), .B1(
        n17081), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16792) );
  AOI211_X1 U20077 ( .C1(n16785), .C2(n16784), .A(n16783), .B(n18931), .ZN(
        n16789) );
  AOI21_X1 U20078 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16787), .A(n16786), .ZN(
        n16788) );
  AOI211_X1 U20079 ( .C1(n16790), .C2(n19009), .A(n16789), .B(n16788), .ZN(
        n16791) );
  OAI211_X1 U20080 ( .C1(n19009), .C2(n16793), .A(n16792), .B(n16791), .ZN(
        P3_U2642) );
  AND2_X1 U20081 ( .A1(n17128), .A2(n16794), .ZN(n16820) );
  AOI22_X1 U20082 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16820), .B1(n17081), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16803) );
  INV_X1 U20083 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19008) );
  INV_X1 U20084 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19005) );
  AOI21_X1 U20085 ( .B1(n19008), .B2(n19005), .A(n16813), .ZN(n16801) );
  AOI211_X1 U20086 ( .C1(n17716), .C2(n16796), .A(n16795), .B(n18931), .ZN(
        n16799) );
  AOI211_X1 U20087 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16809), .A(n16797), .B(
        n17126), .ZN(n16798) );
  AOI211_X1 U20088 ( .C1(n16801), .C2(n16800), .A(n16799), .B(n16798), .ZN(
        n16802) );
  OAI211_X1 U20089 ( .C1(n16804), .C2(n17116), .A(n16803), .B(n16802), .ZN(
        P3_U2643) );
  AOI211_X1 U20090 ( .C1(n16806), .C2(n16805), .A(n9860), .B(n18931), .ZN(
        n16808) );
  INV_X1 U20091 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17738) );
  OAI22_X1 U20092 ( .A1(n17738), .A2(n17116), .B1(n17127), .B2(n16810), .ZN(
        n16807) );
  AOI211_X1 U20093 ( .C1(n16820), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16808), 
        .B(n16807), .ZN(n16812) );
  OAI211_X1 U20094 ( .C1(n16815), .C2(n16810), .A(n17115), .B(n16809), .ZN(
        n16811) );
  OAI211_X1 U20095 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16813), .A(n16812), 
        .B(n16811), .ZN(P3_U2644) );
  AOI22_X1 U20096 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17081), .B1(n16814), 
        .B2(n19003), .ZN(n16822) );
  AOI211_X1 U20097 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16831), .A(n16815), .B(
        n17126), .ZN(n16819) );
  AOI211_X1 U20098 ( .C1(n17748), .C2(n16817), .A(n16816), .B(n18931), .ZN(
        n16818) );
  AOI211_X1 U20099 ( .C1(n16820), .C2(P3_REIP_REG_26__SCAN_IN), .A(n16819), 
        .B(n16818), .ZN(n16821) );
  OAI211_X1 U20100 ( .C1(n10091), .C2(n17116), .A(n16822), .B(n16821), .ZN(
        P3_U2645) );
  INV_X1 U20101 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16834) );
  OAI21_X1 U20102 ( .B1(n17114), .B2(n16835), .A(n17128), .ZN(n16855) );
  OAI21_X1 U20103 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17120), .A(n16855), 
        .ZN(n16830) );
  AOI211_X1 U20104 ( .C1(n16825), .C2(n16824), .A(n16823), .B(n18931), .ZN(
        n16829) );
  INV_X1 U20105 ( .A(n17120), .ZN(n17109) );
  NAND2_X1 U20106 ( .A1(n17109), .A2(n16826), .ZN(n16827) );
  OAI22_X1 U20107 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16827), .B1(n17135), 
        .B2(n17127), .ZN(n16828) );
  AOI211_X1 U20108 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16830), .A(n16829), 
        .B(n16828), .ZN(n16833) );
  OAI211_X1 U20109 ( .C1(n16840), .C2(n17135), .A(n17115), .B(n16831), .ZN(
        n16832) );
  OAI211_X1 U20110 ( .C1(n17116), .C2(n16834), .A(n16833), .B(n16832), .ZN(
        P3_U2646) );
  INV_X1 U20111 ( .A(n16835), .ZN(n16837) );
  NOR2_X1 U20112 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17120), .ZN(n16836) );
  AOI22_X1 U20113 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17091), .B1(
        n16837), .B2(n16836), .ZN(n16844) );
  AOI211_X1 U20114 ( .C1(n17772), .C2(n16839), .A(n16838), .B(n18931), .ZN(
        n16842) );
  AOI211_X1 U20115 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16849), .A(n16840), .B(
        n17126), .ZN(n16841) );
  AOI211_X1 U20116 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17081), .A(n16842), .B(
        n16841), .ZN(n16843) );
  OAI211_X1 U20117 ( .C1(n18999), .C2(n16855), .A(n16844), .B(n16843), .ZN(
        P3_U2647) );
  INV_X1 U20118 ( .A(n16890), .ZN(n16845) );
  NAND2_X1 U20119 ( .A1(n16845), .A2(n16942), .ZN(n16904) );
  NOR2_X1 U20120 ( .A1(n16846), .A2(n16904), .ZN(n16873) );
  NAND2_X1 U20121 ( .A1(n16864), .A2(n16873), .ZN(n16856) );
  INV_X1 U20122 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18998) );
  AOI211_X1 U20123 ( .C1(n17788), .C2(n16848), .A(n16847), .B(n18931), .ZN(
        n16853) );
  OAI211_X1 U20124 ( .C1(n16857), .C2(n16851), .A(n17115), .B(n16849), .ZN(
        n16850) );
  OAI21_X1 U20125 ( .B1(n16851), .B2(n17127), .A(n16850), .ZN(n16852) );
  AOI211_X1 U20126 ( .C1(n17091), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16853), .B(n16852), .ZN(n16854) );
  OAI221_X1 U20127 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n16856), .C1(n18998), 
        .C2(n16855), .A(n16854), .ZN(P3_U2648) );
  AOI211_X1 U20128 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16874), .A(n16857), .B(
        n17126), .ZN(n16858) );
  AOI21_X1 U20129 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17081), .A(n16858), .ZN(
        n16868) );
  NAND2_X1 U20130 ( .A1(n16859), .A2(n17130), .ZN(n16889) );
  INV_X1 U20131 ( .A(n16889), .ZN(n16923) );
  INV_X1 U20132 ( .A(n17128), .ZN(n16924) );
  AOI21_X1 U20133 ( .B1(n16860), .B2(n16923), .A(n16924), .ZN(n16879) );
  AOI211_X1 U20134 ( .C1(n17804), .C2(n16862), .A(n16861), .B(n18931), .ZN(
        n16866) );
  INV_X1 U20135 ( .A(n16873), .ZN(n16863) );
  AOI211_X1 U20136 ( .C1(n18995), .C2(n18993), .A(n16864), .B(n16863), .ZN(
        n16865) );
  AOI211_X1 U20137 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16879), .A(n16866), 
        .B(n16865), .ZN(n16867) );
  OAI211_X1 U20138 ( .C1(n16869), .C2(n17116), .A(n16868), .B(n16867), .ZN(
        P3_U2649) );
  AOI22_X1 U20139 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17091), .B1(
        n17081), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16878) );
  AOI211_X1 U20140 ( .C1(n17810), .C2(n16871), .A(n16870), .B(n18931), .ZN(
        n16872) );
  AOI221_X1 U20141 ( .B1(n16879), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16873), 
        .C2(n18993), .A(n16872), .ZN(n16877) );
  OAI211_X1 U20142 ( .C1(n16883), .C2(n16875), .A(n17115), .B(n16874), .ZN(
        n16876) );
  NAND3_X1 U20143 ( .A1(n16878), .A2(n16877), .A3(n16876), .ZN(P3_U2650) );
  INV_X1 U20144 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18992) );
  INV_X1 U20145 ( .A(n16879), .ZN(n16888) );
  AOI211_X1 U20146 ( .C1(n17828), .C2(n16881), .A(n16880), .B(n18931), .ZN(
        n16882) );
  AOI21_X1 U20147 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17081), .A(n16882), .ZN(
        n16887) );
  INV_X1 U20148 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18989) );
  INV_X1 U20149 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18987) );
  NOR4_X1 U20150 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18989), .A3(n18987), 
        .A4(n16904), .ZN(n16885) );
  AOI211_X1 U20151 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16897), .A(n16883), .B(
        n17126), .ZN(n16884) );
  AOI211_X1 U20152 ( .C1(n17091), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16885), .B(n16884), .ZN(n16886) );
  OAI211_X1 U20153 ( .C1(n18992), .C2(n16888), .A(n16887), .B(n16886), .ZN(
        P3_U2651) );
  NOR2_X1 U20154 ( .A1(n16890), .A2(n16889), .ZN(n16915) );
  AOI21_X1 U20155 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16915), .A(n16924), 
        .ZN(n16909) );
  NOR2_X1 U20156 ( .A1(n18987), .A2(n16904), .ZN(n16892) );
  INV_X1 U20157 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16893) );
  OAI22_X1 U20158 ( .A1(n16893), .A2(n17116), .B1(n17127), .B2(n16898), .ZN(
        n16891) );
  AOI221_X1 U20159 ( .B1(n16909), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16892), 
        .C2(n18989), .A(n16891), .ZN(n16901) );
  NOR2_X1 U20160 ( .A1(n18077), .A2(n17835), .ZN(n17834) );
  NAND2_X1 U20161 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17834), .ZN(
        n16902) );
  INV_X1 U20162 ( .A(n16937), .ZN(n16928) );
  AOI21_X1 U20163 ( .B1(n17045), .B2(n16902), .A(n16928), .ZN(n16896) );
  AOI21_X1 U20164 ( .B1(n16893), .B2(n16902), .A(n17802), .ZN(n16894) );
  INV_X1 U20165 ( .A(n16894), .ZN(n17838) );
  AOI21_X1 U20166 ( .B1(n16896), .B2(n17838), .A(n18931), .ZN(n16895) );
  OAI21_X1 U20167 ( .B1(n16896), .B2(n17838), .A(n16895), .ZN(n16900) );
  OAI211_X1 U20168 ( .C1(n16905), .C2(n16898), .A(n17115), .B(n16897), .ZN(
        n16899) );
  NAND4_X1 U20169 ( .A1(n16901), .A2(n9975), .A3(n16900), .A4(n16899), .ZN(
        P3_U2652) );
  INV_X1 U20170 ( .A(n17834), .ZN(n16912) );
  AOI21_X1 U20171 ( .B1(n17045), .B2(n16912), .A(n16928), .ZN(n16903) );
  OAI21_X1 U20172 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17834), .A(
        n16902), .ZN(n17847) );
  XNOR2_X1 U20173 ( .A(n16903), .B(n17847), .ZN(n16911) );
  NAND2_X1 U20174 ( .A1(n18987), .A2(n16904), .ZN(n16908) );
  AOI211_X1 U20175 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16920), .A(n16905), .B(
        n17126), .ZN(n16907) );
  INV_X1 U20176 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17850) );
  OAI22_X1 U20177 ( .A1(n17850), .A2(n17116), .B1(n17127), .B2(n17274), .ZN(
        n16906) );
  AOI211_X1 U20178 ( .C1(n16909), .C2(n16908), .A(n16907), .B(n16906), .ZN(
        n16910) );
  OAI211_X1 U20179 ( .C1(n18931), .C2(n16911), .A(n16910), .B(n9975), .ZN(
        P3_U2653) );
  NOR2_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18077), .ZN(
        n17087) );
  AOI21_X1 U20181 ( .B1(n9966), .B2(n17087), .A(n9840), .ZN(n16913) );
  AND2_X1 U20182 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9966), .ZN(
        n16926) );
  OAI21_X1 U20183 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16926), .A(
        n16912), .ZN(n17868) );
  XOR2_X1 U20184 ( .A(n16913), .B(n17868), .Z(n16914) );
  OAI21_X1 U20185 ( .B1(n18931), .B2(n16914), .A(n18388), .ZN(n16919) );
  AND3_X1 U20186 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n16942), .ZN(n16917) );
  NOR2_X1 U20187 ( .A1(n16924), .A2(n16915), .ZN(n16916) );
  MUX2_X1 U20188 ( .A(n16917), .B(n16916), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16918) );
  AOI211_X1 U20189 ( .C1(n17091), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16919), .B(n16918), .ZN(n16922) );
  OAI211_X1 U20190 ( .C1(n16925), .C2(n17278), .A(n17115), .B(n16920), .ZN(
        n16921) );
  OAI211_X1 U20191 ( .C1(n17278), .C2(n17127), .A(n16922), .B(n16921), .ZN(
        P3_U2654) );
  NAND2_X1 U20192 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16942), .ZN(n16935) );
  INV_X1 U20193 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18983) );
  INV_X1 U20194 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18981) );
  NOR2_X1 U20195 ( .A1(n16924), .A2(n16923), .ZN(n16951) );
  AOI21_X1 U20196 ( .B1(n16942), .B2(n18981), .A(n16951), .ZN(n16934) );
  AOI211_X1 U20197 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16943), .A(n16925), .B(
        n17126), .ZN(n16932) );
  INV_X1 U20198 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16929) );
  AOI21_X1 U20199 ( .B1(n16929), .B2(n16936), .A(n16926), .ZN(n17873) );
  INV_X1 U20200 ( .A(n17873), .ZN(n16927) );
  AOI221_X1 U20201 ( .B1(n16937), .B2(n17873), .C1(n16928), .C2(n16927), .A(
        n9832), .ZN(n16930) );
  OAI22_X1 U20202 ( .A1(n17057), .A2(n16930), .B1(n16929), .B2(n17116), .ZN(
        n16931) );
  AOI211_X1 U20203 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17081), .A(n16932), .B(
        n16931), .ZN(n16933) );
  OAI221_X1 U20204 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16935), .C1(n18983), 
        .C2(n16934), .A(n16933), .ZN(P3_U2655) );
  INV_X1 U20205 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17887) );
  NAND2_X1 U20206 ( .A1(n17045), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17117) );
  NAND2_X1 U20207 ( .A1(n17076), .A2(n17117), .ZN(n17119) );
  AOI21_X1 U20208 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17045), .A(
        n17119), .ZN(n16939) );
  OAI21_X1 U20209 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17872), .A(
        n16936), .ZN(n17883) );
  OAI21_X1 U20210 ( .B1(n18931), .B2(n16937), .A(n17883), .ZN(n16938) );
  OAI21_X1 U20211 ( .B1(n16939), .B2(n17883), .A(n16938), .ZN(n16940) );
  OAI211_X1 U20212 ( .C1(n17887), .C2(n17116), .A(n16940), .B(n18388), .ZN(
        n16941) );
  AOI221_X1 U20213 ( .B1(n16951), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16942), 
        .C2(n18981), .A(n16941), .ZN(n16945) );
  OAI211_X1 U20214 ( .C1(n16949), .C2(n17272), .A(n17115), .B(n16943), .ZN(
        n16944) );
  OAI211_X1 U20215 ( .C1(n17272), .C2(n17127), .A(n16945), .B(n16944), .ZN(
        P3_U2656) );
  NAND2_X1 U20216 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17927), .ZN(
        n17913) );
  INV_X1 U20217 ( .A(n17913), .ZN(n16972) );
  AND2_X1 U20218 ( .A1(n17916), .A2(n16972), .ZN(n16958) );
  INV_X1 U20219 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17052) );
  AOI21_X1 U20220 ( .B1(n16958), .B2(n17052), .A(n9840), .ZN(n16947) );
  INV_X1 U20221 ( .A(n17872), .ZN(n16946) );
  OAI21_X1 U20222 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16958), .A(
        n16946), .ZN(n17896) );
  XNOR2_X1 U20223 ( .A(n16947), .B(n17896), .ZN(n16948) );
  AOI22_X1 U20224 ( .A1(n17081), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n17076), 
        .B2(n16948), .ZN(n16955) );
  AOI211_X1 U20225 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16963), .A(n16949), .B(
        n17126), .ZN(n16950) );
  AOI21_X1 U20226 ( .B1(n17091), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16950), .ZN(n16954) );
  NOR3_X1 U20227 ( .A1(n17120), .A2(n18977), .A3(n16960), .ZN(n16952) );
  OAI21_X1 U20228 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16952), .A(n16951), 
        .ZN(n16953) );
  NAND4_X1 U20229 ( .A1(n16955), .A2(n16954), .A3(n9975), .A4(n16953), .ZN(
        P3_U2657) );
  NAND2_X1 U20230 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16972), .ZN(
        n16956) );
  AOI21_X1 U20231 ( .B1(n17914), .B2(n16956), .A(n16958), .ZN(n17918) );
  NAND2_X1 U20232 ( .A1(n17045), .A2(n17076), .ZN(n16957) );
  AOI211_X1 U20233 ( .C1(n16958), .C2(n17052), .A(n17918), .B(n16957), .ZN(
        n16969) );
  OAI21_X1 U20234 ( .B1(n17914), .B2(n9840), .A(n17918), .ZN(n16959) );
  OAI22_X1 U20235 ( .A1(n17127), .A2(n16964), .B1(n17119), .B2(n16959), .ZN(
        n16968) );
  OR2_X1 U20236 ( .A1(n17120), .A2(n16960), .ZN(n16962) );
  NOR2_X1 U20237 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17120), .ZN(n16975) );
  OAI21_X1 U20238 ( .B1(n16976), .B2(n17120), .A(n17130), .ZN(n16983) );
  NOR2_X1 U20239 ( .A1(n16975), .A2(n16983), .ZN(n16961) );
  MUX2_X1 U20240 ( .A(n16962), .B(n16961), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n16966) );
  OAI211_X1 U20241 ( .C1(n16970), .C2(n16964), .A(n17115), .B(n16963), .ZN(
        n16965) );
  OAI211_X1 U20242 ( .C1(n17116), .C2(n17914), .A(n16966), .B(n16965), .ZN(
        n16967) );
  OR4_X1 U20243 ( .A1(n9832), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        P3_U2658) );
  AOI211_X1 U20244 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16985), .A(n16970), .B(
        n17126), .ZN(n16971) );
  AOI21_X1 U20245 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17081), .A(n16971), .ZN(
        n16979) );
  AOI22_X1 U20246 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16972), .B1(
        n17913), .B2(n17932), .ZN(n17928) );
  AOI21_X1 U20247 ( .B1(n17927), .B2(n17087), .A(n16764), .ZN(n16973) );
  XOR2_X1 U20248 ( .A(n17928), .B(n16973), .Z(n16974) );
  AOI22_X1 U20249 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17091), .B1(
        n17076), .B2(n16974), .ZN(n16978) );
  AOI22_X1 U20250 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16983), .B1(n16976), 
        .B2(n16975), .ZN(n16977) );
  NAND4_X1 U20251 ( .A1(n16979), .A2(n16978), .A3(n16977), .A4(n9975), .ZN(
        P3_U2659) );
  NAND2_X1 U20252 ( .A1(n17109), .A2(n17027), .ZN(n17028) );
  NAND4_X1 U20253 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .A4(n17048), .ZN(n17001) );
  OAI21_X1 U20254 ( .B1(n16980), .B2(n17001), .A(n18973), .ZN(n16984) );
  OAI22_X1 U20255 ( .A1(n16981), .A2(n17116), .B1(n17127), .B2(n16986), .ZN(
        n16982) );
  AOI21_X1 U20256 ( .B1(n16984), .B2(n16983), .A(n16982), .ZN(n16992) );
  OAI211_X1 U20257 ( .C1(n16995), .C2(n16986), .A(n17115), .B(n16985), .ZN(
        n16991) );
  INV_X1 U20258 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16994) );
  INV_X1 U20259 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17986) );
  INV_X1 U20260 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18002) );
  NOR2_X1 U20261 ( .A1(n17981), .A2(n18002), .ZN(n17984) );
  NAND2_X1 U20262 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17984), .ZN(
        n17030) );
  NOR2_X1 U20263 ( .A1(n17986), .A2(n17030), .ZN(n17020) );
  NAND2_X1 U20264 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17020), .ZN(
        n17006) );
  NOR2_X1 U20265 ( .A1(n16994), .A2(n17006), .ZN(n16993) );
  INV_X1 U20266 ( .A(n16993), .ZN(n16987) );
  OAI21_X1 U20267 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16987), .A(
        n17045), .ZN(n16989) );
  OAI21_X1 U20268 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16993), .A(
        n17913), .ZN(n17941) );
  AOI21_X1 U20269 ( .B1(n16989), .B2(n17941), .A(n18931), .ZN(n16988) );
  OAI21_X1 U20270 ( .B1(n16989), .B2(n17941), .A(n16988), .ZN(n16990) );
  NAND4_X1 U20271 ( .A1(n16992), .A2(n9975), .A3(n16991), .A4(n16990), .ZN(
        P3_U2660) );
  AOI22_X1 U20272 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17091), .B1(
        n17081), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n17005) );
  AOI21_X1 U20273 ( .B1(n16994), .B2(n17006), .A(n16993), .ZN(n17964) );
  INV_X1 U20274 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17957) );
  NAND3_X1 U20275 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17984), .A3(
        n17087), .ZN(n17007) );
  OAI21_X1 U20276 ( .B1(n17957), .B2(n17007), .A(n17045), .ZN(n17008) );
  XNOR2_X1 U20277 ( .A(n17964), .B(n17008), .ZN(n16998) );
  AOI211_X1 U20278 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16996), .A(n16995), .B(
        n17126), .ZN(n16997) );
  AOI211_X1 U20279 ( .C1(n17076), .C2(n16998), .A(n9832), .B(n16997), .ZN(
        n17004) );
  AOI21_X1 U20280 ( .B1(n16999), .B2(n17109), .A(n17114), .ZN(n17000) );
  INV_X1 U20281 ( .A(n17000), .ZN(n17024) );
  NOR2_X1 U20282 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17001), .ZN(n17016) );
  OAI21_X1 U20283 ( .B1(n17024), .B2(n17016), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n17003) );
  INV_X1 U20284 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18969) );
  OR3_X1 U20285 ( .A1(n18969), .A2(n17001), .A3(P3_REIP_REG_10__SCAN_IN), .ZN(
        n17002) );
  NAND4_X1 U20286 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17002), .ZN(
        P3_U2661) );
  OAI21_X1 U20287 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17020), .A(
        n17006), .ZN(n17970) );
  INV_X1 U20288 ( .A(n17970), .ZN(n17009) );
  OAI22_X1 U20289 ( .A1(n17009), .A2(n17008), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17007), .ZN(n17012) );
  INV_X1 U20290 ( .A(n17010), .ZN(n17014) );
  NAND2_X1 U20291 ( .A1(n17115), .A2(n17014), .ZN(n17019) );
  NAND2_X1 U20292 ( .A1(n17076), .A2(n9840), .ZN(n17103) );
  OAI22_X1 U20293 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17019), .B1(n17103), .B2(
        n17970), .ZN(n17011) );
  AOI211_X1 U20294 ( .C1(n17076), .C2(n17012), .A(n9832), .B(n17011), .ZN(
        n17018) );
  AOI221_X1 U20295 ( .B1(n17126), .B2(n17127), .C1(n17014), .C2(n17127), .A(
        n17013), .ZN(n17015) );
  AOI211_X1 U20296 ( .C1(n17024), .C2(P3_REIP_REG_9__SCAN_IN), .A(n17016), .B(
        n17015), .ZN(n17017) );
  OAI211_X1 U20297 ( .C1(n17957), .C2(n17116), .A(n17018), .B(n17017), .ZN(
        P3_U2662) );
  AOI21_X1 U20298 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17036), .A(n17019), .ZN(
        n17023) );
  AOI21_X1 U20299 ( .B1(n17984), .B2(n17087), .A(n9840), .ZN(n17031) );
  AOI21_X1 U20300 ( .B1(n17986), .B2(n17030), .A(n17020), .ZN(n17988) );
  XNOR2_X1 U20301 ( .A(n17031), .B(n17988), .ZN(n17021) );
  OAI21_X1 U20302 ( .B1(n18931), .B2(n17021), .A(n18388), .ZN(n17022) );
  AOI211_X1 U20303 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17081), .A(n17023), .B(
        n17022), .ZN(n17026) );
  INV_X1 U20304 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18965) );
  INV_X1 U20305 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18963) );
  NOR2_X1 U20306 ( .A1(n18965), .A2(n18963), .ZN(n17029) );
  OAI221_X1 U20307 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n17029), .C1(
        P3_REIP_REG_8__SCAN_IN), .C2(n17048), .A(n17024), .ZN(n17025) );
  OAI211_X1 U20308 ( .C1(n17116), .C2(n17986), .A(n17026), .B(n17025), .ZN(
        P3_U2663) );
  OAI21_X1 U20309 ( .B1(n17027), .B2(n17120), .A(n17130), .ZN(n17060) );
  AOI211_X1 U20310 ( .C1(n18965), .C2(n18963), .A(n17029), .B(n17028), .ZN(
        n17035) );
  INV_X1 U20311 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18019) );
  NAND2_X1 U20312 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18015), .ZN(
        n17053) );
  NOR2_X1 U20313 ( .A1(n18019), .A2(n17053), .ZN(n17042) );
  OAI21_X1 U20314 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17042), .A(
        n17030), .ZN(n18006) );
  INV_X1 U20315 ( .A(n18006), .ZN(n17032) );
  INV_X1 U20316 ( .A(n17087), .ZN(n17099) );
  OAI21_X1 U20317 ( .B1(n17981), .B2(n17099), .A(n17045), .ZN(n17043) );
  OAI221_X1 U20318 ( .B1(n17032), .B2(n17031), .C1(n18006), .C2(n17043), .A(
        n17076), .ZN(n17033) );
  OAI211_X1 U20319 ( .C1(n17127), .C2(n17037), .A(n18388), .B(n17033), .ZN(
        n17034) );
  AOI211_X1 U20320 ( .C1(n17060), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17035), .B(
        n17034), .ZN(n17039) );
  OAI211_X1 U20321 ( .C1(n17040), .C2(n17037), .A(n17115), .B(n17036), .ZN(
        n17038) );
  OAI211_X1 U20322 ( .C1(n17116), .C2(n18002), .A(n17039), .B(n17038), .ZN(
        P3_U2664) );
  AOI211_X1 U20323 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17061), .A(n17040), .B(
        n17126), .ZN(n17041) );
  AOI21_X1 U20324 ( .B1(n17091), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17041), .ZN(n17051) );
  AOI21_X1 U20325 ( .B1(n18019), .B2(n17053), .A(n17042), .ZN(n18022) );
  NOR3_X1 U20326 ( .A1(n18022), .A2(n18931), .A3(n17043), .ZN(n17047) );
  INV_X1 U20327 ( .A(n18022), .ZN(n17044) );
  AOI211_X1 U20328 ( .C1(n17045), .C2(n17053), .A(n17044), .B(n17119), .ZN(
        n17046) );
  AOI211_X1 U20329 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17081), .A(n17047), .B(
        n17046), .ZN(n17050) );
  AOI22_X1 U20330 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17060), .B1(n17048), 
        .B2(n18963), .ZN(n17049) );
  NAND4_X1 U20331 ( .A1(n17051), .A2(n17050), .A3(n17049), .A4(n9975), .ZN(
        P3_U2665) );
  OR2_X1 U20332 ( .A1(n17120), .A2(n17065), .ZN(n17083) );
  OAI21_X1 U20333 ( .B1(n18959), .B2(n17083), .A(n18962), .ZN(n17059) );
  NOR2_X1 U20334 ( .A1(n18077), .A2(n18024), .ZN(n17069) );
  AOI21_X1 U20335 ( .B1(n17069), .B2(n17052), .A(n9840), .ZN(n17070) );
  OAI21_X1 U20336 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17069), .A(
        n17053), .ZN(n18032) );
  OAI21_X1 U20337 ( .B1(n17070), .B2(n18032), .A(n18388), .ZN(n17054) );
  AOI21_X1 U20338 ( .B1(n17070), .B2(n18032), .A(n17054), .ZN(n17056) );
  OAI22_X1 U20339 ( .A1(n17057), .A2(n17056), .B1(n17055), .B2(n17116), .ZN(
        n17058) );
  AOI21_X1 U20340 ( .B1(n17060), .B2(n17059), .A(n17058), .ZN(n17063) );
  OAI211_X1 U20341 ( .C1(n17066), .C2(n17064), .A(n17115), .B(n17061), .ZN(
        n17062) );
  OAI211_X1 U20342 ( .C1(n17064), .C2(n17127), .A(n17063), .B(n17062), .ZN(
        P3_U2666) );
  AOI21_X1 U20343 ( .B1(n17109), .B2(n17065), .A(n17114), .ZN(n17084) );
  AOI211_X1 U20344 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17092), .A(n17066), .B(
        n17126), .ZN(n17080) );
  NAND2_X1 U20345 ( .A1(n17068), .A2(n17067), .ZN(n19099) );
  INV_X1 U20346 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17073) );
  NAND2_X1 U20347 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18045), .ZN(
        n17085) );
  AOI21_X1 U20348 ( .B1(n17073), .B2(n17085), .A(n17069), .ZN(n18046) );
  INV_X1 U20349 ( .A(n17070), .ZN(n17071) );
  NAND2_X1 U20350 ( .A1(n18045), .A2(n17073), .ZN(n18042) );
  OAI22_X1 U20351 ( .A1(n18046), .A2(n17071), .B1(n17099), .B2(n18042), .ZN(
        n17075) );
  INV_X1 U20352 ( .A(n18046), .ZN(n17072) );
  OAI22_X1 U20353 ( .A1(n17073), .A2(n17116), .B1(n17072), .B2(n17103), .ZN(
        n17074) );
  AOI211_X1 U20354 ( .C1(n17076), .C2(n17075), .A(n9832), .B(n17074), .ZN(
        n17077) );
  OAI221_X1 U20355 ( .B1(n19099), .B2(n9828), .C1(n19099), .C2(n17078), .A(
        n17077), .ZN(n17079) );
  AOI211_X1 U20356 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17081), .A(n17080), .B(
        n17079), .ZN(n17082) );
  OAI221_X1 U20357 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17083), .C1(n18959), 
        .C2(n17084), .A(n17082), .ZN(P3_U2667) );
  INV_X1 U20358 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U20359 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17108) );
  AOI221_X1 U20360 ( .B1(n17120), .B2(n18957), .C1(n17108), .C2(n18957), .A(
        n17084), .ZN(n17090) );
  NAND2_X1 U20361 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17096) );
  INV_X1 U20362 ( .A(n17085), .ZN(n17086) );
  AOI21_X1 U20363 ( .B1(n18054), .B2(n17096), .A(n17086), .ZN(n18056) );
  AOI21_X1 U20364 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17087), .A(
        n9840), .ZN(n17097) );
  XNOR2_X1 U20365 ( .A(n18056), .B(n17097), .ZN(n17088) );
  OAI22_X1 U20366 ( .A1(n18931), .A2(n17088), .B1(n19099), .B2(n19032), .ZN(
        n17089) );
  AOI211_X1 U20367 ( .C1(n17091), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n17090), .B(n17089), .ZN(n17094) );
  OAI211_X1 U20368 ( .C1(n17095), .C2(n17441), .A(n17115), .B(n17092), .ZN(
        n17093) );
  OAI211_X1 U20369 ( .C1(n17441), .C2(n17127), .A(n17094), .B(n17093), .ZN(
        P3_U2668) );
  NAND2_X1 U20370 ( .A1(n17458), .A2(n17452), .ZN(n17112) );
  AOI211_X1 U20371 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17112), .A(n17095), .B(
        n17126), .ZN(n17107) );
  OAI21_X1 U20372 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17096), .ZN(n18067) );
  INV_X1 U20373 ( .A(n18067), .ZN(n17100) );
  INV_X1 U20374 ( .A(n17097), .ZN(n17098) );
  AOI211_X1 U20375 ( .C1(n17100), .C2(n17099), .A(n18931), .B(n17098), .ZN(
        n17106) );
  INV_X1 U20376 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17102) );
  NAND2_X1 U20377 ( .A1(n18879), .A2(n13184), .ZN(n18873) );
  NAND2_X1 U20378 ( .A1(n17101), .A2(n18873), .ZN(n19043) );
  OAI22_X1 U20379 ( .A1(n17127), .A2(n17102), .B1(n19043), .B2(n19099), .ZN(
        n17105) );
  INV_X1 U20380 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18955) );
  OAI22_X1 U20381 ( .A1(n18955), .A2(n17130), .B1(n18067), .B2(n17103), .ZN(
        n17104) );
  NOR4_X1 U20382 ( .A1(n17107), .A2(n17106), .A3(n17105), .A4(n17104), .ZN(
        n17111) );
  OAI211_X1 U20383 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17109), .B(n17108), .ZN(n17110) );
  OAI211_X1 U20384 ( .C1(n17116), .C2(n18071), .A(n17111), .B(n17110), .ZN(
        P3_U2669) );
  INV_X1 U20385 ( .A(n17112), .ZN(n17113) );
  NOR2_X1 U20386 ( .A1(n17113), .A2(n17447), .ZN(n17450) );
  AOI22_X1 U20387 ( .A1(n17115), .A2(n17450), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n17114), .ZN(n17125) );
  OAI21_X1 U20388 ( .B1(n17117), .B2(n18931), .A(n17116), .ZN(n17123) );
  NAND2_X1 U20389 ( .A1(n18879), .A2(n17118), .ZN(n19048) );
  OAI22_X1 U20390 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17119), .B1(
        n19099), .B2(n19048), .ZN(n17122) );
  OAI22_X1 U20391 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17120), .B1(n17127), 
        .B2(n17452), .ZN(n17121) );
  AOI211_X1 U20392 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17123), .A(
        n17122), .B(n17121), .ZN(n17124) );
  NAND2_X1 U20393 ( .A1(n17125), .A2(n17124), .ZN(P3_U2670) );
  NAND2_X1 U20394 ( .A1(n17127), .A2(n17126), .ZN(n17129) );
  AOI22_X1 U20395 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17129), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17128), .ZN(n17132) );
  NAND3_X1 U20396 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19095), .A3(
        n17130), .ZN(n17131) );
  OAI211_X1 U20397 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n19099), .A(
        n17132), .B(n17131), .ZN(P3_U2671) );
  INV_X1 U20398 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17133) );
  NOR2_X1 U20399 ( .A1(n17133), .A2(n17258), .ZN(n17214) );
  INV_X1 U20400 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17178) );
  NAND4_X1 U20401 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17134)
         );
  NOR3_X1 U20402 ( .A1(n17178), .A2(n17135), .A3(n17134), .ZN(n17136) );
  NAND4_X1 U20403 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17171), .A3(n17214), 
        .A4(n17136), .ZN(n17139) );
  NOR2_X1 U20404 ( .A1(n17140), .A2(n17139), .ZN(n17166) );
  NAND2_X1 U20405 ( .A1(n17451), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17138) );
  NAND2_X1 U20406 ( .A1(n17166), .A2(n17577), .ZN(n17137) );
  OAI22_X1 U20407 ( .A1(n17166), .A2(n17138), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17137), .ZN(P3_U2672) );
  NAND2_X1 U20408 ( .A1(n17140), .A2(n17139), .ZN(n17141) );
  NAND2_X1 U20409 ( .A1(n17141), .A2(n17451), .ZN(n17165) );
  AOI22_X1 U20410 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17142) );
  OAI21_X1 U20411 ( .B1(n17396), .B2(n17143), .A(n17142), .ZN(n17153) );
  AOI22_X1 U20412 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17417), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17151) );
  OAI22_X1 U20413 ( .A1(n10408), .A2(n17144), .B1(n15787), .B2(n18667), .ZN(
        n17149) );
  AOI22_X1 U20414 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17359), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20415 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9830), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n13106), .ZN(n17146) );
  AOI22_X1 U20416 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9965), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n9829), .ZN(n17145) );
  NAND3_X1 U20417 ( .A1(n17147), .A2(n17146), .A3(n17145), .ZN(n17148) );
  AOI211_X1 U20418 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n17318), .A(
        n17149), .B(n17148), .ZN(n17150) );
  OAI211_X1 U20419 ( .C1(n9885), .C2(n18454), .A(n17151), .B(n17150), .ZN(
        n17152) );
  AOI211_X1 U20420 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n17153), .B(n17152), .ZN(n17164) );
  AOI22_X1 U20421 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17163) );
  INV_X1 U20422 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20423 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20424 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17154) );
  OAI211_X1 U20425 ( .C1(n9828), .C2(n17331), .A(n17155), .B(n17154), .ZN(
        n17161) );
  AOI22_X1 U20426 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20427 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20428 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U20429 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n17156) );
  NAND4_X1 U20430 ( .A1(n17159), .A2(n17158), .A3(n17157), .A4(n17156), .ZN(
        n17160) );
  AOI211_X1 U20431 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17161), .B(n17160), .ZN(n17162) );
  OAI211_X1 U20432 ( .C1(n13155), .C2(n18850), .A(n17163), .B(n17162), .ZN(
        n17168) );
  NAND2_X1 U20433 ( .A1(n17169), .A2(n17168), .ZN(n17167) );
  XNOR2_X1 U20434 ( .A(n17164), .B(n17167), .ZN(n17468) );
  OAI22_X1 U20435 ( .A1(n17166), .A2(n17165), .B1(n17468), .B2(n17451), .ZN(
        P3_U2673) );
  OAI21_X1 U20436 ( .B1(n17169), .B2(n17168), .A(n17167), .ZN(n17473) );
  NOR2_X1 U20437 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17182), .ZN(n17170) );
  AOI22_X1 U20438 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17172), .B1(n17171), 
        .B2(n17170), .ZN(n17173) );
  OAI21_X1 U20439 ( .B1(n17473), .B2(n17451), .A(n17173), .ZN(P3_U2674) );
  OAI21_X1 U20440 ( .B1(n17179), .B2(n17175), .A(n17174), .ZN(n17482) );
  NAND3_X1 U20441 ( .A1(n17182), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17451), 
        .ZN(n17176) );
  OAI221_X1 U20442 ( .B1(n17182), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17451), 
        .C2(n17482), .A(n17176), .ZN(P3_U2676) );
  OAI21_X1 U20443 ( .B1(n17178), .B2(n17456), .A(n17177), .ZN(n17181) );
  AOI21_X1 U20444 ( .B1(n17180), .B2(n17184), .A(n17179), .ZN(n17483) );
  AOI22_X1 U20445 ( .A1(n17182), .A2(n17181), .B1(n17483), .B2(n17456), .ZN(
        n17183) );
  INV_X1 U20446 ( .A(n17183), .ZN(P3_U2677) );
  AOI21_X1 U20447 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17451), .A(n17192), .ZN(
        n17186) );
  OAI21_X1 U20448 ( .B1(n17188), .B2(n17185), .A(n17184), .ZN(n17490) );
  OAI22_X1 U20449 ( .A1(n17187), .A2(n17186), .B1(n17490), .B2(n17451), .ZN(
        P3_U2678) );
  AOI21_X1 U20450 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17451), .A(n17198), .ZN(
        n17191) );
  AOI21_X1 U20451 ( .B1(n17189), .B2(n17194), .A(n17188), .ZN(n17491) );
  INV_X1 U20452 ( .A(n17491), .ZN(n17190) );
  OAI22_X1 U20453 ( .A1(n17192), .A2(n17191), .B1(n17190), .B2(n17451), .ZN(
        P3_U2679) );
  INV_X1 U20454 ( .A(n17193), .ZN(n17213) );
  AOI21_X1 U20455 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17451), .A(n17213), .ZN(
        n17197) );
  OAI21_X1 U20456 ( .B1(n17196), .B2(n17195), .A(n17194), .ZN(n17500) );
  OAI22_X1 U20457 ( .A1(n17198), .A2(n17197), .B1(n17500), .B2(n17451), .ZN(
        P3_U2680) );
  AOI21_X1 U20458 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17451), .A(n17199), .ZN(
        n17212) );
  AOI22_X1 U20459 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17210) );
  INV_X1 U20460 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20461 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20462 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17200) );
  OAI211_X1 U20463 ( .C1(n9828), .C2(n17202), .A(n17201), .B(n17200), .ZN(
        n17208) );
  AOI22_X1 U20464 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20465 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20466 ( .A1(n17359), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U20467 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n17203) );
  NAND4_X1 U20468 ( .A1(n17206), .A2(n17205), .A3(n17204), .A4(n17203), .ZN(
        n17207) );
  AOI211_X1 U20469 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17208), .B(n17207), .ZN(n17209) );
  OAI211_X1 U20470 ( .C1(n10419), .C2(n18446), .A(n17210), .B(n17209), .ZN(
        n17501) );
  INV_X1 U20471 ( .A(n17501), .ZN(n17211) );
  OAI22_X1 U20472 ( .A1(n17213), .A2(n17212), .B1(n17211), .B2(n17451), .ZN(
        P3_U2681) );
  NOR2_X1 U20473 ( .A1(n17456), .A2(n17214), .ZN(n17243) );
  AOI22_X1 U20474 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17215) );
  OAI21_X1 U20475 ( .B1(n17328), .B2(n17216), .A(n17215), .ZN(n17227) );
  AOI22_X1 U20476 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17225) );
  INV_X1 U20477 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20478 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17217) );
  OAI21_X1 U20479 ( .B1(n9828), .B2(n17218), .A(n17217), .ZN(n17223) );
  AOI22_X1 U20480 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20481 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17219) );
  OAI211_X1 U20482 ( .C1(n9846), .C2(n17221), .A(n17220), .B(n17219), .ZN(
        n17222) );
  AOI211_X1 U20483 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17223), .B(n17222), .ZN(n17224) );
  OAI211_X1 U20484 ( .C1(n10419), .C2(n18441), .A(n17225), .B(n17224), .ZN(
        n17226) );
  AOI211_X1 U20485 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n17227), .B(n17226), .ZN(n17508) );
  INV_X1 U20486 ( .A(n17508), .ZN(n17228) );
  AOI22_X1 U20487 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17243), .B1(n17456), 
        .B2(n17228), .ZN(n17229) );
  OAI21_X1 U20488 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17230), .A(n17229), .ZN(
        P3_U2682) );
  AOI22_X1 U20489 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20490 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17231) );
  OAI21_X1 U20491 ( .B1(n17415), .B2(n17343), .A(n17231), .ZN(n17240) );
  AOI22_X1 U20492 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17311), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20493 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17233) );
  AOI22_X1 U20494 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17232) );
  OAI211_X1 U20495 ( .C1(n9828), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        n17235) );
  AOI21_X1 U20496 ( .B1(n17318), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17235), .ZN(n17236) );
  OAI211_X1 U20497 ( .C1(n17238), .C2(n17346), .A(n17237), .B(n17236), .ZN(
        n17239) );
  AOI211_X1 U20498 ( .C1(n13275), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n17240), .B(n17239), .ZN(n17241) );
  OAI211_X1 U20499 ( .C1(n10419), .C2(n18435), .A(n17242), .B(n17241), .ZN(
        n17512) );
  INV_X1 U20500 ( .A(n17512), .ZN(n17246) );
  OAI21_X1 U20501 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17244), .A(n17243), .ZN(
        n17245) );
  OAI21_X1 U20502 ( .B1(n17246), .B2(n17451), .A(n17245), .ZN(P3_U2683) );
  AOI22_X1 U20503 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17247) );
  OAI21_X1 U20504 ( .B1(n17396), .B2(n17248), .A(n17247), .ZN(n17257) );
  AOI22_X1 U20505 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17255) );
  OAI22_X1 U20506 ( .A1(n9885), .A2(n18827), .B1(n10419), .B2(n18429), .ZN(
        n17253) );
  AOI22_X1 U20507 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17359), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20508 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20509 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17249) );
  NAND3_X1 U20510 ( .A1(n17251), .A2(n17250), .A3(n17249), .ZN(n17252) );
  AOI211_X1 U20511 ( .C1(n17318), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17253), .B(n17252), .ZN(n17254) );
  OAI211_X1 U20512 ( .C1(n15787), .C2(n18626), .A(n17255), .B(n17254), .ZN(
        n17256) );
  AOI211_X1 U20513 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17257), .B(n17256), .ZN(n17521) );
  OAI21_X1 U20514 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17260), .A(n17258), .ZN(
        n17259) );
  AOI22_X1 U20515 ( .A1(n17456), .A2(n17521), .B1(n17259), .B2(n17451), .ZN(
        P3_U2684) );
  OR2_X1 U20516 ( .A1(n17274), .A2(n17260), .ZN(n17276) );
  INV_X1 U20517 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U20518 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13106), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17261) );
  OAI21_X1 U20519 ( .B1(n17344), .B2(n17378), .A(n17261), .ZN(n17271) );
  AOI22_X1 U20520 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17269) );
  OAI22_X1 U20521 ( .A1(n10419), .A2(n18424), .B1(n9876), .B2(n17262), .ZN(
        n17267) );
  AOI22_X1 U20522 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U20523 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20524 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17263) );
  NAND3_X1 U20525 ( .A1(n17265), .A2(n17264), .A3(n17263), .ZN(n17266) );
  AOI211_X1 U20526 ( .C1(n17417), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17267), .B(n17266), .ZN(n17268) );
  OAI211_X1 U20527 ( .C1(n15787), .C2(n18623), .A(n17269), .B(n17268), .ZN(
        n17270) );
  AOI211_X1 U20528 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17271), .B(n17270), .ZN(n17525) );
  INV_X1 U20529 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17273) );
  NAND2_X1 U20530 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17325), .ZN(n17321) );
  NOR2_X1 U20531 ( .A1(n17272), .A2(n17321), .ZN(n17293) );
  NAND2_X1 U20532 ( .A1(n17577), .A2(n17293), .ZN(n17307) );
  NOR2_X1 U20533 ( .A1(n17273), .A2(n17307), .ZN(n17277) );
  NAND3_X1 U20534 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17277), .A3(n17274), 
        .ZN(n17275) );
  OAI221_X1 U20535 ( .B1(n17456), .B2(n17276), .C1(n17451), .C2(n17525), .A(
        n17275), .ZN(P3_U2685) );
  NOR2_X1 U20536 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17277), .ZN(n17292) );
  AOI211_X1 U20537 ( .C1(n17577), .C2(n17279), .A(n17278), .B(n17437), .ZN(
        n17291) );
  AOI22_X1 U20538 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17280) );
  OAI21_X1 U20539 ( .B1(n17328), .B2(n17406), .A(n17280), .ZN(n17290) );
  AOI22_X1 U20540 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17288) );
  OAI22_X1 U20541 ( .A1(n17377), .A2(n18649), .B1(n9876), .B2(n17397), .ZN(
        n17286) );
  AOI22_X1 U20542 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U20543 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20544 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17282) );
  NAND3_X1 U20545 ( .A1(n17284), .A2(n17283), .A3(n17282), .ZN(n17285) );
  AOI211_X1 U20546 ( .C1(n15772), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n17286), .B(n17285), .ZN(n17287) );
  OAI211_X1 U20547 ( .C1(n10419), .C2(n18419), .A(n17288), .B(n17287), .ZN(
        n17289) );
  AOI211_X1 U20548 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n17290), .B(n17289), .ZN(n17531) );
  OAI22_X1 U20549 ( .A1(n17292), .A2(n17291), .B1(n17531), .B2(n17451), .ZN(
        P3_U2686) );
  NOR2_X1 U20550 ( .A1(n17456), .A2(n17293), .ZN(n17322) );
  AOI22_X1 U20551 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20552 ( .B1(n17377), .B2(n18646), .A(n17294), .ZN(n17304) );
  INV_X1 U20553 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18618) );
  AOI22_X1 U20554 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20555 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17318), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U20556 ( .B1(n10419), .B2(n18415), .A(n17295), .ZN(n17300) );
  AOI22_X1 U20557 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20558 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17296) );
  OAI211_X1 U20559 ( .C1(n17298), .C2(n17413), .A(n17297), .B(n17296), .ZN(
        n17299) );
  AOI211_X1 U20560 ( .C1(n9965), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17300), .B(n17299), .ZN(n17301) );
  OAI211_X1 U20561 ( .C1(n15787), .C2(n18618), .A(n17302), .B(n17301), .ZN(
        n17303) );
  AOI211_X1 U20562 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17304), .B(n17303), .ZN(n17538) );
  INV_X1 U20563 ( .A(n17538), .ZN(n17305) );
  AOI22_X1 U20564 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17322), .B1(n17456), 
        .B2(n17305), .ZN(n17306) );
  OAI21_X1 U20565 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17307), .A(n17306), .ZN(
        P3_U2687) );
  AOI22_X1 U20566 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n13106), .ZN(n17320) );
  INV_X1 U20567 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20568 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17417), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20569 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17359), .B1(
        n17412), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17308) );
  OAI211_X1 U20570 ( .C1(n9828), .C2(n17310), .A(n17309), .B(n17308), .ZN(
        n17317) );
  AOI22_X1 U20571 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20572 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20573 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n9830), .ZN(n17313) );
  NAND2_X1 U20574 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n17312) );
  NAND4_X1 U20575 ( .A1(n17315), .A2(n17314), .A3(n17313), .A4(n17312), .ZN(
        n17316) );
  AOI211_X1 U20576 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n17318), .A(
        n17317), .B(n17316), .ZN(n17319) );
  OAI211_X1 U20577 ( .C1(n18862), .C2(n10419), .A(n17320), .B(n17319), .ZN(
        n17540) );
  INV_X1 U20578 ( .A(n17540), .ZN(n17324) );
  INV_X1 U20579 ( .A(n17321), .ZN(n17341) );
  OAI21_X1 U20580 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17341), .A(n17322), .ZN(
        n17323) );
  OAI21_X1 U20581 ( .B1(n17324), .B2(n17451), .A(n17323), .ZN(P3_U2688) );
  AOI22_X1 U20582 ( .A1(n17577), .A2(n17325), .B1(P3_EBX_REG_14__SCAN_IN), 
        .B2(n17451), .ZN(n17340) );
  AOI22_X1 U20583 ( .A1(n15772), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17359), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20584 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17326) );
  OAI21_X1 U20585 ( .B1(n17328), .B2(n17327), .A(n17326), .ZN(n17336) );
  AOI22_X1 U20586 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20587 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20588 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17329) );
  OAI211_X1 U20589 ( .C1(n9846), .C2(n17331), .A(n17330), .B(n17329), .ZN(
        n17332) );
  AOI21_X1 U20590 ( .B1(n9829), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17332), .ZN(n17333) );
  OAI211_X1 U20591 ( .C1(n10419), .C2(n18850), .A(n17334), .B(n17333), .ZN(
        n17335) );
  AOI211_X1 U20592 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17336), .B(n17335), .ZN(n17337) );
  OAI211_X1 U20593 ( .C1(n17396), .C2(n18446), .A(n17338), .B(n17337), .ZN(
        n17544) );
  INV_X1 U20594 ( .A(n17544), .ZN(n17339) );
  OAI22_X1 U20595 ( .A1(n17341), .A2(n17340), .B1(n17339), .B2(n17451), .ZN(
        P3_U2689) );
  NAND2_X1 U20596 ( .A1(n17577), .A2(n17375), .ZN(n17357) );
  AOI22_X1 U20597 ( .A1(n17363), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17342) );
  OAI21_X1 U20598 ( .B1(n17344), .B2(n17343), .A(n17342), .ZN(n17355) );
  AOI22_X1 U20599 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20600 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17345) );
  OAI21_X1 U20601 ( .B1(n9846), .B2(n17346), .A(n17345), .ZN(n17351) );
  AOI22_X1 U20602 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20603 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17347) );
  OAI211_X1 U20604 ( .C1(n9828), .C2(n17349), .A(n17348), .B(n17347), .ZN(
        n17350) );
  AOI211_X1 U20605 ( .C1(n9829), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17351), .B(n17350), .ZN(n17352) );
  OAI211_X1 U20606 ( .C1(n10419), .C2(n18834), .A(n17353), .B(n17352), .ZN(
        n17354) );
  AOI211_X1 U20607 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17355), .B(n17354), .ZN(n17553) );
  NAND3_X1 U20608 ( .A1(n17357), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17451), 
        .ZN(n17356) );
  OAI221_X1 U20609 ( .B1(n17357), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17451), 
        .C2(n17553), .A(n17356), .ZN(P3_U2691) );
  INV_X1 U20610 ( .A(n17389), .ZN(n17358) );
  OAI21_X1 U20611 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17358), .A(n17451), .ZN(
        n17374) );
  AOI22_X1 U20612 ( .A1(n13275), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17359), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20613 ( .B1(n17377), .B2(n18626), .A(n17361), .ZN(n17373) );
  INV_X1 U20614 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U20615 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17370) );
  OAI22_X1 U20616 ( .A1(n9846), .A2(n17362), .B1(n10419), .B2(n18827), .ZN(
        n17368) );
  AOI22_X1 U20617 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20618 ( .A1(n17398), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20619 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17364) );
  NAND3_X1 U20620 ( .A1(n17366), .A2(n17365), .A3(n17364), .ZN(n17367) );
  AOI211_X1 U20621 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17368), .B(n17367), .ZN(n17369) );
  OAI211_X1 U20622 ( .C1(n15787), .C2(n17371), .A(n17370), .B(n17369), .ZN(
        n17372) );
  AOI211_X1 U20623 ( .C1(n17376), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17373), .B(n17372), .ZN(n17557) );
  OAI22_X1 U20624 ( .A1(n17375), .A2(n17374), .B1(n17557), .B2(n17451), .ZN(
        P3_U2692) );
  AOI22_X1 U20625 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20626 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17412), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17387) );
  OAI22_X1 U20627 ( .A1(n17396), .A2(n18424), .B1(n10419), .B2(n18820), .ZN(
        n17385) );
  OAI22_X1 U20628 ( .A1(n15787), .A2(n17378), .B1(n17377), .B2(n18623), .ZN(
        n17379) );
  AOI21_X1 U20629 ( .B1(n9965), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(n17379), .ZN(n17383) );
  AOI22_X1 U20630 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20631 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20632 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9829), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17380) );
  NAND4_X1 U20633 ( .A1(n17383), .A2(n17382), .A3(n17381), .A4(n17380), .ZN(
        n17384) );
  AOI211_X1 U20634 ( .C1(n17394), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17385), .B(n17384), .ZN(n17386) );
  NAND3_X1 U20635 ( .A1(n17388), .A2(n17387), .A3(n17386), .ZN(n17561) );
  INV_X1 U20636 ( .A(n17561), .ZN(n17391) );
  OAI21_X1 U20637 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17410), .A(n17389), .ZN(
        n17390) );
  AOI22_X1 U20638 ( .A1(n17456), .A2(n17391), .B1(n17390), .B2(n17451), .ZN(
        P3_U2693) );
  NOR3_X1 U20639 ( .A1(n17437), .A2(n17436), .A3(n17392), .ZN(n17393) );
  OAI21_X1 U20640 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17393), .A(n17451), .ZN(
        n17409) );
  AOI22_X1 U20641 ( .A1(n13106), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20642 ( .B1(n17396), .B2(n18419), .A(n17395), .ZN(n17408) );
  AOI22_X1 U20643 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15772), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17405) );
  OAI22_X1 U20644 ( .A1(n13155), .A2(n17397), .B1(n10419), .B2(n18813), .ZN(
        n17403) );
  AOI22_X1 U20645 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20646 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17398), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20647 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17399) );
  NAND3_X1 U20648 ( .A1(n17401), .A2(n17400), .A3(n17399), .ZN(n17402) );
  AOI211_X1 U20649 ( .C1(n9835), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17403), .B(n17402), .ZN(n17404) );
  OAI211_X1 U20650 ( .C1(n17298), .C2(n17406), .A(n17405), .B(n17404), .ZN(
        n17407) );
  AOI211_X1 U20651 ( .C1(n17412), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17408), .B(n17407), .ZN(n17567) );
  OAI22_X1 U20652 ( .A1(n17410), .A2(n17409), .B1(n17567), .B2(n17451), .ZN(
        P3_U2694) );
  NOR2_X1 U20653 ( .A1(n17436), .A2(n17453), .ZN(n17443) );
  NAND2_X1 U20654 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17443), .ZN(n17438) );
  INV_X1 U20655 ( .A(n17438), .ZN(n17433) );
  AND2_X1 U20656 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17433), .ZN(n17435) );
  NAND2_X1 U20657 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17435), .ZN(n17431) );
  AOI22_X1 U20658 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20659 ( .A1(n17412), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17363), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20660 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9965), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17426) );
  OAI22_X1 U20661 ( .A1(n17415), .A2(n17414), .B1(n9876), .B2(n17413), .ZN(
        n17424) );
  AOI22_X1 U20662 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17416), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20663 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20664 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17420) );
  NAND2_X1 U20665 ( .A1(n17318), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17419) );
  NAND4_X1 U20666 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17423) );
  AOI211_X1 U20667 ( .C1(n15772), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17424), .B(n17423), .ZN(n17425) );
  NAND4_X1 U20668 ( .A1(n17428), .A2(n17427), .A3(n17426), .A4(n17425), .ZN(
        n17572) );
  INV_X1 U20669 ( .A(n17572), .ZN(n17430) );
  NAND3_X1 U20670 ( .A1(n17431), .A2(P3_EBX_REG_8__SCAN_IN), .A3(n17451), .ZN(
        n17429) );
  OAI221_X1 U20671 ( .B1(n17431), .B2(P3_EBX_REG_8__SCAN_IN), .C1(n17451), 
        .C2(n17430), .A(n17429), .ZN(P3_U2695) );
  OAI211_X1 U20672 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17435), .A(n17431), .B(
        n17451), .ZN(n17432) );
  OAI21_X1 U20673 ( .B1(n17451), .B2(n18454), .A(n17432), .ZN(P3_U2696) );
  AOI21_X1 U20674 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17451), .A(n17433), .ZN(
        n17434) );
  OAI22_X1 U20675 ( .A1(n17435), .A2(n17434), .B1(n18446), .B2(n17451), .ZN(
        P3_U2697) );
  NOR2_X1 U20676 ( .A1(n17437), .A2(n17436), .ZN(n17439) );
  OAI21_X1 U20677 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17439), .A(n17438), .ZN(
        n17440) );
  AOI22_X1 U20678 ( .A1(n17456), .A2(n18441), .B1(n17440), .B2(n17451), .ZN(
        P3_U2698) );
  INV_X1 U20679 ( .A(n17453), .ZN(n17455) );
  NAND3_X1 U20680 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17447), .A3(n17455), .ZN(
        n17444) );
  NOR2_X1 U20681 ( .A1(n17441), .A2(n17444), .ZN(n17446) );
  AOI21_X1 U20682 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17451), .A(n17446), .ZN(
        n17442) );
  OAI22_X1 U20683 ( .A1(n17443), .A2(n17442), .B1(n18435), .B2(n17451), .ZN(
        P3_U2699) );
  INV_X1 U20684 ( .A(n17444), .ZN(n17449) );
  AOI21_X1 U20685 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17451), .A(n17449), .ZN(
        n17445) );
  OAI22_X1 U20686 ( .A1(n17446), .A2(n17445), .B1(n18429), .B2(n17451), .ZN(
        P3_U2700) );
  AOI22_X1 U20687 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17451), .B1(n17447), .B2(
        n17455), .ZN(n17448) );
  OAI22_X1 U20688 ( .A1(n17449), .A2(n17448), .B1(n18424), .B2(n17451), .ZN(
        P3_U2701) );
  INV_X1 U20689 ( .A(n17450), .ZN(n17454) );
  OAI222_X1 U20690 ( .A1(n17454), .A2(n17453), .B1(n17452), .B2(n17459), .C1(
        n18419), .C2(n17451), .ZN(P3_U2702) );
  AOI22_X1 U20691 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17456), .B1(
        n17455), .B2(n17458), .ZN(n17457) );
  OAI21_X1 U20692 ( .B1(n17459), .B2(n17458), .A(n17457), .ZN(P3_U2703) );
  INV_X1 U20693 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17675) );
  INV_X1 U20694 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17671) );
  INV_X1 U20695 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17667) );
  INV_X1 U20696 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17713) );
  INV_X1 U20697 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17695) );
  INV_X1 U20698 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17681) );
  INV_X1 U20699 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17689) );
  INV_X1 U20700 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17687) );
  INV_X1 U20701 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17685) );
  INV_X1 U20702 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17683) );
  NOR4_X1 U20703 ( .A1(n17689), .A2(n17687), .A3(n17685), .A4(n17683), .ZN(
        n17461) );
  INV_X1 U20704 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17708) );
  INV_X1 U20705 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17706) );
  INV_X1 U20706 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17704) );
  INV_X1 U20707 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17701) );
  NOR4_X1 U20708 ( .A1(n17708), .A2(n17706), .A3(n17704), .A4(n17701), .ZN(
        n17462) );
  INV_X1 U20709 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17662) );
  INV_X1 U20710 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17660) );
  NAND2_X1 U20711 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17478), .ZN(n17475) );
  NAND3_X1 U20712 ( .A1(n17596), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17466), 
        .ZN(n17465) );
  NOR2_X2 U20713 ( .A1(n17463), .A2(n17596), .ZN(n17532) );
  NAND2_X1 U20714 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17532), .ZN(n17464) );
  OAI211_X1 U20715 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17466), .A(n17465), .B(
        n17464), .ZN(P3_U2704) );
  NOR2_X2 U20716 ( .A1(n18437), .A2(n17596), .ZN(n17533) );
  AOI22_X1 U20717 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17532), .ZN(n17467) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17532), .ZN(n17472) );
  AOI211_X1 U20719 ( .C1(n17675), .C2(n17475), .A(n17469), .B(n17516), .ZN(
        n17470) );
  INV_X1 U20720 ( .A(n17470), .ZN(n17471) );
  OAI211_X1 U20721 ( .C1(n17473), .C2(n17607), .A(n17472), .B(n17471), .ZN(
        P3_U2706) );
  INV_X1 U20722 ( .A(n17532), .ZN(n17507) );
  AOI22_X1 U20723 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17533), .B1(n17573), .B2(
        n17474), .ZN(n17477) );
  OAI211_X1 U20724 ( .C1(n17478), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17596), .B(
        n17475), .ZN(n17476) );
  OAI211_X1 U20725 ( .C1(n17507), .C2(n18431), .A(n17477), .B(n17476), .ZN(
        P3_U2707) );
  AOI22_X1 U20726 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17532), .ZN(n17481) );
  AOI211_X1 U20727 ( .C1(n17671), .C2(n17484), .A(n17478), .B(n17516), .ZN(
        n17479) );
  INV_X1 U20728 ( .A(n17479), .ZN(n17480) );
  OAI211_X1 U20729 ( .C1(n17482), .C2(n17607), .A(n17481), .B(n17480), .ZN(
        P3_U2708) );
  AOI22_X1 U20730 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17533), .B1(n17573), .B2(
        n17483), .ZN(n17486) );
  OAI211_X1 U20731 ( .C1(n9881), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17596), .B(
        n17484), .ZN(n17485) );
  OAI211_X1 U20732 ( .C1(n17507), .C2(n19530), .A(n17486), .B(n17485), .ZN(
        P3_U2709) );
  AOI22_X1 U20733 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17532), .ZN(n17489) );
  AOI211_X1 U20734 ( .C1(n17667), .C2(n17492), .A(n9881), .B(n17516), .ZN(
        n17487) );
  INV_X1 U20735 ( .A(n17487), .ZN(n17488) );
  OAI211_X1 U20736 ( .C1(n17490), .C2(n17607), .A(n17489), .B(n17488), .ZN(
        P3_U2710) );
  AOI22_X1 U20737 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17533), .B1(n17573), .B2(
        n17491), .ZN(n17495) );
  OAI211_X1 U20738 ( .C1(n17493), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17596), .B(
        n17492), .ZN(n17494) );
  OAI211_X1 U20739 ( .C1(n17507), .C2(n18409), .A(n17495), .B(n17494), .ZN(
        P3_U2711) );
  AOI22_X1 U20740 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17532), .ZN(n17499) );
  OAI211_X1 U20741 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17497), .A(n17596), .B(
        n17496), .ZN(n17498) );
  OAI211_X1 U20742 ( .C1(n17500), .C2(n17607), .A(n17499), .B(n17498), .ZN(
        P3_U2712) );
  INV_X1 U20743 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17656) );
  INV_X1 U20744 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17652) );
  NAND2_X1 U20745 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17526), .ZN(n17522) );
  NAND2_X1 U20746 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17517), .ZN(n17511) );
  NAND2_X1 U20747 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17662), .ZN(n17506) );
  AOI22_X1 U20748 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17532), .B1(n17573), .B2(
        n17501), .ZN(n17505) );
  NAND2_X1 U20749 ( .A1(n17596), .A2(n17511), .ZN(n17515) );
  OAI21_X1 U20750 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17502), .A(n17515), .ZN(
        n17503) );
  AOI22_X1 U20751 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17533), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17503), .ZN(n17504) );
  OAI211_X1 U20752 ( .C1(n17511), .C2(n17506), .A(n17505), .B(n17504), .ZN(
        P3_U2713) );
  OAI22_X1 U20753 ( .A1(n17508), .A2(n17607), .B1(n15192), .B2(n17507), .ZN(
        n17509) );
  AOI21_X1 U20754 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17533), .A(n17509), .ZN(
        n17510) );
  OAI221_X1 U20755 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17511), .C1(n17660), 
        .C2(n17515), .A(n17510), .ZN(P3_U2714) );
  INV_X1 U20756 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U20757 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17532), .B1(n17573), .B2(
        n17512), .ZN(n17514) );
  AOI22_X1 U20758 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17533), .B1(n17517), .B2(
        n17658), .ZN(n17513) );
  OAI211_X1 U20759 ( .C1(n17658), .C2(n17515), .A(n17514), .B(n17513), .ZN(
        P3_U2715) );
  AOI22_X1 U20760 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17532), .ZN(n17520) );
  AOI211_X1 U20761 ( .C1(n17656), .C2(n17522), .A(n17517), .B(n17516), .ZN(
        n17518) );
  INV_X1 U20762 ( .A(n17518), .ZN(n17519) );
  OAI211_X1 U20763 ( .C1(n17521), .C2(n17607), .A(n17520), .B(n17519), .ZN(
        P3_U2716) );
  AOI22_X1 U20764 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17532), .ZN(n17524) );
  OAI211_X1 U20765 ( .C1(n17526), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17596), .B(
        n17522), .ZN(n17523) );
  OAI211_X1 U20766 ( .C1(n17525), .C2(n17607), .A(n17524), .B(n17523), .ZN(
        P3_U2717) );
  AOI22_X1 U20767 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17532), .ZN(n17530) );
  INV_X1 U20768 ( .A(n17534), .ZN(n17528) );
  INV_X1 U20769 ( .A(n17526), .ZN(n17527) );
  OAI211_X1 U20770 ( .C1(n17528), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17596), .B(
        n17527), .ZN(n17529) );
  OAI211_X1 U20771 ( .C1(n17531), .C2(n17607), .A(n17530), .B(n17529), .ZN(
        P3_U2718) );
  AOI22_X1 U20772 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17533), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17532), .ZN(n17537) );
  OAI211_X1 U20773 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17535), .A(n17596), .B(
        n17534), .ZN(n17536) );
  OAI211_X1 U20774 ( .C1(n17538), .C2(n17607), .A(n17537), .B(n17536), .ZN(
        P3_U2719) );
  OR2_X1 U20775 ( .A1(n18449), .A2(n17539), .ZN(n17542) );
  NAND2_X1 U20776 ( .A1(n17596), .A2(n17539), .ZN(n17546) );
  AOI22_X1 U20777 ( .A1(n17573), .A2(n17540), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17605), .ZN(n17541) );
  OAI221_X1 U20778 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17542), .C1(n17713), 
        .C2(n17546), .A(n17541), .ZN(P3_U2720) );
  NAND2_X1 U20779 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17543) );
  NAND2_X1 U20780 ( .A1(n17577), .A2(n17576), .ZN(n17565) );
  NAND2_X1 U20781 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17564), .ZN(n17552) );
  NOR2_X1 U20782 ( .A1(n17704), .A2(n17552), .ZN(n17555) );
  NAND2_X1 U20783 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17555), .ZN(n17547) );
  AOI22_X1 U20784 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17605), .B1(n17573), .B2(
        n17544), .ZN(n17545) );
  OAI221_X1 U20785 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17547), .C1(n17708), 
        .C2(n17546), .A(n17545), .ZN(P3_U2721) );
  INV_X1 U20786 ( .A(n17547), .ZN(n17550) );
  AOI21_X1 U20787 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17596), .A(n17555), .ZN(
        n17549) );
  OAI222_X1 U20788 ( .A1(n17601), .A2(n17551), .B1(n17550), .B2(n17549), .C1(
        n17607), .C2(n17548), .ZN(P3_U2722) );
  INV_X1 U20789 ( .A(n17552), .ZN(n17559) );
  AOI21_X1 U20790 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17596), .A(n17559), .ZN(
        n17554) );
  OAI222_X1 U20791 ( .A1(n17601), .A2(n17556), .B1(n17555), .B2(n17554), .C1(
        n17607), .C2(n17553), .ZN(P3_U2723) );
  AOI21_X1 U20792 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17596), .A(n17564), .ZN(
        n17558) );
  OAI222_X1 U20793 ( .A1(n17601), .A2(n17560), .B1(n17559), .B2(n17558), .C1(
        n17607), .C2(n17557), .ZN(P3_U2724) );
  INV_X1 U20794 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17697) );
  NOR2_X1 U20795 ( .A1(n17697), .A2(n17565), .ZN(n17569) );
  OAI21_X1 U20796 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17569), .A(n17596), .ZN(
        n17563) );
  AOI22_X1 U20797 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17605), .B1(n17573), .B2(
        n17561), .ZN(n17562) );
  OAI21_X1 U20798 ( .B1(n17564), .B2(n17563), .A(n17562), .ZN(P3_U2725) );
  INV_X1 U20799 ( .A(n17565), .ZN(n17566) );
  AOI21_X1 U20800 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17596), .A(n17566), .ZN(
        n17568) );
  OAI222_X1 U20801 ( .A1(n17601), .A2(n17570), .B1(n17569), .B2(n17568), .C1(
        n17607), .C2(n17567), .ZN(P3_U2726) );
  INV_X1 U20802 ( .A(n17571), .ZN(n17580) );
  OAI21_X1 U20803 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17580), .A(n17596), .ZN(
        n17575) );
  AOI22_X1 U20804 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17605), .B1(n17573), .B2(
        n17572), .ZN(n17574) );
  OAI21_X1 U20805 ( .B1(n17576), .B2(n17575), .A(n17574), .ZN(P3_U2727) );
  INV_X1 U20806 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17691) );
  NAND2_X1 U20807 ( .A1(n17577), .A2(n17602), .ZN(n17594) );
  NAND2_X1 U20808 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17600), .ZN(n17587) );
  NOR2_X1 U20809 ( .A1(n17687), .A2(n17587), .ZN(n17590) );
  NAND2_X1 U20810 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17590), .ZN(n17581) );
  NOR2_X1 U20811 ( .A1(n17691), .A2(n17581), .ZN(n17582) );
  AOI21_X1 U20812 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17596), .A(n17582), .ZN(
        n17579) );
  OAI222_X1 U20813 ( .A1(n17601), .A2(n18447), .B1(n17580), .B2(n17579), .C1(
        n17607), .C2(n17578), .ZN(P3_U2728) );
  INV_X1 U20814 ( .A(n17581), .ZN(n17586) );
  AOI21_X1 U20815 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17596), .A(n17586), .ZN(
        n17583) );
  INV_X1 U20816 ( .A(n18008), .ZN(n18009) );
  OAI222_X1 U20817 ( .A1(n17601), .A2(n18442), .B1(n17583), .B2(n17582), .C1(
        n17607), .C2(n18009), .ZN(P3_U2729) );
  AOI21_X1 U20818 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17596), .A(n17590), .ZN(
        n17585) );
  OAI222_X1 U20819 ( .A1(n18436), .A2(n17601), .B1(n17586), .B2(n17585), .C1(
        n17607), .C2(n17584), .ZN(P3_U2730) );
  INV_X1 U20820 ( .A(n17587), .ZN(n17593) );
  AOI21_X1 U20821 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17596), .A(n17593), .ZN(
        n17589) );
  OAI222_X1 U20822 ( .A1(n18430), .A2(n17601), .B1(n17590), .B2(n17589), .C1(
        n17607), .C2(n17588), .ZN(P3_U2731) );
  AOI21_X1 U20823 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17596), .A(n17600), .ZN(
        n17592) );
  OAI222_X1 U20824 ( .A1(n18425), .A2(n17601), .B1(n17593), .B2(n17592), .C1(
        n17607), .C2(n17591), .ZN(P3_U2732) );
  INV_X1 U20825 ( .A(n17594), .ZN(n17595) );
  AOI21_X1 U20826 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17596), .A(n17595), .ZN(
        n17599) );
  INV_X1 U20827 ( .A(n17597), .ZN(n17598) );
  OAI222_X1 U20828 ( .A1(n18420), .A2(n17601), .B1(n17600), .B2(n17599), .C1(
        n17607), .C2(n17598), .ZN(P3_U2733) );
  AOI21_X1 U20829 ( .B1(n17681), .B2(n17603), .A(n17602), .ZN(n17604) );
  AOI22_X1 U20830 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17605), .B1(n17604), .B2(
        n17596), .ZN(n17606) );
  OAI21_X1 U20831 ( .B1(n17608), .B2(n17607), .A(n17606), .ZN(P3_U2734) );
  NOR2_X4 U20832 ( .A1(n19079), .A2(n17611), .ZN(n17644) );
  AND2_X1 U20833 ( .A1(n17644), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20834 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U20835 ( .A1(n19079), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17644), .ZN(n17612) );
  OAI21_X1 U20836 ( .B1(n17677), .B2(n17627), .A(n17612), .ZN(P3_U2737) );
  AOI22_X1 U20837 ( .A1(n19079), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17613) );
  OAI21_X1 U20838 ( .B1(n17675), .B2(n17627), .A(n17613), .ZN(P3_U2738) );
  INV_X1 U20839 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U20840 ( .A1(n19079), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17614) );
  OAI21_X1 U20841 ( .B1(n17673), .B2(n17627), .A(n17614), .ZN(P3_U2739) );
  AOI22_X1 U20842 ( .A1(n19079), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U20843 ( .B1(n17671), .B2(n17627), .A(n17615), .ZN(P3_U2740) );
  AOI22_X1 U20844 ( .A1(n19079), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17616) );
  OAI21_X1 U20845 ( .B1(n10198), .B2(n17627), .A(n17616), .ZN(P3_U2741) );
  AOI22_X1 U20846 ( .A1(n19079), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17617) );
  OAI21_X1 U20847 ( .B1(n17667), .B2(n17627), .A(n17617), .ZN(P3_U2742) );
  AOI22_X1 U20848 ( .A1(n19079), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17618) );
  OAI21_X1 U20849 ( .B1(n10197), .B2(n17627), .A(n17618), .ZN(P3_U2743) );
  INV_X1 U20850 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U20851 ( .A1(n19079), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20852 ( .B1(n17664), .B2(n17627), .A(n17619), .ZN(P3_U2744) );
  AOI22_X1 U20853 ( .A1(n19079), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17620) );
  OAI21_X1 U20854 ( .B1(n17662), .B2(n17627), .A(n17620), .ZN(P3_U2745) );
  AOI22_X1 U20855 ( .A1(n17637), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17621) );
  OAI21_X1 U20856 ( .B1(n17660), .B2(n17627), .A(n17621), .ZN(P3_U2746) );
  AOI22_X1 U20857 ( .A1(n17637), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17622) );
  OAI21_X1 U20858 ( .B1(n17658), .B2(n17627), .A(n17622), .ZN(P3_U2747) );
  AOI22_X1 U20859 ( .A1(n17637), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17623) );
  OAI21_X1 U20860 ( .B1(n17656), .B2(n17627), .A(n17623), .ZN(P3_U2748) );
  INV_X1 U20861 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U20862 ( .A1(n17637), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17624) );
  OAI21_X1 U20863 ( .B1(n17654), .B2(n17627), .A(n17624), .ZN(P3_U2749) );
  AOI22_X1 U20864 ( .A1(n17637), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17625) );
  OAI21_X1 U20865 ( .B1(n17652), .B2(n17627), .A(n17625), .ZN(P3_U2750) );
  INV_X1 U20866 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U20867 ( .A1(n17637), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U20868 ( .B1(n17650), .B2(n17627), .A(n17626), .ZN(P3_U2751) );
  AOI22_X1 U20869 ( .A1(n17637), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17628) );
  OAI21_X1 U20870 ( .B1(n17713), .B2(n17646), .A(n17628), .ZN(P3_U2752) );
  AOI22_X1 U20871 ( .A1(n17637), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17629) );
  OAI21_X1 U20872 ( .B1(n17708), .B2(n17646), .A(n17629), .ZN(P3_U2753) );
  AOI22_X1 U20873 ( .A1(n17637), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17630) );
  OAI21_X1 U20874 ( .B1(n17706), .B2(n17646), .A(n17630), .ZN(P3_U2754) );
  AOI22_X1 U20875 ( .A1(n17637), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17631) );
  OAI21_X1 U20876 ( .B1(n17704), .B2(n17646), .A(n17631), .ZN(P3_U2755) );
  AOI22_X1 U20877 ( .A1(n19079), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17632) );
  OAI21_X1 U20878 ( .B1(n17701), .B2(n17646), .A(n17632), .ZN(P3_U2756) );
  INV_X1 U20879 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U20880 ( .A1(n19079), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17633) );
  OAI21_X1 U20881 ( .B1(n17699), .B2(n17646), .A(n17633), .ZN(P3_U2757) );
  AOI22_X1 U20882 ( .A1(n19079), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17634) );
  OAI21_X1 U20883 ( .B1(n17697), .B2(n17646), .A(n17634), .ZN(P3_U2758) );
  AOI22_X1 U20884 ( .A1(n19079), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17635) );
  OAI21_X1 U20885 ( .B1(n17695), .B2(n17646), .A(n17635), .ZN(P3_U2759) );
  INV_X1 U20886 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U20887 ( .A1(n19079), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17636) );
  OAI21_X1 U20888 ( .B1(n17693), .B2(n17646), .A(n17636), .ZN(P3_U2760) );
  AOI22_X1 U20889 ( .A1(n17637), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17638) );
  OAI21_X1 U20890 ( .B1(n17691), .B2(n17646), .A(n17638), .ZN(P3_U2761) );
  AOI22_X1 U20891 ( .A1(n19079), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17639) );
  OAI21_X1 U20892 ( .B1(n17689), .B2(n17646), .A(n17639), .ZN(P3_U2762) );
  AOI22_X1 U20893 ( .A1(n19079), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17640) );
  OAI21_X1 U20894 ( .B1(n17687), .B2(n17646), .A(n17640), .ZN(P3_U2763) );
  AOI22_X1 U20895 ( .A1(n19079), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17641) );
  OAI21_X1 U20896 ( .B1(n17685), .B2(n17646), .A(n17641), .ZN(P3_U2764) );
  AOI22_X1 U20897 ( .A1(n19079), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17642) );
  OAI21_X1 U20898 ( .B1(n17683), .B2(n17646), .A(n17642), .ZN(P3_U2765) );
  AOI22_X1 U20899 ( .A1(n19079), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17643) );
  OAI21_X1 U20900 ( .B1(n17681), .B2(n17646), .A(n17643), .ZN(P3_U2766) );
  AOI22_X1 U20901 ( .A1(n19079), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17644), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17645) );
  OAI21_X1 U20902 ( .B1(n17679), .B2(n17646), .A(n17645), .ZN(P3_U2767) );
  INV_X1 U20903 ( .A(n17647), .ZN(n18915) );
  AOI22_X1 U20904 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17710), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17709), .ZN(n17649) );
  OAI21_X1 U20905 ( .B1(n17650), .B2(n17712), .A(n17649), .ZN(P3_U2768) );
  AOI22_X1 U20906 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17709), .ZN(n17651) );
  OAI21_X1 U20907 ( .B1(n17652), .B2(n17712), .A(n17651), .ZN(P3_U2769) );
  AOI22_X1 U20908 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17709), .ZN(n17653) );
  OAI21_X1 U20909 ( .B1(n17654), .B2(n17712), .A(n17653), .ZN(P3_U2770) );
  AOI22_X1 U20910 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17709), .ZN(n17655) );
  OAI21_X1 U20911 ( .B1(n17656), .B2(n17712), .A(n17655), .ZN(P3_U2771) );
  AOI22_X1 U20912 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17709), .ZN(n17657) );
  OAI21_X1 U20913 ( .B1(n17658), .B2(n17712), .A(n17657), .ZN(P3_U2772) );
  AOI22_X1 U20914 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17709), .ZN(n17659) );
  OAI21_X1 U20915 ( .B1(n17660), .B2(n17712), .A(n17659), .ZN(P3_U2773) );
  AOI22_X1 U20916 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17709), .ZN(n17661) );
  OAI21_X1 U20917 ( .B1(n17662), .B2(n17712), .A(n17661), .ZN(P3_U2774) );
  AOI22_X1 U20918 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17709), .ZN(n17663) );
  OAI21_X1 U20919 ( .B1(n17664), .B2(n17712), .A(n17663), .ZN(P3_U2775) );
  AOI22_X1 U20920 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17709), .ZN(n17665) );
  OAI21_X1 U20921 ( .B1(n10197), .B2(n17712), .A(n17665), .ZN(P3_U2776) );
  AOI22_X1 U20922 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17709), .ZN(n17666) );
  OAI21_X1 U20923 ( .B1(n17667), .B2(n17712), .A(n17666), .ZN(P3_U2777) );
  AOI22_X1 U20924 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17709), .ZN(n17668) );
  OAI21_X1 U20925 ( .B1(n10198), .B2(n17712), .A(n17668), .ZN(P3_U2778) );
  AOI22_X1 U20926 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17669), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17709), .ZN(n17670) );
  OAI21_X1 U20927 ( .B1(n17671), .B2(n17712), .A(n17670), .ZN(P3_U2779) );
  AOI22_X1 U20928 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17710), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17709), .ZN(n17672) );
  OAI21_X1 U20929 ( .B1(n17673), .B2(n17712), .A(n17672), .ZN(P3_U2780) );
  AOI22_X1 U20930 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17710), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17709), .ZN(n17674) );
  OAI21_X1 U20931 ( .B1(n17675), .B2(n17712), .A(n17674), .ZN(P3_U2781) );
  AOI22_X1 U20932 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17710), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17709), .ZN(n17676) );
  OAI21_X1 U20933 ( .B1(n17677), .B2(n17712), .A(n17676), .ZN(P3_U2782) );
  AOI22_X1 U20934 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17709), .ZN(n17678) );
  OAI21_X1 U20935 ( .B1(n17679), .B2(n17712), .A(n17678), .ZN(P3_U2783) );
  AOI22_X1 U20936 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17709), .ZN(n17680) );
  OAI21_X1 U20937 ( .B1(n17681), .B2(n17712), .A(n17680), .ZN(P3_U2784) );
  AOI22_X1 U20938 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17709), .ZN(n17682) );
  OAI21_X1 U20939 ( .B1(n17683), .B2(n17712), .A(n17682), .ZN(P3_U2785) );
  AOI22_X1 U20940 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17702), .ZN(n17684) );
  OAI21_X1 U20941 ( .B1(n17685), .B2(n17712), .A(n17684), .ZN(P3_U2786) );
  AOI22_X1 U20942 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17702), .ZN(n17686) );
  OAI21_X1 U20943 ( .B1(n17687), .B2(n17712), .A(n17686), .ZN(P3_U2787) );
  AOI22_X1 U20944 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17702), .ZN(n17688) );
  OAI21_X1 U20945 ( .B1(n17689), .B2(n17712), .A(n17688), .ZN(P3_U2788) );
  AOI22_X1 U20946 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17702), .ZN(n17690) );
  OAI21_X1 U20947 ( .B1(n17691), .B2(n17712), .A(n17690), .ZN(P3_U2789) );
  AOI22_X1 U20948 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17702), .ZN(n17692) );
  OAI21_X1 U20949 ( .B1(n17693), .B2(n17712), .A(n17692), .ZN(P3_U2790) );
  AOI22_X1 U20950 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17702), .ZN(n17694) );
  OAI21_X1 U20951 ( .B1(n17695), .B2(n17712), .A(n17694), .ZN(P3_U2791) );
  AOI22_X1 U20952 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17702), .ZN(n17696) );
  OAI21_X1 U20953 ( .B1(n17697), .B2(n17712), .A(n17696), .ZN(P3_U2792) );
  AOI22_X1 U20954 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17702), .ZN(n17698) );
  OAI21_X1 U20955 ( .B1(n17699), .B2(n17712), .A(n17698), .ZN(P3_U2793) );
  AOI22_X1 U20956 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17702), .ZN(n17700) );
  OAI21_X1 U20957 ( .B1(n17701), .B2(n17712), .A(n17700), .ZN(P3_U2794) );
  AOI22_X1 U20958 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17702), .ZN(n17703) );
  OAI21_X1 U20959 ( .B1(n17704), .B2(n17712), .A(n17703), .ZN(P3_U2795) );
  AOI22_X1 U20960 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17709), .ZN(n17705) );
  OAI21_X1 U20961 ( .B1(n17706), .B2(n17712), .A(n17705), .ZN(P3_U2796) );
  AOI22_X1 U20962 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17709), .ZN(n17707) );
  OAI21_X1 U20963 ( .B1(n17708), .B2(n17712), .A(n17707), .ZN(P3_U2797) );
  AOI22_X1 U20964 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17710), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17709), .ZN(n17711) );
  OAI21_X1 U20965 ( .B1(n17713), .B2(n17712), .A(n17711), .ZN(P3_U2798) );
  OAI21_X1 U20966 ( .B1(n17714), .B2(n18936), .A(n18083), .ZN(n17715) );
  AOI21_X1 U20967 ( .B1(n17982), .B2(n17726), .A(n17715), .ZN(n17751) );
  OAI21_X1 U20968 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17823), .A(
        n17751), .ZN(n17737) );
  AOI22_X1 U20969 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17737), .B1(
        n17929), .B2(n17716), .ZN(n17730) );
  NOR2_X1 U20970 ( .A1(n17911), .A2(n17999), .ZN(n17829) );
  INV_X1 U20971 ( .A(n17717), .ZN(n18093) );
  INV_X1 U20972 ( .A(n18095), .ZN(n17718) );
  OAI22_X1 U20973 ( .A1(n18093), .A2(n17992), .B1(n17718), .B2(n18088), .ZN(
        n17753) );
  NOR2_X1 U20974 ( .A1(n18097), .A2(n17753), .ZN(n17720) );
  NOR3_X1 U20975 ( .A1(n17829), .A2(n17720), .A3(n17719), .ZN(n17724) );
  NAND2_X1 U20976 ( .A1(n9832), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17729) );
  NOR2_X1 U20977 ( .A1(n17875), .A2(n17726), .ZN(n17739) );
  OAI211_X1 U20978 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17739), .B(n17727), .ZN(n17728) );
  INV_X1 U20979 ( .A(n17731), .ZN(n17733) );
  NAND2_X1 U20980 ( .A1(n17733), .A2(n17732), .ZN(n17734) );
  XNOR2_X1 U20981 ( .A(n15863), .B(n17734), .ZN(n18101) );
  OAI22_X1 U20982 ( .A1(n18388), .A2(n19005), .B1(n17884), .B2(n17735), .ZN(
        n17736) );
  AOI221_X1 U20983 ( .B1(n17739), .B2(n17738), .C1(n17737), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17736), .ZN(n17743) );
  INV_X1 U20984 ( .A(n17794), .ZN(n17746) );
  NOR2_X1 U20985 ( .A1(n17740), .A2(n17746), .ZN(n17741) );
  AOI22_X1 U20986 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17753), .B1(
        n17741), .B2(n18097), .ZN(n17742) );
  OAI211_X1 U20987 ( .C1(n18101), .C2(n17978), .A(n17743), .B(n17742), .ZN(
        P3_U2803) );
  AOI21_X1 U20988 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17745), .A(
        n17744), .ZN(n18110) );
  NOR2_X1 U20989 ( .A1(n18104), .A2(n17746), .ZN(n17754) );
  AOI21_X1 U20990 ( .B1(n18741), .B2(n17747), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17750) );
  OAI21_X1 U20991 ( .B1(n17929), .B2(n17858), .A(n17748), .ZN(n17749) );
  NAND2_X1 U20992 ( .A1(n9832), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18108) );
  OAI211_X1 U20993 ( .C1(n17751), .C2(n17750), .A(n17749), .B(n18108), .ZN(
        n17752) );
  AOI221_X1 U20994 ( .B1(n17754), .B2(n18105), .C1(n17753), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17752), .ZN(n17755) );
  OAI21_X1 U20995 ( .B1(n18110), .B2(n17978), .A(n17755), .ZN(P3_U2804) );
  OAI21_X1 U20996 ( .B1(n17951), .B2(n17757), .A(n17756), .ZN(n17758) );
  XNOR2_X1 U20997 ( .A(n17758), .B(n18119), .ZN(n18124) );
  NAND2_X1 U20998 ( .A1(n18741), .A2(n17760), .ZN(n17791) );
  OAI211_X1 U20999 ( .C1(n17759), .C2(n18936), .A(n18083), .B(n17791), .ZN(
        n17786) );
  NOR2_X1 U21000 ( .A1(n17875), .A2(n17760), .ZN(n17776) );
  OAI211_X1 U21001 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17776), .B(n17761), .ZN(n17762) );
  NAND2_X1 U21002 ( .A1(n9832), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18122) );
  OAI211_X1 U21003 ( .C1(n17884), .C2(n17763), .A(n17762), .B(n18122), .ZN(
        n17764) );
  AOI21_X1 U21004 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17786), .A(
        n17764), .ZN(n17769) );
  AOI21_X1 U21005 ( .B1(n18119), .B2(n17766), .A(n17765), .ZN(n18115) );
  XNOR2_X1 U21006 ( .A(n17767), .B(n18119), .ZN(n18116) );
  AOI22_X1 U21007 ( .A1(n17911), .A2(n18115), .B1(n17999), .B2(n18116), .ZN(
        n17768) );
  OAI211_X1 U21008 ( .C1(n17978), .C2(n18124), .A(n17769), .B(n17768), .ZN(
        P3_U2805) );
  AOI21_X1 U21009 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17771), .A(
        n17770), .ZN(n18139) );
  INV_X1 U21010 ( .A(n17772), .ZN(n17773) );
  OAI22_X1 U21011 ( .A1(n18388), .A2(n18999), .B1(n17884), .B2(n17773), .ZN(
        n17774) );
  AOI221_X1 U21012 ( .B1(n17776), .B2(n17775), .C1(n17786), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17774), .ZN(n17779) );
  INV_X1 U21013 ( .A(n18129), .ZN(n17777) );
  OAI22_X1 U21014 ( .A1(n18131), .A2(n17992), .B1(n17777), .B2(n18088), .ZN(
        n17793) );
  NOR2_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18133), .ZN(
        n18125) );
  AOI22_X1 U21016 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17793), .B1(
        n17794), .B2(n18125), .ZN(n17778) );
  OAI211_X1 U21017 ( .C1(n18139), .C2(n17978), .A(n17779), .B(n17778), .ZN(
        P3_U2806) );
  INV_X1 U21018 ( .A(n17780), .ZN(n17797) );
  AOI22_X1 U21019 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17951), .B1(
        n17781), .B2(n17798), .ZN(n17782) );
  NAND2_X1 U21020 ( .A1(n17780), .A2(n17782), .ZN(n17783) );
  XNOR2_X1 U21021 ( .A(n17783), .B(n18133), .ZN(n18146) );
  AOI21_X1 U21022 ( .B1(n17858), .B2(n17784), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17785) );
  INV_X1 U21023 ( .A(n17785), .ZN(n17787) );
  AOI22_X1 U21024 ( .A1(n17929), .A2(n17788), .B1(n17787), .B2(n17786), .ZN(
        n17789) );
  NAND2_X1 U21025 ( .A1(n9832), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18145) );
  OAI211_X1 U21026 ( .C1(n17791), .C2(n17790), .A(n17789), .B(n18145), .ZN(
        n17792) );
  AOI221_X1 U21027 ( .B1(n17794), .B2(n18133), .C1(n17793), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17792), .ZN(n17795) );
  OAI21_X1 U21028 ( .B1(n17978), .B2(n18146), .A(n17795), .ZN(P3_U2807) );
  INV_X1 U21029 ( .A(n18149), .ZN(n18166) );
  NOR2_X1 U21030 ( .A1(n18166), .A2(n17796), .ZN(n17801) );
  INV_X1 U21031 ( .A(n17801), .ZN(n18158) );
  AOI221_X1 U21032 ( .B1(n17799), .B2(n17798), .C1(n18158), .C2(n17798), .A(
        n17797), .ZN(n17800) );
  XNOR2_X1 U21033 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17800), .ZN(
        n18164) );
  NOR2_X1 U21034 ( .A1(n17882), .A2(n18158), .ZN(n17808) );
  NOR2_X1 U21035 ( .A1(n18157), .A2(n18088), .ZN(n17890) );
  AOI21_X1 U21036 ( .B1(n17911), .B2(n18218), .A(n17890), .ZN(n17881) );
  OAI21_X1 U21037 ( .B1(n17829), .B2(n17801), .A(n17881), .ZN(n17819) );
  NOR2_X1 U21038 ( .A1(n17802), .A2(n18936), .ZN(n17803) );
  OAI21_X1 U21039 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17823), .A(
        n17826), .ZN(n17813) );
  NOR2_X1 U21040 ( .A1(n17875), .A2(n17805), .ZN(n17815) );
  OAI211_X1 U21041 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17815), .B(n17806), .ZN(n17807) );
  NAND2_X1 U21042 ( .A1(n18156), .A2(n17809), .ZN(n18172) );
  INV_X1 U21043 ( .A(n17882), .ZN(n17865) );
  NAND2_X1 U21044 ( .A1(n18149), .A2(n17865), .ZN(n17846) );
  INV_X1 U21045 ( .A(n17810), .ZN(n17811) );
  OAI22_X1 U21046 ( .A1(n18388), .A2(n18993), .B1(n17884), .B2(n17811), .ZN(
        n17812) );
  AOI221_X1 U21047 ( .B1(n17815), .B2(n17814), .C1(n17813), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17812), .ZN(n17821) );
  NOR3_X1 U21048 ( .A1(n17951), .A2(n18147), .A3(n17816), .ZN(n17840) );
  INV_X1 U21049 ( .A(n17854), .ZN(n17841) );
  AOI22_X1 U21050 ( .A1(n18156), .A2(n17840), .B1(n17841), .B2(n17817), .ZN(
        n17818) );
  XNOR2_X1 U21051 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17818), .ZN(
        n18167) );
  AOI22_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17819), .B1(
        n17989), .B2(n18167), .ZN(n17820) );
  OAI211_X1 U21053 ( .C1(n18172), .C2(n17846), .A(n17821), .B(n17820), .ZN(
        P3_U2809) );
  NAND2_X1 U21054 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17822), .ZN(
        n18181) );
  AOI21_X1 U21055 ( .B1(n17824), .B2(n18741), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17825) );
  OAI22_X1 U21056 ( .A1(n17826), .A2(n17825), .B1(n18388), .B2(n18992), .ZN(
        n17827) );
  AOI221_X1 U21057 ( .B1(n17929), .B2(n17828), .C1(n17858), .C2(n17828), .A(
        n17827), .ZN(n17833) );
  NOR2_X1 U21058 ( .A1(n18166), .A2(n17830), .ZN(n18150) );
  OAI21_X1 U21059 ( .B1(n17829), .B2(n18150), .A(n17881), .ZN(n17843) );
  OAI221_X1 U21060 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17853), 
        .C1(n17830), .C2(n17840), .A(n17780), .ZN(n17831) );
  XNOR2_X1 U21061 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17831), .ZN(
        n18173) );
  AOI22_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17843), .B1(
        n17989), .B2(n18173), .ZN(n17832) );
  OAI211_X1 U21063 ( .C1(n17846), .C2(n18181), .A(n17833), .B(n17832), .ZN(
        P3_U2810) );
  AOI21_X1 U21064 ( .B1(n17982), .B2(n17835), .A(n18055), .ZN(n17861) );
  OAI21_X1 U21065 ( .B1(n17834), .B2(n18936), .A(n17861), .ZN(n17849) );
  NAND2_X1 U21066 ( .A1(n9832), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18184) );
  NOR2_X1 U21067 ( .A1(n17875), .A2(n17835), .ZN(n17851) );
  OAI211_X1 U21068 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17851), .B(n17836), .ZN(n17837) );
  OAI211_X1 U21069 ( .C1(n17884), .C2(n17838), .A(n18184), .B(n17837), .ZN(
        n17839) );
  AOI21_X1 U21070 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17849), .A(
        n17839), .ZN(n17845) );
  AOI21_X1 U21071 ( .B1(n17853), .B2(n17841), .A(n17840), .ZN(n17842) );
  XNOR2_X1 U21072 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17842), .ZN(
        n18182) );
  AOI22_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17843), .B1(
        n17989), .B2(n18182), .ZN(n17844) );
  OAI211_X1 U21074 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17846), .A(
        n17845), .B(n17844), .ZN(P3_U2811) );
  NAND2_X1 U21075 ( .A1(n17852), .A2(n18147), .ZN(n18202) );
  OAI22_X1 U21076 ( .A1(n18388), .A2(n18987), .B1(n17884), .B2(n17847), .ZN(
        n17848) );
  AOI221_X1 U21077 ( .B1(n17851), .B2(n17850), .C1(n17849), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17848), .ZN(n17857) );
  OAI21_X1 U21078 ( .B1(n17852), .B2(n17882), .A(n17881), .ZN(n17864) );
  AOI21_X1 U21079 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15863), .A(
        n17853), .ZN(n17855) );
  XNOR2_X1 U21080 ( .A(n17855), .B(n17854), .ZN(n18198) );
  AOI22_X1 U21081 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17864), .B1(
        n17989), .B2(n18198), .ZN(n17856) );
  OAI211_X1 U21082 ( .C1(n17882), .C2(n18202), .A(n17857), .B(n17856), .ZN(
        P3_U2812) );
  OAI21_X1 U21083 ( .B1(n17860), .B2(n18203), .A(n17859), .ZN(n18207) );
  AOI21_X1 U21084 ( .B1(n9966), .B2(n18741), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17862) );
  INV_X1 U21085 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18986) );
  OAI22_X1 U21086 ( .A1(n17862), .A2(n17861), .B1(n9975), .B2(n18986), .ZN(
        n17863) );
  AOI21_X1 U21087 ( .B1(n17989), .B2(n18207), .A(n17863), .ZN(n17867) );
  OAI221_X1 U21088 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17865), .A(n17864), .ZN(
        n17866) );
  OAI211_X1 U21089 ( .C1(n9826), .C2(n17868), .A(n17867), .B(n17866), .ZN(
        P3_U2813) );
  NAND3_X1 U21090 ( .A1(n15863), .A2(n18189), .A3(n17869), .ZN(n17967) );
  OAI21_X1 U21091 ( .B1(n18148), .B2(n17967), .A(n17870), .ZN(n17871) );
  XNOR2_X1 U21092 ( .A(n17871), .B(n18216), .ZN(n18213) );
  AOI21_X1 U21093 ( .B1(n17982), .B2(n17874), .A(n18055), .ZN(n17898) );
  OAI21_X1 U21094 ( .B1(n17872), .B2(n18936), .A(n17898), .ZN(n17886) );
  AOI22_X1 U21095 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17886), .B1(
        n17929), .B2(n17873), .ZN(n17878) );
  NOR2_X1 U21096 ( .A1(n17875), .A2(n17874), .ZN(n17888) );
  OAI211_X1 U21097 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17888), .B(n17876), .ZN(n17877) );
  OAI211_X1 U21098 ( .C1(n18983), .C2(n9975), .A(n17878), .B(n17877), .ZN(
        n17879) );
  AOI21_X1 U21099 ( .B1(n17989), .B2(n18213), .A(n17879), .ZN(n17880) );
  OAI221_X1 U21100 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17882), 
        .C1(n18216), .C2(n17881), .A(n17880), .ZN(P3_U2814) );
  AOI21_X1 U21101 ( .B1(n17900), .B2(n18271), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18226) );
  NAND2_X1 U21102 ( .A1(n17911), .A2(n18218), .ZN(n17893) );
  OAI22_X1 U21103 ( .A1(n18388), .A2(n18981), .B1(n17884), .B2(n17883), .ZN(
        n17885) );
  AOI221_X1 U21104 ( .B1(n17888), .B2(n17887), .C1(n17886), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17885), .ZN(n17892) );
  INV_X1 U21105 ( .A(n17910), .ZN(n18233) );
  NOR2_X1 U21106 ( .A1(n18233), .A2(n17967), .ZN(n17905) );
  NAND2_X1 U21107 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15850), .ZN(
        n17904) );
  OAI221_X1 U21108 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17906), 
        .C1(n17903), .C2(n17905), .A(n17904), .ZN(n17889) );
  XNOR2_X1 U21109 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17889), .ZN(
        n18227) );
  NAND4_X1 U21110 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17910), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n17947), .ZN(n17894) );
  NAND2_X1 U21111 ( .A1(n18231), .A2(n17894), .ZN(n18222) );
  AOI22_X1 U21112 ( .A1(n17989), .A2(n18227), .B1(n17890), .B2(n18222), .ZN(
        n17891) );
  OAI211_X1 U21113 ( .C1(n18226), .C2(n17893), .A(n17892), .B(n17891), .ZN(
        P3_U2815) );
  NAND2_X1 U21114 ( .A1(n17910), .A2(n17947), .ZN(n18249) );
  NOR2_X1 U21115 ( .A1(n15850), .A2(n18249), .ZN(n17895) );
  OAI21_X1 U21116 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17895), .A(
        n17894), .ZN(n18246) );
  AND2_X1 U21117 ( .A1(n18741), .A2(n17927), .ZN(n17943) );
  AOI21_X1 U21118 ( .B1(n17916), .B2(n17943), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17897) );
  OAI22_X1 U21119 ( .A1(n17898), .A2(n17897), .B1(n9826), .B2(n17896), .ZN(
        n17899) );
  AOI21_X1 U21120 ( .B1(n9832), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17899), .ZN(
        n17909) );
  INV_X1 U21121 ( .A(n17900), .ZN(n18219) );
  NOR2_X1 U21122 ( .A1(n17902), .A2(n18219), .ZN(n17901) );
  AOI221_X1 U21123 ( .B1(n18237), .B2(n17903), .C1(n17902), .C2(n17903), .A(
        n17901), .ZN(n18235) );
  OAI21_X1 U21124 ( .B1(n17906), .B2(n17905), .A(n17904), .ZN(n17907) );
  XNOR2_X1 U21125 ( .A(n17907), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18242) );
  AOI22_X1 U21126 ( .A1(n17911), .A2(n18235), .B1(n17989), .B2(n18242), .ZN(
        n17908) );
  OAI211_X1 U21127 ( .C1(n18088), .C2(n18246), .A(n17909), .B(n17908), .ZN(
        P3_U2816) );
  NAND2_X1 U21128 ( .A1(n18271), .A2(n17910), .ZN(n18247) );
  AOI22_X1 U21129 ( .A1(n17911), .A2(n18247), .B1(n17999), .B2(n18249), .ZN(
        n17937) );
  NOR2_X1 U21130 ( .A1(n18388), .A2(n18977), .ZN(n18255) );
  OAI211_X1 U21131 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17927), .B(n17926), .ZN(n17915) );
  OAI21_X1 U21132 ( .B1(n17927), .B2(n18044), .A(n18936), .ZN(n17912) );
  AOI21_X1 U21133 ( .B1(n17913), .B2(n17912), .A(n18055), .ZN(n17931) );
  OAI22_X1 U21134 ( .A1(n17916), .A2(n17915), .B1(n17931), .B2(n17914), .ZN(
        n17917) );
  AOI211_X1 U21135 ( .C1(n17929), .C2(n17918), .A(n18255), .B(n17917), .ZN(
        n17923) );
  OAI22_X1 U21136 ( .A1(n15863), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17952), .B2(n18233), .ZN(n17919) );
  OAI21_X1 U21137 ( .B1(n15863), .B2(n17924), .A(n17919), .ZN(n17920) );
  XOR2_X1 U21138 ( .A(n17920), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18258) );
  INV_X1 U21139 ( .A(n18258), .ZN(n17921) );
  NOR2_X1 U21140 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18233), .ZN(
        n18256) );
  AOI22_X1 U21141 ( .A1(n17989), .A2(n17921), .B1(n18256), .B2(n17974), .ZN(
        n17922) );
  OAI211_X1 U21142 ( .C1(n17937), .C2(n15850), .A(n17923), .B(n17922), .ZN(
        P3_U2817) );
  OAI21_X1 U21143 ( .B1(n18260), .B2(n17967), .A(n10045), .ZN(n17925) );
  XNOR2_X1 U21144 ( .A(n17925), .B(n18267), .ZN(n18259) );
  INV_X1 U21145 ( .A(n17974), .ZN(n17946) );
  NOR3_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17946), .A3(
        n18260), .ZN(n17935) );
  NAND2_X1 U21147 ( .A1(n17927), .A2(n17926), .ZN(n17933) );
  AOI22_X1 U21148 ( .A1(n9832), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n17929), 
        .B2(n17928), .ZN(n17930) );
  OAI221_X1 U21149 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17933), .C1(
        n17932), .C2(n17931), .A(n17930), .ZN(n17934) );
  AOI211_X1 U21150 ( .C1(n17989), .C2(n18259), .A(n17935), .B(n17934), .ZN(
        n17936) );
  OAI21_X1 U21151 ( .B1(n17937), .B2(n18267), .A(n17936), .ZN(P3_U2818) );
  INV_X1 U21152 ( .A(n18276), .ZN(n17955) );
  OAI21_X1 U21153 ( .B1(n17967), .B2(n17955), .A(n17938), .ZN(n17939) );
  XNOR2_X1 U21154 ( .A(n17939), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18281) );
  NOR2_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17955), .ZN(
        n18268) );
  NOR2_X1 U21156 ( .A1(n9975), .A2(n18973), .ZN(n17945) );
  NAND3_X1 U21157 ( .A1(n18741), .A2(n18015), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18003) );
  NOR2_X1 U21158 ( .A1(n17940), .A2(n18003), .ZN(n17959) );
  AOI21_X1 U21159 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18078), .A(
        n17959), .ZN(n17942) );
  OAI22_X1 U21160 ( .A1(n17943), .A2(n17942), .B1(n9826), .B2(n17941), .ZN(
        n17944) );
  AOI211_X1 U21161 ( .C1(n18268), .C2(n17974), .A(n17945), .B(n17944), .ZN(
        n17949) );
  NOR2_X1 U21162 ( .A1(n18276), .A2(n17946), .ZN(n17956) );
  OAI22_X1 U21163 ( .A1(n18271), .A2(n17992), .B1(n18088), .B2(n17947), .ZN(
        n17975) );
  OAI21_X1 U21164 ( .B1(n17956), .B2(n17975), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17948) );
  OAI211_X1 U21165 ( .C1(n18281), .C2(n17978), .A(n17949), .B(n17948), .ZN(
        P3_U2819) );
  OAI221_X1 U21166 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17966), .C1(
        n18290), .C2(n17967), .A(n17950), .ZN(n17954) );
  NAND4_X1 U21167 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17952), .A3(
        n17951), .A4(n18290), .ZN(n17953) );
  OAI211_X1 U21168 ( .C1(n17967), .C2(n17955), .A(n17954), .B(n17953), .ZN(
        n18289) );
  INV_X1 U21169 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18971) );
  NOR2_X1 U21170 ( .A1(n9975), .A2(n18971), .ZN(n17963) );
  NOR2_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17961) );
  AOI21_X1 U21172 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17975), .A(
        n17956), .ZN(n17960) );
  NAND2_X1 U21173 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17983) );
  NOR3_X1 U21174 ( .A1(n17983), .A2(n17957), .A3(n18003), .ZN(n17972) );
  AOI21_X1 U21175 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18078), .A(
        n17972), .ZN(n17958) );
  OAI22_X1 U21176 ( .A1(n17961), .A2(n17960), .B1(n17959), .B2(n17958), .ZN(
        n17962) );
  AOI211_X1 U21177 ( .C1(n17964), .C2(n9825), .A(n17963), .B(n17962), .ZN(
        n17965) );
  OAI21_X1 U21178 ( .B1(n17978), .B2(n18289), .A(n17965), .ZN(P3_U2820) );
  NAND2_X1 U21179 ( .A1(n17967), .A2(n17966), .ZN(n17968) );
  XNOR2_X1 U21180 ( .A(n17968), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18300) );
  NOR2_X1 U21181 ( .A1(n17983), .A2(n18003), .ZN(n17969) );
  AOI21_X1 U21182 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18078), .A(
        n17969), .ZN(n17971) );
  OAI22_X1 U21183 ( .A1(n17972), .A2(n17971), .B1(n9826), .B2(n17970), .ZN(
        n17973) );
  AOI21_X1 U21184 ( .B1(n9832), .B2(P3_REIP_REG_9__SCAN_IN), .A(n17973), .ZN(
        n17977) );
  AOI22_X1 U21185 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17975), .B1(
        n17974), .B2(n18290), .ZN(n17976) );
  OAI211_X1 U21186 ( .C1(n18300), .C2(n17978), .A(n17977), .B(n17976), .ZN(
        P3_U2821) );
  AOI21_X1 U21187 ( .B1(n17980), .B2(n18319), .A(n17979), .ZN(n18303) );
  AOI21_X1 U21188 ( .B1(n17982), .B2(n17981), .A(n18055), .ZN(n18001) );
  OAI211_X1 U21189 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17984), .A(
        n18741), .B(n17983), .ZN(n17985) );
  NAND2_X1 U21190 ( .A1(n9832), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18317) );
  OAI211_X1 U21191 ( .C1(n18001), .C2(n17986), .A(n17985), .B(n18317), .ZN(
        n17987) );
  AOI21_X1 U21192 ( .B1(n17999), .B2(n18303), .A(n17987), .ZN(n17991) );
  AOI21_X1 U21193 ( .B1(n15863), .B2(n18312), .A(n9941), .ZN(n18314) );
  AOI22_X1 U21194 ( .A1(n17989), .A2(n18314), .B1(n17988), .B2(n9825), .ZN(
        n17990) );
  OAI211_X1 U21195 ( .C1(n17992), .C2(n18312), .A(n17991), .B(n17990), .ZN(
        P3_U2822) );
  AOI21_X1 U21196 ( .B1(n18301), .B2(n17994), .A(n17993), .ZN(n18320) );
  OAI21_X1 U21197 ( .B1(n17997), .B2(n17996), .A(n17995), .ZN(n17998) );
  XNOR2_X1 U21198 ( .A(n17998), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18321) );
  AOI22_X1 U21199 ( .A1(n17999), .A2(n18321), .B1(n9832), .B2(
        P3_REIP_REG_7__SCAN_IN), .ZN(n18000) );
  OAI221_X1 U21200 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18003), .C1(
        n18002), .C2(n18001), .A(n18000), .ZN(n18004) );
  AOI21_X1 U21201 ( .B1(n18076), .B2(n18320), .A(n18004), .ZN(n18005) );
  OAI21_X1 U21202 ( .B1(n9826), .B2(n18006), .A(n18005), .ZN(P3_U2823) );
  AOI22_X1 U21203 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18009), .B1(
        n18008), .B2(n18007), .ZN(n18014) );
  AOI22_X1 U21204 ( .A1(n18012), .A2(n18029), .B1(n18011), .B2(n18010), .ZN(
        n18013) );
  XNOR2_X1 U21205 ( .A(n18014), .B(n18013), .ZN(n18338) );
  NAND2_X1 U21206 ( .A1(n18741), .A2(n18015), .ZN(n18020) );
  NAND2_X1 U21207 ( .A1(n18078), .A2(n18020), .ZN(n18035) );
  AOI21_X1 U21208 ( .B1(n9954), .B2(n18017), .A(n18016), .ZN(n18335) );
  AOI22_X1 U21209 ( .A1(n18076), .A2(n18335), .B1(n9832), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18018) );
  OAI221_X1 U21210 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18020), .C1(
        n18019), .C2(n18035), .A(n18018), .ZN(n18021) );
  AOI21_X1 U21211 ( .B1(n18022), .B2(n9825), .A(n18021), .ZN(n18023) );
  OAI21_X1 U21212 ( .B1(n18338), .B2(n18088), .A(n18023), .ZN(P3_U2824) );
  INV_X1 U21213 ( .A(n18024), .ZN(n18025) );
  AOI21_X1 U21214 ( .B1(n18025), .B2(n18083), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18036) );
  AOI21_X1 U21215 ( .B1(n18028), .B2(n18027), .A(n18026), .ZN(n18344) );
  NOR2_X1 U21216 ( .A1(n9975), .A2(n18962), .ZN(n18343) );
  OAI21_X1 U21217 ( .B1(n18031), .B2(n18030), .A(n18029), .ZN(n18346) );
  OAI22_X1 U21218 ( .A1(n9826), .A2(n18032), .B1(n18088), .B2(n18346), .ZN(
        n18033) );
  AOI211_X1 U21219 ( .C1(n18076), .C2(n18344), .A(n18343), .B(n18033), .ZN(
        n18034) );
  OAI21_X1 U21220 ( .B1(n18036), .B2(n18035), .A(n18034), .ZN(P3_U2825) );
  OAI21_X1 U21221 ( .B1(n18039), .B2(n18038), .A(n18037), .ZN(n18355) );
  AOI21_X1 U21222 ( .B1(n18041), .B2(n18040), .A(n9962), .ZN(n18353) );
  OAI22_X1 U21223 ( .A1(n9975), .A2(n18959), .B1(n18797), .B2(n18042), .ZN(
        n18043) );
  AOI21_X1 U21224 ( .B1(n18076), .B2(n18353), .A(n18043), .ZN(n18048) );
  OAI21_X1 U21225 ( .B1(n18045), .B2(n18044), .A(n18083), .ZN(n18058) );
  AOI22_X1 U21226 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18058), .B1(
        n18046), .B2(n9825), .ZN(n18047) );
  OAI211_X1 U21227 ( .C1(n18088), .C2(n18355), .A(n18048), .B(n18047), .ZN(
        P3_U2826) );
  OAI21_X1 U21228 ( .B1(n18051), .B2(n18050), .A(n18049), .ZN(n18364) );
  AOI21_X1 U21229 ( .B1(n18358), .B2(n18053), .A(n18052), .ZN(n18356) );
  AOI22_X1 U21230 ( .A1(n18076), .A2(n18356), .B1(n9832), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18060) );
  OAI21_X1 U21231 ( .B1(n18055), .B2(n18071), .A(n18054), .ZN(n18057) );
  AOI22_X1 U21232 ( .A1(n18058), .A2(n18057), .B1(n18056), .B2(n9825), .ZN(
        n18059) );
  OAI211_X1 U21233 ( .C1(n18088), .C2(n18364), .A(n18060), .B(n18059), .ZN(
        P3_U2827) );
  AOI21_X1 U21234 ( .B1(n18063), .B2(n18062), .A(n18061), .ZN(n18375) );
  NOR2_X1 U21235 ( .A1(n18388), .A2(n18955), .ZN(n18374) );
  OAI21_X1 U21236 ( .B1(n18066), .B2(n18065), .A(n18064), .ZN(n18370) );
  OAI22_X1 U21237 ( .A1(n9826), .A2(n18067), .B1(n18088), .B2(n18370), .ZN(
        n18069) );
  AOI211_X1 U21238 ( .C1(n18076), .C2(n18375), .A(n18374), .B(n18069), .ZN(
        n18070) );
  OAI221_X1 U21239 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18797), .C1(
        n18071), .C2(n18083), .A(n18070), .ZN(P3_U2828) );
  AOI21_X1 U21240 ( .B1(n18073), .B2(n18081), .A(n18072), .ZN(n18387) );
  AOI21_X1 U21241 ( .B1(n18075), .B2(n18082), .A(n18074), .ZN(n18382) );
  AOI22_X1 U21242 ( .A1(n18076), .A2(n18382), .B1(n9832), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18080) );
  AOI22_X1 U21243 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18078), .B1(
        n9825), .B2(n18077), .ZN(n18079) );
  OAI211_X1 U21244 ( .C1(n18387), .C2(n18088), .A(n18080), .B(n18079), .ZN(
        P3_U2829) );
  NAND2_X1 U21245 ( .A1(n18082), .A2(n18081), .ZN(n18087) );
  INV_X1 U21246 ( .A(n18087), .ZN(n18396) );
  NAND3_X1 U21247 ( .A1(n19042), .A2(n18936), .A3(n18083), .ZN(n18084) );
  AOI22_X1 U21248 ( .A1(n9832), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18084), .ZN(n18085) );
  OAI221_X1 U21249 ( .B1(n18396), .B2(n18088), .C1(n18087), .C2(n18086), .A(
        n18085), .ZN(P3_U2830) );
  NAND2_X1 U21250 ( .A1(n9832), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18100) );
  INV_X1 U21251 ( .A(n18126), .ZN(n18103) );
  NOR3_X1 U21252 ( .A1(n18105), .A2(n18104), .A3(n18103), .ZN(n18098) );
  NAND2_X1 U21253 ( .A1(n18882), .A2(n9820), .ZN(n18090) );
  INV_X1 U21254 ( .A(n18192), .ZN(n18305) );
  OAI221_X1 U21255 ( .B1(n18307), .B2(n18112), .C1(n18307), .C2(n18127), .A(
        n18305), .ZN(n18113) );
  AOI211_X1 U21256 ( .C1(n18091), .C2(n18090), .A(n18089), .B(n18113), .ZN(
        n18092) );
  OAI21_X1 U21257 ( .B1(n18093), .B2(n18313), .A(n18092), .ZN(n18094) );
  AOI21_X1 U21258 ( .B1(n18868), .B2(n18095), .A(n18094), .ZN(n18102) );
  NAND2_X1 U21259 ( .A1(n18102), .A2(n18328), .ZN(n18096) );
  OAI221_X1 U21260 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18098), 
        .C1(n18097), .C2(n18096), .A(n9975), .ZN(n18099) );
  OAI211_X1 U21261 ( .C1(n18101), .C2(n18299), .A(n18100), .B(n18099), .ZN(
        P3_U2835) );
  INV_X1 U21262 ( .A(n18102), .ZN(n18107) );
  OAI22_X1 U21263 ( .A1(n18105), .A2(n18392), .B1(n18104), .B2(n18103), .ZN(
        n18106) );
  AOI22_X1 U21264 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18384), .B1(
        n18107), .B2(n18106), .ZN(n18109) );
  OAI211_X1 U21265 ( .C1(n18110), .C2(n18299), .A(n18109), .B(n18108), .ZN(
        P3_U2836) );
  NAND2_X1 U21266 ( .A1(n18111), .A2(n18112), .ZN(n18120) );
  AOI21_X1 U21267 ( .B1(n18112), .B2(n18132), .A(n10174), .ZN(n18114) );
  NOR2_X1 U21268 ( .A1(n18114), .A2(n18113), .ZN(n18118) );
  AOI22_X1 U21269 ( .A1(n18868), .A2(n18116), .B1(n18248), .B2(n18115), .ZN(
        n18117) );
  OAI221_X1 U21270 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18120), 
        .C1(n18119), .C2(n18118), .A(n18117), .ZN(n18121) );
  AOI22_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18384), .B1(
        n18328), .B2(n18121), .ZN(n18123) );
  OAI211_X1 U21272 ( .C1(n18124), .C2(n18299), .A(n18123), .B(n18122), .ZN(
        P3_U2837) );
  AOI22_X1 U21273 ( .A1(n9832), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18126), 
        .B2(n18125), .ZN(n18138) );
  OAI21_X1 U21274 ( .B1(n18307), .B2(n18127), .A(n18305), .ZN(n18128) );
  AOI211_X1 U21275 ( .C1(n18868), .C2(n18129), .A(n18384), .B(n18128), .ZN(
        n18130) );
  OAI21_X1 U21276 ( .B1(n18131), .B2(n18313), .A(n18130), .ZN(n18136) );
  NOR2_X1 U21277 ( .A1(n18132), .A2(n10174), .ZN(n18134) );
  NOR3_X1 U21278 ( .A1(n18134), .A2(n18133), .A3(n18136), .ZN(n18135) );
  NOR2_X1 U21279 ( .A1(n18135), .A2(n9832), .ZN(n18141) );
  OAI211_X1 U21280 ( .C1(n18309), .C2(n18136), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18141), .ZN(n18137) );
  OAI211_X1 U21281 ( .C1(n18139), .C2(n18299), .A(n18138), .B(n18137), .ZN(
        P3_U2838) );
  NOR2_X1 U21282 ( .A1(n18384), .A2(n18140), .ZN(n18143) );
  OAI221_X1 U21283 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18143), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18142), .A(n18141), .ZN(
        n18144) );
  OAI211_X1 U21284 ( .C1(n18146), .C2(n18299), .A(n18145), .B(n18144), .ZN(
        P3_U2839) );
  AOI22_X1 U21285 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18384), .B1(
        n9832), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n18163) );
  OR3_X1 U21286 ( .A1(n18197), .A2(n18147), .A3(n18193), .ZN(n18154) );
  NAND2_X1 U21287 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18209), .ZN(
        n18292) );
  NOR2_X1 U21288 ( .A1(n18148), .A2(n18292), .ZN(n18211) );
  AOI21_X1 U21289 ( .B1(n18149), .B2(n18211), .A(n18882), .ZN(n18153) );
  INV_X1 U21290 ( .A(n18150), .ZN(n18174) );
  OAI21_X1 U21291 ( .B1(n18191), .B2(n18174), .A(n18874), .ZN(n18151) );
  INV_X1 U21292 ( .A(n18151), .ZN(n18152) );
  AOI211_X1 U21293 ( .C1(n18890), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        n18176) );
  NAND2_X1 U21294 ( .A1(n10170), .A2(n18313), .ZN(n18269) );
  NAND2_X1 U21295 ( .A1(n18158), .A2(n18269), .ZN(n18155) );
  OAI211_X1 U21296 ( .C1(n18308), .C2(n18156), .A(n18176), .B(n18155), .ZN(
        n18169) );
  NOR2_X1 U21297 ( .A1(n18157), .A2(n10170), .ZN(n18223) );
  AOI21_X1 U21298 ( .B1(n18248), .B2(n18218), .A(n18223), .ZN(n18168) );
  OAI211_X1 U21299 ( .C1(n18308), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18168), .ZN(n18161) );
  OAI22_X1 U21300 ( .A1(n18159), .A2(n18392), .B1(n18165), .B2(n18158), .ZN(
        n18160) );
  OAI21_X1 U21301 ( .B1(n18169), .B2(n18161), .A(n18160), .ZN(n18162) );
  OAI211_X1 U21302 ( .C1(n18164), .C2(n18299), .A(n18163), .B(n18162), .ZN(
        P3_U2840) );
  AOI22_X1 U21303 ( .A1(n9832), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18315), 
        .B2(n18167), .ZN(n18171) );
  NAND2_X1 U21304 ( .A1(n18328), .A2(n18168), .ZN(n18212) );
  OAI211_X1 U21305 ( .C1(n18212), .C2(n18169), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n9975), .ZN(n18170) );
  OAI211_X1 U21306 ( .C1(n18172), .C2(n18186), .A(n18171), .B(n18170), .ZN(
        P3_U2841) );
  AOI22_X1 U21307 ( .A1(n9832), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18315), 
        .B2(n18173), .ZN(n18180) );
  AOI21_X1 U21308 ( .B1(n18174), .B2(n18269), .A(n18212), .ZN(n18175) );
  AOI21_X1 U21309 ( .B1(n18176), .B2(n18175), .A(n9832), .ZN(n18183) );
  NOR3_X1 U21310 ( .A1(n18383), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n18177), .ZN(n18178) );
  OAI21_X1 U21311 ( .B1(n18183), .B2(n18178), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18179) );
  OAI211_X1 U21312 ( .C1(n18181), .C2(n18186), .A(n18180), .B(n18179), .ZN(
        P3_U2842) );
  AOI22_X1 U21313 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18183), .B1(
        n18315), .B2(n18182), .ZN(n18185) );
  OAI211_X1 U21314 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18186), .A(
        n18185), .B(n18184), .ZN(P3_U2843) );
  OAI22_X1 U21315 ( .A1(n18304), .A2(n10174), .B1(n18187), .B2(n18366), .ZN(
        n18357) );
  NAND2_X1 U21316 ( .A1(n18189), .A2(n18324), .ZN(n18261) );
  AOI21_X1 U21317 ( .B1(n18262), .B2(n18261), .A(n18392), .ZN(n18291) );
  NAND2_X1 U21318 ( .A1(n18190), .A2(n18291), .ZN(n18217) );
  NOR3_X1 U21319 ( .A1(n18192), .A2(n18191), .A3(n18216), .ZN(n18195) );
  NOR2_X1 U21320 ( .A1(n18197), .A2(n18193), .ZN(n18194) );
  OAI22_X1 U21321 ( .A1(n18307), .A2(n18195), .B1(n18194), .B2(n10174), .ZN(
        n18196) );
  AOI211_X1 U21322 ( .C1(n18197), .C2(n18269), .A(n18212), .B(n18196), .ZN(
        n18204) );
  AOI221_X1 U21323 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18204), 
        .C1(n18307), .C2(n18204), .A(n9832), .ZN(n18199) );
  AOI22_X1 U21324 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18199), .B1(
        n18315), .B2(n18198), .ZN(n18201) );
  NAND2_X1 U21325 ( .A1(n9832), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18200) );
  OAI211_X1 U21326 ( .C1(n18202), .C2(n18217), .A(n18201), .B(n18200), .ZN(
        P3_U2844) );
  NOR3_X1 U21327 ( .A1(n9832), .A2(n18204), .A3(n18203), .ZN(n18206) );
  NOR3_X1 U21328 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18216), .A3(
        n18217), .ZN(n18205) );
  AOI211_X1 U21329 ( .C1(n18315), .C2(n18207), .A(n18206), .B(n18205), .ZN(
        n18208) );
  OAI21_X1 U21330 ( .B1(n9975), .B2(n18986), .A(n18208), .ZN(P3_U2845) );
  NOR2_X1 U21331 ( .A1(n9820), .A2(n18209), .ZN(n18250) );
  INV_X1 U21332 ( .A(n18250), .ZN(n18293) );
  OAI21_X1 U21333 ( .B1(n18270), .B2(n10174), .A(n18293), .ZN(n18232) );
  AOI21_X1 U21334 ( .B1(n18219), .B2(n18283), .A(n18232), .ZN(n18210) );
  OAI211_X1 U21335 ( .C1(n18211), .C2(n18882), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18210), .ZN(n18221) );
  OAI221_X1 U21336 ( .B1(n18212), .B2(n18309), .C1(n18212), .C2(n18221), .A(
        n9975), .ZN(n18215) );
  AOI22_X1 U21337 ( .A1(n9832), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18315), 
        .B2(n18213), .ZN(n18214) );
  OAI221_X1 U21338 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18217), 
        .C1(n18216), .C2(n18215), .A(n18214), .ZN(P3_U2846) );
  NAND2_X1 U21339 ( .A1(n18248), .A2(n18218), .ZN(n18225) );
  OAI21_X1 U21340 ( .B1(n18219), .B2(n18261), .A(n18231), .ZN(n18220) );
  AOI22_X1 U21341 ( .A1(n18223), .A2(n18222), .B1(n18221), .B2(n18220), .ZN(
        n18224) );
  OAI21_X1 U21342 ( .B1(n18226), .B2(n18225), .A(n18224), .ZN(n18228) );
  AOI22_X1 U21343 ( .A1(n18328), .A2(n18228), .B1(n18315), .B2(n18227), .ZN(
        n18230) );
  NAND2_X1 U21344 ( .A1(n9832), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18229) );
  OAI211_X1 U21345 ( .C1(n18371), .C2(n18231), .A(n18230), .B(n18229), .ZN(
        P3_U2847) );
  AOI22_X1 U21346 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18384), .B1(
        n9832), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18245) );
  AOI221_X1 U21347 ( .B1(n18233), .B2(n18892), .C1(n18292), .C2(n18892), .A(
        n18232), .ZN(n18252) );
  AOI22_X1 U21348 ( .A1(n18890), .A2(n18233), .B1(n18874), .B2(n18237), .ZN(
        n18234) );
  OAI211_X1 U21349 ( .C1(n18383), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18252), .B(n18234), .ZN(n18236) );
  AOI22_X1 U21350 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18236), .B1(
        n18248), .B2(n18235), .ZN(n18241) );
  INV_X1 U21351 ( .A(n18237), .ZN(n18239) );
  INV_X1 U21352 ( .A(n18261), .ZN(n18238) );
  NAND3_X1 U21353 ( .A1(n18239), .A2(n17903), .A3(n18238), .ZN(n18240) );
  NAND2_X1 U21354 ( .A1(n18241), .A2(n18240), .ZN(n18243) );
  AOI22_X1 U21355 ( .A1(n18328), .A2(n18243), .B1(n18315), .B2(n18242), .ZN(
        n18244) );
  OAI211_X1 U21356 ( .C1(n18395), .C2(n18246), .A(n18245), .B(n18244), .ZN(
        P3_U2848) );
  AOI22_X1 U21357 ( .A1(n18868), .A2(n18249), .B1(n18248), .B2(n18247), .ZN(
        n18251) );
  OAI21_X1 U21358 ( .B1(n18250), .B2(n18260), .A(n18283), .ZN(n18277) );
  NAND3_X1 U21359 ( .A1(n18252), .A2(n18251), .A3(n18277), .ZN(n18263) );
  AOI211_X1 U21360 ( .C1(n18267), .C2(n18283), .A(n18392), .B(n18263), .ZN(
        n18253) );
  NOR3_X1 U21361 ( .A1(n9832), .A2(n18253), .A3(n15850), .ZN(n18254) );
  AOI211_X1 U21362 ( .C1(n18256), .C2(n18291), .A(n18255), .B(n18254), .ZN(
        n18257) );
  OAI21_X1 U21363 ( .B1(n18299), .B2(n18258), .A(n18257), .ZN(P3_U2849) );
  AOI22_X1 U21364 ( .A1(n9832), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18315), 
        .B2(n18259), .ZN(n18266) );
  AOI21_X1 U21365 ( .B1(n18262), .B2(n18261), .A(n18260), .ZN(n18264) );
  OAI221_X1 U21366 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18264), 
        .C1(n18267), .C2(n18263), .A(n18328), .ZN(n18265) );
  OAI211_X1 U21367 ( .C1(n18371), .C2(n18267), .A(n18266), .B(n18265), .ZN(
        P3_U2850) );
  AOI22_X1 U21368 ( .A1(n9832), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18291), 
        .B2(n18268), .ZN(n18280) );
  INV_X1 U21369 ( .A(n18269), .ZN(n18275) );
  OAI22_X1 U21370 ( .A1(n18271), .A2(n18313), .B1(n18270), .B2(n10174), .ZN(
        n18272) );
  AOI211_X1 U21371 ( .C1(n18868), .C2(n18273), .A(n18392), .B(n18272), .ZN(
        n18294) );
  OAI21_X1 U21372 ( .B1(n18290), .B2(n18292), .A(n18892), .ZN(n18274) );
  OAI211_X1 U21373 ( .C1(n18276), .C2(n18275), .A(n18294), .B(n18274), .ZN(
        n18286) );
  OAI21_X1 U21374 ( .B1(n18882), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18277), .ZN(n18278) );
  OAI211_X1 U21375 ( .C1(n18286), .C2(n18278), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9975), .ZN(n18279) );
  OAI211_X1 U21376 ( .C1(n18281), .C2(n18299), .A(n18280), .B(n18279), .ZN(
        P3_U2851) );
  NOR2_X1 U21377 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18290), .ZN(
        n18282) );
  AOI22_X1 U21378 ( .A1(n9832), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18291), 
        .B2(n18282), .ZN(n18288) );
  INV_X1 U21379 ( .A(n18283), .ZN(n18284) );
  OAI21_X1 U21380 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18284), .A(
        n18293), .ZN(n18285) );
  OAI211_X1 U21381 ( .C1(n18286), .C2(n18285), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n9975), .ZN(n18287) );
  OAI211_X1 U21382 ( .C1(n18299), .C2(n18289), .A(n18288), .B(n18287), .ZN(
        P3_U2852) );
  AOI22_X1 U21383 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n9832), .B1(n18291), .B2(
        n18290), .ZN(n18298) );
  INV_X1 U21384 ( .A(n18292), .ZN(n18295) );
  OAI211_X1 U21385 ( .C1(n18882), .C2(n18295), .A(n18294), .B(n18293), .ZN(
        n18296) );
  NAND3_X1 U21386 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n9975), .A3(
        n18296), .ZN(n18297) );
  OAI211_X1 U21387 ( .C1(n18300), .C2(n18299), .A(n18298), .B(n18297), .ZN(
        P3_U2853) );
  NOR2_X1 U21388 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18301), .ZN(
        n18302) );
  AOI22_X1 U21389 ( .A1(n18868), .A2(n18303), .B1(n18324), .B2(n18302), .ZN(
        n18311) );
  INV_X1 U21390 ( .A(n18366), .ZN(n18306) );
  NAND2_X1 U21391 ( .A1(n18890), .A2(n18304), .ZN(n18365) );
  OAI211_X1 U21392 ( .C1(n18307), .C2(n18306), .A(n18365), .B(n18305), .ZN(
        n18369) );
  AOI21_X1 U21393 ( .B1(n18309), .B2(n18329), .A(n18369), .ZN(n18330) );
  OAI211_X1 U21394 ( .C1(n18308), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18330), .ZN(n18323) );
  NAND3_X1 U21395 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18309), .A3(
        n18323), .ZN(n18310) );
  OAI211_X1 U21396 ( .C1(n18313), .C2(n18312), .A(n18311), .B(n18310), .ZN(
        n18316) );
  AOI22_X1 U21397 ( .A1(n18328), .A2(n18316), .B1(n18315), .B2(n18314), .ZN(
        n18318) );
  OAI211_X1 U21398 ( .C1(n18371), .C2(n18319), .A(n18318), .B(n18317), .ZN(
        P3_U2854) );
  AOI22_X1 U21399 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18384), .B1(
        n9832), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18327) );
  AOI22_X1 U21400 ( .A1(n18322), .A2(n18321), .B1(n18391), .B2(n18320), .ZN(
        n18326) );
  OAI211_X1 U21401 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18324), .A(
        n18328), .B(n18323), .ZN(n18325) );
  NAND3_X1 U21402 ( .A1(n18327), .A2(n18326), .A3(n18325), .ZN(P3_U2855) );
  NAND2_X1 U21403 ( .A1(n18328), .A2(n18357), .ZN(n18339) );
  NOR2_X1 U21404 ( .A1(n18329), .A2(n18339), .ZN(n18333) );
  INV_X1 U21405 ( .A(n18330), .ZN(n18331) );
  OAI21_X1 U21406 ( .B1(n18392), .B2(n18331), .A(n18388), .ZN(n18332) );
  INV_X1 U21407 ( .A(n18332), .ZN(n18340) );
  MUX2_X1 U21408 ( .A(n18333), .B(n18340), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n18334) );
  AOI21_X1 U21409 ( .B1(n18391), .B2(n18335), .A(n18334), .ZN(n18337) );
  NAND2_X1 U21410 ( .A1(n9832), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18336) );
  OAI211_X1 U21411 ( .C1(n18338), .C2(n18395), .A(n18337), .B(n18336), .ZN(
        P3_U2856) );
  OR2_X1 U21412 ( .A1(n18358), .A2(n18339), .ZN(n18349) );
  NOR2_X1 U21413 ( .A1(n18348), .A2(n18349), .ZN(n18341) );
  MUX2_X1 U21414 ( .A(n18341), .B(n18340), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18342) );
  AOI211_X1 U21415 ( .C1(n18391), .C2(n18344), .A(n18343), .B(n18342), .ZN(
        n18345) );
  OAI21_X1 U21416 ( .B1(n18395), .B2(n18346), .A(n18345), .ZN(P3_U2857) );
  NOR2_X1 U21417 ( .A1(n9975), .A2(n18959), .ZN(n18352) );
  OR2_X1 U21418 ( .A1(n18358), .A2(n18369), .ZN(n18360) );
  AOI21_X1 U21419 ( .B1(n18347), .B2(n18360), .A(n18384), .ZN(n18350) );
  AOI22_X1 U21420 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18350), .B1(
        n18349), .B2(n18348), .ZN(n18351) );
  AOI211_X1 U21421 ( .C1(n18391), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        n18354) );
  OAI21_X1 U21422 ( .B1(n18395), .B2(n18355), .A(n18354), .ZN(P3_U2858) );
  AOI22_X1 U21423 ( .A1(n9832), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18391), .B2(
        n18356), .ZN(n18363) );
  INV_X1 U21424 ( .A(n18357), .ZN(n18359) );
  AOI21_X1 U21425 ( .B1(n18359), .B2(n18358), .A(n18392), .ZN(n18361) );
  AOI22_X1 U21426 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18384), .B1(
        n18361), .B2(n18360), .ZN(n18362) );
  OAI211_X1 U21427 ( .C1(n18395), .C2(n18364), .A(n18363), .B(n18362), .ZN(
        P3_U2859) );
  NOR2_X1 U21428 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18874), .ZN(
        n18379) );
  INV_X1 U21429 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19041) );
  OAI211_X1 U21430 ( .C1(n18379), .C2(n19041), .A(n18372), .B(n18365), .ZN(
        n18368) );
  NOR3_X1 U21431 ( .A1(n10174), .A2(n19059), .A3(n18366), .ZN(n18367) );
  AOI21_X1 U21432 ( .B1(n18369), .B2(n18368), .A(n18367), .ZN(n18377) );
  OAI22_X1 U21433 ( .A1(n18372), .A2(n18371), .B1(n18395), .B2(n18370), .ZN(
        n18373) );
  AOI211_X1 U21434 ( .C1(n18391), .C2(n18375), .A(n18374), .B(n18373), .ZN(
        n18376) );
  OAI21_X1 U21435 ( .B1(n18377), .B2(n18392), .A(n18376), .ZN(P3_U2860) );
  NOR2_X1 U21436 ( .A1(n9975), .A2(n19063), .ZN(n18381) );
  NOR3_X1 U21437 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18379), .A3(
        n18378), .ZN(n18380) );
  AOI211_X1 U21438 ( .C1(n18391), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        n18386) );
  NOR3_X1 U21439 ( .A1(n18383), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18392), .ZN(n18389) );
  OAI21_X1 U21440 ( .B1(n18384), .B2(n18389), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18385) );
  OAI211_X1 U21441 ( .C1(n18387), .C2(n18395), .A(n18386), .B(n18385), .ZN(
        P3_U2861) );
  INV_X1 U21442 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19069) );
  NOR2_X1 U21443 ( .A1(n9975), .A2(n19069), .ZN(n18390) );
  AOI211_X1 U21444 ( .C1(n18391), .C2(n18396), .A(n18390), .B(n18389), .ZN(
        n18394) );
  OAI211_X1 U21445 ( .C1(n18874), .C2(n18392), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n9975), .ZN(n18393) );
  OAI211_X1 U21446 ( .C1(n18396), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        P3_U2862) );
  OAI211_X1 U21447 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18397), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18922)
         );
  INV_X1 U21448 ( .A(n18398), .ZN(n18455) );
  OAI21_X1 U21449 ( .B1(n18400), .B2(n19077), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18399) );
  OAI221_X1 U21450 ( .B1(n18400), .B2(n18922), .C1(n18400), .C2(n18455), .A(
        n18399), .ZN(P3_U2863) );
  INV_X1 U21451 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18589) );
  NOR2_X1 U21452 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18589), .ZN(
        n18712) );
  NOR2_X1 U21453 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18903), .ZN(
        n18592) );
  NOR2_X1 U21454 ( .A1(n18712), .A2(n18592), .ZN(n18402) );
  OAI22_X1 U21455 ( .A1(n18403), .A2(n18589), .B1(n18402), .B2(n18401), .ZN(
        P3_U2866) );
  NOR2_X1 U21456 ( .A1(n18405), .A2(n18404), .ZN(P3_U2867) );
  NOR2_X1 U21457 ( .A1(n18897), .A2(n19031), .ZN(n18407) );
  INV_X1 U21458 ( .A(n18406), .ZN(n18588) );
  NAND2_X1 U21459 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18588), .ZN(
        n18798) );
  NOR2_X1 U21460 ( .A1(n18897), .A2(n18798), .ZN(n18845) );
  INV_X1 U21461 ( .A(n18845), .ZN(n18841) );
  INV_X1 U21462 ( .A(n18841), .ZN(n18855) );
  NAND2_X1 U21463 ( .A1(n18898), .A2(n18897), .ZN(n18899) );
  NAND2_X1 U21464 ( .A1(n18903), .A2(n18589), .ZN(n18496) );
  NOR2_X1 U21465 ( .A1(n18899), .A2(n18496), .ZN(n18515) );
  OAI21_X1 U21466 ( .B1(n18855), .B2(n18511), .A(n18765), .ZN(n18475) );
  NOR2_X1 U21467 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18898), .ZN(
        n18668) );
  NOR2_X1 U21468 ( .A1(n18897), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18643) );
  NOR2_X1 U21469 ( .A1(n18668), .A2(n18643), .ZN(n18716) );
  OR3_X1 U21470 ( .A1(n18589), .A2(n18903), .A3(n18716), .ZN(n18761) );
  OAI22_X1 U21471 ( .A1(n18407), .A2(n18475), .B1(n18797), .B2(n18761), .ZN(
        n18453) );
  NAND3_X1 U21472 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18668), .ZN(n18794) );
  AND2_X1 U21473 ( .A1(n18741), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18801) );
  AND2_X1 U21474 ( .A1(n18765), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18800) );
  OAI21_X1 U21475 ( .B1(n18855), .B2(n18511), .A(n18926), .ZN(n18408) );
  INV_X1 U21476 ( .A(n18408), .ZN(n18448) );
  AOI22_X1 U21477 ( .A1(n18767), .A2(n18801), .B1(n18800), .B2(n18448), .ZN(
        n18414) );
  NAND3_X1 U21478 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18898), .ZN(n18796) );
  INV_X1 U21479 ( .A(n18796), .ZN(n18739) );
  NAND2_X1 U21480 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18739), .ZN(
        n18763) );
  INV_X1 U21481 ( .A(n18763), .ZN(n18858) );
  NOR2_X2 U21482 ( .A1(n18409), .A2(n18797), .ZN(n18803) );
  NOR2_X1 U21483 ( .A1(n18411), .A2(n18410), .ZN(n18450) );
  NAND2_X1 U21484 ( .A1(n18450), .A2(n18412), .ZN(n18770) );
  INV_X1 U21485 ( .A(n18770), .ZN(n18802) );
  AOI22_X1 U21486 ( .A1(n18858), .A2(n18803), .B1(n18802), .B2(n18515), .ZN(
        n18413) );
  OAI211_X1 U21487 ( .C1(n18415), .C2(n18453), .A(n18414), .B(n18413), .ZN(
        P3_U2868) );
  AND2_X1 U21488 ( .A1(n18741), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18808) );
  AND2_X1 U21489 ( .A1(n18765), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18807) );
  AOI22_X1 U21490 ( .A1(n18767), .A2(n18808), .B1(n18807), .B2(n18448), .ZN(
        n18418) );
  NOR2_X2 U21491 ( .A1(n19525), .A2(n18797), .ZN(n18810) );
  NAND2_X1 U21492 ( .A1(n18450), .A2(n18416), .ZN(n18773) );
  INV_X1 U21493 ( .A(n18773), .ZN(n18809) );
  AOI22_X1 U21494 ( .A1(n18858), .A2(n18810), .B1(n18809), .B2(n18515), .ZN(
        n18417) );
  OAI211_X1 U21495 ( .C1(n18419), .C2(n18453), .A(n18418), .B(n18417), .ZN(
        P3_U2869) );
  AND2_X1 U21496 ( .A1(n18741), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18815) );
  NOR2_X2 U21497 ( .A1(n18565), .A2(n18420), .ZN(n18814) );
  AOI22_X1 U21498 ( .A1(n18767), .A2(n18815), .B1(n18814), .B2(n18448), .ZN(
        n18423) );
  NOR2_X2 U21499 ( .A1(n19530), .A2(n18797), .ZN(n18817) );
  NAND2_X1 U21500 ( .A1(n18450), .A2(n18421), .ZN(n18776) );
  INV_X1 U21501 ( .A(n18776), .ZN(n18816) );
  AOI22_X1 U21502 ( .A1(n18858), .A2(n18817), .B1(n18816), .B2(n18515), .ZN(
        n18422) );
  OAI211_X1 U21503 ( .C1(n18424), .C2(n18453), .A(n18423), .B(n18422), .ZN(
        P3_U2870) );
  NOR2_X2 U21504 ( .A1(n18797), .A2(n14030), .ZN(n18824) );
  NOR2_X2 U21505 ( .A1(n18565), .A2(n18425), .ZN(n18821) );
  AOI22_X1 U21506 ( .A1(n18767), .A2(n18824), .B1(n18821), .B2(n18448), .ZN(
        n18428) );
  AND2_X1 U21507 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18741), .ZN(n18822) );
  NAND2_X1 U21508 ( .A1(n18450), .A2(n18426), .ZN(n18779) );
  INV_X1 U21509 ( .A(n18779), .ZN(n18823) );
  AOI22_X1 U21510 ( .A1(n18858), .A2(n18822), .B1(n18823), .B2(n18515), .ZN(
        n18427) );
  OAI211_X1 U21511 ( .C1(n18429), .C2(n18453), .A(n18428), .B(n18427), .ZN(
        P3_U2871) );
  NOR2_X2 U21512 ( .A1(n18797), .A2(n19539), .ZN(n18831) );
  NOR2_X2 U21513 ( .A1(n18565), .A2(n18430), .ZN(n18828) );
  AOI22_X1 U21514 ( .A1(n18767), .A2(n18831), .B1(n18828), .B2(n18448), .ZN(
        n18434) );
  NOR2_X2 U21515 ( .A1(n18431), .A2(n18797), .ZN(n18829) );
  NAND2_X1 U21516 ( .A1(n18450), .A2(n18432), .ZN(n18782) );
  INV_X1 U21517 ( .A(n18782), .ZN(n18830) );
  AOI22_X1 U21518 ( .A1(n18858), .A2(n18829), .B1(n18830), .B2(n18515), .ZN(
        n18433) );
  OAI211_X1 U21519 ( .C1(n18435), .C2(n18453), .A(n18434), .B(n18433), .ZN(
        P3_U2872) );
  NOR2_X2 U21520 ( .A1(n19546), .A2(n18797), .ZN(n18837) );
  NOR2_X2 U21521 ( .A1(n18565), .A2(n18436), .ZN(n18835) );
  AOI22_X1 U21522 ( .A1(n18858), .A2(n18837), .B1(n18835), .B2(n18448), .ZN(
        n18440) );
  NOR2_X2 U21523 ( .A1(n18797), .A2(n15192), .ZN(n18836) );
  NAND2_X1 U21524 ( .A1(n18450), .A2(n18437), .ZN(n18842) );
  INV_X1 U21525 ( .A(n18842), .ZN(n18438) );
  AOI22_X1 U21526 ( .A1(n18767), .A2(n18836), .B1(n18438), .B2(n18515), .ZN(
        n18439) );
  OAI211_X1 U21527 ( .C1(n18441), .C2(n18453), .A(n18440), .B(n18439), .ZN(
        P3_U2873) );
  AND2_X1 U21528 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18741), .ZN(n18847) );
  NOR2_X2 U21529 ( .A1(n18442), .A2(n18565), .ZN(n18843) );
  AOI22_X1 U21530 ( .A1(n18767), .A2(n18847), .B1(n18843), .B2(n18448), .ZN(
        n18445) );
  NOR2_X2 U21531 ( .A1(n19553), .A2(n18797), .ZN(n18844) );
  NAND2_X1 U21532 ( .A1(n18450), .A2(n18443), .ZN(n18787) );
  INV_X1 U21533 ( .A(n18787), .ZN(n18846) );
  AOI22_X1 U21534 ( .A1(n18858), .A2(n18844), .B1(n18846), .B2(n18515), .ZN(
        n18444) );
  OAI211_X1 U21535 ( .C1(n18446), .C2(n18453), .A(n18445), .B(n18444), .ZN(
        P3_U2874) );
  NOR2_X2 U21536 ( .A1(n18797), .A2(n19561), .ZN(n18853) );
  NOR2_X2 U21537 ( .A1(n18447), .A2(n18565), .ZN(n18852) );
  AOI22_X1 U21538 ( .A1(n18858), .A2(n18853), .B1(n18852), .B2(n18448), .ZN(
        n18452) );
  AND2_X1 U21539 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18741), .ZN(n18857) );
  NAND2_X1 U21540 ( .A1(n18450), .A2(n18449), .ZN(n18793) );
  INV_X1 U21541 ( .A(n18793), .ZN(n18856) );
  AOI22_X1 U21542 ( .A1(n18767), .A2(n18857), .B1(n18856), .B2(n18515), .ZN(
        n18451) );
  OAI211_X1 U21543 ( .C1(n18454), .C2(n18453), .A(n18452), .B(n18451), .ZN(
        P3_U2875) );
  INV_X1 U21544 ( .A(n18496), .ZN(n18497) );
  NAND2_X1 U21545 ( .A1(n18643), .A2(n18497), .ZN(n18498) );
  NAND2_X1 U21546 ( .A1(n18898), .A2(n18926), .ZN(n18642) );
  NOR2_X1 U21547 ( .A1(n18496), .A2(n18642), .ZN(n18471) );
  AOI22_X1 U21548 ( .A1(n18800), .A2(n18471), .B1(n18801), .B2(n18855), .ZN(
        n18458) );
  INV_X1 U21549 ( .A(n18798), .ZN(n18456) );
  NAND2_X1 U21550 ( .A1(n18765), .A2(n18455), .ZN(n18795) );
  NOR2_X1 U21551 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18795), .ZN(
        n18544) );
  AOI22_X1 U21552 ( .A1(n18741), .A2(n18456), .B1(n18497), .B2(n18544), .ZN(
        n18472) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18472), .B1(
        n18767), .B2(n18803), .ZN(n18457) );
  OAI211_X1 U21554 ( .C1(n18770), .C2(n18498), .A(n18458), .B(n18457), .ZN(
        P3_U2876) );
  AOI22_X1 U21555 ( .A1(n18808), .A2(n18855), .B1(n18807), .B2(n18471), .ZN(
        n18460) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18472), .B1(
        n18767), .B2(n18810), .ZN(n18459) );
  OAI211_X1 U21557 ( .C1(n18773), .C2(n18498), .A(n18460), .B(n18459), .ZN(
        P3_U2877) );
  AOI22_X1 U21558 ( .A1(n18814), .A2(n18471), .B1(n18815), .B2(n18855), .ZN(
        n18462) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18472), .B1(
        n18767), .B2(n18817), .ZN(n18461) );
  OAI211_X1 U21560 ( .C1(n18776), .C2(n18498), .A(n18462), .B(n18461), .ZN(
        P3_U2878) );
  AOI22_X1 U21561 ( .A1(n18767), .A2(n18822), .B1(n18821), .B2(n18471), .ZN(
        n18464) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18472), .B1(
        n18824), .B2(n18845), .ZN(n18463) );
  OAI211_X1 U21563 ( .C1(n18779), .C2(n18498), .A(n18464), .B(n18463), .ZN(
        P3_U2879) );
  AOI22_X1 U21564 ( .A1(n18767), .A2(n18829), .B1(n18828), .B2(n18471), .ZN(
        n18466) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18472), .B1(
        n18831), .B2(n18845), .ZN(n18465) );
  OAI211_X1 U21566 ( .C1(n18782), .C2(n18498), .A(n18466), .B(n18465), .ZN(
        P3_U2880) );
  AOI22_X1 U21567 ( .A1(n18835), .A2(n18471), .B1(n18836), .B2(n18855), .ZN(
        n18468) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18472), .B1(
        n18767), .B2(n18837), .ZN(n18467) );
  OAI211_X1 U21569 ( .C1(n18842), .C2(n18498), .A(n18468), .B(n18467), .ZN(
        P3_U2881) );
  AOI22_X1 U21570 ( .A1(n18767), .A2(n18844), .B1(n18843), .B2(n18471), .ZN(
        n18470) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18472), .B1(
        n18847), .B2(n18845), .ZN(n18469) );
  OAI211_X1 U21572 ( .C1(n18787), .C2(n18498), .A(n18470), .B(n18469), .ZN(
        P3_U2882) );
  AOI22_X1 U21573 ( .A1(n18857), .A2(n18855), .B1(n18852), .B2(n18471), .ZN(
        n18474) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18472), .B1(
        n18767), .B2(n18853), .ZN(n18473) );
  OAI211_X1 U21575 ( .C1(n18793), .C2(n18498), .A(n18474), .B(n18473), .ZN(
        P3_U2883) );
  NAND2_X1 U21576 ( .A1(n18668), .A2(n18497), .ZN(n18495) );
  INV_X1 U21577 ( .A(n18926), .ZN(n18799) );
  AOI21_X1 U21578 ( .B1(n18498), .B2(n18495), .A(n18799), .ZN(n18491) );
  AOI22_X1 U21579 ( .A1(n18803), .A2(n18855), .B1(n18800), .B2(n18491), .ZN(
        n18478) );
  INV_X1 U21580 ( .A(n18495), .ZN(n18561) );
  AOI21_X1 U21581 ( .B1(n18498), .B2(n18495), .A(n18565), .ZN(n18520) );
  NOR2_X1 U21582 ( .A1(n18762), .A2(n18475), .ZN(n18476) );
  OAI22_X1 U21583 ( .A1(n18561), .A2(n19031), .B1(n18520), .B2(n18476), .ZN(
        n18492) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18492), .B1(
        n18801), .B2(n18515), .ZN(n18477) );
  OAI211_X1 U21585 ( .C1(n18770), .C2(n18495), .A(n18478), .B(n18477), .ZN(
        P3_U2884) );
  AOI22_X1 U21586 ( .A1(n18808), .A2(n18511), .B1(n18807), .B2(n18491), .ZN(
        n18480) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18492), .B1(
        n18810), .B2(n18855), .ZN(n18479) );
  OAI211_X1 U21588 ( .C1(n18773), .C2(n18495), .A(n18480), .B(n18479), .ZN(
        P3_U2885) );
  AOI22_X1 U21589 ( .A1(n18814), .A2(n18491), .B1(n18815), .B2(n18511), .ZN(
        n18482) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18492), .B1(
        n18817), .B2(n18855), .ZN(n18481) );
  OAI211_X1 U21591 ( .C1(n18776), .C2(n18495), .A(n18482), .B(n18481), .ZN(
        P3_U2886) );
  AOI22_X1 U21592 ( .A1(n18824), .A2(n18511), .B1(n18821), .B2(n18491), .ZN(
        n18484) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18492), .B1(
        n18822), .B2(n18855), .ZN(n18483) );
  OAI211_X1 U21594 ( .C1(n18779), .C2(n18495), .A(n18484), .B(n18483), .ZN(
        P3_U2887) );
  AOI22_X1 U21595 ( .A1(n18829), .A2(n18855), .B1(n18828), .B2(n18491), .ZN(
        n18486) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18492), .B1(
        n18831), .B2(n18511), .ZN(n18485) );
  OAI211_X1 U21597 ( .C1(n18782), .C2(n18495), .A(n18486), .B(n18485), .ZN(
        P3_U2888) );
  AOI22_X1 U21598 ( .A1(n18835), .A2(n18491), .B1(n18836), .B2(n18511), .ZN(
        n18488) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18492), .B1(
        n18837), .B2(n18845), .ZN(n18487) );
  OAI211_X1 U21600 ( .C1(n18842), .C2(n18495), .A(n18488), .B(n18487), .ZN(
        P3_U2889) );
  AOI22_X1 U21601 ( .A1(n18844), .A2(n18855), .B1(n18843), .B2(n18491), .ZN(
        n18490) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18492), .B1(
        n18847), .B2(n18511), .ZN(n18489) );
  OAI211_X1 U21603 ( .C1(n18787), .C2(n18495), .A(n18490), .B(n18489), .ZN(
        P3_U2890) );
  AOI22_X1 U21604 ( .A1(n18852), .A2(n18491), .B1(n18853), .B2(n18855), .ZN(
        n18494) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18492), .B1(
        n18857), .B2(n18515), .ZN(n18493) );
  OAI211_X1 U21606 ( .C1(n18793), .C2(n18495), .A(n18494), .B(n18493), .ZN(
        P3_U2891) );
  NOR2_X1 U21607 ( .A1(n18898), .A2(n18496), .ZN(n18545) );
  NAND2_X1 U21608 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18545), .ZN(
        n18519) );
  AND2_X1 U21609 ( .A1(n18926), .A2(n18545), .ZN(n18514) );
  AOI22_X1 U21610 ( .A1(n18803), .A2(n18511), .B1(n18800), .B2(n18514), .ZN(
        n18500) );
  AOI21_X1 U21611 ( .B1(n18898), .B2(n18762), .A(n18795), .ZN(n18591) );
  NAND2_X1 U21612 ( .A1(n18497), .A2(n18591), .ZN(n18516) );
  INV_X1 U21613 ( .A(n18498), .ZN(n18538) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18516), .B1(
        n18801), .B2(n18538), .ZN(n18499) );
  OAI211_X1 U21615 ( .C1(n18770), .C2(n18519), .A(n18500), .B(n18499), .ZN(
        P3_U2892) );
  AOI22_X1 U21616 ( .A1(n18810), .A2(n18511), .B1(n18807), .B2(n18514), .ZN(
        n18502) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18516), .B1(
        n18808), .B2(n18538), .ZN(n18501) );
  OAI211_X1 U21618 ( .C1(n18773), .C2(n18519), .A(n18502), .B(n18501), .ZN(
        P3_U2893) );
  AOI22_X1 U21619 ( .A1(n18814), .A2(n18514), .B1(n18815), .B2(n18538), .ZN(
        n18504) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18516), .B1(
        n18817), .B2(n18511), .ZN(n18503) );
  OAI211_X1 U21621 ( .C1(n18776), .C2(n18519), .A(n18504), .B(n18503), .ZN(
        P3_U2894) );
  AOI22_X1 U21622 ( .A1(n18821), .A2(n18514), .B1(n18822), .B2(n18511), .ZN(
        n18506) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18516), .B1(
        n18824), .B2(n18538), .ZN(n18505) );
  OAI211_X1 U21624 ( .C1(n18779), .C2(n18519), .A(n18506), .B(n18505), .ZN(
        P3_U2895) );
  AOI22_X1 U21625 ( .A1(n18831), .A2(n18538), .B1(n18828), .B2(n18514), .ZN(
        n18508) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18516), .B1(
        n18829), .B2(n18511), .ZN(n18507) );
  OAI211_X1 U21627 ( .C1(n18782), .C2(n18519), .A(n18508), .B(n18507), .ZN(
        P3_U2896) );
  AOI22_X1 U21628 ( .A1(n18835), .A2(n18514), .B1(n18836), .B2(n18538), .ZN(
        n18510) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18516), .B1(
        n18837), .B2(n18511), .ZN(n18509) );
  OAI211_X1 U21630 ( .C1(n18842), .C2(n18519), .A(n18510), .B(n18509), .ZN(
        P3_U2897) );
  AOI22_X1 U21631 ( .A1(n18844), .A2(n18511), .B1(n18843), .B2(n18514), .ZN(
        n18513) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18516), .B1(
        n18847), .B2(n18538), .ZN(n18512) );
  OAI211_X1 U21633 ( .C1(n18787), .C2(n18519), .A(n18513), .B(n18512), .ZN(
        P3_U2898) );
  AOI22_X1 U21634 ( .A1(n18857), .A2(n18538), .B1(n18852), .B2(n18514), .ZN(
        n18518) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18516), .B1(
        n18853), .B2(n18515), .ZN(n18517) );
  OAI211_X1 U21636 ( .C1(n18793), .C2(n18519), .A(n18518), .B(n18517), .ZN(
        P3_U2899) );
  INV_X1 U21637 ( .A(n18592), .ZN(n18543) );
  NOR2_X2 U21638 ( .A1(n18899), .A2(n18543), .ZN(n18607) );
  INV_X1 U21639 ( .A(n18607), .ZN(n18542) );
  NOR2_X1 U21640 ( .A1(n18582), .A2(n18607), .ZN(n18566) );
  NOR2_X1 U21641 ( .A1(n18799), .A2(n18566), .ZN(n18537) );
  AOI22_X1 U21642 ( .A1(n18800), .A2(n18537), .B1(n18801), .B2(n18561), .ZN(
        n18524) );
  INV_X1 U21643 ( .A(n18520), .ZN(n18521) );
  OAI22_X1 U21644 ( .A1(n18566), .A2(n18565), .B1(n18762), .B2(n18521), .ZN(
        n18522) );
  OAI21_X1 U21645 ( .B1(n18607), .B2(n19031), .A(n18522), .ZN(n18539) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18539), .B1(
        n18803), .B2(n18538), .ZN(n18523) );
  OAI211_X1 U21647 ( .C1(n18770), .C2(n18542), .A(n18524), .B(n18523), .ZN(
        P3_U2900) );
  AOI22_X1 U21648 ( .A1(n18808), .A2(n18561), .B1(n18807), .B2(n18537), .ZN(
        n18526) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18539), .B1(
        n18810), .B2(n18538), .ZN(n18525) );
  OAI211_X1 U21650 ( .C1(n18773), .C2(n18542), .A(n18526), .B(n18525), .ZN(
        P3_U2901) );
  AOI22_X1 U21651 ( .A1(n18817), .A2(n18538), .B1(n18814), .B2(n18537), .ZN(
        n18528) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18539), .B1(
        n18815), .B2(n18561), .ZN(n18527) );
  OAI211_X1 U21653 ( .C1(n18776), .C2(n18542), .A(n18528), .B(n18527), .ZN(
        P3_U2902) );
  AOI22_X1 U21654 ( .A1(n18824), .A2(n18561), .B1(n18821), .B2(n18537), .ZN(
        n18530) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18539), .B1(
        n18822), .B2(n18538), .ZN(n18529) );
  OAI211_X1 U21656 ( .C1(n18779), .C2(n18542), .A(n18530), .B(n18529), .ZN(
        P3_U2903) );
  AOI22_X1 U21657 ( .A1(n18831), .A2(n18561), .B1(n18828), .B2(n18537), .ZN(
        n18532) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18539), .B1(
        n18829), .B2(n18538), .ZN(n18531) );
  OAI211_X1 U21659 ( .C1(n18782), .C2(n18542), .A(n18532), .B(n18531), .ZN(
        P3_U2904) );
  AOI22_X1 U21660 ( .A1(n18837), .A2(n18538), .B1(n18835), .B2(n18537), .ZN(
        n18534) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18539), .B1(
        n18836), .B2(n18561), .ZN(n18533) );
  OAI211_X1 U21662 ( .C1(n18842), .C2(n18542), .A(n18534), .B(n18533), .ZN(
        P3_U2905) );
  AOI22_X1 U21663 ( .A1(n18847), .A2(n18561), .B1(n18843), .B2(n18537), .ZN(
        n18536) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18539), .B1(
        n18844), .B2(n18538), .ZN(n18535) );
  OAI211_X1 U21665 ( .C1(n18787), .C2(n18542), .A(n18536), .B(n18535), .ZN(
        P3_U2906) );
  AOI22_X1 U21666 ( .A1(n18857), .A2(n18561), .B1(n18852), .B2(n18537), .ZN(
        n18541) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18539), .B1(
        n18853), .B2(n18538), .ZN(n18540) );
  OAI211_X1 U21668 ( .C1(n18793), .C2(n18542), .A(n18541), .B(n18540), .ZN(
        P3_U2907) );
  NAND2_X1 U21669 ( .A1(n18643), .A2(n18592), .ZN(n18590) );
  NOR2_X1 U21670 ( .A1(n18543), .A2(n18642), .ZN(n18560) );
  AOI22_X1 U21671 ( .A1(n18800), .A2(n18560), .B1(n18801), .B2(n18582), .ZN(
        n18547) );
  AOI22_X1 U21672 ( .A1(n18741), .A2(n18545), .B1(n18592), .B2(n18544), .ZN(
        n18562) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18562), .B1(
        n18803), .B2(n18561), .ZN(n18546) );
  OAI211_X1 U21674 ( .C1(n18770), .C2(n18590), .A(n18547), .B(n18546), .ZN(
        P3_U2908) );
  AOI22_X1 U21675 ( .A1(n18808), .A2(n18582), .B1(n18807), .B2(n18560), .ZN(
        n18549) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18562), .B1(
        n18810), .B2(n18561), .ZN(n18548) );
  OAI211_X1 U21677 ( .C1(n18773), .C2(n18590), .A(n18549), .B(n18548), .ZN(
        P3_U2909) );
  AOI22_X1 U21678 ( .A1(n18814), .A2(n18560), .B1(n18815), .B2(n18582), .ZN(
        n18551) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18562), .B1(
        n18817), .B2(n18561), .ZN(n18550) );
  OAI211_X1 U21680 ( .C1(n18776), .C2(n18590), .A(n18551), .B(n18550), .ZN(
        P3_U2910) );
  AOI22_X1 U21681 ( .A1(n18821), .A2(n18560), .B1(n18822), .B2(n18561), .ZN(
        n18553) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18562), .B1(
        n18824), .B2(n18582), .ZN(n18552) );
  OAI211_X1 U21683 ( .C1(n18779), .C2(n18590), .A(n18553), .B(n18552), .ZN(
        P3_U2911) );
  AOI22_X1 U21684 ( .A1(n18829), .A2(n18561), .B1(n18828), .B2(n18560), .ZN(
        n18555) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18562), .B1(
        n18831), .B2(n18582), .ZN(n18554) );
  OAI211_X1 U21686 ( .C1(n18782), .C2(n18590), .A(n18555), .B(n18554), .ZN(
        P3_U2912) );
  AOI22_X1 U21687 ( .A1(n18835), .A2(n18560), .B1(n18836), .B2(n18582), .ZN(
        n18557) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18562), .B1(
        n18837), .B2(n18561), .ZN(n18556) );
  OAI211_X1 U21689 ( .C1(n18842), .C2(n18590), .A(n18557), .B(n18556), .ZN(
        P3_U2913) );
  AOI22_X1 U21690 ( .A1(n18844), .A2(n18561), .B1(n18843), .B2(n18560), .ZN(
        n18559) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18562), .B1(
        n18847), .B2(n18582), .ZN(n18558) );
  OAI211_X1 U21692 ( .C1(n18787), .C2(n18590), .A(n18559), .B(n18558), .ZN(
        P3_U2914) );
  AOI22_X1 U21693 ( .A1(n18857), .A2(n18582), .B1(n18852), .B2(n18560), .ZN(
        n18564) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18562), .B1(
        n18853), .B2(n18561), .ZN(n18563) );
  OAI211_X1 U21695 ( .C1(n18793), .C2(n18590), .A(n18564), .B(n18563), .ZN(
        P3_U2915) );
  NAND2_X1 U21696 ( .A1(n18668), .A2(n18592), .ZN(n18587) );
  AOI21_X1 U21697 ( .B1(n18590), .B2(n18587), .A(n18799), .ZN(n18583) );
  AOI22_X1 U21698 ( .A1(n18803), .A2(n18582), .B1(n18800), .B2(n18583), .ZN(
        n18569) );
  AOI21_X1 U21699 ( .B1(n18590), .B2(n18587), .A(n18565), .ZN(n18613) );
  NOR2_X1 U21700 ( .A1(n18566), .A2(n18797), .ZN(n18567) );
  OAI22_X1 U21701 ( .A1(n18663), .A2(n19031), .B1(n18613), .B2(n18567), .ZN(
        n18584) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18584), .B1(
        n18801), .B2(n18607), .ZN(n18568) );
  OAI211_X1 U21703 ( .C1(n18770), .C2(n18587), .A(n18569), .B(n18568), .ZN(
        P3_U2916) );
  AOI22_X1 U21704 ( .A1(n18808), .A2(n18607), .B1(n18807), .B2(n18583), .ZN(
        n18571) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18584), .B1(
        n18810), .B2(n18582), .ZN(n18570) );
  OAI211_X1 U21706 ( .C1(n18773), .C2(n18587), .A(n18571), .B(n18570), .ZN(
        P3_U2917) );
  AOI22_X1 U21707 ( .A1(n18814), .A2(n18583), .B1(n18815), .B2(n18607), .ZN(
        n18573) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18584), .B1(
        n18817), .B2(n18582), .ZN(n18572) );
  OAI211_X1 U21709 ( .C1(n18776), .C2(n18587), .A(n18573), .B(n18572), .ZN(
        P3_U2918) );
  AOI22_X1 U21710 ( .A1(n18824), .A2(n18607), .B1(n18821), .B2(n18583), .ZN(
        n18575) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18584), .B1(
        n18822), .B2(n18582), .ZN(n18574) );
  OAI211_X1 U21712 ( .C1(n18779), .C2(n18587), .A(n18575), .B(n18574), .ZN(
        P3_U2919) );
  AOI22_X1 U21713 ( .A1(n18829), .A2(n18582), .B1(n18828), .B2(n18583), .ZN(
        n18577) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18584), .B1(
        n18831), .B2(n18607), .ZN(n18576) );
  OAI211_X1 U21715 ( .C1(n18782), .C2(n18587), .A(n18577), .B(n18576), .ZN(
        P3_U2920) );
  AOI22_X1 U21716 ( .A1(n18837), .A2(n18582), .B1(n18835), .B2(n18583), .ZN(
        n18579) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18584), .B1(
        n18836), .B2(n18607), .ZN(n18578) );
  OAI211_X1 U21718 ( .C1(n18842), .C2(n18587), .A(n18579), .B(n18578), .ZN(
        P3_U2921) );
  AOI22_X1 U21719 ( .A1(n18847), .A2(n18607), .B1(n18843), .B2(n18583), .ZN(
        n18581) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18584), .B1(
        n18844), .B2(n18582), .ZN(n18580) );
  OAI211_X1 U21721 ( .C1(n18787), .C2(n18587), .A(n18581), .B(n18580), .ZN(
        P3_U2922) );
  AOI22_X1 U21722 ( .A1(n18852), .A2(n18583), .B1(n18853), .B2(n18582), .ZN(
        n18586) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18584), .B1(
        n18857), .B2(n18607), .ZN(n18585) );
  OAI211_X1 U21724 ( .C1(n18793), .C2(n18587), .A(n18586), .B(n18585), .ZN(
        P3_U2923) );
  NAND2_X1 U21725 ( .A1(n18589), .A2(n18588), .ZN(n18641) );
  NOR2_X2 U21726 ( .A1(n18897), .A2(n18641), .ZN(n18686) );
  INV_X1 U21727 ( .A(n18686), .ZN(n18612) );
  NOR2_X1 U21728 ( .A1(n18799), .A2(n18641), .ZN(n18608) );
  INV_X1 U21729 ( .A(n18590), .ZN(n18634) );
  AOI22_X1 U21730 ( .A1(n18800), .A2(n18608), .B1(n18801), .B2(n18634), .ZN(
        n18594) );
  NAND2_X1 U21731 ( .A1(n18592), .A2(n18591), .ZN(n18609) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18609), .B1(
        n18803), .B2(n18607), .ZN(n18593) );
  OAI211_X1 U21733 ( .C1(n18770), .C2(n18612), .A(n18594), .B(n18593), .ZN(
        P3_U2924) );
  AOI22_X1 U21734 ( .A1(n18808), .A2(n18634), .B1(n18807), .B2(n18608), .ZN(
        n18596) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18609), .B1(
        n18810), .B2(n18607), .ZN(n18595) );
  OAI211_X1 U21736 ( .C1(n18773), .C2(n18612), .A(n18596), .B(n18595), .ZN(
        P3_U2925) );
  AOI22_X1 U21737 ( .A1(n18817), .A2(n18607), .B1(n18814), .B2(n18608), .ZN(
        n18598) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18609), .B1(
        n18815), .B2(n18634), .ZN(n18597) );
  OAI211_X1 U21739 ( .C1(n18776), .C2(n18612), .A(n18598), .B(n18597), .ZN(
        P3_U2926) );
  AOI22_X1 U21740 ( .A1(n18821), .A2(n18608), .B1(n18822), .B2(n18607), .ZN(
        n18600) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18609), .B1(
        n18824), .B2(n18634), .ZN(n18599) );
  OAI211_X1 U21742 ( .C1(n18779), .C2(n18612), .A(n18600), .B(n18599), .ZN(
        P3_U2927) );
  AOI22_X1 U21743 ( .A1(n18829), .A2(n18607), .B1(n18828), .B2(n18608), .ZN(
        n18602) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18609), .B1(
        n18831), .B2(n18634), .ZN(n18601) );
  OAI211_X1 U21745 ( .C1(n18782), .C2(n18612), .A(n18602), .B(n18601), .ZN(
        P3_U2928) );
  AOI22_X1 U21746 ( .A1(n18835), .A2(n18608), .B1(n18836), .B2(n18634), .ZN(
        n18604) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18609), .B1(
        n18837), .B2(n18607), .ZN(n18603) );
  OAI211_X1 U21748 ( .C1(n18842), .C2(n18612), .A(n18604), .B(n18603), .ZN(
        P3_U2929) );
  AOI22_X1 U21749 ( .A1(n18847), .A2(n18634), .B1(n18843), .B2(n18608), .ZN(
        n18606) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18609), .B1(
        n18844), .B2(n18607), .ZN(n18605) );
  OAI211_X1 U21751 ( .C1(n18787), .C2(n18612), .A(n18606), .B(n18605), .ZN(
        P3_U2930) );
  AOI22_X1 U21752 ( .A1(n18852), .A2(n18608), .B1(n18853), .B2(n18607), .ZN(
        n18611) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18609), .B1(
        n18857), .B2(n18634), .ZN(n18610) );
  OAI211_X1 U21754 ( .C1(n18793), .C2(n18612), .A(n18611), .B(n18610), .ZN(
        P3_U2931) );
  INV_X1 U21755 ( .A(n18712), .ZN(n18692) );
  NOR2_X2 U21756 ( .A1(n18899), .A2(n18692), .ZN(n18708) );
  INV_X1 U21757 ( .A(n18708), .ZN(n18639) );
  NAND2_X1 U21758 ( .A1(n18612), .A2(n18639), .ZN(n18615) );
  AOI22_X1 U21759 ( .A1(n18765), .A2(n18615), .B1(n18713), .B2(n18613), .ZN(
        n18614) );
  AOI21_X1 U21760 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18639), .A(n18614), 
        .ZN(n18627) );
  INV_X1 U21761 ( .A(n18615), .ZN(n18670) );
  NOR2_X1 U21762 ( .A1(n18799), .A2(n18670), .ZN(n18635) );
  AOI22_X1 U21763 ( .A1(n18800), .A2(n18635), .B1(n18801), .B2(n18663), .ZN(
        n18617) );
  AOI22_X1 U21764 ( .A1(n18803), .A2(n18634), .B1(n18802), .B2(n18708), .ZN(
        n18616) );
  OAI211_X1 U21765 ( .C1(n18627), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2932) );
  AOI22_X1 U21766 ( .A1(n18810), .A2(n18634), .B1(n18807), .B2(n18635), .ZN(
        n18620) );
  INV_X1 U21767 ( .A(n18627), .ZN(n18636) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18636), .B1(
        n18808), .B2(n18663), .ZN(n18619) );
  OAI211_X1 U21769 ( .C1(n18773), .C2(n18639), .A(n18620), .B(n18619), .ZN(
        P3_U2933) );
  AOI22_X1 U21770 ( .A1(n18817), .A2(n18634), .B1(n18814), .B2(n18635), .ZN(
        n18622) );
  AOI22_X1 U21771 ( .A1(n18816), .A2(n18708), .B1(n18815), .B2(n18663), .ZN(
        n18621) );
  OAI211_X1 U21772 ( .C1(n18627), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        P3_U2934) );
  AOI22_X1 U21773 ( .A1(n18824), .A2(n18663), .B1(n18821), .B2(n18635), .ZN(
        n18625) );
  AOI22_X1 U21774 ( .A1(n18823), .A2(n18708), .B1(n18822), .B2(n18634), .ZN(
        n18624) );
  OAI211_X1 U21775 ( .C1(n18627), .C2(n18626), .A(n18625), .B(n18624), .ZN(
        P3_U2935) );
  AOI22_X1 U21776 ( .A1(n18829), .A2(n18634), .B1(n18828), .B2(n18635), .ZN(
        n18629) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18636), .B1(
        n18831), .B2(n18663), .ZN(n18628) );
  OAI211_X1 U21778 ( .C1(n18782), .C2(n18639), .A(n18629), .B(n18628), .ZN(
        P3_U2936) );
  AOI22_X1 U21779 ( .A1(n18837), .A2(n18634), .B1(n18835), .B2(n18635), .ZN(
        n18631) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18636), .B1(
        n18836), .B2(n18663), .ZN(n18630) );
  OAI211_X1 U21781 ( .C1(n18842), .C2(n18639), .A(n18631), .B(n18630), .ZN(
        P3_U2937) );
  AOI22_X1 U21782 ( .A1(n18844), .A2(n18634), .B1(n18843), .B2(n18635), .ZN(
        n18633) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18636), .B1(
        n18847), .B2(n18663), .ZN(n18632) );
  OAI211_X1 U21784 ( .C1(n18787), .C2(n18639), .A(n18633), .B(n18632), .ZN(
        P3_U2938) );
  AOI22_X1 U21785 ( .A1(n18852), .A2(n18635), .B1(n18853), .B2(n18634), .ZN(
        n18638) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18636), .B1(
        n18857), .B2(n18663), .ZN(n18637) );
  OAI211_X1 U21787 ( .C1(n18793), .C2(n18639), .A(n18638), .B(n18637), .ZN(
        P3_U2939) );
  NAND2_X1 U21788 ( .A1(n18712), .A2(n18898), .ZN(n18640) );
  OAI22_X1 U21789 ( .A1(n18797), .A2(n18641), .B1(n18795), .B2(n18640), .ZN(
        n18666) );
  NOR2_X1 U21790 ( .A1(n18692), .A2(n18642), .ZN(n18662) );
  AOI22_X1 U21791 ( .A1(n18800), .A2(n18662), .B1(n18801), .B2(n18686), .ZN(
        n18645) );
  NAND2_X1 U21792 ( .A1(n18712), .A2(n18643), .ZN(n18669) );
  AOI22_X1 U21793 ( .A1(n18803), .A2(n18663), .B1(n18802), .B2(n18733), .ZN(
        n18644) );
  OAI211_X1 U21794 ( .C1(n18646), .C2(n18666), .A(n18645), .B(n18644), .ZN(
        P3_U2940) );
  AOI22_X1 U21795 ( .A1(n18808), .A2(n18686), .B1(n18807), .B2(n18662), .ZN(
        n18648) );
  AOI22_X1 U21796 ( .A1(n18809), .A2(n18733), .B1(n18810), .B2(n18663), .ZN(
        n18647) );
  OAI211_X1 U21797 ( .C1(n18649), .C2(n18666), .A(n18648), .B(n18647), .ZN(
        P3_U2941) );
  AOI22_X1 U21798 ( .A1(n18814), .A2(n18662), .B1(n18815), .B2(n18686), .ZN(
        n18651) );
  INV_X1 U21799 ( .A(n18666), .ZN(n18659) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18659), .B1(
        n18817), .B2(n18663), .ZN(n18650) );
  OAI211_X1 U21801 ( .C1(n18776), .C2(n18669), .A(n18651), .B(n18650), .ZN(
        P3_U2942) );
  AOI22_X1 U21802 ( .A1(n18821), .A2(n18662), .B1(n18822), .B2(n18663), .ZN(
        n18653) );
  AOI22_X1 U21803 ( .A1(n18824), .A2(n18686), .B1(n18823), .B2(n18733), .ZN(
        n18652) );
  OAI211_X1 U21804 ( .C1(n18654), .C2(n18666), .A(n18653), .B(n18652), .ZN(
        P3_U2943) );
  AOI22_X1 U21805 ( .A1(n18829), .A2(n18663), .B1(n18828), .B2(n18662), .ZN(
        n18656) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18659), .B1(
        n18831), .B2(n18686), .ZN(n18655) );
  OAI211_X1 U21807 ( .C1(n18782), .C2(n18669), .A(n18656), .B(n18655), .ZN(
        P3_U2944) );
  AOI22_X1 U21808 ( .A1(n18837), .A2(n18663), .B1(n18835), .B2(n18662), .ZN(
        n18658) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18659), .B1(
        n18836), .B2(n18686), .ZN(n18657) );
  OAI211_X1 U21810 ( .C1(n18842), .C2(n18669), .A(n18658), .B(n18657), .ZN(
        P3_U2945) );
  AOI22_X1 U21811 ( .A1(n18844), .A2(n18663), .B1(n18843), .B2(n18662), .ZN(
        n18661) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18659), .B1(
        n18847), .B2(n18686), .ZN(n18660) );
  OAI211_X1 U21813 ( .C1(n18787), .C2(n18669), .A(n18661), .B(n18660), .ZN(
        P3_U2946) );
  AOI22_X1 U21814 ( .A1(n18857), .A2(n18686), .B1(n18852), .B2(n18662), .ZN(
        n18665) );
  AOI22_X1 U21815 ( .A1(n18856), .A2(n18733), .B1(n18853), .B2(n18663), .ZN(
        n18664) );
  OAI211_X1 U21816 ( .C1(n18667), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2947) );
  NAND2_X1 U21817 ( .A1(n18668), .A2(n18712), .ZN(n18691) );
  AOI21_X1 U21818 ( .B1(n18669), .B2(n18691), .A(n18799), .ZN(n18687) );
  AOI22_X1 U21819 ( .A1(n18800), .A2(n18687), .B1(n18801), .B2(n18708), .ZN(
        n18673) );
  OAI211_X1 U21820 ( .C1(n18670), .C2(n18762), .A(n18669), .B(n18691), .ZN(
        n18671) );
  OAI211_X1 U21821 ( .C1(n18757), .C2(n19031), .A(n18765), .B(n18671), .ZN(
        n18688) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18688), .B1(
        n18803), .B2(n18686), .ZN(n18672) );
  OAI211_X1 U21823 ( .C1(n18770), .C2(n18691), .A(n18673), .B(n18672), .ZN(
        P3_U2948) );
  AOI22_X1 U21824 ( .A1(n18808), .A2(n18708), .B1(n18807), .B2(n18687), .ZN(
        n18675) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18688), .B1(
        n18810), .B2(n18686), .ZN(n18674) );
  OAI211_X1 U21826 ( .C1(n18773), .C2(n18691), .A(n18675), .B(n18674), .ZN(
        P3_U2949) );
  AOI22_X1 U21827 ( .A1(n18817), .A2(n18686), .B1(n18814), .B2(n18687), .ZN(
        n18677) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18688), .B1(
        n18815), .B2(n18708), .ZN(n18676) );
  OAI211_X1 U21829 ( .C1(n18776), .C2(n18691), .A(n18677), .B(n18676), .ZN(
        P3_U2950) );
  AOI22_X1 U21830 ( .A1(n18824), .A2(n18708), .B1(n18821), .B2(n18687), .ZN(
        n18679) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18688), .B1(
        n18822), .B2(n18686), .ZN(n18678) );
  OAI211_X1 U21832 ( .C1(n18779), .C2(n18691), .A(n18679), .B(n18678), .ZN(
        P3_U2951) );
  AOI22_X1 U21833 ( .A1(n18831), .A2(n18708), .B1(n18828), .B2(n18687), .ZN(
        n18681) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18688), .B1(
        n18829), .B2(n18686), .ZN(n18680) );
  OAI211_X1 U21835 ( .C1(n18782), .C2(n18691), .A(n18681), .B(n18680), .ZN(
        P3_U2952) );
  AOI22_X1 U21836 ( .A1(n18837), .A2(n18686), .B1(n18835), .B2(n18687), .ZN(
        n18683) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18688), .B1(
        n18836), .B2(n18708), .ZN(n18682) );
  OAI211_X1 U21838 ( .C1(n18842), .C2(n18691), .A(n18683), .B(n18682), .ZN(
        P3_U2953) );
  AOI22_X1 U21839 ( .A1(n18847), .A2(n18708), .B1(n18843), .B2(n18687), .ZN(
        n18685) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18688), .B1(
        n18844), .B2(n18686), .ZN(n18684) );
  OAI211_X1 U21841 ( .C1(n18787), .C2(n18691), .A(n18685), .B(n18684), .ZN(
        P3_U2954) );
  AOI22_X1 U21842 ( .A1(n18852), .A2(n18687), .B1(n18853), .B2(n18686), .ZN(
        n18690) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18688), .B1(
        n18857), .B2(n18708), .ZN(n18689) );
  OAI211_X1 U21844 ( .C1(n18793), .C2(n18691), .A(n18690), .B(n18689), .ZN(
        P3_U2955) );
  NOR2_X1 U21845 ( .A1(n18898), .A2(n18692), .ZN(n18740) );
  NAND2_X1 U21846 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18740), .ZN(
        n18714) );
  AND2_X1 U21847 ( .A1(n18926), .A2(n18740), .ZN(n18707) );
  AOI22_X1 U21848 ( .A1(n18800), .A2(n18707), .B1(n18801), .B2(n18733), .ZN(
        n18694) );
  INV_X1 U21849 ( .A(n18795), .ZN(n18738) );
  OAI211_X1 U21850 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18741), .A(
        n18738), .B(n18712), .ZN(n18709) );
  AOI22_X1 U21851 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18709), .B1(
        n18803), .B2(n18708), .ZN(n18693) );
  OAI211_X1 U21852 ( .C1(n18714), .C2(n18770), .A(n18694), .B(n18693), .ZN(
        P3_U2956) );
  AOI22_X1 U21853 ( .A1(n18810), .A2(n18708), .B1(n18807), .B2(n18707), .ZN(
        n18696) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18709), .B1(
        n18808), .B2(n18733), .ZN(n18695) );
  OAI211_X1 U21855 ( .C1(n18714), .C2(n18773), .A(n18696), .B(n18695), .ZN(
        P3_U2957) );
  AOI22_X1 U21856 ( .A1(n18814), .A2(n18707), .B1(n18815), .B2(n18733), .ZN(
        n18698) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18709), .B1(
        n18817), .B2(n18708), .ZN(n18697) );
  OAI211_X1 U21858 ( .C1(n18714), .C2(n18776), .A(n18698), .B(n18697), .ZN(
        P3_U2958) );
  AOI22_X1 U21859 ( .A1(n18824), .A2(n18733), .B1(n18821), .B2(n18707), .ZN(
        n18700) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18709), .B1(
        n18822), .B2(n18708), .ZN(n18699) );
  OAI211_X1 U21861 ( .C1(n18714), .C2(n18779), .A(n18700), .B(n18699), .ZN(
        P3_U2959) );
  AOI22_X1 U21862 ( .A1(n18831), .A2(n18733), .B1(n18828), .B2(n18707), .ZN(
        n18702) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18709), .B1(
        n18829), .B2(n18708), .ZN(n18701) );
  OAI211_X1 U21864 ( .C1(n18714), .C2(n18782), .A(n18702), .B(n18701), .ZN(
        P3_U2960) );
  AOI22_X1 U21865 ( .A1(n18837), .A2(n18708), .B1(n18835), .B2(n18707), .ZN(
        n18704) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18709), .B1(
        n18836), .B2(n18733), .ZN(n18703) );
  OAI211_X1 U21867 ( .C1(n18714), .C2(n18842), .A(n18704), .B(n18703), .ZN(
        P3_U2961) );
  AOI22_X1 U21868 ( .A1(n18844), .A2(n18708), .B1(n18843), .B2(n18707), .ZN(
        n18706) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18709), .B1(
        n18847), .B2(n18733), .ZN(n18705) );
  OAI211_X1 U21870 ( .C1(n18714), .C2(n18787), .A(n18706), .B(n18705), .ZN(
        P3_U2962) );
  AOI22_X1 U21871 ( .A1(n18857), .A2(n18733), .B1(n18852), .B2(n18707), .ZN(
        n18711) );
  AOI22_X1 U21872 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18709), .B1(
        n18853), .B2(n18708), .ZN(n18710) );
  OAI211_X1 U21873 ( .C1(n18714), .C2(n18793), .A(n18711), .B(n18710), .ZN(
        P3_U2963) );
  NOR2_X2 U21874 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18796), .ZN(
        n18854) );
  INV_X1 U21875 ( .A(n18854), .ZN(n18737) );
  NAND2_X1 U21876 ( .A1(n18713), .A2(n18712), .ZN(n18715) );
  INV_X1 U21877 ( .A(n18714), .ZN(n18789) );
  NOR2_X1 U21878 ( .A1(n18854), .A2(n18789), .ZN(n18764) );
  OAI21_X1 U21879 ( .B1(n18716), .B2(n18715), .A(n18764), .ZN(n18717) );
  OAI211_X1 U21880 ( .C1(n18854), .C2(n19031), .A(n18765), .B(n18717), .ZN(
        n18734) );
  NOR2_X1 U21881 ( .A1(n18799), .A2(n18764), .ZN(n18732) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18734), .B1(
        n18800), .B2(n18732), .ZN(n18719) );
  AOI22_X1 U21883 ( .A1(n18803), .A2(n18733), .B1(n18801), .B2(n18757), .ZN(
        n18718) );
  OAI211_X1 U21884 ( .C1(n18737), .C2(n18770), .A(n18719), .B(n18718), .ZN(
        P3_U2964) );
  AOI22_X1 U21885 ( .A1(n18810), .A2(n18733), .B1(n18807), .B2(n18732), .ZN(
        n18721) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18734), .B1(
        n18808), .B2(n18757), .ZN(n18720) );
  OAI211_X1 U21887 ( .C1(n18737), .C2(n18773), .A(n18721), .B(n18720), .ZN(
        P3_U2965) );
  AOI22_X1 U21888 ( .A1(n18814), .A2(n18732), .B1(n18815), .B2(n18757), .ZN(
        n18723) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18734), .B1(
        n18817), .B2(n18733), .ZN(n18722) );
  OAI211_X1 U21890 ( .C1(n18737), .C2(n18776), .A(n18723), .B(n18722), .ZN(
        P3_U2966) );
  AOI22_X1 U21891 ( .A1(n18821), .A2(n18732), .B1(n18822), .B2(n18733), .ZN(
        n18725) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18734), .B1(
        n18824), .B2(n18757), .ZN(n18724) );
  OAI211_X1 U21893 ( .C1(n18737), .C2(n18779), .A(n18725), .B(n18724), .ZN(
        P3_U2967) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18734), .B1(
        n18828), .B2(n18732), .ZN(n18727) );
  AOI22_X1 U21895 ( .A1(n18829), .A2(n18733), .B1(n18831), .B2(n18757), .ZN(
        n18726) );
  OAI211_X1 U21896 ( .C1(n18737), .C2(n18782), .A(n18727), .B(n18726), .ZN(
        P3_U2968) );
  AOI22_X1 U21897 ( .A1(n18835), .A2(n18732), .B1(n18836), .B2(n18757), .ZN(
        n18729) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18734), .B1(
        n18837), .B2(n18733), .ZN(n18728) );
  OAI211_X1 U21899 ( .C1(n18737), .C2(n18842), .A(n18729), .B(n18728), .ZN(
        P3_U2969) );
  AOI22_X1 U21900 ( .A1(n18844), .A2(n18733), .B1(n18843), .B2(n18732), .ZN(
        n18731) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18734), .B1(
        n18847), .B2(n18757), .ZN(n18730) );
  OAI211_X1 U21902 ( .C1(n18737), .C2(n18787), .A(n18731), .B(n18730), .ZN(
        P3_U2970) );
  AOI22_X1 U21903 ( .A1(n18857), .A2(n18757), .B1(n18852), .B2(n18732), .ZN(
        n18736) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18734), .B1(
        n18853), .B2(n18733), .ZN(n18735) );
  OAI211_X1 U21905 ( .C1(n18737), .C2(n18793), .A(n18736), .B(n18735), .ZN(
        P3_U2971) );
  NOR2_X1 U21906 ( .A1(n18799), .A2(n18796), .ZN(n18756) );
  AOI22_X1 U21907 ( .A1(n18789), .A2(n18801), .B1(n18800), .B2(n18756), .ZN(
        n18743) );
  AOI22_X1 U21908 ( .A1(n18741), .A2(n18740), .B1(n18739), .B2(n18738), .ZN(
        n18758) );
  AOI22_X1 U21909 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18758), .B1(
        n18803), .B2(n18757), .ZN(n18742) );
  OAI211_X1 U21910 ( .C1(n18763), .C2(n18770), .A(n18743), .B(n18742), .ZN(
        P3_U2972) );
  AOI22_X1 U21911 ( .A1(n18810), .A2(n18757), .B1(n18807), .B2(n18756), .ZN(
        n18745) );
  AOI22_X1 U21912 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18758), .B1(
        n18789), .B2(n18808), .ZN(n18744) );
  OAI211_X1 U21913 ( .C1(n18763), .C2(n18773), .A(n18745), .B(n18744), .ZN(
        P3_U2973) );
  AOI22_X1 U21914 ( .A1(n18789), .A2(n18815), .B1(n18814), .B2(n18756), .ZN(
        n18747) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18758), .B1(
        n18817), .B2(n18757), .ZN(n18746) );
  OAI211_X1 U21916 ( .C1(n18763), .C2(n18776), .A(n18747), .B(n18746), .ZN(
        P3_U2974) );
  AOI22_X1 U21917 ( .A1(n18789), .A2(n18824), .B1(n18821), .B2(n18756), .ZN(
        n18749) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18758), .B1(
        n18822), .B2(n18757), .ZN(n18748) );
  OAI211_X1 U21919 ( .C1(n18763), .C2(n18779), .A(n18749), .B(n18748), .ZN(
        P3_U2975) );
  AOI22_X1 U21920 ( .A1(n18829), .A2(n18757), .B1(n18828), .B2(n18756), .ZN(
        n18751) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18758), .B1(
        n18789), .B2(n18831), .ZN(n18750) );
  OAI211_X1 U21922 ( .C1(n18763), .C2(n18782), .A(n18751), .B(n18750), .ZN(
        P3_U2976) );
  AOI22_X1 U21923 ( .A1(n18789), .A2(n18836), .B1(n18835), .B2(n18756), .ZN(
        n18753) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18758), .B1(
        n18837), .B2(n18757), .ZN(n18752) );
  OAI211_X1 U21925 ( .C1(n18763), .C2(n18842), .A(n18753), .B(n18752), .ZN(
        P3_U2977) );
  AOI22_X1 U21926 ( .A1(n18844), .A2(n18757), .B1(n18843), .B2(n18756), .ZN(
        n18755) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18758), .B1(
        n18789), .B2(n18847), .ZN(n18754) );
  OAI211_X1 U21928 ( .C1(n18763), .C2(n18787), .A(n18755), .B(n18754), .ZN(
        P3_U2978) );
  AOI22_X1 U21929 ( .A1(n18789), .A2(n18857), .B1(n18852), .B2(n18756), .ZN(
        n18760) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18758), .B1(
        n18853), .B2(n18757), .ZN(n18759) );
  OAI211_X1 U21931 ( .C1(n18763), .C2(n18793), .A(n18760), .B(n18759), .ZN(
        P3_U2979) );
  NOR2_X1 U21932 ( .A1(n18799), .A2(n18761), .ZN(n18788) );
  AOI22_X1 U21933 ( .A1(n18854), .A2(n18801), .B1(n18800), .B2(n18788), .ZN(
        n18769) );
  AOI221_X1 U21934 ( .B1(n18764), .B2(n18763), .C1(n18762), .C2(n18763), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18766) );
  OAI21_X1 U21935 ( .B1(n18767), .B2(n18766), .A(n18765), .ZN(n18790) );
  AOI22_X1 U21936 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18790), .B1(
        n18789), .B2(n18803), .ZN(n18768) );
  OAI211_X1 U21937 ( .C1(n18794), .C2(n18770), .A(n18769), .B(n18768), .ZN(
        P3_U2980) );
  AOI22_X1 U21938 ( .A1(n18789), .A2(n18810), .B1(n18788), .B2(n18807), .ZN(
        n18772) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18790), .B1(
        n18854), .B2(n18808), .ZN(n18771) );
  OAI211_X1 U21940 ( .C1(n18794), .C2(n18773), .A(n18772), .B(n18771), .ZN(
        P3_U2981) );
  AOI22_X1 U21941 ( .A1(n18854), .A2(n18815), .B1(n18788), .B2(n18814), .ZN(
        n18775) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18790), .B1(
        n18789), .B2(n18817), .ZN(n18774) );
  OAI211_X1 U21943 ( .C1(n18794), .C2(n18776), .A(n18775), .B(n18774), .ZN(
        P3_U2982) );
  AOI22_X1 U21944 ( .A1(n18789), .A2(n18822), .B1(n18788), .B2(n18821), .ZN(
        n18778) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18790), .B1(
        n18854), .B2(n18824), .ZN(n18777) );
  OAI211_X1 U21946 ( .C1(n18794), .C2(n18779), .A(n18778), .B(n18777), .ZN(
        P3_U2983) );
  AOI22_X1 U21947 ( .A1(n18854), .A2(n18831), .B1(n18788), .B2(n18828), .ZN(
        n18781) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18790), .B1(
        n18789), .B2(n18829), .ZN(n18780) );
  OAI211_X1 U21949 ( .C1(n18794), .C2(n18782), .A(n18781), .B(n18780), .ZN(
        P3_U2984) );
  AOI22_X1 U21950 ( .A1(n18854), .A2(n18836), .B1(n18788), .B2(n18835), .ZN(
        n18784) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18790), .B1(
        n18789), .B2(n18837), .ZN(n18783) );
  OAI211_X1 U21952 ( .C1(n18794), .C2(n18842), .A(n18784), .B(n18783), .ZN(
        P3_U2985) );
  AOI22_X1 U21953 ( .A1(n18789), .A2(n18844), .B1(n18788), .B2(n18843), .ZN(
        n18786) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18790), .B1(
        n18854), .B2(n18847), .ZN(n18785) );
  OAI211_X1 U21955 ( .C1(n18794), .C2(n18787), .A(n18786), .B(n18785), .ZN(
        P3_U2986) );
  AOI22_X1 U21956 ( .A1(n18789), .A2(n18853), .B1(n18788), .B2(n18852), .ZN(
        n18792) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18790), .B1(
        n18854), .B2(n18857), .ZN(n18791) );
  OAI211_X1 U21958 ( .C1(n18794), .C2(n18793), .A(n18792), .B(n18791), .ZN(
        P3_U2987) );
  OAI22_X1 U21959 ( .A1(n18797), .A2(n18796), .B1(n18798), .B2(n18795), .ZN(
        n18861) );
  NOR2_X1 U21960 ( .A1(n18799), .A2(n18798), .ZN(n18851) );
  AOI22_X1 U21961 ( .A1(n18858), .A2(n18801), .B1(n18800), .B2(n18851), .ZN(
        n18805) );
  AOI22_X1 U21962 ( .A1(n18854), .A2(n18803), .B1(n18802), .B2(n18845), .ZN(
        n18804) );
  OAI211_X1 U21963 ( .C1(n18806), .C2(n18861), .A(n18805), .B(n18804), .ZN(
        P3_U2988) );
  AOI22_X1 U21964 ( .A1(n18858), .A2(n18808), .B1(n18807), .B2(n18851), .ZN(
        n18812) );
  AOI22_X1 U21965 ( .A1(n18854), .A2(n18810), .B1(n18809), .B2(n18845), .ZN(
        n18811) );
  OAI211_X1 U21966 ( .C1(n18813), .C2(n18861), .A(n18812), .B(n18811), .ZN(
        P3_U2989) );
  AOI22_X1 U21967 ( .A1(n18858), .A2(n18815), .B1(n18814), .B2(n18851), .ZN(
        n18819) );
  AOI22_X1 U21968 ( .A1(n18854), .A2(n18817), .B1(n18816), .B2(n18845), .ZN(
        n18818) );
  OAI211_X1 U21969 ( .C1(n18820), .C2(n18861), .A(n18819), .B(n18818), .ZN(
        P3_U2990) );
  AOI22_X1 U21970 ( .A1(n18854), .A2(n18822), .B1(n18821), .B2(n18851), .ZN(
        n18826) );
  AOI22_X1 U21971 ( .A1(n18858), .A2(n18824), .B1(n18823), .B2(n18845), .ZN(
        n18825) );
  OAI211_X1 U21972 ( .C1(n18827), .C2(n18861), .A(n18826), .B(n18825), .ZN(
        P3_U2991) );
  AOI22_X1 U21973 ( .A1(n18854), .A2(n18829), .B1(n18828), .B2(n18851), .ZN(
        n18833) );
  AOI22_X1 U21974 ( .A1(n18858), .A2(n18831), .B1(n18830), .B2(n18845), .ZN(
        n18832) );
  OAI211_X1 U21975 ( .C1(n18834), .C2(n18861), .A(n18833), .B(n18832), .ZN(
        P3_U2992) );
  AOI22_X1 U21976 ( .A1(n18858), .A2(n18836), .B1(n18835), .B2(n18851), .ZN(
        n18840) );
  INV_X1 U21977 ( .A(n18861), .ZN(n18838) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18838), .B1(
        n18854), .B2(n18837), .ZN(n18839) );
  OAI211_X1 U21979 ( .C1(n18842), .C2(n18841), .A(n18840), .B(n18839), .ZN(
        P3_U2993) );
  AOI22_X1 U21980 ( .A1(n18854), .A2(n18844), .B1(n18843), .B2(n18851), .ZN(
        n18849) );
  AOI22_X1 U21981 ( .A1(n18858), .A2(n18847), .B1(n18846), .B2(n18845), .ZN(
        n18848) );
  OAI211_X1 U21982 ( .C1(n18850), .C2(n18861), .A(n18849), .B(n18848), .ZN(
        P3_U2994) );
  AOI22_X1 U21983 ( .A1(n18854), .A2(n18853), .B1(n18852), .B2(n18851), .ZN(
        n18860) );
  AOI22_X1 U21984 ( .A1(n18858), .A2(n18857), .B1(n18856), .B2(n18855), .ZN(
        n18859) );
  OAI211_X1 U21985 ( .C1(n18862), .C2(n18861), .A(n18860), .B(n18859), .ZN(
        P3_U2995) );
  OAI22_X1 U21986 ( .A1(n18866), .A2(n18865), .B1(n18864), .B2(n18863), .ZN(
        n18867) );
  AOI221_X1 U21987 ( .B1(n18890), .B2(n18869), .C1(n18868), .C2(n18869), .A(
        n18867), .ZN(n19075) );
  AOI211_X1 U21988 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18901), .A(
        n18871), .B(n18870), .ZN(n18913) );
  INV_X1 U21989 ( .A(n18901), .ZN(n18891) );
  AOI21_X1 U21990 ( .B1(n18880), .B2(n18874), .A(n18878), .ZN(n18872) );
  NOR2_X1 U21991 ( .A1(n19037), .A2(n19036), .ZN(n18877) );
  INV_X1 U21992 ( .A(n18873), .ZN(n18875) );
  NOR2_X1 U21993 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18874), .ZN(
        n18895) );
  OAI22_X1 U21994 ( .A1(n18875), .A2(n10174), .B1(n18895), .B2(n18880), .ZN(
        n19033) );
  AOI21_X1 U21995 ( .B1(n19033), .B2(n18891), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18876) );
  AOI21_X1 U21996 ( .B1(n18891), .B2(n18877), .A(n18876), .ZN(n18910) );
  AOI21_X1 U21997 ( .B1(n19055), .B2(n18883), .A(n18878), .ZN(n18888) );
  NAND2_X1 U21998 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18879), .ZN(
        n18887) );
  OAI211_X1 U21999 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18881), .B(n18880), .ZN(
        n18886) );
  NOR2_X1 U22000 ( .A1(n18882), .A2(n13107), .ZN(n18884) );
  OAI211_X1 U22001 ( .C1(n18884), .C2(n18883), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n13184), .ZN(n18885) );
  OAI211_X1 U22002 ( .C1(n18888), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        n18889) );
  AOI21_X1 U22003 ( .B1(n18890), .B2(n19043), .A(n18889), .ZN(n19045) );
  AOI22_X1 U22004 ( .A1(n18901), .A2(n13184), .B1(n19045), .B2(n18891), .ZN(
        n18904) );
  OAI22_X1 U22005 ( .A1(n18896), .A2(n19048), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18895), .ZN(n19053) );
  OAI21_X1 U22006 ( .B1(n18901), .B2(n18900), .A(n18899), .ZN(n18902) );
  AOI222_X1 U22007 ( .A1(n18903), .A2(n18904), .B1(n18903), .B2(n18902), .C1(
        n18904), .C2(n18902), .ZN(n18906) );
  INV_X1 U22008 ( .A(n18904), .ZN(n18905) );
  OAI221_X1 U22009 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18906), .A(n18905), .ZN(
        n18909) );
  NOR2_X1 U22010 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18908) );
  INV_X1 U22011 ( .A(n18906), .ZN(n18907) );
  OAI21_X1 U22012 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18911), .ZN(n18912) );
  NOR2_X1 U22013 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19085), .ZN(n18924) );
  NOR2_X1 U22014 ( .A1(n18925), .A2(n18926), .ZN(n18918) );
  NAND2_X1 U22015 ( .A1(n18938), .A2(n19079), .ZN(n18930) );
  INV_X1 U22016 ( .A(n18930), .ZN(n18916) );
  AOI211_X1 U22017 ( .C1(n19056), .C2(n19087), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18916), .ZN(n18917) );
  AOI211_X1 U22018 ( .C1(n18920), .C2(n18919), .A(n18918), .B(n18917), .ZN(
        n18921) );
  OAI221_X1 U22019 ( .B1(n18923), .B2(n18927), .C1(n18923), .C2(n18922), .A(
        n18921), .ZN(P3_U2996) );
  NAND3_X1 U22020 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18924), .ZN(n18933) );
  INV_X1 U22021 ( .A(n18925), .ZN(n18928) );
  NAND3_X1 U22022 ( .A1(n18928), .A2(n18927), .A3(n18926), .ZN(n18929) );
  NAND4_X1 U22023 ( .A1(n18931), .A2(n18930), .A3(n18933), .A4(n18929), .ZN(
        P3_U2997) );
  OAI21_X1 U22024 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18932), .ZN(n18935) );
  INV_X1 U22025 ( .A(n18933), .ZN(n18934) );
  AOI21_X1 U22026 ( .B1(n18936), .B2(n18935), .A(n18934), .ZN(P3_U2998) );
  AND2_X1 U22027 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19024), .ZN(
        P3_U2999) );
  AND2_X1 U22028 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19024), .ZN(
        P3_U3000) );
  AND2_X1 U22029 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18937), .ZN(
        P3_U3001) );
  AND2_X1 U22030 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18937), .ZN(
        P3_U3002) );
  AND2_X1 U22031 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18937), .ZN(
        P3_U3003) );
  AND2_X1 U22032 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18937), .ZN(
        P3_U3004) );
  AND2_X1 U22033 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18937), .ZN(
        P3_U3005) );
  AND2_X1 U22034 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18937), .ZN(
        P3_U3006) );
  AND2_X1 U22035 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18937), .ZN(
        P3_U3007) );
  AND2_X1 U22036 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18937), .ZN(
        P3_U3008) );
  AND2_X1 U22037 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18937), .ZN(
        P3_U3009) );
  AND2_X1 U22038 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18937), .ZN(
        P3_U3010) );
  AND2_X1 U22039 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18937), .ZN(
        P3_U3011) );
  AND2_X1 U22040 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18937), .ZN(
        P3_U3012) );
  AND2_X1 U22041 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18937), .ZN(
        P3_U3013) );
  AND2_X1 U22042 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18937), .ZN(
        P3_U3014) );
  AND2_X1 U22043 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18937), .ZN(
        P3_U3015) );
  AND2_X1 U22044 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18937), .ZN(
        P3_U3016) );
  AND2_X1 U22045 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18937), .ZN(
        P3_U3017) );
  AND2_X1 U22046 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18937), .ZN(
        P3_U3018) );
  AND2_X1 U22047 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18937), .ZN(
        P3_U3019) );
  AND2_X1 U22048 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18937), .ZN(
        P3_U3020) );
  AND2_X1 U22049 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18937), .ZN(P3_U3021) );
  AND2_X1 U22050 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19024), .ZN(P3_U3022) );
  AND2_X1 U22051 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19024), .ZN(P3_U3023) );
  AND2_X1 U22052 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19024), .ZN(P3_U3024) );
  AND2_X1 U22053 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19024), .ZN(P3_U3025) );
  AND2_X1 U22054 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19024), .ZN(P3_U3026) );
  AND2_X1 U22055 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19024), .ZN(P3_U3027) );
  AND2_X1 U22056 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19024), .ZN(P3_U3028) );
  INV_X1 U22057 ( .A(HOLD), .ZN(n21329) );
  NOR2_X1 U22058 ( .A1(n18953), .A2(n21329), .ZN(n18948) );
  INV_X1 U22059 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18941) );
  AOI211_X1 U22060 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n18948), .B(
        n18941), .ZN(n18940) );
  NAND2_X1 U22061 ( .A1(n18938), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18946) );
  AND2_X1 U22062 ( .A1(n18946), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18952) );
  AOI21_X1 U22063 ( .B1(NA), .B2(n18939), .A(n18953), .ZN(n18945) );
  OAI22_X1 U22064 ( .A1(n19092), .A2(n18940), .B1(n18952), .B2(n18945), .ZN(
        P3_U3029) );
  NOR2_X1 U22065 ( .A1(n18948), .A2(n18941), .ZN(n18943) );
  AND2_X1 U22066 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n18942) );
  AOI22_X1 U22067 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18943), .B1(n18942), 
        .B2(n18953), .ZN(n18944) );
  NAND3_X1 U22068 ( .A1(n18944), .A2(n19082), .A3(n18946), .ZN(P3_U3030) );
  INV_X1 U22069 ( .A(n18945), .ZN(n18951) );
  OAI22_X1 U22070 ( .A1(NA), .A2(n18946), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18947) );
  OAI22_X1 U22071 ( .A1(n18948), .A2(n18947), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18949) );
  OAI22_X1 U22072 ( .A1(n18952), .A2(n18951), .B1(n18950), .B2(n18949), .ZN(
        P3_U3031) );
  OAI222_X1 U22073 ( .A1(n19063), .A2(n19015), .B1(n18954), .B2(n19092), .C1(
        n18955), .C2(n19011), .ZN(P3_U3032) );
  OAI222_X1 U22074 ( .A1(n19011), .A2(n18957), .B1(n18956), .B2(n19092), .C1(
        n18955), .C2(n19015), .ZN(P3_U3033) );
  OAI222_X1 U22075 ( .A1(n19011), .A2(n18959), .B1(n18958), .B2(n19092), .C1(
        n18957), .C2(n19015), .ZN(P3_U3034) );
  OAI222_X1 U22076 ( .A1(n19011), .A2(n18962), .B1(n18960), .B2(n19092), .C1(
        n18959), .C2(n19015), .ZN(P3_U3035) );
  OAI222_X1 U22077 ( .A1(n18962), .A2(n19015), .B1(n18961), .B2(n19092), .C1(
        n18963), .C2(n19011), .ZN(P3_U3036) );
  OAI222_X1 U22078 ( .A1(n19011), .A2(n18965), .B1(n18964), .B2(n19092), .C1(
        n18963), .C2(n19015), .ZN(P3_U3037) );
  INV_X1 U22079 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18968) );
  OAI222_X1 U22080 ( .A1(n19011), .A2(n18968), .B1(n18966), .B2(n19092), .C1(
        n18965), .C2(n19015), .ZN(P3_U3038) );
  OAI222_X1 U22081 ( .A1(n18968), .A2(n19015), .B1(n18967), .B2(n19092), .C1(
        n18969), .C2(n19011), .ZN(P3_U3039) );
  OAI222_X1 U22082 ( .A1(n19011), .A2(n18971), .B1(n18970), .B2(n19092), .C1(
        n18969), .C2(n19015), .ZN(P3_U3040) );
  OAI222_X1 U22083 ( .A1(n19011), .A2(n18973), .B1(n18972), .B2(n19092), .C1(
        n18971), .C2(n19015), .ZN(P3_U3041) );
  INV_X1 U22084 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18975) );
  OAI222_X1 U22085 ( .A1(n19011), .A2(n18975), .B1(n18974), .B2(n19092), .C1(
        n18973), .C2(n19015), .ZN(P3_U3042) );
  OAI222_X1 U22086 ( .A1(n19011), .A2(n18977), .B1(n18976), .B2(n19092), .C1(
        n18975), .C2(n19015), .ZN(P3_U3043) );
  OAI222_X1 U22087 ( .A1(n19011), .A2(n18980), .B1(n18978), .B2(n19092), .C1(
        n18977), .C2(n19015), .ZN(P3_U3044) );
  OAI222_X1 U22088 ( .A1(n18980), .A2(n19015), .B1(n18979), .B2(n19092), .C1(
        n18981), .C2(n19011), .ZN(P3_U3045) );
  OAI222_X1 U22089 ( .A1(n19011), .A2(n18983), .B1(n18982), .B2(n19092), .C1(
        n18981), .C2(n19015), .ZN(P3_U3046) );
  OAI222_X1 U22090 ( .A1(n19011), .A2(n18986), .B1(n18984), .B2(n19092), .C1(
        n18983), .C2(n19015), .ZN(P3_U3047) );
  OAI222_X1 U22091 ( .A1(n18986), .A2(n19015), .B1(n18985), .B2(n19092), .C1(
        n18987), .C2(n19011), .ZN(P3_U3048) );
  OAI222_X1 U22092 ( .A1(n19011), .A2(n18989), .B1(n18988), .B2(n19092), .C1(
        n18987), .C2(n19015), .ZN(P3_U3049) );
  OAI222_X1 U22093 ( .A1(n19011), .A2(n18992), .B1(n18990), .B2(n19092), .C1(
        n18989), .C2(n19015), .ZN(P3_U3050) );
  OAI222_X1 U22094 ( .A1(n18992), .A2(n19015), .B1(n18991), .B2(n19092), .C1(
        n18993), .C2(n19011), .ZN(P3_U3051) );
  OAI222_X1 U22095 ( .A1(n19011), .A2(n18995), .B1(n18994), .B2(n19092), .C1(
        n18993), .C2(n19015), .ZN(P3_U3052) );
  OAI222_X1 U22096 ( .A1(n19011), .A2(n18998), .B1(n18996), .B2(n19092), .C1(
        n18995), .C2(n19015), .ZN(P3_U3053) );
  OAI222_X1 U22097 ( .A1(n18998), .A2(n19015), .B1(n18997), .B2(n19092), .C1(
        n18999), .C2(n19011), .ZN(P3_U3054) );
  INV_X1 U22098 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19001) );
  OAI222_X1 U22099 ( .A1(n19011), .A2(n19001), .B1(n19000), .B2(n19092), .C1(
        n18999), .C2(n19015), .ZN(P3_U3055) );
  OAI222_X1 U22100 ( .A1(n19011), .A2(n19003), .B1(n19002), .B2(n19092), .C1(
        n19001), .C2(n19015), .ZN(P3_U3056) );
  OAI222_X1 U22101 ( .A1(n19011), .A2(n19005), .B1(n19004), .B2(n19092), .C1(
        n19003), .C2(n19015), .ZN(P3_U3057) );
  OAI222_X1 U22102 ( .A1(n19011), .A2(n19008), .B1(n19006), .B2(n19092), .C1(
        n19005), .C2(n19015), .ZN(P3_U3058) );
  OAI222_X1 U22103 ( .A1(n19008), .A2(n19015), .B1(n19007), .B2(n19092), .C1(
        n19009), .C2(n19011), .ZN(P3_U3059) );
  OAI222_X1 U22104 ( .A1(n19011), .A2(n19014), .B1(n19010), .B2(n19092), .C1(
        n19009), .C2(n19015), .ZN(P3_U3060) );
  INV_X1 U22105 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19013) );
  OAI222_X1 U22106 ( .A1(n19015), .A2(n19014), .B1(n19013), .B2(n19092), .C1(
        n19012), .C2(n19011), .ZN(P3_U3061) );
  INV_X1 U22107 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19016) );
  AOI22_X1 U22108 ( .A1(n19092), .A2(n19017), .B1(n19016), .B2(n19093), .ZN(
        P3_U3274) );
  INV_X1 U22109 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19065) );
  INV_X1 U22110 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19018) );
  AOI22_X1 U22111 ( .A1(n19092), .A2(n19065), .B1(n19018), .B2(n19093), .ZN(
        P3_U3275) );
  INV_X1 U22112 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19019) );
  AOI22_X1 U22113 ( .A1(n19092), .A2(n19020), .B1(n19019), .B2(n19093), .ZN(
        P3_U3276) );
  INV_X1 U22114 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19071) );
  INV_X1 U22115 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19021) );
  AOI22_X1 U22116 ( .A1(n19092), .A2(n19071), .B1(n19021), .B2(n19093), .ZN(
        P3_U3277) );
  INV_X1 U22117 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19023) );
  INV_X1 U22118 ( .A(n19025), .ZN(n19022) );
  AOI21_X1 U22119 ( .B1(n19024), .B2(n19023), .A(n19022), .ZN(P3_U3280) );
  OAI21_X1 U22120 ( .B1(n19027), .B2(n19026), .A(n19025), .ZN(P3_U3281) );
  INV_X1 U22121 ( .A(n19028), .ZN(n19030) );
  OAI221_X1 U22122 ( .B1(n19031), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19031), 
        .C2(n19030), .A(n19029), .ZN(P3_U3282) );
  INV_X1 U22123 ( .A(n19032), .ZN(n19035) );
  NOR2_X1 U22124 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19095), .ZN(
        n19034) );
  AOI22_X1 U22125 ( .A1(n19056), .A2(n19035), .B1(n19034), .B2(n19033), .ZN(
        n19039) );
  AOI21_X1 U22126 ( .B1(n19058), .B2(n19036), .A(n19062), .ZN(n19038) );
  OAI22_X1 U22127 ( .A1(n19062), .A2(n19039), .B1(n19038), .B2(n19037), .ZN(
        P3_U3285) );
  AOI22_X1 U22128 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19041), .B2(n19040), .ZN(
        n19049) );
  NOR2_X1 U22129 ( .A1(n19042), .A2(n19059), .ZN(n19050) );
  INV_X1 U22130 ( .A(n19056), .ZN(n19044) );
  OAI22_X1 U22131 ( .A1(n19045), .A2(n19095), .B1(n19044), .B2(n19043), .ZN(
        n19046) );
  AOI21_X1 U22132 ( .B1(n19049), .B2(n19050), .A(n19046), .ZN(n19047) );
  AOI22_X1 U22133 ( .A1(n19062), .A2(n13184), .B1(n19047), .B2(n19060), .ZN(
        P3_U3288) );
  INV_X1 U22134 ( .A(n19048), .ZN(n19052) );
  INV_X1 U22135 ( .A(n19049), .ZN(n19051) );
  AOI222_X1 U22136 ( .A1(n19053), .A2(n19058), .B1(n19056), .B2(n19052), .C1(
        n19051), .C2(n19050), .ZN(n19054) );
  AOI22_X1 U22137 ( .A1(n19062), .A2(n19055), .B1(n19054), .B2(n19060), .ZN(
        P3_U3289) );
  AOI222_X1 U22138 ( .A1(n19059), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19058), 
        .B2(n19057), .C1(n13107), .C2(n19056), .ZN(n19061) );
  AOI22_X1 U22139 ( .A1(n19062), .A2(n13107), .B1(n19061), .B2(n19060), .ZN(
        P3_U3290) );
  AOI21_X1 U22140 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19064) );
  AOI22_X1 U22141 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19064), .B2(n19063), .ZN(n19066) );
  AOI22_X1 U22142 ( .A1(n19067), .A2(n19066), .B1(n19065), .B2(n19070), .ZN(
        P3_U3292) );
  NOR2_X1 U22143 ( .A1(n19070), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19068) );
  AOI22_X1 U22144 ( .A1(n19071), .A2(n19070), .B1(n19069), .B2(n19068), .ZN(
        P3_U3293) );
  INV_X1 U22145 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19072) );
  AOI22_X1 U22146 ( .A1(n19092), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19072), 
        .B2(n19093), .ZN(P3_U3294) );
  INV_X1 U22147 ( .A(n19073), .ZN(n19076) );
  NAND2_X1 U22148 ( .A1(n19076), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19074) );
  OAI21_X1 U22149 ( .B1(n19076), .B2(n19075), .A(n19074), .ZN(P3_U3295) );
  AOI22_X1 U22150 ( .A1(n19085), .A2(n19079), .B1(n19078), .B2(n19077), .ZN(
        n19080) );
  AND2_X1 U22151 ( .A1(n19097), .A2(n19080), .ZN(n19091) );
  INV_X1 U22152 ( .A(n19081), .ZN(n19096) );
  AOI21_X1 U22153 ( .B1(n19084), .B2(n19083), .A(n19082), .ZN(n19086) );
  OAI211_X1 U22154 ( .C1(n19096), .C2(n19086), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19085), .ZN(n19088) );
  AOI21_X1 U22155 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19088), .A(n19087), 
        .ZN(n19090) );
  NAND2_X1 U22156 ( .A1(n19091), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19089) );
  OAI21_X1 U22157 ( .B1(n19091), .B2(n19090), .A(n19089), .ZN(P3_U3296) );
  OAI22_X1 U22158 ( .A1(n19093), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19092), .ZN(n19094) );
  INV_X1 U22159 ( .A(n19094), .ZN(P3_U3297) );
  OAI21_X1 U22160 ( .B1(n19095), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19097), 
        .ZN(n19100) );
  OAI22_X1 U22161 ( .A1(n19100), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19097), 
        .B2(n19096), .ZN(n19098) );
  INV_X1 U22162 ( .A(n19098), .ZN(P3_U3298) );
  OAI21_X1 U22163 ( .B1(n19100), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19099), 
        .ZN(n19101) );
  INV_X1 U22164 ( .A(n19101), .ZN(P3_U3299) );
  INV_X1 U22165 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19102) );
  INV_X1 U22166 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20098) );
  NAND2_X1 U22167 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20098), .ZN(n20090) );
  AOI22_X1 U22168 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20090), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20083), .ZN(n20161) );
  OAI21_X1 U22169 ( .B1(n20083), .B2(n19102), .A(n20081), .ZN(P2_U2815) );
  INV_X1 U22170 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19104) );
  OAI22_X1 U22171 ( .A1(n20214), .A2(n19104), .B1(n20218), .B2(n19103), .ZN(
        P2_U2816) );
  AOI21_X1 U22172 ( .B1(n20083), .B2(n20098), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19105) );
  AOI22_X1 U22173 ( .A1(n20148), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19105), 
        .B2(n20230), .ZN(P2_U2817) );
  OAI21_X1 U22174 ( .B1(n20091), .B2(BS16), .A(n20161), .ZN(n20159) );
  OAI21_X1 U22175 ( .B1(n20161), .B2(n12714), .A(n20159), .ZN(P2_U2818) );
  NOR2_X1 U22176 ( .A1(n19107), .A2(n19106), .ZN(n20208) );
  INV_X1 U22177 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19109) );
  OAI21_X1 U22178 ( .B1(n20208), .B2(n19109), .A(n19108), .ZN(P2_U2819) );
  NOR4_X1 U22179 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19113) );
  NOR4_X1 U22180 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19112) );
  NOR4_X1 U22181 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19111) );
  NOR4_X1 U22182 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19110) );
  NAND4_X1 U22183 ( .A1(n19113), .A2(n19112), .A3(n19111), .A4(n19110), .ZN(
        n19119) );
  NOR4_X1 U22184 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19117) );
  AOI211_X1 U22185 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19116) );
  NOR4_X1 U22186 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19115) );
  NOR4_X1 U22187 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19114) );
  NAND4_X1 U22188 ( .A1(n19117), .A2(n19116), .A3(n19115), .A4(n19114), .ZN(
        n19118) );
  NOR2_X1 U22189 ( .A1(n19119), .A2(n19118), .ZN(n19126) );
  INV_X1 U22190 ( .A(n19126), .ZN(n19125) );
  NOR2_X1 U22191 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19125), .ZN(n19120) );
  INV_X1 U22192 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20157) );
  AOI22_X1 U22193 ( .A1(n19120), .A2(n19341), .B1(n19125), .B2(n20157), .ZN(
        P2_U2820) );
  OR3_X1 U22194 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19124) );
  INV_X1 U22195 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U22196 ( .A1(n19120), .A2(n19124), .B1(n19125), .B2(n20155), .ZN(
        P2_U2821) );
  INV_X1 U22197 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20160) );
  NAND2_X1 U22198 ( .A1(n19120), .A2(n20160), .ZN(n19123) );
  OAI21_X1 U22199 ( .B1(n19341), .B2(n20099), .A(n19126), .ZN(n19121) );
  OAI21_X1 U22200 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19126), .A(n19121), 
        .ZN(n19122) );
  OAI221_X1 U22201 ( .B1(n19123), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19123), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19122), .ZN(P2_U2822) );
  INV_X1 U22202 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20153) );
  OAI221_X1 U22203 ( .B1(n19126), .B2(n20153), .C1(n19125), .C2(n19124), .A(
        n19123), .ZN(P2_U2823) );
  INV_X1 U22204 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20128) );
  OAI22_X1 U22205 ( .A1(n19127), .A2(n19353), .B1(n20128), .B2(n19342), .ZN(
        n19131) );
  INV_X1 U22206 ( .A(n19128), .ZN(n19129) );
  OAI22_X1 U22207 ( .A1(n19129), .A2(n19328), .B1(n14130), .B2(n19343), .ZN(
        n19130) );
  AOI211_X1 U22208 ( .C1(n19132), .C2(n19333), .A(n19131), .B(n19130), .ZN(
        n19137) );
  OAI211_X1 U22209 ( .C1(n19135), .C2(n19134), .A(n19303), .B(n19133), .ZN(
        n19136) );
  OAI211_X1 U22210 ( .C1(n19349), .C2(n19138), .A(n19137), .B(n19136), .ZN(
        P2_U2834) );
  INV_X1 U22211 ( .A(n19143), .ZN(n19140) );
  AOI22_X1 U22212 ( .A1(n19335), .A2(n19140), .B1(n19346), .B2(n19139), .ZN(
        n19150) );
  INV_X1 U22213 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19141) );
  OAI22_X1 U22214 ( .A1(n19141), .A2(n19353), .B1(n20126), .B2(n19342), .ZN(
        n19147) );
  OAI21_X1 U22215 ( .B1(n19144), .B2(n19143), .A(n19142), .ZN(n19145) );
  OAI22_X1 U22216 ( .A1(n19343), .A2(n14129), .B1(n19358), .B2(n19145), .ZN(
        n19146) );
  AOI211_X1 U22217 ( .C1(n19148), .C2(n19290), .A(n19147), .B(n19146), .ZN(
        n19149) );
  OAI211_X1 U22218 ( .C1(n19151), .C2(n19340), .A(n19150), .B(n19149), .ZN(
        P2_U2835) );
  NAND2_X1 U22219 ( .A1(n9843), .A2(n19152), .ZN(n19153) );
  XOR2_X1 U22220 ( .A(n19154), .B(n19153), .Z(n19162) );
  AOI22_X1 U22221 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19324), .ZN(n19155) );
  OAI21_X1 U22222 ( .B1(n19156), .B2(n19328), .A(n19155), .ZN(n19157) );
  AOI211_X1 U22223 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19323), .A(n19310), 
        .B(n19157), .ZN(n19161) );
  AOI22_X1 U22224 ( .A1(n19159), .A2(n19290), .B1(n19158), .B2(n19333), .ZN(
        n19160) );
  OAI211_X1 U22225 ( .C1(n19339), .C2(n19162), .A(n19161), .B(n19160), .ZN(
        P2_U2836) );
  OAI21_X1 U22226 ( .B1(n20123), .B2(n19342), .A(n19294), .ZN(n19165) );
  OAI22_X1 U22227 ( .A1(n19163), .A2(n19328), .B1(n11175), .B2(n19343), .ZN(
        n19164) );
  AOI211_X1 U22228 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19324), .A(
        n19165), .B(n19164), .ZN(n19171) );
  NOR2_X1 U22229 ( .A1(n19315), .A2(n19166), .ZN(n19179) );
  XNOR2_X1 U22230 ( .A(n19179), .B(n19167), .ZN(n19168) );
  AOI22_X1 U22231 ( .A1(n19169), .A2(n19290), .B1(n19303), .B2(n19168), .ZN(
        n19170) );
  OAI211_X1 U22232 ( .C1(n19172), .C2(n19340), .A(n19171), .B(n19170), .ZN(
        P2_U2837) );
  AOI22_X1 U22233 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19324), .ZN(n19173) );
  OAI211_X1 U22234 ( .C1(n20121), .C2(n19342), .A(n19173), .B(n19294), .ZN(
        n19176) );
  OAI22_X1 U22235 ( .A1(n19352), .A2(n19180), .B1(n19174), .B2(n19328), .ZN(
        n19175) );
  AOI211_X1 U22236 ( .C1(n19177), .C2(n19290), .A(n19176), .B(n19175), .ZN(
        n19183) );
  INV_X1 U22237 ( .A(n19178), .ZN(n19181) );
  OAI211_X1 U22238 ( .C1(n19181), .C2(n19180), .A(n19303), .B(n19179), .ZN(
        n19182) );
  OAI211_X1 U22239 ( .C1(n19340), .C2(n19184), .A(n19183), .B(n19182), .ZN(
        P2_U2838) );
  OAI21_X1 U22240 ( .B1(n20119), .B2(n19342), .A(n19294), .ZN(n19188) );
  INV_X1 U22241 ( .A(n19185), .ZN(n19186) );
  OAI22_X1 U22242 ( .A1(n19186), .A2(n19328), .B1(n14145), .B2(n19343), .ZN(
        n19187) );
  AOI211_X1 U22243 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19324), .A(
        n19188), .B(n19187), .ZN(n19195) );
  NOR2_X1 U22244 ( .A1(n19315), .A2(n19189), .ZN(n19191) );
  XNOR2_X1 U22245 ( .A(n19191), .B(n19190), .ZN(n19192) );
  AOI22_X1 U22246 ( .A1(n19193), .A2(n19290), .B1(n19303), .B2(n19192), .ZN(
        n19194) );
  OAI211_X1 U22247 ( .C1(n19196), .C2(n19340), .A(n19195), .B(n19194), .ZN(
        P2_U2839) );
  NAND2_X1 U22248 ( .A1(n15010), .A2(n19197), .ZN(n19199) );
  XOR2_X1 U22249 ( .A(n19199), .B(n19198), .Z(n19207) );
  INV_X1 U22250 ( .A(n19200), .ZN(n19201) );
  AOI22_X1 U22251 ( .A1(n19201), .A2(n19346), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19324), .ZN(n19202) );
  OAI211_X1 U22252 ( .C1(n20117), .C2(n19342), .A(n19202), .B(n19294), .ZN(
        n19205) );
  OAI22_X1 U22253 ( .A1(n19203), .A2(n19349), .B1(n19372), .B2(n19340), .ZN(
        n19204) );
  AOI211_X1 U22254 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19325), .A(n19205), .B(
        n19204), .ZN(n19206) );
  OAI21_X1 U22255 ( .B1(n19207), .B2(n19339), .A(n19206), .ZN(P2_U2840) );
  AOI22_X1 U22256 ( .A1(n19208), .A2(n19346), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19325), .ZN(n19209) );
  OAI211_X1 U22257 ( .C1(n13965), .C2(n19342), .A(n19209), .B(n19294), .ZN(
        n19210) );
  AOI21_X1 U22258 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19324), .A(
        n19210), .ZN(n19216) );
  OR2_X1 U22259 ( .A1(n19315), .A2(n19211), .ZN(n19217) );
  XOR2_X1 U22260 ( .A(n19217), .B(n19212), .Z(n19213) );
  AOI22_X1 U22261 ( .A1(n19214), .A2(n19290), .B1(n19303), .B2(n19213), .ZN(
        n19215) );
  OAI211_X1 U22262 ( .C1(n19374), .C2(n19340), .A(n19216), .B(n19215), .ZN(
        P2_U2841) );
  AOI211_X1 U22263 ( .C1(n19226), .C2(n19218), .A(n19339), .B(n19217), .ZN(
        n19225) );
  NAND2_X1 U22264 ( .A1(n19219), .A2(n19346), .ZN(n19223) );
  AOI22_X1 U22265 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19324), .ZN(n19220) );
  OAI211_X1 U22266 ( .C1(n19342), .C2(n13957), .A(n19220), .B(n19294), .ZN(
        n19221) );
  INV_X1 U22267 ( .A(n19221), .ZN(n19222) );
  NAND2_X1 U22268 ( .A1(n19223), .A2(n19222), .ZN(n19224) );
  NOR2_X1 U22269 ( .A1(n19225), .A2(n19224), .ZN(n19228) );
  AOI22_X1 U22270 ( .A1(n19226), .A2(n19335), .B1(n19375), .B2(n19333), .ZN(
        n19227) );
  OAI211_X1 U22271 ( .C1(n19229), .C2(n19349), .A(n19228), .B(n19227), .ZN(
        P2_U2842) );
  AOI22_X1 U22272 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19324), .ZN(n19230) );
  OAI21_X1 U22273 ( .B1(n19231), .B2(n19328), .A(n19230), .ZN(n19232) );
  AOI211_X1 U22274 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19323), .A(n19310), 
        .B(n19232), .ZN(n19239) );
  NOR2_X1 U22275 ( .A1(n19315), .A2(n19233), .ZN(n19235) );
  XNOR2_X1 U22276 ( .A(n19235), .B(n19234), .ZN(n19236) );
  AOI22_X1 U22277 ( .A1(n19237), .A2(n19290), .B1(n19303), .B2(n19236), .ZN(
        n19238) );
  OAI211_X1 U22278 ( .C1(n19378), .C2(n19340), .A(n19239), .B(n19238), .ZN(
        P2_U2843) );
  AOI22_X1 U22279 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19324), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n19325), .ZN(n19240) );
  OAI21_X1 U22280 ( .B1(n19241), .B2(n19328), .A(n19240), .ZN(n19242) );
  AOI211_X1 U22281 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19323), .A(n19310), 
        .B(n19242), .ZN(n19249) );
  NOR2_X1 U22282 ( .A1(n19315), .A2(n19243), .ZN(n19245) );
  XNOR2_X1 U22283 ( .A(n19245), .B(n19244), .ZN(n19246) );
  AOI22_X1 U22284 ( .A1(n19247), .A2(n19290), .B1(n19303), .B2(n19246), .ZN(
        n19248) );
  OAI211_X1 U22285 ( .C1(n19383), .C2(n19340), .A(n19249), .B(n19248), .ZN(
        P2_U2845) );
  AOI22_X1 U22286 ( .A1(n19250), .A2(n19346), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19325), .ZN(n19251) );
  OAI21_X1 U22287 ( .B1(n19252), .B2(n19353), .A(n19251), .ZN(n19253) );
  AOI211_X1 U22288 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19323), .A(n19310), .B(
        n19253), .ZN(n19259) );
  NAND2_X1 U22289 ( .A1(n15010), .A2(n19254), .ZN(n19255) );
  XNOR2_X1 U22290 ( .A(n19256), .B(n19255), .ZN(n19257) );
  AOI22_X1 U22291 ( .A1(n19386), .A2(n19333), .B1(n19303), .B2(n19257), .ZN(
        n19258) );
  OAI211_X1 U22292 ( .C1(n19260), .C2(n19349), .A(n19259), .B(n19258), .ZN(
        P2_U2846) );
  INV_X1 U22293 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U22294 ( .A1(n19261), .A2(n19346), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19325), .ZN(n19262) );
  OAI211_X1 U22295 ( .C1(n20108), .C2(n19342), .A(n19262), .B(n19294), .ZN(
        n19263) );
  AOI21_X1 U22296 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19324), .A(
        n19263), .ZN(n19270) );
  NOR2_X1 U22297 ( .A1(n19315), .A2(n19264), .ZN(n19266) );
  XNOR2_X1 U22298 ( .A(n19266), .B(n19265), .ZN(n19268) );
  AOI22_X1 U22299 ( .A1(n19303), .A2(n19268), .B1(n19290), .B2(n19267), .ZN(
        n19269) );
  OAI211_X1 U22300 ( .C1(n19340), .C2(n19390), .A(n19270), .B(n19269), .ZN(
        P2_U2847) );
  AOI22_X1 U22301 ( .A1(n19271), .A2(n19346), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19325), .ZN(n19272) );
  OAI21_X1 U22302 ( .B1(n19273), .B2(n19353), .A(n19272), .ZN(n19274) );
  AOI211_X1 U22303 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n19323), .A(n19310), .B(
        n19274), .ZN(n19280) );
  NAND2_X1 U22304 ( .A1(n9843), .A2(n19275), .ZN(n19276) );
  XNOR2_X1 U22305 ( .A(n19277), .B(n19276), .ZN(n19278) );
  AOI22_X1 U22306 ( .A1(n19303), .A2(n19278), .B1(n19333), .B2(n19392), .ZN(
        n19279) );
  OAI211_X1 U22307 ( .C1(n19349), .C2(n19281), .A(n19280), .B(n19279), .ZN(
        P2_U2848) );
  NOR2_X1 U22308 ( .A1(n19315), .A2(n19282), .ZN(n19284) );
  XOR2_X1 U22309 ( .A(n19284), .B(n19283), .Z(n19293) );
  AOI22_X1 U22310 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19324), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n19325), .ZN(n19285) );
  OAI21_X1 U22311 ( .B1(n19286), .B2(n19328), .A(n19285), .ZN(n19287) );
  AOI211_X1 U22312 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19323), .A(n19310), .B(
        n19287), .ZN(n19292) );
  INV_X1 U22313 ( .A(n19288), .ZN(n19394) );
  AOI22_X1 U22314 ( .A1(n19333), .A2(n19394), .B1(n19290), .B2(n19289), .ZN(
        n19291) );
  OAI211_X1 U22315 ( .C1(n19339), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U2849) );
  OAI21_X1 U22316 ( .B1(n12476), .B2(n19342), .A(n19294), .ZN(n19298) );
  OAI22_X1 U22317 ( .A1(n19296), .A2(n19328), .B1(n19295), .B2(n19353), .ZN(
        n19297) );
  AOI211_X1 U22318 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19325), .A(n19298), .B(
        n19297), .ZN(n19305) );
  NAND2_X1 U22319 ( .A1(n9843), .A2(n19299), .ZN(n19300) );
  XNOR2_X1 U22320 ( .A(n19301), .B(n19300), .ZN(n19302) );
  AOI22_X1 U22321 ( .A1(n19303), .A2(n19302), .B1(n19333), .B2(n19397), .ZN(
        n19304) );
  OAI211_X1 U22322 ( .C1(n19349), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P2_U2850) );
  INV_X1 U22323 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19307) );
  OAI22_X1 U22324 ( .A1(n19308), .A2(n19328), .B1(n19353), .B2(n19307), .ZN(
        n19309) );
  AOI211_X1 U22325 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19323), .A(n19310), .B(
        n19309), .ZN(n19322) );
  AOI22_X1 U22326 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19325), .B1(n19333), .B2(
        n19404), .ZN(n19321) );
  OAI22_X1 U22327 ( .A1(n19405), .A2(n19312), .B1(n19311), .B2(n19349), .ZN(
        n19313) );
  INV_X1 U22328 ( .A(n19313), .ZN(n19320) );
  INV_X1 U22329 ( .A(n19499), .ZN(n19318) );
  NOR2_X1 U22330 ( .A1(n19315), .A2(n19314), .ZN(n19317) );
  AOI21_X1 U22331 ( .B1(n19318), .B2(n19317), .A(n19339), .ZN(n19316) );
  OAI21_X1 U22332 ( .B1(n19318), .B2(n19317), .A(n19316), .ZN(n19319) );
  NAND4_X1 U22333 ( .A1(n19322), .A2(n19321), .A3(n19320), .A4(n19319), .ZN(
        P2_U2851) );
  NAND2_X1 U22334 ( .A1(n19323), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19327) );
  AOI22_X1 U22335 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19325), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19324), .ZN(n19326) );
  OAI211_X1 U22336 ( .C1(n19329), .C2(n19328), .A(n19327), .B(n19326), .ZN(
        n19332) );
  NOR2_X1 U22337 ( .A1(n19330), .A2(n19349), .ZN(n19331) );
  AOI211_X1 U22338 ( .C1(n19333), .C2(n20188), .A(n19332), .B(n19331), .ZN(
        n19337) );
  AOI22_X1 U22339 ( .A1(n19335), .A2(n19334), .B1(n19356), .B2(n20184), .ZN(
        n19336) );
  OAI211_X1 U22340 ( .C1(n19339), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P2_U2854) );
  OAI22_X1 U22341 ( .A1(n19342), .A2(n19341), .B1(n19340), .B2(n19398), .ZN(
        n19345) );
  NOR2_X1 U22342 ( .A1(n19343), .A2(n12390), .ZN(n19344) );
  AOI211_X1 U22343 ( .C1(n19347), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        n19348) );
  OAI21_X1 U22344 ( .B1(n19350), .B2(n19349), .A(n19348), .ZN(n19355) );
  INV_X1 U22345 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19351) );
  AOI21_X1 U22346 ( .B1(n19353), .B2(n19352), .A(n19351), .ZN(n19354) );
  AOI211_X1 U22347 ( .C1(n19356), .C2(n19582), .A(n19355), .B(n19354), .ZN(
        n19357) );
  OAI21_X1 U22348 ( .B1(n19359), .B2(n19358), .A(n19357), .ZN(P2_U2855) );
  AOI22_X1 U22349 ( .A1(n19361), .A2(n19428), .B1(n19360), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19364) );
  AOI22_X1 U22350 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19362), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19427), .ZN(n19363) );
  NAND2_X1 U22351 ( .A1(n19364), .A2(n19363), .ZN(P2_U2888) );
  INV_X1 U22352 ( .A(n19367), .ZN(n19370) );
  INV_X1 U22353 ( .A(n19368), .ZN(n19369) );
  OAI222_X1 U22354 ( .A1(n12641), .A2(n19391), .B1(n19372), .B2(n19389), .C1(
        n19371), .C2(n19434), .ZN(P2_U2904) );
  INV_X1 U22355 ( .A(n19434), .ZN(n19384) );
  AOI22_X1 U22356 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19427), .B1(n19480), 
        .B2(n19384), .ZN(n19373) );
  OAI21_X1 U22357 ( .B1(n19389), .B2(n19374), .A(n19373), .ZN(P2_U2905) );
  INV_X1 U22358 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19448) );
  AOI22_X1 U22359 ( .A1(n19375), .A2(n19396), .B1(n19478), .B2(n19384), .ZN(
        n19376) );
  OAI21_X1 U22360 ( .B1(n19391), .B2(n19448), .A(n19376), .ZN(P2_U2906) );
  INV_X1 U22361 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19450) );
  OAI222_X1 U22362 ( .A1(n19450), .A2(n19391), .B1(n19378), .B2(n19389), .C1(
        n19434), .C2(n19377), .ZN(P2_U2907) );
  AOI22_X1 U22363 ( .A1(n19380), .A2(n19396), .B1(n19379), .B2(n19384), .ZN(
        n19381) );
  OAI21_X1 U22364 ( .B1(n19391), .B2(n19452), .A(n19381), .ZN(P2_U2908) );
  INV_X1 U22365 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19454) );
  OAI222_X1 U22366 ( .A1(n19454), .A2(n19391), .B1(n19383), .B2(n19389), .C1(
        n19434), .C2(n19382), .ZN(P2_U2909) );
  AOI22_X1 U22367 ( .A1(n19386), .A2(n19396), .B1(n19385), .B2(n19384), .ZN(
        n19387) );
  OAI21_X1 U22368 ( .B1(n19391), .B2(n19456), .A(n19387), .ZN(P2_U2910) );
  INV_X1 U22369 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19458) );
  OAI222_X1 U22370 ( .A1(n19458), .A2(n19391), .B1(n19390), .B2(n19389), .C1(
        n19434), .C2(n19388), .ZN(P2_U2911) );
  AOI22_X1 U22371 ( .A1(n19392), .A2(n19396), .B1(P2_EAX_REG_7__SCAN_IN), .B2(
        n19427), .ZN(n19393) );
  OAI21_X1 U22372 ( .B1(n19567), .B2(n19434), .A(n19393), .ZN(P2_U2912) );
  AOI22_X1 U22373 ( .A1(n19394), .A2(n19396), .B1(P2_EAX_REG_6__SCAN_IN), .B2(
        n19427), .ZN(n19395) );
  OAI21_X1 U22374 ( .B1(n19555), .B2(n19434), .A(n19395), .ZN(P2_U2913) );
  AOI22_X1 U22375 ( .A1(n19397), .A2(n19396), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19427), .ZN(n19403) );
  XOR2_X1 U22376 ( .A(n20179), .B(n20174), .Z(n19418) );
  XNOR2_X1 U22377 ( .A(n19667), .B(n20188), .ZN(n19423) );
  INV_X1 U22378 ( .A(n19398), .ZN(n19431) );
  NAND2_X1 U22379 ( .A1(n19582), .A2(n19431), .ZN(n19430) );
  NAND2_X1 U22380 ( .A1(n19423), .A2(n19430), .ZN(n19422) );
  OAI21_X1 U22381 ( .B1(n20188), .B2(n20184), .A(n19422), .ZN(n19417) );
  NAND2_X1 U22382 ( .A1(n19418), .A2(n19417), .ZN(n19416) );
  OAI21_X1 U22383 ( .B1(n20174), .B2(n20179), .A(n19416), .ZN(n19411) );
  XNOR2_X1 U22384 ( .A(n19583), .B(n20166), .ZN(n19412) );
  NAND2_X1 U22385 ( .A1(n19411), .A2(n19412), .ZN(n19410) );
  OAI21_X1 U22386 ( .B1(n20166), .B2(n20167), .A(n19410), .ZN(n19400) );
  NAND2_X1 U22387 ( .A1(n19400), .A2(n19399), .ZN(n19406) );
  INV_X1 U22388 ( .A(n19405), .ZN(n19401) );
  NAND3_X1 U22389 ( .A1(n19406), .A2(n19401), .A3(n19429), .ZN(n19402) );
  OAI211_X1 U22390 ( .C1(n19549), .C2(n19434), .A(n19403), .B(n19402), .ZN(
        P2_U2914) );
  AOI22_X1 U22391 ( .A1(n19428), .A2(n19404), .B1(n19427), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19409) );
  XNOR2_X1 U22392 ( .A(n19406), .B(n19405), .ZN(n19407) );
  NAND2_X1 U22393 ( .A1(n19407), .A2(n19429), .ZN(n19408) );
  OAI211_X1 U22394 ( .C1(n19542), .C2(n19434), .A(n19409), .B(n19408), .ZN(
        P2_U2915) );
  AOI22_X1 U22395 ( .A1(n19428), .A2(n20166), .B1(n19427), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19415) );
  OAI21_X1 U22396 ( .B1(n19412), .B2(n19411), .A(n19410), .ZN(n19413) );
  NAND2_X1 U22397 ( .A1(n19413), .A2(n19429), .ZN(n19414) );
  OAI211_X1 U22398 ( .C1(n19535), .C2(n19434), .A(n19415), .B(n19414), .ZN(
        P2_U2916) );
  AOI22_X1 U22399 ( .A1(n19428), .A2(n20179), .B1(n19427), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19421) );
  OAI21_X1 U22400 ( .B1(n19418), .B2(n19417), .A(n19416), .ZN(n19419) );
  NAND2_X1 U22401 ( .A1(n19419), .A2(n19429), .ZN(n19420) );
  OAI211_X1 U22402 ( .C1(n19531), .C2(n19434), .A(n19421), .B(n19420), .ZN(
        P2_U2917) );
  AOI22_X1 U22403 ( .A1(n19428), .A2(n20188), .B1(n19427), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19426) );
  OAI21_X1 U22404 ( .B1(n19423), .B2(n19430), .A(n19422), .ZN(n19424) );
  NAND2_X1 U22405 ( .A1(n19424), .A2(n19429), .ZN(n19425) );
  OAI211_X1 U22406 ( .C1(n19526), .C2(n19434), .A(n19426), .B(n19425), .ZN(
        P2_U2918) );
  AOI22_X1 U22407 ( .A1(n19428), .A2(n19431), .B1(n19427), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19433) );
  OAI211_X1 U22408 ( .C1(n19582), .C2(n19431), .A(n19430), .B(n19429), .ZN(
        n19432) );
  OAI211_X1 U22409 ( .C1(n19435), .C2(n19434), .A(n19433), .B(n19432), .ZN(
        P2_U2919) );
  NOR2_X1 U22410 ( .A1(n19443), .A2(n19436), .ZN(P2_U2920) );
  INV_X1 U22411 ( .A(n19437), .ZN(n19440) );
  AOI22_X1 U22412 ( .A1(n19440), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19474), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19438) );
  OAI21_X1 U22413 ( .B1(n19439), .B2(n19443), .A(n19438), .ZN(P2_U2921) );
  AOI22_X1 U22414 ( .A1(n19440), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19474), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19441) );
  OAI21_X1 U22415 ( .B1(n19443), .B2(n19442), .A(n19441), .ZN(P2_U2922) );
  AOI22_X1 U22416 ( .A1(n19474), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19444) );
  OAI21_X1 U22417 ( .B1(n12641), .B2(n19476), .A(n19444), .ZN(P2_U2936) );
  INV_X1 U22418 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19446) );
  AOI22_X1 U22419 ( .A1(n19474), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22420 ( .B1(n19446), .B2(n19476), .A(n19445), .ZN(P2_U2937) );
  AOI22_X1 U22421 ( .A1(n19474), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19447) );
  OAI21_X1 U22422 ( .B1(n19448), .B2(n19476), .A(n19447), .ZN(P2_U2938) );
  AOI22_X1 U22423 ( .A1(n19474), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19449) );
  OAI21_X1 U22424 ( .B1(n19450), .B2(n19476), .A(n19449), .ZN(P2_U2939) );
  AOI22_X1 U22425 ( .A1(n19474), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19451) );
  OAI21_X1 U22426 ( .B1(n19452), .B2(n19476), .A(n19451), .ZN(P2_U2940) );
  AOI22_X1 U22427 ( .A1(n19474), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19453) );
  OAI21_X1 U22428 ( .B1(n19454), .B2(n19476), .A(n19453), .ZN(P2_U2941) );
  AOI22_X1 U22429 ( .A1(n19474), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19455) );
  OAI21_X1 U22430 ( .B1(n19456), .B2(n19476), .A(n19455), .ZN(P2_U2942) );
  AOI22_X1 U22431 ( .A1(n19474), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19457) );
  OAI21_X1 U22432 ( .B1(n19458), .B2(n19476), .A(n19457), .ZN(P2_U2943) );
  INV_X1 U22433 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19460) );
  AOI22_X1 U22434 ( .A1(n19474), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19459) );
  OAI21_X1 U22435 ( .B1(n19460), .B2(n19476), .A(n19459), .ZN(P2_U2944) );
  INV_X1 U22436 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19462) );
  AOI22_X1 U22437 ( .A1(n19474), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19461) );
  OAI21_X1 U22438 ( .B1(n19462), .B2(n19476), .A(n19461), .ZN(P2_U2945) );
  INV_X1 U22439 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19464) );
  AOI22_X1 U22440 ( .A1(n19474), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19463) );
  OAI21_X1 U22441 ( .B1(n19464), .B2(n19476), .A(n19463), .ZN(P2_U2946) );
  INV_X1 U22442 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19466) );
  AOI22_X1 U22443 ( .A1(n19474), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19465) );
  OAI21_X1 U22444 ( .B1(n19466), .B2(n19476), .A(n19465), .ZN(P2_U2947) );
  INV_X1 U22445 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19468) );
  AOI22_X1 U22446 ( .A1(n19474), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19467) );
  OAI21_X1 U22447 ( .B1(n19468), .B2(n19476), .A(n19467), .ZN(P2_U2948) );
  INV_X1 U22448 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19470) );
  AOI22_X1 U22449 ( .A1(n19474), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19469) );
  OAI21_X1 U22450 ( .B1(n19470), .B2(n19476), .A(n19469), .ZN(P2_U2949) );
  INV_X1 U22451 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19472) );
  AOI22_X1 U22452 ( .A1(n19474), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19471) );
  OAI21_X1 U22453 ( .B1(n19472), .B2(n19476), .A(n19471), .ZN(P2_U2950) );
  INV_X1 U22454 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19477) );
  AOI22_X1 U22455 ( .A1(n19474), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19473), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19475) );
  OAI21_X1 U22456 ( .B1(n19477), .B2(n19476), .A(n19475), .ZN(P2_U2951) );
  AOI22_X1 U22457 ( .A1(n19487), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19479) );
  NAND2_X1 U22458 ( .A1(n19481), .A2(n19478), .ZN(n19484) );
  NAND2_X1 U22459 ( .A1(n19479), .A2(n19484), .ZN(P2_U2965) );
  AOI22_X1 U22460 ( .A1(n19487), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19482) );
  NAND2_X1 U22461 ( .A1(n19481), .A2(n19480), .ZN(n19488) );
  NAND2_X1 U22462 ( .A1(n19482), .A2(n19488), .ZN(P2_U2966) );
  AOI22_X1 U22463 ( .A1(n19487), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19483), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19485) );
  NAND2_X1 U22464 ( .A1(n19485), .A2(n19484), .ZN(P2_U2980) );
  AOI22_X1 U22465 ( .A1(n19487), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19489) );
  NAND2_X1 U22466 ( .A1(n19489), .A2(n19488), .ZN(P2_U2981) );
  AOI22_X1 U22467 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19490), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19310), .ZN(n19498) );
  INV_X1 U22468 ( .A(n19491), .ZN(n19492) );
  OAI22_X1 U22469 ( .A1(n19494), .A2(n19493), .B1(n19492), .B2(n19501), .ZN(
        n19495) );
  AOI21_X1 U22470 ( .B1(n19510), .B2(n19496), .A(n19495), .ZN(n19497) );
  OAI211_X1 U22471 ( .C1(n19503), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        P2_U3010) );
  INV_X1 U22472 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19513) );
  OAI22_X1 U22473 ( .A1(n19503), .A2(n19502), .B1(n19501), .B2(n19500), .ZN(
        n19508) );
  AND3_X1 U22474 ( .A1(n19506), .A2(n19505), .A3(n19504), .ZN(n19507) );
  AOI211_X1 U22475 ( .C1(n19510), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        n19512) );
  OAI211_X1 U22476 ( .C1(n19514), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3012) );
  NAND2_X1 U22477 ( .A1(n19573), .A2(n20190), .ZN(n19579) );
  NOR2_X1 U22478 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19579), .ZN(
        n19566) );
  AOI22_X1 U22479 ( .A1(n19946), .A2(n20066), .B1(n20016), .B2(n19566), .ZN(
        n19524) );
  AOI21_X1 U22480 ( .B1(n20059), .B2(n19604), .A(n12714), .ZN(n19515) );
  NOR2_X1 U22481 ( .A1(n19515), .A2(n19973), .ZN(n19519) );
  INV_X1 U22482 ( .A(n19516), .ZN(n19520) );
  AOI21_X1 U22483 ( .B1(n19520), .B2(n12466), .A(n20169), .ZN(n19517) );
  AOI21_X1 U22484 ( .B1(n19519), .B2(n20020), .A(n19517), .ZN(n19518) );
  OAI21_X1 U22485 ( .B1(n19518), .B2(n19566), .A(n19975), .ZN(n19569) );
  INV_X1 U22486 ( .A(n20020), .ZN(n20062) );
  OAI21_X1 U22487 ( .B1(n20062), .B2(n19566), .A(n19519), .ZN(n19522) );
  OAI21_X1 U22488 ( .B1(n19520), .B2(n19566), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19521) );
  NAND2_X1 U22489 ( .A1(n19522), .A2(n19521), .ZN(n19568) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19569), .B1(
        n13458), .B2(n19568), .ZN(n19523) );
  OAI211_X1 U22491 ( .C1(n19949), .C2(n19604), .A(n19524), .B(n19523), .ZN(
        P2_U3048) );
  AOI22_X1 U22492 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19559), .ZN(n20033) );
  OAI22_X2 U22493 ( .A1(n19525), .A2(n19560), .B1(n20439), .B2(n19562), .ZN(
        n20030) );
  NOR2_X2 U22494 ( .A1(n9839), .A2(n19564), .ZN(n20029) );
  AOI22_X1 U22495 ( .A1(n20030), .A2(n20066), .B1(n20029), .B2(n19566), .ZN(
        n19529) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19569), .B1(
        n19527), .B2(n19568), .ZN(n19528) );
  OAI211_X1 U22497 ( .C1(n20033), .C2(n19604), .A(n19529), .B(n19528), .ZN(
        P2_U3049) );
  OAI22_X2 U22498 ( .A1(n20445), .A2(n19562), .B1(n19530), .B2(n19560), .ZN(
        n20035) );
  AOI22_X1 U22499 ( .A1(n20035), .A2(n20066), .B1(n9818), .B2(n19566), .ZN(
        n19534) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19569), .B1(
        n19532), .B2(n19568), .ZN(n19533) );
  OAI211_X1 U22501 ( .C1(n20038), .C2(n19604), .A(n19534), .B(n19533), .ZN(
        P2_U3050) );
  AOI22_X1 U22502 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19559), .ZN(n20043) );
  NOR2_X2 U22503 ( .A1(n10014), .A2(n19564), .ZN(n20039) );
  AOI22_X1 U22504 ( .A1(n19988), .A2(n20066), .B1(n20039), .B2(n19566), .ZN(
        n19538) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19569), .B1(
        n19536), .B2(n19568), .ZN(n19537) );
  OAI211_X1 U22506 ( .C1(n19991), .C2(n19604), .A(n19538), .B(n19537), .ZN(
        P2_U3051) );
  AOI22_X1 U22507 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19559), .ZN(n19995) );
  NOR2_X2 U22508 ( .A1(n19541), .A2(n19564), .ZN(n20044) );
  AOI22_X1 U22509 ( .A1(n20045), .A2(n20066), .B1(n20044), .B2(n19566), .ZN(
        n19545) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19569), .B1(
        n19543), .B2(n19568), .ZN(n19544) );
  OAI211_X1 U22511 ( .C1(n20048), .C2(n19604), .A(n19545), .B(n19544), .ZN(
        P2_U3052) );
  AOI22_X1 U22512 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19558), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19559), .ZN(n20052) );
  AOI22_X1 U22513 ( .A1(n20049), .A2(n20066), .B1(n19548), .B2(n19566), .ZN(
        n19552) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19569), .B1(
        n19550), .B2(n19568), .ZN(n19551) );
  OAI211_X1 U22515 ( .C1(n20052), .C2(n19604), .A(n19552), .B(n19551), .ZN(
        P2_U3053) );
  OAI22_X2 U22516 ( .A1(n19553), .A2(n19560), .B1(n20470), .B2(n19562), .ZN(
        n20055) );
  NOR2_X2 U22517 ( .A1(n19554), .A2(n19564), .ZN(n20053) );
  AOI22_X1 U22518 ( .A1(n20055), .A2(n20066), .B1(n20053), .B2(n19566), .ZN(
        n19557) );
  NOR2_X2 U22519 ( .A1(n19555), .A2(n20019), .ZN(n20054) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19569), .B1(
        n20054), .B2(n19568), .ZN(n19556) );
  OAI211_X1 U22521 ( .C1(n20060), .C2(n19604), .A(n19557), .B(n19556), .ZN(
        P2_U3054) );
  AOI22_X1 U22522 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19559), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19558), .ZN(n20010) );
  NOR2_X2 U22523 ( .A1(n19565), .A2(n19564), .ZN(n20061) );
  AOI22_X1 U22524 ( .A1(n20005), .A2(n20066), .B1(n20061), .B2(n19566), .ZN(
        n19571) );
  NOR2_X2 U22525 ( .A1(n19567), .A2(n20019), .ZN(n20063) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19569), .B1(
        n20063), .B2(n19568), .ZN(n19570) );
  OAI211_X1 U22527 ( .C1(n20010), .C2(n19604), .A(n19571), .B(n19570), .ZN(
        P2_U3055) );
  INV_X1 U22528 ( .A(n20075), .ZN(n19576) );
  INV_X1 U22529 ( .A(n19572), .ZN(n19575) );
  INV_X1 U22530 ( .A(n19573), .ZN(n19635) );
  NOR2_X1 U22531 ( .A1(n19574), .A2(n19635), .ZN(n19599) );
  NOR3_X1 U22532 ( .A1(n19575), .A2(n19599), .A3(n20013), .ZN(n19578) );
  AOI211_X2 U22533 ( .C1(n19579), .C2(n20013), .A(n19576), .B(n19578), .ZN(
        n19600) );
  AOI22_X1 U22534 ( .A1(n19600), .A2(n13458), .B1(n20016), .B2(n19599), .ZN(
        n19586) );
  NAND2_X1 U22535 ( .A1(n19583), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19759) );
  INV_X1 U22536 ( .A(n19759), .ZN(n19577) );
  NAND2_X1 U22537 ( .A1(n19577), .A2(n19584), .ZN(n19580) );
  AOI21_X1 U22538 ( .B1(n19580), .B2(n19579), .A(n19578), .ZN(n19581) );
  OAI211_X1 U22539 ( .C1(n19599), .C2(n12466), .A(n19581), .B(n19975), .ZN(
        n19601) );
  NAND2_X1 U22540 ( .A1(n19584), .A2(n19763), .ZN(n19608) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n20025), .ZN(n19585) );
  OAI211_X1 U22542 ( .C1(n20028), .C2(n19604), .A(n19586), .B(n19585), .ZN(
        P2_U3056) );
  AOI22_X1 U22543 ( .A1(n19600), .A2(n19527), .B1(n20029), .B2(n19599), .ZN(
        n19588) );
  INV_X1 U22544 ( .A(n20033), .ZN(n19911) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n19911), .ZN(n19587) );
  OAI211_X1 U22546 ( .C1(n19914), .C2(n19604), .A(n19588), .B(n19587), .ZN(
        P2_U3057) );
  INV_X1 U22547 ( .A(n20035), .ZN(n19918) );
  AOI22_X1 U22548 ( .A1(n19600), .A2(n19532), .B1(n9818), .B2(n19599), .ZN(
        n19590) );
  INV_X1 U22549 ( .A(n20038), .ZN(n19915) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n19915), .ZN(n19589) );
  OAI211_X1 U22551 ( .C1(n19918), .C2(n19604), .A(n19590), .B(n19589), .ZN(
        P2_U3058) );
  AOI22_X1 U22552 ( .A1(n19600), .A2(n19536), .B1(n20039), .B2(n19599), .ZN(
        n19592) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n20040), .ZN(n19591) );
  OAI211_X1 U22554 ( .C1(n20043), .C2(n19604), .A(n19592), .B(n19591), .ZN(
        P2_U3059) );
  AOI22_X1 U22555 ( .A1(n19600), .A2(n19543), .B1(n20044), .B2(n19599), .ZN(
        n19594) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n19992), .ZN(n19593) );
  OAI211_X1 U22557 ( .C1(n19995), .C2(n19604), .A(n19594), .B(n19593), .ZN(
        P2_U3060) );
  AOI22_X1 U22558 ( .A1(n19600), .A2(n19550), .B1(n19548), .B2(n19599), .ZN(
        n19596) );
  INV_X1 U22559 ( .A(n20052), .ZN(n19923) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n19923), .ZN(n19595) );
  OAI211_X1 U22561 ( .C1(n19926), .C2(n19604), .A(n19596), .B(n19595), .ZN(
        P2_U3061) );
  INV_X1 U22562 ( .A(n20055), .ZN(n20002) );
  AOI22_X1 U22563 ( .A1(n19600), .A2(n20054), .B1(n20053), .B2(n19599), .ZN(
        n19598) );
  INV_X1 U22564 ( .A(n20060), .ZN(n19998) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n19998), .ZN(n19597) );
  OAI211_X1 U22566 ( .C1(n20002), .C2(n19604), .A(n19598), .B(n19597), .ZN(
        P2_U3062) );
  INV_X1 U22567 ( .A(n20005), .ZN(n20071) );
  AOI22_X1 U22568 ( .A1(n19600), .A2(n20063), .B1(n20061), .B2(n19599), .ZN(
        n19603) );
  INV_X1 U22569 ( .A(n20010), .ZN(n20065) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19601), .B1(
        n19630), .B2(n20065), .ZN(n19602) );
  OAI211_X1 U22571 ( .C1(n20071), .C2(n19604), .A(n19603), .B(n19602), .ZN(
        P2_U3063) );
  INV_X1 U22572 ( .A(n13805), .ZN(n19607) );
  NOR2_X1 U22573 ( .A1(n19836), .A2(n19635), .ZN(n19628) );
  OAI21_X1 U22574 ( .B1(n19607), .B2(n19628), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  NOR2_X1 U22575 ( .A1(n19839), .A2(n19635), .ZN(n19609) );
  INV_X1 U22576 ( .A(n19609), .ZN(n19605) );
  NAND2_X1 U22577 ( .A1(n19606), .A2(n19605), .ZN(n19629) );
  AOI22_X1 U22578 ( .A1(n19629), .A2(n13458), .B1(n20016), .B2(n19628), .ZN(
        n19615) );
  AOI21_X1 U22579 ( .B1(n19607), .B2(n12466), .A(n19628), .ZN(n19612) );
  AOI21_X1 U22580 ( .B1(n19666), .B2(n19608), .A(n12714), .ZN(n19610) );
  NOR2_X1 U22581 ( .A1(n19610), .A2(n19609), .ZN(n19611) );
  MUX2_X1 U22582 ( .A(n19612), .B(n19611), .S(n20169), .Z(n19613) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19946), .ZN(n19614) );
  OAI211_X1 U22584 ( .C1(n19949), .C2(n19666), .A(n19615), .B(n19614), .ZN(
        P2_U3064) );
  AOI22_X1 U22585 ( .A1(n19629), .A2(n19527), .B1(n20029), .B2(n19628), .ZN(
        n19617) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20030), .ZN(n19616) );
  OAI211_X1 U22587 ( .C1(n20033), .C2(n19666), .A(n19617), .B(n19616), .ZN(
        P2_U3065) );
  AOI22_X1 U22588 ( .A1(n19629), .A2(n19532), .B1(n9818), .B2(n19628), .ZN(
        n19619) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20035), .ZN(n19618) );
  OAI211_X1 U22590 ( .C1(n20038), .C2(n19666), .A(n19619), .B(n19618), .ZN(
        P2_U3066) );
  AOI22_X1 U22591 ( .A1(n19629), .A2(n19536), .B1(n20039), .B2(n19628), .ZN(
        n19621) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n19988), .ZN(n19620) );
  OAI211_X1 U22593 ( .C1(n19991), .C2(n19666), .A(n19621), .B(n19620), .ZN(
        P2_U3067) );
  AOI22_X1 U22594 ( .A1(n19629), .A2(n19543), .B1(n20044), .B2(n19628), .ZN(
        n19623) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20045), .ZN(n19622) );
  OAI211_X1 U22596 ( .C1(n20048), .C2(n19666), .A(n19623), .B(n19622), .ZN(
        P2_U3068) );
  AOI22_X1 U22597 ( .A1(n19629), .A2(n19550), .B1(n19548), .B2(n19628), .ZN(
        n19625) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20049), .ZN(n19624) );
  OAI211_X1 U22599 ( .C1(n20052), .C2(n19666), .A(n19625), .B(n19624), .ZN(
        P2_U3069) );
  AOI22_X1 U22600 ( .A1(n19629), .A2(n20054), .B1(n20053), .B2(n19628), .ZN(
        n19627) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20055), .ZN(n19626) );
  OAI211_X1 U22602 ( .C1(n20060), .C2(n19666), .A(n19627), .B(n19626), .ZN(
        P2_U3070) );
  AOI22_X1 U22603 ( .A1(n19629), .A2(n20063), .B1(n20061), .B2(n19628), .ZN(
        n19633) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19631), .B1(
        n19630), .B2(n20005), .ZN(n19632) );
  OAI211_X1 U22605 ( .C1(n20010), .C2(n19666), .A(n19633), .B(n19632), .ZN(
        P2_U3071) );
  NOR2_X1 U22606 ( .A1(n19865), .A2(n19635), .ZN(n19661) );
  AOI22_X1 U22607 ( .A1(n20025), .A2(n19693), .B1(n20016), .B2(n19661), .ZN(
        n19646) );
  INV_X1 U22608 ( .A(n20162), .ZN(n19634) );
  OAI21_X1 U22609 ( .B1(n19634), .B2(n19759), .A(n20169), .ZN(n19644) );
  NOR2_X1 U22610 ( .A1(n20190), .A2(n19635), .ZN(n19640) );
  INV_X1 U22611 ( .A(n19636), .ZN(n19641) );
  OAI21_X1 U22612 ( .B1(n19641), .B2(n20013), .A(n12466), .ZN(n19638) );
  INV_X1 U22613 ( .A(n19661), .ZN(n19637) );
  AOI21_X1 U22614 ( .B1(n19638), .B2(n19637), .A(n20019), .ZN(n19639) );
  OAI21_X1 U22615 ( .B1(n19644), .B2(n19640), .A(n19639), .ZN(n19663) );
  INV_X1 U22616 ( .A(n19640), .ZN(n19643) );
  OAI21_X1 U22617 ( .B1(n19641), .B2(n19661), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19642) );
  OAI21_X1 U22618 ( .B1(n19644), .B2(n19643), .A(n19642), .ZN(n19662) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19663), .B1(
        n13458), .B2(n19662), .ZN(n19645) );
  OAI211_X1 U22620 ( .C1(n20028), .C2(n19666), .A(n19646), .B(n19645), .ZN(
        P2_U3072) );
  AOI22_X1 U22621 ( .A1(n19911), .A2(n19693), .B1(n19661), .B2(n20029), .ZN(
        n19648) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19663), .B1(
        n19527), .B2(n19662), .ZN(n19647) );
  OAI211_X1 U22623 ( .C1(n19914), .C2(n19666), .A(n19648), .B(n19647), .ZN(
        P2_U3073) );
  AOI22_X1 U22624 ( .A1(n19915), .A2(n19693), .B1(n19661), .B2(n9818), .ZN(
        n19650) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19663), .B1(
        n19532), .B2(n19662), .ZN(n19649) );
  OAI211_X1 U22626 ( .C1(n19918), .C2(n19666), .A(n19650), .B(n19649), .ZN(
        P2_U3074) );
  AOI22_X1 U22627 ( .A1(n20040), .A2(n19693), .B1(n19661), .B2(n20039), .ZN(
        n19652) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19663), .B1(
        n19536), .B2(n19662), .ZN(n19651) );
  OAI211_X1 U22629 ( .C1(n20043), .C2(n19666), .A(n19652), .B(n19651), .ZN(
        P2_U3075) );
  INV_X1 U22630 ( .A(n19693), .ZN(n19660) );
  INV_X1 U22631 ( .A(n19666), .ZN(n19657) );
  AOI22_X1 U22632 ( .A1(n20045), .A2(n19657), .B1(n19661), .B2(n20044), .ZN(
        n19654) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19663), .B1(
        n19543), .B2(n19662), .ZN(n19653) );
  OAI211_X1 U22634 ( .C1(n20048), .C2(n19660), .A(n19654), .B(n19653), .ZN(
        P2_U3076) );
  AOI22_X1 U22635 ( .A1(n19923), .A2(n19693), .B1(n19661), .B2(n19548), .ZN(
        n19656) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19663), .B1(
        n19550), .B2(n19662), .ZN(n19655) );
  OAI211_X1 U22637 ( .C1(n19926), .C2(n19666), .A(n19656), .B(n19655), .ZN(
        P2_U3077) );
  AOI22_X1 U22638 ( .A1(n20055), .A2(n19657), .B1(n19661), .B2(n20053), .ZN(
        n19659) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19663), .B1(
        n20054), .B2(n19662), .ZN(n19658) );
  OAI211_X1 U22640 ( .C1(n20060), .C2(n19660), .A(n19659), .B(n19658), .ZN(
        P2_U3078) );
  AOI22_X1 U22641 ( .A1(n20065), .A2(n19693), .B1(n19661), .B2(n20061), .ZN(
        n19665) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19663), .B1(
        n20063), .B2(n19662), .ZN(n19664) );
  OAI211_X1 U22643 ( .C1(n20071), .C2(n19666), .A(n19665), .B(n19664), .ZN(
        P2_U3079) );
  INV_X1 U22644 ( .A(n19668), .ZN(n19670) );
  NOR2_X1 U22645 ( .A1(n19670), .A2(n19669), .ZN(n19907) );
  NAND2_X1 U22646 ( .A1(n19907), .A2(n10685), .ZN(n19675) );
  NAND3_X1 U22647 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n10685), .A3(
        n20190), .ZN(n19703) );
  NOR2_X1 U22648 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19703), .ZN(
        n19691) );
  OAI21_X1 U22649 ( .B1(n19672), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19671) );
  OAI21_X1 U22650 ( .B1(n19675), .B2(n19973), .A(n19671), .ZN(n19692) );
  AOI22_X1 U22651 ( .A1(n19692), .A2(n13458), .B1(n20016), .B2(n19691), .ZN(
        n19678) );
  OAI21_X1 U22652 ( .B1(n19693), .B2(n19717), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19674) );
  AOI211_X1 U22653 ( .C1(n19672), .C2(n12466), .A(n20169), .B(n19691), .ZN(
        n19673) );
  AOI211_X1 U22654 ( .C1(n19675), .C2(n19674), .A(n20019), .B(n19673), .ZN(
        n19676) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19946), .ZN(n19677) );
  OAI211_X1 U22656 ( .C1(n19949), .C2(n19724), .A(n19678), .B(n19677), .ZN(
        P2_U3080) );
  AOI22_X1 U22657 ( .A1(n19692), .A2(n19527), .B1(n20029), .B2(n19691), .ZN(
        n19680) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20030), .ZN(n19679) );
  OAI211_X1 U22659 ( .C1(n20033), .C2(n19724), .A(n19680), .B(n19679), .ZN(
        P2_U3081) );
  AOI22_X1 U22660 ( .A1(n19692), .A2(n19532), .B1(n9818), .B2(n19691), .ZN(
        n19682) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20035), .ZN(n19681) );
  OAI211_X1 U22662 ( .C1(n20038), .C2(n19724), .A(n19682), .B(n19681), .ZN(
        P2_U3082) );
  AOI22_X1 U22663 ( .A1(n19692), .A2(n19536), .B1(n20039), .B2(n19691), .ZN(
        n19684) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19988), .ZN(n19683) );
  OAI211_X1 U22665 ( .C1(n19991), .C2(n19724), .A(n19684), .B(n19683), .ZN(
        P2_U3083) );
  AOI22_X1 U22666 ( .A1(n19692), .A2(n19543), .B1(n20044), .B2(n19691), .ZN(
        n19686) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20045), .ZN(n19685) );
  OAI211_X1 U22668 ( .C1(n20048), .C2(n19724), .A(n19686), .B(n19685), .ZN(
        P2_U3084) );
  AOI22_X1 U22669 ( .A1(n19692), .A2(n19550), .B1(n19548), .B2(n19691), .ZN(
        n19688) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20049), .ZN(n19687) );
  OAI211_X1 U22671 ( .C1(n20052), .C2(n19724), .A(n19688), .B(n19687), .ZN(
        P2_U3085) );
  AOI22_X1 U22672 ( .A1(n19692), .A2(n20054), .B1(n20053), .B2(n19691), .ZN(
        n19690) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20055), .ZN(n19689) );
  OAI211_X1 U22674 ( .C1(n20060), .C2(n19724), .A(n19690), .B(n19689), .ZN(
        P2_U3086) );
  AOI22_X1 U22675 ( .A1(n19692), .A2(n20063), .B1(n20061), .B2(n19691), .ZN(
        n19696) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n20005), .ZN(n19695) );
  OAI211_X1 U22677 ( .C1(n20010), .C2(n19724), .A(n19696), .B(n19695), .ZN(
        P2_U3087) );
  NOR2_X1 U22678 ( .A1(n20199), .A2(n19703), .ZN(n19727) );
  AOI22_X1 U22679 ( .A1(n20025), .A2(n19747), .B1(n20016), .B2(n19727), .ZN(
        n19706) );
  OAI21_X1 U22680 ( .B1(n19759), .B2(n19935), .A(n20169), .ZN(n19704) );
  INV_X1 U22681 ( .A(n19703), .ZN(n19700) );
  INV_X1 U22682 ( .A(n19697), .ZN(n19701) );
  OAI21_X1 U22683 ( .B1(n19701), .B2(n20013), .A(n12466), .ZN(n19698) );
  INV_X1 U22684 ( .A(n19727), .ZN(n19732) );
  AOI21_X1 U22685 ( .B1(n19698), .B2(n19732), .A(n20019), .ZN(n19699) );
  OAI21_X1 U22686 ( .B1(n19704), .B2(n19700), .A(n19699), .ZN(n19721) );
  OAI21_X1 U22687 ( .B1(n19701), .B2(n19727), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19702) );
  OAI21_X1 U22688 ( .B1(n19704), .B2(n19703), .A(n19702), .ZN(n19720) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19721), .B1(
        n13458), .B2(n19720), .ZN(n19705) );
  OAI211_X1 U22690 ( .C1(n20028), .C2(n19724), .A(n19706), .B(n19705), .ZN(
        P2_U3088) );
  AOI22_X1 U22691 ( .A1(n19911), .A2(n19747), .B1(n20029), .B2(n19727), .ZN(
        n19708) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19721), .B1(
        n19527), .B2(n19720), .ZN(n19707) );
  OAI211_X1 U22693 ( .C1(n19914), .C2(n19724), .A(n19708), .B(n19707), .ZN(
        P2_U3089) );
  AOI22_X1 U22694 ( .A1(n20035), .A2(n19717), .B1(n9818), .B2(n19727), .ZN(
        n19710) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19721), .B1(
        n19532), .B2(n19720), .ZN(n19709) );
  OAI211_X1 U22696 ( .C1(n20038), .C2(n19755), .A(n19710), .B(n19709), .ZN(
        P2_U3090) );
  AOI22_X1 U22697 ( .A1(n19988), .A2(n19717), .B1(n20039), .B2(n19727), .ZN(
        n19712) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19721), .B1(
        n19536), .B2(n19720), .ZN(n19711) );
  OAI211_X1 U22699 ( .C1(n19991), .C2(n19755), .A(n19712), .B(n19711), .ZN(
        P2_U3091) );
  AOI22_X1 U22700 ( .A1(n19992), .A2(n19747), .B1(n20044), .B2(n19727), .ZN(
        n19714) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19721), .B1(
        n19543), .B2(n19720), .ZN(n19713) );
  OAI211_X1 U22702 ( .C1(n19995), .C2(n19724), .A(n19714), .B(n19713), .ZN(
        P2_U3092) );
  AOI22_X1 U22703 ( .A1(n19923), .A2(n19747), .B1(n19548), .B2(n19727), .ZN(
        n19716) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19721), .B1(
        n19550), .B2(n19720), .ZN(n19715) );
  OAI211_X1 U22705 ( .C1(n19926), .C2(n19724), .A(n19716), .B(n19715), .ZN(
        P2_U3093) );
  AOI22_X1 U22706 ( .A1(n20055), .A2(n19717), .B1(n20053), .B2(n19727), .ZN(
        n19719) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19721), .B1(
        n20054), .B2(n19720), .ZN(n19718) );
  OAI211_X1 U22708 ( .C1(n20060), .C2(n19755), .A(n19719), .B(n19718), .ZN(
        P2_U3094) );
  AOI22_X1 U22709 ( .A1(n20065), .A2(n19747), .B1(n20061), .B2(n19727), .ZN(
        n19723) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19721), .B1(
        n20063), .B2(n19720), .ZN(n19722) );
  OAI211_X1 U22711 ( .C1(n20071), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3095) );
  NOR2_X1 U22712 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20012), .ZN(
        n19762) );
  NAND2_X1 U22713 ( .A1(n20199), .A2(n19762), .ZN(n19730) );
  NAND3_X1 U22714 ( .A1(n19726), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19730), 
        .ZN(n19733) );
  INV_X1 U22715 ( .A(n19730), .ZN(n19750) );
  NOR2_X1 U22716 ( .A1(n19727), .A2(n19750), .ZN(n19728) );
  OAI21_X1 U22717 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19728), .A(n20013), 
        .ZN(n19729) );
  AOI22_X1 U22718 ( .A1(n19751), .A2(n13458), .B1(n20016), .B2(n19750), .ZN(
        n19736) );
  OAI21_X1 U22719 ( .B1(n19747), .B2(n19772), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19731) );
  OAI221_X1 U22720 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19732), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19731), .A(n19730), .ZN(n19734) );
  NAND3_X1 U22721 ( .A1(n19734), .A2(n19975), .A3(n19733), .ZN(n19752) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19752), .B1(
        n19747), .B2(n19946), .ZN(n19735) );
  OAI211_X1 U22723 ( .C1(n19949), .C2(n19783), .A(n19736), .B(n19735), .ZN(
        P2_U3096) );
  AOI22_X1 U22724 ( .A1(n19751), .A2(n19527), .B1(n20029), .B2(n19750), .ZN(
        n19738) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19752), .B1(
        n19747), .B2(n20030), .ZN(n19737) );
  OAI211_X1 U22726 ( .C1(n20033), .C2(n19783), .A(n19738), .B(n19737), .ZN(
        P2_U3097) );
  AOI22_X1 U22727 ( .A1(n19751), .A2(n19532), .B1(n9818), .B2(n19750), .ZN(
        n19740) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19752), .B1(
        n19772), .B2(n19915), .ZN(n19739) );
  OAI211_X1 U22729 ( .C1(n19918), .C2(n19755), .A(n19740), .B(n19739), .ZN(
        P2_U3098) );
  AOI22_X1 U22730 ( .A1(n19751), .A2(n19536), .B1(n20039), .B2(n19750), .ZN(
        n19742) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19752), .B1(
        n19772), .B2(n20040), .ZN(n19741) );
  OAI211_X1 U22732 ( .C1(n20043), .C2(n19755), .A(n19742), .B(n19741), .ZN(
        P2_U3099) );
  AOI22_X1 U22733 ( .A1(n19751), .A2(n19543), .B1(n20044), .B2(n19750), .ZN(
        n19744) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19752), .B1(
        n19772), .B2(n19992), .ZN(n19743) );
  OAI211_X1 U22735 ( .C1(n19995), .C2(n19755), .A(n19744), .B(n19743), .ZN(
        P2_U3100) );
  AOI22_X1 U22736 ( .A1(n19751), .A2(n19550), .B1(n19548), .B2(n19750), .ZN(
        n19746) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19752), .B1(
        n19772), .B2(n19923), .ZN(n19745) );
  OAI211_X1 U22738 ( .C1(n19926), .C2(n19755), .A(n19746), .B(n19745), .ZN(
        P2_U3101) );
  AOI22_X1 U22739 ( .A1(n19751), .A2(n20054), .B1(n20053), .B2(n19750), .ZN(
        n19749) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19752), .B1(
        n19747), .B2(n20055), .ZN(n19748) );
  OAI211_X1 U22741 ( .C1(n20060), .C2(n19783), .A(n19749), .B(n19748), .ZN(
        P2_U3102) );
  AOI22_X1 U22742 ( .A1(n19751), .A2(n20063), .B1(n20061), .B2(n19750), .ZN(
        n19754) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19752), .B1(
        n19772), .B2(n20065), .ZN(n19753) );
  OAI211_X1 U22744 ( .C1(n20071), .C2(n19755), .A(n19754), .B(n19753), .ZN(
        P2_U3103) );
  INV_X1 U22745 ( .A(n19762), .ZN(n19758) );
  INV_X1 U22746 ( .A(n19760), .ZN(n19756) );
  NOR2_X1 U22747 ( .A1(n20199), .A2(n19758), .ZN(n19791) );
  OAI21_X1 U22748 ( .B1(n19756), .B2(n19791), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19757) );
  OAI21_X1 U22749 ( .B1(n19758), .B2(n19973), .A(n19757), .ZN(n19779) );
  AOI22_X1 U22750 ( .A1(n19779), .A2(n13458), .B1(n20016), .B2(n19791), .ZN(
        n19765) );
  NOR2_X1 U22751 ( .A1(n19759), .A2(n19968), .ZN(n20170) );
  INV_X1 U22752 ( .A(n19791), .ZN(n19788) );
  OAI211_X1 U22753 ( .C1(n19760), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19973), 
        .B(n19788), .ZN(n19761) );
  OAI211_X1 U22754 ( .C1(n20170), .C2(n19762), .A(n19975), .B(n19761), .ZN(
        n19780) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n20025), .ZN(n19764) );
  OAI211_X1 U22756 ( .C1(n20028), .C2(n19783), .A(n19765), .B(n19764), .ZN(
        P2_U3104) );
  AOI22_X1 U22757 ( .A1(n19779), .A2(n19527), .B1(n20029), .B2(n19791), .ZN(
        n19767) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n19911), .ZN(n19766) );
  OAI211_X1 U22759 ( .C1(n19914), .C2(n19783), .A(n19767), .B(n19766), .ZN(
        P2_U3105) );
  AOI22_X1 U22760 ( .A1(n19779), .A2(n19532), .B1(n9818), .B2(n19791), .ZN(
        n19769) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n19915), .ZN(n19768) );
  OAI211_X1 U22762 ( .C1(n19918), .C2(n19783), .A(n19769), .B(n19768), .ZN(
        P2_U3106) );
  AOI22_X1 U22763 ( .A1(n19779), .A2(n19536), .B1(n20039), .B2(n19791), .ZN(
        n19771) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19780), .B1(
        n19772), .B2(n19988), .ZN(n19770) );
  OAI211_X1 U22765 ( .C1(n19991), .C2(n19805), .A(n19771), .B(n19770), .ZN(
        P2_U3107) );
  AOI22_X1 U22766 ( .A1(n19779), .A2(n19543), .B1(n20044), .B2(n19791), .ZN(
        n19774) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19780), .B1(
        n19772), .B2(n20045), .ZN(n19773) );
  OAI211_X1 U22768 ( .C1(n20048), .C2(n19805), .A(n19774), .B(n19773), .ZN(
        P2_U3108) );
  AOI22_X1 U22769 ( .A1(n19779), .A2(n19550), .B1(n19548), .B2(n19791), .ZN(
        n19776) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n19923), .ZN(n19775) );
  OAI211_X1 U22771 ( .C1(n19926), .C2(n19783), .A(n19776), .B(n19775), .ZN(
        P2_U3109) );
  AOI22_X1 U22772 ( .A1(n19779), .A2(n20054), .B1(n20053), .B2(n19791), .ZN(
        n19778) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n19998), .ZN(n19777) );
  OAI211_X1 U22774 ( .C1(n20002), .C2(n19783), .A(n19778), .B(n19777), .ZN(
        P2_U3110) );
  AOI22_X1 U22775 ( .A1(n19779), .A2(n20063), .B1(n20061), .B2(n19791), .ZN(
        n19782) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19780), .B1(
        n19811), .B2(n20065), .ZN(n19781) );
  OAI211_X1 U22777 ( .C1(n20071), .C2(n19783), .A(n19782), .B(n19781), .ZN(
        P2_U3111) );
  NOR2_X1 U22778 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19784), .ZN(
        n19810) );
  AOI22_X1 U22779 ( .A1(n19946), .A2(n19811), .B1(n20016), .B2(n19810), .ZN(
        n19796) );
  NAND2_X1 U22780 ( .A1(n19805), .A2(n19826), .ZN(n19785) );
  AOI21_X1 U22781 ( .B1(n19785), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19973), 
        .ZN(n19790) );
  INV_X1 U22782 ( .A(n19786), .ZN(n19792) );
  OAI21_X1 U22783 ( .B1(n19792), .B2(n20013), .A(n12466), .ZN(n19787) );
  AOI21_X1 U22784 ( .B1(n19790), .B2(n19788), .A(n19787), .ZN(n19789) );
  OAI21_X1 U22785 ( .B1(n19810), .B2(n19789), .A(n19975), .ZN(n19813) );
  OAI21_X1 U22786 ( .B1(n19810), .B2(n19791), .A(n19790), .ZN(n19794) );
  OAI21_X1 U22787 ( .B1(n19792), .B2(n19810), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19793) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19813), .B1(
        n13458), .B2(n19812), .ZN(n19795) );
  OAI211_X1 U22789 ( .C1(n19949), .C2(n19826), .A(n19796), .B(n19795), .ZN(
        P2_U3112) );
  AOI22_X1 U22790 ( .A1(n20030), .A2(n19811), .B1(n19810), .B2(n20029), .ZN(
        n19798) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19527), .ZN(n19797) );
  OAI211_X1 U22792 ( .C1(n20033), .C2(n19826), .A(n19798), .B(n19797), .ZN(
        P2_U3113) );
  AOI22_X1 U22793 ( .A1(n20035), .A2(n19811), .B1(n19810), .B2(n9818), .ZN(
        n19800) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19532), .ZN(n19799) );
  OAI211_X1 U22795 ( .C1(n20038), .C2(n19826), .A(n19800), .B(n19799), .ZN(
        P2_U3114) );
  AOI22_X1 U22796 ( .A1(n20040), .A2(n19829), .B1(n19810), .B2(n20039), .ZN(
        n19802) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19536), .ZN(n19801) );
  OAI211_X1 U22798 ( .C1(n20043), .C2(n19805), .A(n19802), .B(n19801), .ZN(
        P2_U3115) );
  AOI22_X1 U22799 ( .A1(n19992), .A2(n19829), .B1(n19810), .B2(n20044), .ZN(
        n19804) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19543), .ZN(n19803) );
  OAI211_X1 U22801 ( .C1(n19995), .C2(n19805), .A(n19804), .B(n19803), .ZN(
        P2_U3116) );
  AOI22_X1 U22802 ( .A1(n20049), .A2(n19811), .B1(n19810), .B2(n19548), .ZN(
        n19807) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19550), .ZN(n19806) );
  OAI211_X1 U22804 ( .C1(n20052), .C2(n19826), .A(n19807), .B(n19806), .ZN(
        P2_U3117) );
  AOI22_X1 U22805 ( .A1(n20055), .A2(n19811), .B1(n19810), .B2(n20053), .ZN(
        n19809) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n20054), .ZN(n19808) );
  OAI211_X1 U22807 ( .C1(n20060), .C2(n19826), .A(n19809), .B(n19808), .ZN(
        P2_U3118) );
  AOI22_X1 U22808 ( .A1(n20005), .A2(n19811), .B1(n19810), .B2(n20061), .ZN(
        n19815) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n20063), .ZN(n19814) );
  OAI211_X1 U22810 ( .C1(n20010), .C2(n19826), .A(n19815), .B(n19814), .ZN(
        P2_U3119) );
  AOI22_X1 U22811 ( .A1(n19911), .A2(n19859), .B1(n19840), .B2(n20029), .ZN(
        n19817) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19831), .B1(
        n19527), .B2(n19830), .ZN(n19816) );
  OAI211_X1 U22813 ( .C1(n19914), .C2(n19826), .A(n19817), .B(n19816), .ZN(
        P2_U3121) );
  INV_X1 U22814 ( .A(n19859), .ZN(n19834) );
  AOI22_X1 U22815 ( .A1(n20035), .A2(n19829), .B1(n19840), .B2(n9818), .ZN(
        n19819) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19831), .B1(
        n19532), .B2(n19830), .ZN(n19818) );
  OAI211_X1 U22817 ( .C1(n20038), .C2(n19834), .A(n19819), .B(n19818), .ZN(
        P2_U3122) );
  AOI22_X1 U22818 ( .A1(n20040), .A2(n19859), .B1(n19840), .B2(n20039), .ZN(
        n19821) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19831), .B1(
        n19536), .B2(n19830), .ZN(n19820) );
  OAI211_X1 U22820 ( .C1(n20043), .C2(n19826), .A(n19821), .B(n19820), .ZN(
        P2_U3123) );
  AOI22_X1 U22821 ( .A1(n20045), .A2(n19829), .B1(n19840), .B2(n20044), .ZN(
        n19823) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19831), .B1(
        n19543), .B2(n19830), .ZN(n19822) );
  OAI211_X1 U22823 ( .C1(n20048), .C2(n19834), .A(n19823), .B(n19822), .ZN(
        P2_U3124) );
  AOI22_X1 U22824 ( .A1(n19923), .A2(n19859), .B1(n19840), .B2(n19548), .ZN(
        n19825) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19831), .B1(
        n19550), .B2(n19830), .ZN(n19824) );
  OAI211_X1 U22826 ( .C1(n19926), .C2(n19826), .A(n19825), .B(n19824), .ZN(
        P2_U3125) );
  AOI22_X1 U22827 ( .A1(n20055), .A2(n19829), .B1(n19840), .B2(n20053), .ZN(
        n19828) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19831), .B1(
        n20054), .B2(n19830), .ZN(n19827) );
  OAI211_X1 U22829 ( .C1(n20060), .C2(n19834), .A(n19828), .B(n19827), .ZN(
        P2_U3126) );
  AOI22_X1 U22830 ( .A1(n20005), .A2(n19829), .B1(n19840), .B2(n20061), .ZN(
        n19833) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19831), .B1(
        n20063), .B2(n19830), .ZN(n19832) );
  OAI211_X1 U22832 ( .C1(n20010), .C2(n19834), .A(n19833), .B(n19832), .ZN(
        P2_U3127) );
  INV_X1 U22833 ( .A(n13784), .ZN(n19837) );
  NOR2_X1 U22834 ( .A1(n19836), .A2(n19869), .ZN(n19857) );
  OAI21_X1 U22835 ( .B1(n19837), .B2(n19857), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19838) );
  OAI21_X1 U22836 ( .B1(n19869), .B2(n19839), .A(n19838), .ZN(n19858) );
  AOI22_X1 U22837 ( .A1(n19858), .A2(n13458), .B1(n20016), .B2(n19857), .ZN(
        n19844) );
  AOI221_X1 U22838 ( .B1(n19859), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19894), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19840), .ZN(n19841) );
  AOI211_X1 U22839 ( .C1(n13784), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19841), .ZN(n19842) );
  OAI21_X1 U22840 ( .B1(n19842), .B2(n19857), .A(n19975), .ZN(n19860) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n19946), .ZN(n19843) );
  OAI211_X1 U22842 ( .C1(n19949), .C2(n19863), .A(n19844), .B(n19843), .ZN(
        P2_U3128) );
  AOI22_X1 U22843 ( .A1(n19858), .A2(n19527), .B1(n20029), .B2(n19857), .ZN(
        n19846) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20030), .ZN(n19845) );
  OAI211_X1 U22845 ( .C1(n20033), .C2(n19863), .A(n19846), .B(n19845), .ZN(
        P2_U3129) );
  AOI22_X1 U22846 ( .A1(n19858), .A2(n19532), .B1(n9818), .B2(n19857), .ZN(
        n19848) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20035), .ZN(n19847) );
  OAI211_X1 U22848 ( .C1(n20038), .C2(n19863), .A(n19848), .B(n19847), .ZN(
        P2_U3130) );
  AOI22_X1 U22849 ( .A1(n19858), .A2(n19536), .B1(n20039), .B2(n19857), .ZN(
        n19850) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n19988), .ZN(n19849) );
  OAI211_X1 U22851 ( .C1(n19991), .C2(n19863), .A(n19850), .B(n19849), .ZN(
        P2_U3131) );
  AOI22_X1 U22852 ( .A1(n19858), .A2(n19543), .B1(n20044), .B2(n19857), .ZN(
        n19852) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20045), .ZN(n19851) );
  OAI211_X1 U22854 ( .C1(n20048), .C2(n19863), .A(n19852), .B(n19851), .ZN(
        P2_U3132) );
  AOI22_X1 U22855 ( .A1(n19858), .A2(n19550), .B1(n19548), .B2(n19857), .ZN(
        n19854) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20049), .ZN(n19853) );
  OAI211_X1 U22857 ( .C1(n20052), .C2(n19863), .A(n19854), .B(n19853), .ZN(
        P2_U3133) );
  AOI22_X1 U22858 ( .A1(n19858), .A2(n20054), .B1(n20053), .B2(n19857), .ZN(
        n19856) );
  AOI22_X1 U22859 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20055), .ZN(n19855) );
  OAI211_X1 U22860 ( .C1(n20060), .C2(n19863), .A(n19856), .B(n19855), .ZN(
        P2_U3134) );
  AOI22_X1 U22861 ( .A1(n19858), .A2(n20063), .B1(n20061), .B2(n19857), .ZN(
        n19862) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19860), .B1(
        n19859), .B2(n20005), .ZN(n19861) );
  OAI211_X1 U22863 ( .C1(n20010), .C2(n19863), .A(n19862), .B(n19861), .ZN(
        P2_U3135) );
  INV_X1 U22864 ( .A(n19865), .ZN(n19867) );
  INV_X1 U22865 ( .A(n19869), .ZN(n19866) );
  NAND2_X1 U22866 ( .A1(n19867), .A2(n19866), .ZN(n19875) );
  NAND3_X1 U22867 ( .A1(n19868), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19875), 
        .ZN(n19873) );
  NOR2_X1 U22868 ( .A1(n20190), .A2(n19869), .ZN(n19877) );
  INV_X1 U22869 ( .A(n19877), .ZN(n19870) );
  OAI21_X1 U22870 ( .B1(n19870), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20013), 
        .ZN(n19871) );
  AND2_X1 U22871 ( .A1(n19873), .A2(n19871), .ZN(n19893) );
  INV_X1 U22872 ( .A(n19875), .ZN(n19892) );
  AOI22_X1 U22873 ( .A1(n19893), .A2(n13458), .B1(n20016), .B2(n19892), .ZN(
        n19879) );
  INV_X1 U22874 ( .A(n19872), .ZN(n20022) );
  INV_X1 U22875 ( .A(n19873), .ZN(n19874) );
  AOI211_X1 U22876 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19875), .A(n20019), 
        .B(n19874), .ZN(n19876) );
  OAI221_X1 U22877 ( .B1(n19877), .B2(n20162), .C1(n19877), .C2(n20022), .A(
        n19876), .ZN(n19895) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n19946), .ZN(n19878) );
  OAI211_X1 U22879 ( .C1(n19949), .C2(n19934), .A(n19879), .B(n19878), .ZN(
        P2_U3136) );
  AOI22_X1 U22880 ( .A1(n19893), .A2(n19527), .B1(n20029), .B2(n19892), .ZN(
        n19881) );
  AOI22_X1 U22881 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20030), .ZN(n19880) );
  OAI211_X1 U22882 ( .C1(n20033), .C2(n19934), .A(n19881), .B(n19880), .ZN(
        P2_U3137) );
  AOI22_X1 U22883 ( .A1(n19893), .A2(n19532), .B1(n9818), .B2(n19892), .ZN(
        n19883) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20035), .ZN(n19882) );
  OAI211_X1 U22885 ( .C1(n20038), .C2(n19934), .A(n19883), .B(n19882), .ZN(
        P2_U3138) );
  AOI22_X1 U22886 ( .A1(n19893), .A2(n19536), .B1(n20039), .B2(n19892), .ZN(
        n19885) );
  AOI22_X1 U22887 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n19988), .ZN(n19884) );
  OAI211_X1 U22888 ( .C1(n19991), .C2(n19934), .A(n19885), .B(n19884), .ZN(
        P2_U3139) );
  AOI22_X1 U22889 ( .A1(n19893), .A2(n19543), .B1(n20044), .B2(n19892), .ZN(
        n19887) );
  AOI22_X1 U22890 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20045), .ZN(n19886) );
  OAI211_X1 U22891 ( .C1(n20048), .C2(n19934), .A(n19887), .B(n19886), .ZN(
        P2_U3140) );
  AOI22_X1 U22892 ( .A1(n19893), .A2(n19550), .B1(n19548), .B2(n19892), .ZN(
        n19889) );
  AOI22_X1 U22893 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20049), .ZN(n19888) );
  OAI211_X1 U22894 ( .C1(n20052), .C2(n19934), .A(n19889), .B(n19888), .ZN(
        P2_U3141) );
  AOI22_X1 U22895 ( .A1(n19893), .A2(n20054), .B1(n20053), .B2(n19892), .ZN(
        n19891) );
  AOI22_X1 U22896 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20055), .ZN(n19890) );
  OAI211_X1 U22897 ( .C1(n20060), .C2(n19934), .A(n19891), .B(n19890), .ZN(
        P2_U3142) );
  AOI22_X1 U22898 ( .A1(n19893), .A2(n20063), .B1(n20061), .B2(n19892), .ZN(
        n19897) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19895), .B1(
        n19894), .B2(n20005), .ZN(n19896) );
  OAI211_X1 U22900 ( .C1(n20010), .C2(n19934), .A(n19897), .B(n19896), .ZN(
        P2_U3143) );
  INV_X1 U22901 ( .A(n19898), .ZN(n19902) );
  INV_X1 U22902 ( .A(n19907), .ZN(n19901) );
  INV_X1 U22903 ( .A(n19899), .ZN(n19903) );
  NOR3_X1 U22904 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20181), .A3(
        n10685), .ZN(n19945) );
  INV_X1 U22905 ( .A(n19945), .ZN(n19937) );
  NOR2_X1 U22906 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19937), .ZN(
        n19929) );
  OAI21_X1 U22907 ( .B1(n19903), .B2(n19929), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19900) );
  OAI21_X1 U22908 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(n19930) );
  AOI22_X1 U22909 ( .A1(n19930), .A2(n13458), .B1(n20016), .B2(n19929), .ZN(
        n19910) );
  INV_X1 U22910 ( .A(n19958), .ZN(n19967) );
  AOI21_X1 U22911 ( .B1(n19934), .B2(n19967), .A(n12714), .ZN(n19908) );
  OAI21_X1 U22912 ( .B1(n19903), .B2(n20013), .A(n12466), .ZN(n19905) );
  INV_X1 U22913 ( .A(n19929), .ZN(n19904) );
  AOI21_X1 U22914 ( .B1(n19905), .B2(n19904), .A(n20019), .ZN(n19906) );
  OAI211_X1 U22915 ( .C1(n19908), .C2(n19907), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19906), .ZN(n19931) );
  AOI22_X1 U22916 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n20025), .ZN(n19909) );
  OAI211_X1 U22917 ( .C1(n20028), .C2(n19934), .A(n19910), .B(n19909), .ZN(
        P2_U3144) );
  AOI22_X1 U22918 ( .A1(n19930), .A2(n19527), .B1(n20029), .B2(n19929), .ZN(
        n19913) );
  AOI22_X1 U22919 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n19911), .ZN(n19912) );
  OAI211_X1 U22920 ( .C1(n19914), .C2(n19934), .A(n19913), .B(n19912), .ZN(
        P2_U3145) );
  AOI22_X1 U22921 ( .A1(n19930), .A2(n19532), .B1(n9818), .B2(n19929), .ZN(
        n19917) );
  AOI22_X1 U22922 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n19915), .ZN(n19916) );
  OAI211_X1 U22923 ( .C1(n19918), .C2(n19934), .A(n19917), .B(n19916), .ZN(
        P2_U3146) );
  AOI22_X1 U22924 ( .A1(n19930), .A2(n19536), .B1(n20039), .B2(n19929), .ZN(
        n19920) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n20040), .ZN(n19919) );
  OAI211_X1 U22926 ( .C1(n20043), .C2(n19934), .A(n19920), .B(n19919), .ZN(
        P2_U3147) );
  AOI22_X1 U22927 ( .A1(n19930), .A2(n19543), .B1(n20044), .B2(n19929), .ZN(
        n19922) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n19992), .ZN(n19921) );
  OAI211_X1 U22929 ( .C1(n19995), .C2(n19934), .A(n19922), .B(n19921), .ZN(
        P2_U3148) );
  AOI22_X1 U22930 ( .A1(n19930), .A2(n19550), .B1(n19548), .B2(n19929), .ZN(
        n19925) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n19923), .ZN(n19924) );
  OAI211_X1 U22932 ( .C1(n19926), .C2(n19934), .A(n19925), .B(n19924), .ZN(
        P2_U3149) );
  AOI22_X1 U22933 ( .A1(n19930), .A2(n20054), .B1(n20053), .B2(n19929), .ZN(
        n19928) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n19998), .ZN(n19927) );
  OAI211_X1 U22935 ( .C1(n20002), .C2(n19934), .A(n19928), .B(n19927), .ZN(
        P2_U3150) );
  AOI22_X1 U22936 ( .A1(n19930), .A2(n20063), .B1(n20061), .B2(n19929), .ZN(
        n19933) );
  AOI22_X1 U22937 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19931), .B1(
        n19958), .B2(n20065), .ZN(n19932) );
  OAI211_X1 U22938 ( .C1(n20071), .C2(n19934), .A(n19933), .B(n19932), .ZN(
        P2_U3151) );
  OR2_X1 U22939 ( .A1(n19937), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19940) );
  INV_X1 U22940 ( .A(n19938), .ZN(n19939) );
  NAND2_X1 U22941 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19945), .ZN(
        n19942) );
  INV_X1 U22942 ( .A(n19942), .ZN(n19971) );
  NOR3_X1 U22943 ( .A1(n19939), .A2(n19971), .A3(n20013), .ZN(n19941) );
  AOI21_X1 U22944 ( .B1(n20013), .B2(n19940), .A(n19941), .ZN(n19963) );
  AOI22_X1 U22945 ( .A1(n19963), .A2(n13458), .B1(n20016), .B2(n19971), .ZN(
        n19948) );
  AOI211_X1 U22946 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19942), .A(n20019), 
        .B(n19941), .ZN(n19943) );
  OAI221_X1 U22947 ( .B1(n19945), .B2(n19944), .C1(n19945), .C2(n20022), .A(
        n19943), .ZN(n19964) );
  AOI22_X1 U22948 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n19946), .ZN(n19947) );
  OAI211_X1 U22949 ( .C1(n19949), .C2(n20001), .A(n19948), .B(n19947), .ZN(
        P2_U3152) );
  AOI22_X1 U22950 ( .A1(n19963), .A2(n19527), .B1(n20029), .B2(n19971), .ZN(
        n19951) );
  AOI22_X1 U22951 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n20030), .ZN(n19950) );
  OAI211_X1 U22952 ( .C1(n20033), .C2(n20001), .A(n19951), .B(n19950), .ZN(
        P2_U3153) );
  AOI22_X1 U22953 ( .A1(n19963), .A2(n19532), .B1(n9818), .B2(n19971), .ZN(
        n19953) );
  AOI22_X1 U22954 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n20035), .ZN(n19952) );
  OAI211_X1 U22955 ( .C1(n20038), .C2(n20001), .A(n19953), .B(n19952), .ZN(
        P2_U3154) );
  AOI22_X1 U22956 ( .A1(n19963), .A2(n19536), .B1(n20039), .B2(n19971), .ZN(
        n19955) );
  AOI22_X1 U22957 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n19988), .ZN(n19954) );
  OAI211_X1 U22958 ( .C1(n19991), .C2(n20001), .A(n19955), .B(n19954), .ZN(
        P2_U3155) );
  AOI22_X1 U22959 ( .A1(n19963), .A2(n19543), .B1(n20044), .B2(n19971), .ZN(
        n19957) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n20045), .ZN(n19956) );
  OAI211_X1 U22961 ( .C1(n20048), .C2(n20001), .A(n19957), .B(n19956), .ZN(
        P2_U3156) );
  AOI22_X1 U22962 ( .A1(n19963), .A2(n19550), .B1(n19548), .B2(n19971), .ZN(
        n19960) );
  AOI22_X1 U22963 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19964), .B1(
        n19958), .B2(n20049), .ZN(n19959) );
  OAI211_X1 U22964 ( .C1(n20052), .C2(n20001), .A(n19960), .B(n19959), .ZN(
        P2_U3157) );
  AOI22_X1 U22965 ( .A1(n19963), .A2(n20054), .B1(n20053), .B2(n19971), .ZN(
        n19962) );
  AOI22_X1 U22966 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19964), .B1(
        n20004), .B2(n19998), .ZN(n19961) );
  OAI211_X1 U22967 ( .C1(n20002), .C2(n19967), .A(n19962), .B(n19961), .ZN(
        P2_U3158) );
  AOI22_X1 U22968 ( .A1(n19963), .A2(n20063), .B1(n20061), .B2(n19971), .ZN(
        n19966) );
  AOI22_X1 U22969 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19964), .B1(
        n20004), .B2(n20065), .ZN(n19965) );
  OAI211_X1 U22970 ( .C1(n20071), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        P2_U3159) );
  NOR3_X2 U22971 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10685), .A3(
        n20012), .ZN(n20003) );
  AOI22_X1 U22972 ( .A1(n20025), .A2(n20056), .B1(n20016), .B2(n20003), .ZN(
        n19983) );
  NOR2_X1 U22973 ( .A1(n20056), .A2(n20004), .ZN(n19970) );
  OAI21_X1 U22974 ( .B1(n19970), .B2(n12714), .A(n20169), .ZN(n19981) );
  NOR2_X1 U22975 ( .A1(n20003), .A2(n19971), .ZN(n19980) );
  INV_X1 U22976 ( .A(n19980), .ZN(n19976) );
  INV_X1 U22977 ( .A(n20003), .ZN(n19972) );
  OAI211_X1 U22978 ( .C1(n19977), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19973), 
        .B(n19972), .ZN(n19974) );
  OAI211_X1 U22979 ( .C1(n19981), .C2(n19976), .A(n19975), .B(n19974), .ZN(
        n20007) );
  INV_X1 U22980 ( .A(n19977), .ZN(n19978) );
  OAI21_X1 U22981 ( .B1(n19978), .B2(n20003), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19979) );
  AOI22_X1 U22982 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20007), .B1(
        n13458), .B2(n20006), .ZN(n19982) );
  OAI211_X1 U22983 ( .C1(n20028), .C2(n20001), .A(n19983), .B(n19982), .ZN(
        P2_U3160) );
  AOI22_X1 U22984 ( .A1(n20030), .A2(n20004), .B1(n20029), .B2(n20003), .ZN(
        n19985) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20007), .B1(
        n19527), .B2(n20006), .ZN(n19984) );
  OAI211_X1 U22986 ( .C1(n20033), .C2(n20070), .A(n19985), .B(n19984), .ZN(
        P2_U3161) );
  AOI22_X1 U22987 ( .A1(n20035), .A2(n20004), .B1(n9818), .B2(n20003), .ZN(
        n19987) );
  AOI22_X1 U22988 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20007), .B1(
        n19532), .B2(n20006), .ZN(n19986) );
  OAI211_X1 U22989 ( .C1(n20038), .C2(n20070), .A(n19987), .B(n19986), .ZN(
        P2_U3162) );
  AOI22_X1 U22990 ( .A1(n19988), .A2(n20004), .B1(n20039), .B2(n20003), .ZN(
        n19990) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20007), .B1(
        n19536), .B2(n20006), .ZN(n19989) );
  OAI211_X1 U22992 ( .C1(n19991), .C2(n20070), .A(n19990), .B(n19989), .ZN(
        P2_U3163) );
  AOI22_X1 U22993 ( .A1(n19992), .A2(n20056), .B1(n20044), .B2(n20003), .ZN(
        n19994) );
  AOI22_X1 U22994 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20007), .B1(
        n19543), .B2(n20006), .ZN(n19993) );
  OAI211_X1 U22995 ( .C1(n19995), .C2(n20001), .A(n19994), .B(n19993), .ZN(
        P2_U3164) );
  AOI22_X1 U22996 ( .A1(n20049), .A2(n20004), .B1(n20003), .B2(n19548), .ZN(
        n19997) );
  AOI22_X1 U22997 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20007), .B1(
        n19550), .B2(n20006), .ZN(n19996) );
  OAI211_X1 U22998 ( .C1(n20052), .C2(n20070), .A(n19997), .B(n19996), .ZN(
        P2_U3165) );
  AOI22_X1 U22999 ( .A1(n19998), .A2(n20056), .B1(n20053), .B2(n20003), .ZN(
        n20000) );
  AOI22_X1 U23000 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20007), .B1(
        n20054), .B2(n20006), .ZN(n19999) );
  OAI211_X1 U23001 ( .C1(n20002), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3166) );
  AOI22_X1 U23002 ( .A1(n20005), .A2(n20004), .B1(n20061), .B2(n20003), .ZN(
        n20009) );
  AOI22_X1 U23003 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20007), .B1(
        n20063), .B2(n20006), .ZN(n20008) );
  OAI211_X1 U23004 ( .C1(n20010), .C2(n20070), .A(n20009), .B(n20008), .ZN(
        P2_U3167) );
  NAND3_X1 U23005 ( .A1(n20011), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20020), 
        .ZN(n20017) );
  NOR2_X1 U23006 ( .A1(n10685), .A2(n20012), .ZN(n20024) );
  INV_X1 U23007 ( .A(n20024), .ZN(n20014) );
  OAI21_X1 U23008 ( .B1(n20014), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20013), 
        .ZN(n20015) );
  AND2_X1 U23009 ( .A1(n20017), .A2(n20015), .ZN(n20064) );
  AOI22_X1 U23010 ( .A1(n20064), .A2(n13458), .B1(n20062), .B2(n20016), .ZN(
        n20027) );
  INV_X1 U23011 ( .A(n20017), .ZN(n20018) );
  AOI211_X1 U23012 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20020), .A(n20019), 
        .B(n20018), .ZN(n20021) );
  OAI221_X1 U23013 ( .B1(n20024), .B2(n20023), .C1(n20024), .C2(n20022), .A(
        n20021), .ZN(n20067) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20067), .B1(
        n20066), .B2(n20025), .ZN(n20026) );
  OAI211_X1 U23015 ( .C1(n20028), .C2(n20070), .A(n20027), .B(n20026), .ZN(
        P2_U3168) );
  AOI22_X1 U23016 ( .A1(n20064), .A2(n19527), .B1(n20062), .B2(n20029), .ZN(
        n20032) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20067), .B1(
        n20056), .B2(n20030), .ZN(n20031) );
  OAI211_X1 U23018 ( .C1(n20033), .C2(n20059), .A(n20032), .B(n20031), .ZN(
        P2_U3169) );
  AOI22_X1 U23019 ( .A1(n20064), .A2(n19532), .B1(n20062), .B2(n9818), .ZN(
        n20037) );
  AOI22_X1 U23020 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20067), .B1(
        n20056), .B2(n20035), .ZN(n20036) );
  OAI211_X1 U23021 ( .C1(n20038), .C2(n20059), .A(n20037), .B(n20036), .ZN(
        P2_U3170) );
  AOI22_X1 U23022 ( .A1(n20064), .A2(n19536), .B1(n20062), .B2(n20039), .ZN(
        n20042) );
  AOI22_X1 U23023 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20067), .B1(
        n20066), .B2(n20040), .ZN(n20041) );
  OAI211_X1 U23024 ( .C1(n20043), .C2(n20070), .A(n20042), .B(n20041), .ZN(
        P2_U3171) );
  AOI22_X1 U23025 ( .A1(n20064), .A2(n19543), .B1(n20062), .B2(n20044), .ZN(
        n20047) );
  AOI22_X1 U23026 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20067), .B1(
        n20056), .B2(n20045), .ZN(n20046) );
  OAI211_X1 U23027 ( .C1(n20048), .C2(n20059), .A(n20047), .B(n20046), .ZN(
        P2_U3172) );
  AOI22_X1 U23028 ( .A1(n20064), .A2(n19550), .B1(n20062), .B2(n19548), .ZN(
        n20051) );
  AOI22_X1 U23029 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20067), .B1(
        n20056), .B2(n20049), .ZN(n20050) );
  OAI211_X1 U23030 ( .C1(n20052), .C2(n20059), .A(n20051), .B(n20050), .ZN(
        P2_U3173) );
  AOI22_X1 U23031 ( .A1(n20064), .A2(n20054), .B1(n20062), .B2(n20053), .ZN(
        n20058) );
  AOI22_X1 U23032 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20067), .B1(
        n20056), .B2(n20055), .ZN(n20057) );
  OAI211_X1 U23033 ( .C1(n20060), .C2(n20059), .A(n20058), .B(n20057), .ZN(
        P2_U3174) );
  AOI22_X1 U23034 ( .A1(n20064), .A2(n20063), .B1(n20062), .B2(n20061), .ZN(
        n20069) );
  AOI22_X1 U23035 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20067), .B1(
        n20066), .B2(n20065), .ZN(n20068) );
  OAI211_X1 U23036 ( .C1(n20071), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P2_U3175) );
  AOI21_X1 U23037 ( .B1(n20074), .B2(n20073), .A(n20072), .ZN(n20080) );
  OAI211_X1 U23038 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20216), .A(n20076), 
        .B(n20075), .ZN(n20077) );
  OAI22_X1 U23039 ( .A1(n20080), .A2(n20079), .B1(n20078), .B2(n20077), .ZN(
        P2_U3177) );
  AND2_X1 U23040 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20081), .ZN(
        P2_U3179) );
  AND2_X1 U23041 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20081), .ZN(
        P2_U3180) );
  AND2_X1 U23042 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20081), .ZN(
        P2_U3181) );
  AND2_X1 U23043 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20081), .ZN(
        P2_U3182) );
  AND2_X1 U23044 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20081), .ZN(
        P2_U3183) );
  AND2_X1 U23045 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20081), .ZN(
        P2_U3184) );
  AND2_X1 U23046 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20081), .ZN(
        P2_U3185) );
  AND2_X1 U23047 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20081), .ZN(
        P2_U3186) );
  AND2_X1 U23048 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20081), .ZN(
        P2_U3187) );
  AND2_X1 U23049 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20081), .ZN(
        P2_U3188) );
  AND2_X1 U23050 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20081), .ZN(
        P2_U3189) );
  AND2_X1 U23051 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20081), .ZN(
        P2_U3190) );
  AND2_X1 U23052 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20081), .ZN(
        P2_U3191) );
  AND2_X1 U23053 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20081), .ZN(
        P2_U3192) );
  AND2_X1 U23054 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20081), .ZN(
        P2_U3193) );
  AND2_X1 U23055 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20081), .ZN(
        P2_U3194) );
  AND2_X1 U23056 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20081), .ZN(
        P2_U3195) );
  AND2_X1 U23057 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20081), .ZN(
        P2_U3196) );
  AND2_X1 U23058 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20081), .ZN(
        P2_U3197) );
  AND2_X1 U23059 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20081), .ZN(
        P2_U3198) );
  AND2_X1 U23060 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20081), .ZN(
        P2_U3199) );
  AND2_X1 U23061 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20081), .ZN(
        P2_U3200) );
  AND2_X1 U23062 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20081), .ZN(P2_U3201) );
  AND2_X1 U23063 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20081), .ZN(P2_U3202) );
  AND2_X1 U23064 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20081), .ZN(P2_U3203) );
  AND2_X1 U23065 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20081), .ZN(P2_U3204) );
  AND2_X1 U23066 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20081), .ZN(P2_U3205) );
  AND2_X1 U23067 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20081), .ZN(P2_U3206) );
  AND2_X1 U23068 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20081), .ZN(P2_U3207) );
  AND2_X1 U23069 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20081), .ZN(P2_U3208) );
  INV_X1 U23070 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20082) );
  NOR2_X1 U23071 ( .A1(n20216), .A2(n20082), .ZN(n20093) );
  INV_X1 U23072 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20229) );
  NOR3_X1 U23073 ( .A1(n20093), .A2(n20229), .A3(n20083), .ZN(n20087) );
  OAI211_X1 U23074 ( .C1(HOLD), .C2(n20229), .A(n20230), .B(n20084), .ZN(
        n20086) );
  INV_X1 U23075 ( .A(NA), .ZN(n21039) );
  NOR3_X1 U23076 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21039), .ZN(n20095) );
  INV_X1 U23077 ( .A(n20095), .ZN(n20085) );
  OAI211_X1 U23078 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20087), .A(n20086), 
        .B(n20085), .ZN(P2_U3209) );
  AOI21_X1 U23079 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21329), .A(n20098), 
        .ZN(n20092) );
  NOR3_X1 U23080 ( .A1(n20083), .A2(n20092), .A3(n20229), .ZN(n20088) );
  NOR3_X1 U23081 ( .A1(n20224), .A2(n20093), .A3(n20088), .ZN(n20089) );
  OAI21_X1 U23082 ( .B1(n21329), .B2(n20090), .A(n20089), .ZN(P2_U3210) );
  AOI22_X1 U23083 ( .A1(n20091), .A2(n20229), .B1(n20093), .B2(n21039), .ZN(
        n20097) );
  OAI21_X1 U23084 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20096) );
  AOI21_X1 U23085 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20093), .A(n20092), 
        .ZN(n20094) );
  OAI22_X1 U23086 ( .A1(n20097), .A2(n20096), .B1(n20095), .B2(n20094), .ZN(
        P2_U3211) );
  NAND2_X1 U23087 ( .A1(n20148), .A2(n20098), .ZN(n20151) );
  OAI222_X1 U23088 ( .A1(n20145), .A2(n15007), .B1(n20100), .B2(n20148), .C1(
        n20099), .C2(n20146), .ZN(P2_U3212) );
  OAI222_X1 U23089 ( .A1(n20146), .A2(n15007), .B1(n20101), .B2(n20148), .C1(
        n13568), .C2(n20145), .ZN(P2_U3213) );
  OAI222_X1 U23090 ( .A1(n20146), .A2(n13568), .B1(n20102), .B2(n20148), .C1(
        n12532), .C2(n20145), .ZN(P2_U3214) );
  OAI222_X1 U23091 ( .A1(n20151), .A2(n12476), .B1(n20103), .B2(n20148), .C1(
        n12532), .C2(n20146), .ZN(P2_U3215) );
  OAI222_X1 U23092 ( .A1(n20151), .A2(n12535), .B1(n20104), .B2(n20148), .C1(
        n12476), .C2(n20146), .ZN(P2_U3216) );
  INV_X1 U23093 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20106) );
  OAI222_X1 U23094 ( .A1(n20151), .A2(n20106), .B1(n20105), .B2(n20148), .C1(
        n12535), .C2(n20146), .ZN(P2_U3217) );
  OAI222_X1 U23095 ( .A1(n20151), .A2(n20108), .B1(n20107), .B2(n20148), .C1(
        n20106), .C2(n20146), .ZN(P2_U3218) );
  OAI222_X1 U23096 ( .A1(n20151), .A2(n12538), .B1(n20109), .B2(n20148), .C1(
        n20108), .C2(n20146), .ZN(P2_U3219) );
  OAI222_X1 U23097 ( .A1(n20145), .A2(n12543), .B1(n20110), .B2(n20148), .C1(
        n12538), .C2(n20146), .ZN(P2_U3220) );
  OAI222_X1 U23098 ( .A1(n20145), .A2(n20112), .B1(n20111), .B2(n20148), .C1(
        n12543), .C2(n20146), .ZN(P2_U3221) );
  OAI222_X1 U23099 ( .A1(n20145), .A2(n13956), .B1(n20113), .B2(n20148), .C1(
        n20112), .C2(n20146), .ZN(P2_U3222) );
  OAI222_X1 U23100 ( .A1(n20145), .A2(n13957), .B1(n20114), .B2(n20148), .C1(
        n13956), .C2(n20146), .ZN(P2_U3223) );
  OAI222_X1 U23101 ( .A1(n20145), .A2(n13965), .B1(n20115), .B2(n20148), .C1(
        n13957), .C2(n20146), .ZN(P2_U3224) );
  OAI222_X1 U23102 ( .A1(n20145), .A2(n20117), .B1(n20116), .B2(n20148), .C1(
        n13965), .C2(n20146), .ZN(P2_U3225) );
  OAI222_X1 U23103 ( .A1(n20151), .A2(n20119), .B1(n20118), .B2(n20148), .C1(
        n20117), .C2(n20146), .ZN(P2_U3226) );
  OAI222_X1 U23104 ( .A1(n20151), .A2(n20121), .B1(n20120), .B2(n20148), .C1(
        n20119), .C2(n20146), .ZN(P2_U3227) );
  OAI222_X1 U23105 ( .A1(n20151), .A2(n20123), .B1(n20122), .B2(n20148), .C1(
        n20121), .C2(n20146), .ZN(P2_U3228) );
  OAI222_X1 U23106 ( .A1(n20151), .A2(n14022), .B1(n20124), .B2(n20148), .C1(
        n20123), .C2(n20146), .ZN(P2_U3229) );
  OAI222_X1 U23107 ( .A1(n20151), .A2(n20126), .B1(n20125), .B2(n20148), .C1(
        n14022), .C2(n20146), .ZN(P2_U3230) );
  OAI222_X1 U23108 ( .A1(n20151), .A2(n20128), .B1(n20127), .B2(n20148), .C1(
        n20126), .C2(n20146), .ZN(P2_U3231) );
  OAI222_X1 U23109 ( .A1(n20145), .A2(n20130), .B1(n20129), .B2(n20148), .C1(
        n20128), .C2(n20146), .ZN(P2_U3232) );
  OAI222_X1 U23110 ( .A1(n20145), .A2(n15287), .B1(n20131), .B2(n20148), .C1(
        n20130), .C2(n20146), .ZN(P2_U3233) );
  INV_X1 U23111 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20133) );
  OAI222_X1 U23112 ( .A1(n20145), .A2(n20133), .B1(n20132), .B2(n20148), .C1(
        n15287), .C2(n20146), .ZN(P2_U3234) );
  OAI222_X1 U23113 ( .A1(n20145), .A2(n20135), .B1(n20134), .B2(n20148), .C1(
        n20133), .C2(n20146), .ZN(P2_U3235) );
  OAI222_X1 U23114 ( .A1(n20145), .A2(n20137), .B1(n20136), .B2(n20148), .C1(
        n20135), .C2(n20146), .ZN(P2_U3236) );
  OAI222_X1 U23115 ( .A1(n20145), .A2(n20140), .B1(n20138), .B2(n20148), .C1(
        n20137), .C2(n20146), .ZN(P2_U3237) );
  OAI222_X1 U23116 ( .A1(n20146), .A2(n20140), .B1(n20139), .B2(n20148), .C1(
        n20141), .C2(n20145), .ZN(P2_U3238) );
  OAI222_X1 U23117 ( .A1(n20145), .A2(n20143), .B1(n20142), .B2(n20148), .C1(
        n20141), .C2(n20146), .ZN(P2_U3239) );
  OAI222_X1 U23118 ( .A1(n20145), .A2(n20147), .B1(n20144), .B2(n20148), .C1(
        n20143), .C2(n20146), .ZN(P2_U3240) );
  INV_X1 U23119 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20149) );
  OAI222_X1 U23120 ( .A1(n20151), .A2(n20150), .B1(n20149), .B2(n20148), .C1(
        n20147), .C2(n20146), .ZN(P2_U3241) );
  INV_X1 U23121 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20152) );
  AOI22_X1 U23122 ( .A1(n20148), .A2(n20153), .B1(n20152), .B2(n20230), .ZN(
        P2_U3585) );
  MUX2_X1 U23123 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20148), .Z(P2_U3586) );
  INV_X1 U23124 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20154) );
  AOI22_X1 U23125 ( .A1(n20148), .A2(n20155), .B1(n20154), .B2(n20230), .ZN(
        P2_U3587) );
  INV_X1 U23126 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U23127 ( .A1(n20148), .A2(n20157), .B1(n20156), .B2(n20230), .ZN(
        P2_U3588) );
  OAI21_X1 U23128 ( .B1(n20161), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20159), 
        .ZN(n20158) );
  INV_X1 U23129 ( .A(n20158), .ZN(P2_U3591) );
  OAI21_X1 U23130 ( .B1(n20161), .B2(n20160), .A(n20159), .ZN(P2_U3592) );
  AND2_X1 U23131 ( .A1(n20169), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20186) );
  NAND2_X1 U23132 ( .A1(n20162), .A2(n20186), .ZN(n20175) );
  NOR2_X1 U23133 ( .A1(n20163), .A2(n12714), .ZN(n20164) );
  NAND2_X1 U23134 ( .A1(n20184), .A2(n20164), .ZN(n20165) );
  NAND2_X1 U23135 ( .A1(n20165), .A2(n20182), .ZN(n20176) );
  NAND2_X1 U23136 ( .A1(n20175), .A2(n20176), .ZN(n20168) );
  AOI22_X1 U23137 ( .A1(n20168), .A2(n20167), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20166), .ZN(n20172) );
  NAND2_X1 U23138 ( .A1(n20170), .A2(n20169), .ZN(n20171) );
  AND2_X1 U23139 ( .A1(n20172), .A2(n20171), .ZN(n20173) );
  AOI22_X1 U23140 ( .A1(n20197), .A2(n10685), .B1(n20173), .B2(n20198), .ZN(
        P2_U3602) );
  INV_X1 U23141 ( .A(n20174), .ZN(n20177) );
  OAI21_X1 U23142 ( .B1(n20177), .B2(n20176), .A(n20175), .ZN(n20178) );
  AOI21_X1 U23143 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20179), .A(n20178), 
        .ZN(n20180) );
  AOI22_X1 U23144 ( .A1(n20197), .A2(n20181), .B1(n20180), .B2(n20198), .ZN(
        P2_U3603) );
  INV_X1 U23145 ( .A(n20182), .ZN(n20193) );
  NOR2_X1 U23146 ( .A1(n20193), .A2(n20183), .ZN(n20185) );
  MUX2_X1 U23147 ( .A(n20186), .B(n20185), .S(n20184), .Z(n20187) );
  AOI21_X1 U23148 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20188), .A(n20187), 
        .ZN(n20189) );
  AOI22_X1 U23149 ( .A1(n20197), .A2(n20190), .B1(n20189), .B2(n20198), .ZN(
        P2_U3604) );
  OAI22_X1 U23150 ( .A1(n20194), .A2(n20193), .B1(n20192), .B2(n20191), .ZN(
        n20195) );
  AOI21_X1 U23151 ( .B1(n20199), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20195), 
        .ZN(n20196) );
  OAI22_X1 U23152 ( .A1(n20199), .A2(n20198), .B1(n20197), .B2(n20196), .ZN(
        P2_U3605) );
  INV_X1 U23153 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20200) );
  AOI22_X1 U23154 ( .A1(n20148), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20200), 
        .B2(n20230), .ZN(P2_U3608) );
  INV_X1 U23155 ( .A(n20201), .ZN(n20202) );
  AOI22_X1 U23156 ( .A1(n20205), .A2(n20204), .B1(n20203), .B2(n20202), .ZN(
        n20206) );
  NAND2_X1 U23157 ( .A1(n20207), .A2(n20206), .ZN(n20209) );
  MUX2_X1 U23158 ( .A(P2_MORE_REG_SCAN_IN), .B(n20209), .S(n20208), .Z(
        P2_U3609) );
  INV_X1 U23159 ( .A(n20216), .ZN(n20212) );
  OAI22_X1 U23160 ( .A1(n20212), .A2(n20211), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20210), .ZN(n20213) );
  NOR2_X1 U23161 ( .A1(n20214), .A2(n20213), .ZN(n20228) );
  NAND2_X1 U23162 ( .A1(n20218), .A2(n20215), .ZN(n20221) );
  NAND2_X1 U23163 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20216), .ZN(n20220) );
  NOR4_X1 U23164 ( .A1(n20224), .A2(n9838), .A3(n20218), .A4(n20217), .ZN(
        n20219) );
  AOI21_X1 U23165 ( .B1(n20221), .B2(n20220), .A(n20219), .ZN(n20227) );
  AOI211_X1 U23166 ( .C1(n20224), .C2(P2_STATEBS16_REG_SCAN_IN), .A(n9833), 
        .B(n20222), .ZN(n20225) );
  NOR2_X1 U23167 ( .A1(n20228), .A2(n20225), .ZN(n20226) );
  AOI22_X1 U23168 ( .A1(n20229), .A2(n20228), .B1(n20227), .B2(n20226), .ZN(
        P2_U3610) );
  OAI22_X1 U23169 ( .A1(n20230), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20148), .ZN(n20231) );
  INV_X1 U23170 ( .A(n20231), .ZN(P2_U3611) );
  NOR2_X1 U23171 ( .A1(n21036), .A2(n21038), .ZN(n20240) );
  INV_X1 U23172 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20233) );
  INV_X1 U23173 ( .A(n21115), .ZN(n21116) );
  AOI21_X1 U23174 ( .B1(n20240), .B2(n20233), .A(n21116), .ZN(P1_U2802) );
  INV_X1 U23175 ( .A(n20234), .ZN(n20236) );
  OAI21_X1 U23176 ( .B1(n20236), .B2(n20235), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20237) );
  OAI21_X1 U23177 ( .B1(n20238), .B2(n21026), .A(n20237), .ZN(P1_U2803) );
  INV_X1 U23178 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n21347) );
  NOR2_X1 U23179 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20241) );
  NOR2_X1 U23180 ( .A1(n21116), .A2(n20241), .ZN(n20239) );
  AOI22_X1 U23181 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n21116), .B1(n21347), 
        .B2(n20239), .ZN(P1_U2804) );
  NOR2_X1 U23182 ( .A1(n21116), .A2(n20240), .ZN(n21030) );
  OAI21_X1 U23183 ( .B1(BS16), .B2(n20241), .A(n21030), .ZN(n21092) );
  OAI21_X1 U23184 ( .B1(n21030), .B2(n21220), .A(n21092), .ZN(P1_U2805) );
  OAI21_X1 U23185 ( .B1(n20243), .B2(n21311), .A(n20242), .ZN(P1_U2806) );
  NOR4_X1 U23186 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20247) );
  NOR4_X1 U23187 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20246) );
  NOR4_X1 U23188 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20245) );
  NOR4_X1 U23189 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20244) );
  NAND4_X1 U23190 ( .A1(n20247), .A2(n20246), .A3(n20245), .A4(n20244), .ZN(
        n20253) );
  NOR4_X1 U23191 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20251) );
  AOI211_X1 U23192 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20250) );
  NOR4_X1 U23193 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20249) );
  NOR4_X1 U23194 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20248) );
  NAND4_X1 U23195 ( .A1(n20251), .A2(n20250), .A3(n20249), .A4(n20248), .ZN(
        n20252) );
  NOR2_X1 U23196 ( .A1(n20253), .A2(n20252), .ZN(n21103) );
  INV_X1 U23197 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21282) );
  NOR3_X1 U23198 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20255) );
  OAI21_X1 U23199 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20255), .A(n21103), .ZN(
        n20254) );
  OAI21_X1 U23200 ( .B1(n21103), .B2(n21282), .A(n20254), .ZN(P1_U2807) );
  INV_X1 U23201 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21276) );
  NOR2_X1 U23202 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21098) );
  OAI21_X1 U23203 ( .B1(n20255), .B2(n21098), .A(n21103), .ZN(n20256) );
  OAI21_X1 U23204 ( .B1(n21103), .B2(n21276), .A(n20256), .ZN(P1_U2808) );
  NAND2_X1 U23205 ( .A1(n20270), .A2(n20257), .ZN(n20261) );
  INV_X1 U23206 ( .A(n20258), .ZN(n20259) );
  AOI22_X1 U23207 ( .A1(n20288), .A2(n20259), .B1(n20315), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20260) );
  OAI21_X1 U23208 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20261), .A(n20260), .ZN(
        n20262) );
  AOI211_X1 U23209 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20306), .B(n20262), .ZN(n20267) );
  AOI22_X1 U23210 ( .A1(n20265), .A2(n20292), .B1(n20264), .B2(n20263), .ZN(
        n20266) );
  OAI211_X1 U23211 ( .C1(n20268), .C2(n21326), .A(n20267), .B(n20266), .ZN(
        P1_U2831) );
  AOI22_X1 U23212 ( .A1(n20288), .A2(n20269), .B1(n20315), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20274) );
  AND2_X1 U23213 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .ZN(n20280) );
  INV_X1 U23214 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20272) );
  NAND2_X1 U23215 ( .A1(n20270), .A2(n20276), .ZN(n20300) );
  INV_X1 U23216 ( .A(n20300), .ZN(n20271) );
  NAND3_X1 U23217 ( .A1(n20280), .A2(n20272), .A3(n20271), .ZN(n20273) );
  NAND2_X1 U23218 ( .A1(n20274), .A2(n20273), .ZN(n20275) );
  AOI211_X1 U23219 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20306), .B(n20275), .ZN(n20283) );
  OR2_X1 U23220 ( .A1(n20318), .A2(n20276), .ZN(n20278) );
  AND2_X1 U23221 ( .A1(n20278), .A2(n20277), .ZN(n20316) );
  OAI21_X1 U23222 ( .B1(n20280), .B2(n20279), .A(n20316), .ZN(n20293) );
  AOI22_X1 U23223 ( .A1(n20281), .A2(n20292), .B1(n20293), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20282) );
  OAI211_X1 U23224 ( .C1(n20284), .C2(n20324), .A(n20283), .B(n20282), .ZN(
        P1_U2833) );
  INV_X1 U23225 ( .A(n20285), .ZN(n20287) );
  NOR2_X1 U23226 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20300), .ZN(n20286) );
  AOI22_X1 U23227 ( .A1(n20288), .A2(n20287), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20286), .ZN(n20289) );
  OAI21_X1 U23228 ( .B1(n21248), .B2(n20297), .A(n20289), .ZN(n20290) );
  AOI211_X1 U23229 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20306), .B(n20290), .ZN(n20295) );
  AOI22_X1 U23230 ( .A1(n20293), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20292), 
        .B2(n20291), .ZN(n20294) );
  OAI211_X1 U23231 ( .C1(n20296), .C2(n20324), .A(n20295), .B(n20294), .ZN(
        P1_U2834) );
  INV_X1 U23232 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21218) );
  OAI22_X1 U23233 ( .A1(n20316), .A2(n21218), .B1(n21450), .B2(n20297), .ZN(
        n20298) );
  AOI211_X1 U23234 ( .C1(n20307), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20306), .B(n20298), .ZN(n20304) );
  OAI22_X1 U23235 ( .A1(n20300), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20313), 
        .B2(n20299), .ZN(n20301) );
  AOI21_X1 U23236 ( .B1(n20302), .B2(n20321), .A(n20301), .ZN(n20303) );
  OAI211_X1 U23237 ( .C1(n20305), .C2(n20324), .A(n20304), .B(n20303), .ZN(
        P1_U2835) );
  AOI21_X1 U23238 ( .B1(n20307), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20306), .ZN(n20311) );
  NAND2_X1 U23239 ( .A1(n20309), .A2(n20308), .ZN(n20310) );
  OAI211_X1 U23240 ( .C1(n20313), .C2(n20312), .A(n20311), .B(n20310), .ZN(
        n20314) );
  AOI21_X1 U23241 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n20315), .A(n20314), .ZN(
        n20323) );
  INV_X1 U23242 ( .A(n20316), .ZN(n20320) );
  OAI21_X1 U23243 ( .B1(n20318), .B2(n20317), .A(n21265), .ZN(n20319) );
  AOI22_X1 U23244 ( .A1(n20369), .A2(n20321), .B1(n20320), .B2(n20319), .ZN(
        n20322) );
  OAI211_X1 U23245 ( .C1(n20373), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        P1_U2836) );
  AOI22_X1 U23246 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20328), .B1(n15999), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20325) );
  OAI21_X1 U23247 ( .B1(n20327), .B2(n20326), .A(n20325), .ZN(P1_U2921) );
  AOI22_X1 U23248 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20329) );
  OAI21_X1 U23249 ( .B1(n14072), .B2(n20349), .A(n20329), .ZN(P1_U2922) );
  AOI22_X1 U23250 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20330) );
  OAI21_X1 U23251 ( .B1(n14675), .B2(n20349), .A(n20330), .ZN(P1_U2923) );
  AOI22_X1 U23252 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20331) );
  OAI21_X1 U23253 ( .B1(n14053), .B2(n20349), .A(n20331), .ZN(P1_U2924) );
  AOI22_X1 U23254 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20332) );
  OAI21_X1 U23255 ( .B1(n13981), .B2(n20349), .A(n20332), .ZN(P1_U2925) );
  AOI22_X1 U23256 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20333) );
  OAI21_X1 U23257 ( .B1(n13750), .B2(n20349), .A(n20333), .ZN(P1_U2926) );
  AOI22_X1 U23258 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20334) );
  OAI21_X1 U23259 ( .B1(n13728), .B2(n20349), .A(n20334), .ZN(P1_U2927) );
  AOI22_X1 U23260 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20335) );
  OAI21_X1 U23261 ( .B1(n13661), .B2(n20349), .A(n20335), .ZN(P1_U2928) );
  AOI22_X1 U23262 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20336) );
  OAI21_X1 U23263 ( .B1(n20337), .B2(n20349), .A(n20336), .ZN(P1_U2929) );
  AOI22_X1 U23264 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20338) );
  OAI21_X1 U23265 ( .B1(n11632), .B2(n20349), .A(n20338), .ZN(P1_U2930) );
  AOI22_X1 U23266 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20339) );
  OAI21_X1 U23267 ( .B1(n11553), .B2(n20349), .A(n20339), .ZN(P1_U2931) );
  AOI22_X1 U23268 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20340) );
  OAI21_X1 U23269 ( .B1(n20341), .B2(n20349), .A(n20340), .ZN(P1_U2932) );
  AOI22_X1 U23270 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20342) );
  OAI21_X1 U23271 ( .B1(n20343), .B2(n20349), .A(n20342), .ZN(P1_U2933) );
  AOI22_X1 U23272 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20344) );
  OAI21_X1 U23273 ( .B1(n20345), .B2(n20349), .A(n20344), .ZN(P1_U2934) );
  AOI22_X1 U23274 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20346) );
  OAI21_X1 U23275 ( .B1(n20347), .B2(n20349), .A(n20346), .ZN(P1_U2935) );
  AOI22_X1 U23276 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21111), .B1(n15999), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20348) );
  OAI21_X1 U23277 ( .B1(n20350), .B2(n20349), .A(n20348), .ZN(P1_U2936) );
  AOI22_X1 U23278 ( .A1(n20362), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20361), .ZN(n20352) );
  NAND2_X1 U23279 ( .A1(n20352), .A2(n20351), .ZN(P1_U2961) );
  AOI22_X1 U23280 ( .A1(n20362), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20361), .ZN(n20354) );
  NAND2_X1 U23281 ( .A1(n20354), .A2(n20353), .ZN(P1_U2962) );
  AOI22_X1 U23282 ( .A1(n20362), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20361), .ZN(n20356) );
  NAND2_X1 U23283 ( .A1(n20356), .A2(n20355), .ZN(P1_U2963) );
  AOI22_X1 U23284 ( .A1(n20362), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20361), .ZN(n20358) );
  NAND2_X1 U23285 ( .A1(n20358), .A2(n20357), .ZN(P1_U2964) );
  AOI22_X1 U23286 ( .A1(n20362), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20361), .ZN(n20360) );
  NAND2_X1 U23287 ( .A1(n20360), .A2(n20359), .ZN(P1_U2965) );
  AOI22_X1 U23288 ( .A1(n20362), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20361), .ZN(n20364) );
  NAND2_X1 U23289 ( .A1(n20364), .A2(n20363), .ZN(P1_U2966) );
  AOI22_X1 U23290 ( .A1(n20365), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20380), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20372) );
  XOR2_X1 U23291 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n20366), .Z(
        n20367) );
  XNOR2_X1 U23292 ( .A(n20368), .B(n20367), .ZN(n20378) );
  AOI22_X1 U23293 ( .A1(n20378), .A2(n20370), .B1(n14411), .B2(n20369), .ZN(
        n20371) );
  OAI211_X1 U23294 ( .C1(n20374), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P1_U2995) );
  INV_X1 U23295 ( .A(n20375), .ZN(n20376) );
  NOR2_X1 U23296 ( .A1(n20377), .A2(n20376), .ZN(n20394) );
  AOI222_X1 U23297 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20380), .B1(n20404), 
        .B2(n20379), .C1(n20405), .C2(n20378), .ZN(n20384) );
  OAI211_X1 U23298 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20382), .B(n20381), .ZN(n20383) );
  OAI211_X1 U23299 ( .C1(n20394), .C2(n13670), .A(n20384), .B(n20383), .ZN(
        P1_U3027) );
  AOI21_X1 U23300 ( .B1(n20404), .B2(n20386), .A(n20385), .ZN(n20392) );
  OAI22_X1 U23301 ( .A1(n20389), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20388), .B2(n20387), .ZN(n20390) );
  INV_X1 U23302 ( .A(n20390), .ZN(n20391) );
  OAI211_X1 U23303 ( .C1(n20394), .C2(n20393), .A(n20392), .B(n20391), .ZN(
        P1_U3028) );
  AOI21_X1 U23304 ( .B1(n20397), .B2(n20396), .A(n20395), .ZN(n20410) );
  NAND3_X1 U23305 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20399) );
  AOI21_X1 U23306 ( .B1(n20400), .B2(n20399), .A(n20398), .ZN(n20401) );
  AOI211_X1 U23307 ( .C1(n20404), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        n20408) );
  NAND3_X1 U23308 ( .A1(n20406), .A2(n13328), .A3(n20405), .ZN(n20407) );
  AND2_X1 U23309 ( .A1(n20408), .A2(n20407), .ZN(n20409) );
  OAI221_X1 U23310 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20412), .C1(
        n20411), .C2(n20410), .A(n20409), .ZN(P1_U3029) );
  NOR2_X1 U23311 ( .A1(n20414), .A2(n20413), .ZN(P1_U3032) );
  AOI22_X1 U23312 ( .A1(DATAI_16_), .A2(n20477), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20476), .ZN(n20898) );
  INV_X1 U23313 ( .A(n12986), .ZN(n20418) );
  INV_X1 U23314 ( .A(n20476), .ZN(n20469) );
  INV_X1 U23315 ( .A(DATAI_24_), .ZN(n21469) );
  OAI22_X1 U23316 ( .A1(n20421), .A2(n20469), .B1(n21469), .B2(n20468), .ZN(
        n20895) );
  INV_X1 U23317 ( .A(n20895), .ZN(n20980) );
  NAND2_X1 U23318 ( .A1(n20479), .A2(n20423), .ZN(n20840) );
  NAND3_X1 U23319 ( .A1(n20804), .A2(n20764), .A3(n20839), .ZN(n20487) );
  OR2_X1 U23320 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20487), .ZN(
        n20480) );
  OAI22_X1 U23321 ( .A1(n20976), .A2(n20980), .B1(n20840), .B2(n20480), .ZN(
        n20424) );
  INV_X1 U23322 ( .A(n20424), .ZN(n20438) );
  INV_X1 U23323 ( .A(n20425), .ZN(n20711) );
  INV_X1 U23324 ( .A(n20768), .ZN(n20426) );
  NOR2_X1 U23325 ( .A1(n20711), .A2(n20426), .ZN(n20434) );
  NAND2_X1 U23326 ( .A1(n20433), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20930) );
  NAND3_X1 U23327 ( .A1(n20506), .A2(n20842), .A3(n20976), .ZN(n20428) );
  NAND2_X1 U23328 ( .A1(n20842), .A2(n21220), .ZN(n20843) );
  NAND2_X1 U23329 ( .A1(n20428), .A2(n20843), .ZN(n20432) );
  NAND2_X1 U23330 ( .A1(n9928), .A2(n20932), .ZN(n20435) );
  AOI22_X1 U23331 ( .A1(n20432), .A2(n20435), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20480), .ZN(n20430) );
  OAI211_X1 U23332 ( .C1(n20434), .C2(n21028), .A(n20771), .B(n20430), .ZN(
        n20484) );
  NOR2_X2 U23333 ( .A1(n20431), .A2(n20593), .ZN(n20968) );
  INV_X1 U23334 ( .A(n20432), .ZN(n20436) );
  NOR2_X1 U23335 ( .A1(n20433), .A2(n21028), .ZN(n20594) );
  INV_X1 U23336 ( .A(n20594), .ZN(n20774) );
  INV_X1 U23337 ( .A(n20434), .ZN(n20590) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20484), .B1(
        n20968), .B2(n20483), .ZN(n20437) );
  OAI211_X1 U23339 ( .C1(n20898), .C2(n20506), .A(n20438), .B(n20437), .ZN(
        P1_U3033) );
  AOI22_X1 U23340 ( .A1(DATAI_17_), .A2(n20477), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20476), .ZN(n20902) );
  INV_X1 U23341 ( .A(DATAI_25_), .ZN(n21263) );
  OAI22_X1 U23342 ( .A1(n20439), .A2(n20469), .B1(n21263), .B2(n20468), .ZN(
        n20899) );
  INV_X1 U23343 ( .A(n20899), .ZN(n20985) );
  NAND2_X1 U23344 ( .A1(n20479), .A2(n20440), .ZN(n20855) );
  OAI22_X1 U23345 ( .A1(n20976), .A2(n20985), .B1(n20855), .B2(n20480), .ZN(
        n20441) );
  INV_X1 U23346 ( .A(n20441), .ZN(n20444) );
  NOR2_X2 U23347 ( .A1(n20442), .A2(n20593), .ZN(n20981) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20484), .B1(
        n20981), .B2(n20483), .ZN(n20443) );
  OAI211_X1 U23349 ( .C1(n9983), .C2(n20506), .A(n20444), .B(n20443), .ZN(
        P1_U3034) );
  INV_X1 U23350 ( .A(DATAI_26_), .ZN(n21212) );
  OAI22_X1 U23351 ( .A1(n20445), .A2(n20469), .B1(n21212), .B2(n20468), .ZN(
        n20903) );
  INV_X1 U23352 ( .A(n20903), .ZN(n20991) );
  NAND2_X1 U23353 ( .A1(n20479), .A2(n20446), .ZN(n20859) );
  OAI22_X1 U23354 ( .A1(n20976), .A2(n20991), .B1(n20859), .B2(n20480), .ZN(
        n20447) );
  INV_X1 U23355 ( .A(n20447), .ZN(n20450) );
  NOR2_X2 U23356 ( .A1(n20448), .A2(n20593), .ZN(n20986) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20484), .B1(
        n20986), .B2(n20483), .ZN(n20449) );
  OAI211_X1 U23358 ( .C1(n20906), .C2(n20506), .A(n20450), .B(n20449), .ZN(
        P1_U3035) );
  AOI22_X1 U23359 ( .A1(DATAI_19_), .A2(n20477), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20476), .ZN(n20910) );
  INV_X1 U23360 ( .A(DATAI_27_), .ZN(n21287) );
  OAI22_X1 U23361 ( .A1(n20451), .A2(n20469), .B1(n21287), .B2(n20468), .ZN(
        n20907) );
  NAND2_X1 U23362 ( .A1(n20479), .A2(n20452), .ZN(n20863) );
  OAI22_X1 U23363 ( .A1(n20976), .A2(n20997), .B1(n20863), .B2(n20480), .ZN(
        n20453) );
  INV_X1 U23364 ( .A(n20453), .ZN(n20456) );
  NOR2_X2 U23365 ( .A1(n20454), .A2(n20593), .ZN(n20992) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20484), .B1(
        n20992), .B2(n20483), .ZN(n20455) );
  OAI211_X1 U23367 ( .C1(n20910), .C2(n20506), .A(n20456), .B(n20455), .ZN(
        P1_U3036) );
  AOI22_X1 U23368 ( .A1(DATAI_20_), .A2(n20477), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20476), .ZN(n20914) );
  INV_X1 U23369 ( .A(DATAI_28_), .ZN(n21284) );
  OAI22_X1 U23370 ( .A1(n20457), .A2(n20469), .B1(n21284), .B2(n20468), .ZN(
        n20911) );
  INV_X1 U23371 ( .A(n20911), .ZN(n21002) );
  OAI22_X1 U23372 ( .A1(n20976), .A2(n21002), .B1(n20867), .B2(n20480), .ZN(
        n20458) );
  INV_X1 U23373 ( .A(n20458), .ZN(n20461) );
  NOR2_X2 U23374 ( .A1(n20459), .A2(n20593), .ZN(n20998) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20484), .B1(
        n20998), .B2(n20483), .ZN(n20460) );
  OAI211_X1 U23376 ( .C1(n9979), .C2(n20506), .A(n20461), .B(n20460), .ZN(
        P1_U3037) );
  AOI22_X1 U23377 ( .A1(DATAI_21_), .A2(n20477), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20476), .ZN(n20918) );
  INV_X1 U23378 ( .A(DATAI_29_), .ZN(n21274) );
  OAI22_X1 U23379 ( .A1(n20462), .A2(n20469), .B1(n21274), .B2(n20468), .ZN(
        n20915) );
  INV_X1 U23380 ( .A(n20915), .ZN(n21008) );
  NAND2_X1 U23381 ( .A1(n20479), .A2(n20463), .ZN(n20871) );
  OAI22_X1 U23382 ( .A1(n20976), .A2(n21008), .B1(n20871), .B2(n20480), .ZN(
        n20464) );
  INV_X1 U23383 ( .A(n20464), .ZN(n20467) );
  NOR2_X2 U23384 ( .A1(n20465), .A2(n20593), .ZN(n21003) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20484), .B1(
        n21003), .B2(n20483), .ZN(n20466) );
  OAI211_X1 U23386 ( .C1(n20918), .C2(n20506), .A(n20467), .B(n20466), .ZN(
        P1_U3038) );
  INV_X1 U23387 ( .A(DATAI_30_), .ZN(n21211) );
  OAI22_X1 U23388 ( .A1(n20470), .A2(n20469), .B1(n21211), .B2(n20468), .ZN(
        n20919) );
  INV_X1 U23389 ( .A(n20919), .ZN(n21014) );
  NAND2_X1 U23390 ( .A1(n20479), .A2(n20471), .ZN(n20875) );
  OAI22_X1 U23391 ( .A1(n20976), .A2(n21014), .B1(n20875), .B2(n20480), .ZN(
        n20472) );
  INV_X1 U23392 ( .A(n20472), .ZN(n20475) );
  NOR2_X2 U23393 ( .A1(n20473), .A2(n20593), .ZN(n21009) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20484), .B1(
        n21009), .B2(n20483), .ZN(n20474) );
  OAI211_X1 U23395 ( .C1(n20922), .C2(n20506), .A(n20475), .B(n20474), .ZN(
        P1_U3039) );
  AOI22_X1 U23396 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20476), .B1(DATAI_23_), 
        .B2(n20477), .ZN(n20929) );
  AOI22_X1 U23397 ( .A1(DATAI_31_), .A2(n20477), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20476), .ZN(n21024) );
  NAND2_X1 U23398 ( .A1(n20479), .A2(n20478), .ZN(n20880) );
  OAI22_X1 U23399 ( .A1(n20976), .A2(n9977), .B1(n20880), .B2(n20480), .ZN(
        n20481) );
  INV_X1 U23400 ( .A(n20481), .ZN(n20486) );
  NOR2_X2 U23401 ( .A1(n20593), .A2(n20482), .ZN(n21016) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20484), .B1(
        n21016), .B2(n20483), .ZN(n20485) );
  OAI211_X1 U23403 ( .C1(n9981), .C2(n20506), .A(n20486), .B(n20485), .ZN(
        P1_U3040) );
  NOR2_X1 U23404 ( .A1(n20889), .A2(n20487), .ZN(n20508) );
  INV_X1 U23405 ( .A(n20890), .ZN(n20736) );
  AOI21_X1 U23406 ( .B1(n9928), .B2(n20736), .A(n20508), .ZN(n20488) );
  OAI22_X1 U23407 ( .A1(n20488), .A2(n20967), .B1(n20487), .B2(n21028), .ZN(
        n20507) );
  AOI22_X1 U23408 ( .A1(n20969), .A2(n20508), .B1(n20507), .B2(n20968), .ZN(
        n20492) );
  INV_X1 U23409 ( .A(n20487), .ZN(n20490) );
  OAI211_X1 U23410 ( .C1(n20555), .C2(n21220), .A(n20842), .B(n20488), .ZN(
        n20489) );
  OAI211_X1 U23411 ( .C1(n20842), .C2(n20490), .A(n20974), .B(n20489), .ZN(
        n20510) );
  INV_X1 U23412 ( .A(n20548), .ZN(n20503) );
  INV_X1 U23413 ( .A(n20898), .ZN(n20977) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20510), .B1(
        n20503), .B2(n20977), .ZN(n20491) );
  OAI211_X1 U23415 ( .C1(n20980), .C2(n20506), .A(n20492), .B(n20491), .ZN(
        P1_U3041) );
  AOI22_X1 U23416 ( .A1(n20982), .A2(n20508), .B1(n20507), .B2(n20981), .ZN(
        n20494) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20510), .B1(
        n20503), .B2(n9982), .ZN(n20493) );
  OAI211_X1 U23418 ( .C1(n20985), .C2(n20506), .A(n20494), .B(n20493), .ZN(
        P1_U3042) );
  AOI22_X1 U23419 ( .A1(n20987), .A2(n20508), .B1(n20507), .B2(n20986), .ZN(
        n20496) );
  INV_X1 U23420 ( .A(n20506), .ZN(n20509) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20510), .B1(
        n20509), .B2(n20903), .ZN(n20495) );
  OAI211_X1 U23422 ( .C1(n20906), .C2(n20548), .A(n20496), .B(n20495), .ZN(
        P1_U3043) );
  AOI22_X1 U23423 ( .A1(n20993), .A2(n20508), .B1(n20507), .B2(n20992), .ZN(
        n20498) );
  INV_X1 U23424 ( .A(n20910), .ZN(n20994) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20510), .B1(
        n20503), .B2(n20994), .ZN(n20497) );
  OAI211_X1 U23426 ( .C1(n20997), .C2(n20506), .A(n20498), .B(n20497), .ZN(
        P1_U3044) );
  AOI22_X1 U23427 ( .A1(n20999), .A2(n20508), .B1(n20507), .B2(n20998), .ZN(
        n20500) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20510), .B1(
        n20509), .B2(n20911), .ZN(n20499) );
  OAI211_X1 U23429 ( .C1(n9979), .C2(n20548), .A(n20500), .B(n20499), .ZN(
        P1_U3045) );
  AOI22_X1 U23430 ( .A1(n21004), .A2(n20508), .B1(n20507), .B2(n21003), .ZN(
        n20502) );
  INV_X1 U23431 ( .A(n20918), .ZN(n21005) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20510), .B1(
        n20503), .B2(n21005), .ZN(n20501) );
  OAI211_X1 U23433 ( .C1(n21008), .C2(n20506), .A(n20502), .B(n20501), .ZN(
        P1_U3046) );
  AOI22_X1 U23434 ( .A1(n21010), .A2(n20508), .B1(n20507), .B2(n21009), .ZN(
        n20505) );
  INV_X1 U23435 ( .A(n20922), .ZN(n21011) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20510), .B1(
        n20503), .B2(n21011), .ZN(n20504) );
  OAI211_X1 U23437 ( .C1(n21014), .C2(n20506), .A(n20505), .B(n20504), .ZN(
        P1_U3047) );
  AOI22_X1 U23438 ( .A1(n21018), .A2(n20508), .B1(n21016), .B2(n20507), .ZN(
        n20512) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20510), .B1(
        n20509), .B2(n9976), .ZN(n20511) );
  OAI211_X1 U23440 ( .C1(n9981), .C2(n20548), .A(n20512), .B(n20511), .ZN(
        P1_U3048) );
  NAND3_X1 U23441 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20804), .A3(
        n20764), .ZN(n20558) );
  NOR2_X1 U23442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20558), .ZN(
        n20516) );
  INV_X1 U23443 ( .A(n20516), .ZN(n20542) );
  OAI22_X1 U23444 ( .A1(n20548), .A2(n20980), .B1(n20542), .B2(n20840), .ZN(
        n20514) );
  INV_X1 U23445 ( .A(n20514), .ZN(n20523) );
  NAND2_X1 U23446 ( .A1(n20582), .A2(n20548), .ZN(n20515) );
  AOI21_X1 U23447 ( .B1(n20515), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20967), 
        .ZN(n20519) );
  NAND2_X1 U23448 ( .A1(n9928), .A2(n20936), .ZN(n20520) );
  NOR2_X1 U23449 ( .A1(n20516), .A2(n20847), .ZN(n20517) );
  AOI21_X1 U23450 ( .B1(n20519), .B2(n20520), .A(n20517), .ZN(n20518) );
  OR2_X1 U23451 ( .A1(n20768), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20648) );
  NAND2_X1 U23452 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20648), .ZN(n20645) );
  NAND3_X1 U23453 ( .A1(n20771), .A2(n20518), .A3(n20645), .ZN(n20545) );
  INV_X1 U23454 ( .A(n20519), .ZN(n20521) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20545), .B1(
        n20968), .B2(n20544), .ZN(n20522) );
  OAI211_X1 U23456 ( .C1(n20898), .C2(n20582), .A(n20523), .B(n20522), .ZN(
        P1_U3049) );
  OAI22_X1 U23457 ( .A1(n20582), .A2(n9983), .B1(n20855), .B2(n20542), .ZN(
        n20524) );
  INV_X1 U23458 ( .A(n20524), .ZN(n20526) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20545), .B1(
        n20981), .B2(n20544), .ZN(n20525) );
  OAI211_X1 U23460 ( .C1(n20985), .C2(n20548), .A(n20526), .B(n20525), .ZN(
        P1_U3050) );
  OAI22_X1 U23461 ( .A1(n20548), .A2(n20991), .B1(n20542), .B2(n20859), .ZN(
        n20527) );
  INV_X1 U23462 ( .A(n20527), .ZN(n20529) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20545), .B1(
        n20986), .B2(n20544), .ZN(n20528) );
  OAI211_X1 U23464 ( .C1(n20906), .C2(n20582), .A(n20529), .B(n20528), .ZN(
        P1_U3051) );
  OAI22_X1 U23465 ( .A1(n20582), .A2(n20910), .B1(n20542), .B2(n20863), .ZN(
        n20530) );
  INV_X1 U23466 ( .A(n20530), .ZN(n20532) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20545), .B1(
        n20992), .B2(n20544), .ZN(n20531) );
  OAI211_X1 U23468 ( .C1(n20997), .C2(n20548), .A(n20532), .B(n20531), .ZN(
        P1_U3052) );
  OAI22_X1 U23469 ( .A1(n20582), .A2(n9979), .B1(n20542), .B2(n20867), .ZN(
        n20533) );
  INV_X1 U23470 ( .A(n20533), .ZN(n20535) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20545), .B1(
        n20998), .B2(n20544), .ZN(n20534) );
  OAI211_X1 U23472 ( .C1(n21002), .C2(n20548), .A(n20535), .B(n20534), .ZN(
        P1_U3053) );
  OAI22_X1 U23473 ( .A1(n20582), .A2(n20918), .B1(n20542), .B2(n20871), .ZN(
        n20536) );
  INV_X1 U23474 ( .A(n20536), .ZN(n20538) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20545), .B1(
        n21003), .B2(n20544), .ZN(n20537) );
  OAI211_X1 U23476 ( .C1(n21008), .C2(n20548), .A(n20538), .B(n20537), .ZN(
        P1_U3054) );
  OAI22_X1 U23477 ( .A1(n20548), .A2(n21014), .B1(n20542), .B2(n20875), .ZN(
        n20539) );
  INV_X1 U23478 ( .A(n20539), .ZN(n20541) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20545), .B1(
        n21009), .B2(n20544), .ZN(n20540) );
  OAI211_X1 U23480 ( .C1(n20922), .C2(n20582), .A(n20541), .B(n20540), .ZN(
        P1_U3055) );
  OAI22_X1 U23481 ( .A1(n20582), .A2(n9981), .B1(n20542), .B2(n20880), .ZN(
        n20543) );
  INV_X1 U23482 ( .A(n20543), .ZN(n20547) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20545), .B1(
        n21016), .B2(n20544), .ZN(n20546) );
  OAI211_X1 U23484 ( .C1(n9977), .C2(n20548), .A(n20547), .B(n20546), .ZN(
        P1_U3056) );
  INV_X1 U23485 ( .A(n20805), .ZN(n20549) );
  NAND2_X1 U23486 ( .A1(n20549), .A2(n20804), .ZN(n20581) );
  OAI22_X1 U23487 ( .A1(n20596), .A2(n20898), .B1(n20581), .B2(n20840), .ZN(
        n20550) );
  INV_X1 U23488 ( .A(n20550), .ZN(n20562) );
  NOR2_X1 U23489 ( .A1(n20552), .A2(n20551), .ZN(n20963) );
  INV_X1 U23490 ( .A(n20581), .ZN(n20553) );
  AOI21_X1 U23491 ( .B1(n9928), .B2(n20963), .A(n20553), .ZN(n20559) );
  AOI21_X1 U23492 ( .B1(n20555), .B2(n20842), .A(n20554), .ZN(n20560) );
  INV_X1 U23493 ( .A(n20560), .ZN(n20556) );
  AOI22_X1 U23494 ( .A1(n20559), .A2(n20556), .B1(n20967), .B2(n20558), .ZN(
        n20557) );
  NAND2_X1 U23495 ( .A1(n20974), .A2(n20557), .ZN(n20585) );
  OAI22_X1 U23496 ( .A1(n20560), .A2(n20559), .B1(n21028), .B2(n20558), .ZN(
        n20584) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20585), .B1(
        n20968), .B2(n20584), .ZN(n20561) );
  OAI211_X1 U23498 ( .C1(n20980), .C2(n20582), .A(n20562), .B(n20561), .ZN(
        P1_U3057) );
  OAI22_X1 U23499 ( .A1(n20582), .A2(n20985), .B1(n20855), .B2(n20581), .ZN(
        n20563) );
  INV_X1 U23500 ( .A(n20563), .ZN(n20565) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20585), .B1(
        n20981), .B2(n20584), .ZN(n20564) );
  OAI211_X1 U23502 ( .C1(n9983), .C2(n20596), .A(n20565), .B(n20564), .ZN(
        P1_U3058) );
  OAI22_X1 U23503 ( .A1(n20582), .A2(n20991), .B1(n20581), .B2(n20859), .ZN(
        n20566) );
  INV_X1 U23504 ( .A(n20566), .ZN(n20568) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20585), .B1(
        n20986), .B2(n20584), .ZN(n20567) );
  OAI211_X1 U23506 ( .C1(n20906), .C2(n20596), .A(n20568), .B(n20567), .ZN(
        P1_U3059) );
  OAI22_X1 U23507 ( .A1(n20596), .A2(n20910), .B1(n20863), .B2(n20581), .ZN(
        n20569) );
  INV_X1 U23508 ( .A(n20569), .ZN(n20571) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20585), .B1(
        n20992), .B2(n20584), .ZN(n20570) );
  OAI211_X1 U23510 ( .C1(n20997), .C2(n20582), .A(n20571), .B(n20570), .ZN(
        P1_U3060) );
  OAI22_X1 U23511 ( .A1(n20582), .A2(n21002), .B1(n20867), .B2(n20581), .ZN(
        n20572) );
  INV_X1 U23512 ( .A(n20572), .ZN(n20574) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20585), .B1(
        n20998), .B2(n20584), .ZN(n20573) );
  OAI211_X1 U23514 ( .C1(n9979), .C2(n20596), .A(n20574), .B(n20573), .ZN(
        P1_U3061) );
  OAI22_X1 U23515 ( .A1(n20596), .A2(n20918), .B1(n20871), .B2(n20581), .ZN(
        n20575) );
  INV_X1 U23516 ( .A(n20575), .ZN(n20577) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20585), .B1(
        n21003), .B2(n20584), .ZN(n20576) );
  OAI211_X1 U23518 ( .C1(n21008), .C2(n20582), .A(n20577), .B(n20576), .ZN(
        P1_U3062) );
  OAI22_X1 U23519 ( .A1(n20582), .A2(n21014), .B1(n20581), .B2(n20875), .ZN(
        n20578) );
  INV_X1 U23520 ( .A(n20578), .ZN(n20580) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20585), .B1(
        n21009), .B2(n20584), .ZN(n20579) );
  OAI211_X1 U23522 ( .C1(n20922), .C2(n20596), .A(n20580), .B(n20579), .ZN(
        P1_U3063) );
  OAI22_X1 U23523 ( .A1(n20582), .A2(n9977), .B1(n20880), .B2(n20581), .ZN(
        n20583) );
  INV_X1 U23524 ( .A(n20583), .ZN(n20587) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20585), .B1(
        n21016), .B2(n20584), .ZN(n20586) );
  OAI211_X1 U23526 ( .C1(n9981), .C2(n20596), .A(n20587), .B(n20586), .ZN(
        P1_U3064) );
  NAND3_X1 U23527 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20804), .A3(
        n20839), .ZN(n20617) );
  NOR2_X1 U23528 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20617), .ZN(
        n20612) );
  NOR2_X1 U23529 ( .A1(n20845), .A2(n20588), .ZN(n20679) );
  NAND3_X1 U23530 ( .A1(n20679), .A2(n20842), .A3(n20932), .ZN(n20589) );
  OAI21_X1 U23531 ( .B1(n20930), .B2(n20590), .A(n20589), .ZN(n20611) );
  AOI22_X1 U23532 ( .A1(n20969), .A2(n20612), .B1(n20968), .B2(n20611), .ZN(
        n20598) );
  AOI21_X1 U23533 ( .B1(n20596), .B2(n20642), .A(n21220), .ZN(n20591) );
  AOI21_X1 U23534 ( .B1(n20679), .B2(n20932), .A(n20591), .ZN(n20592) );
  NOR2_X1 U23535 ( .A1(n20592), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20595) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20895), .ZN(n20597) );
  OAI211_X1 U23537 ( .C1(n20898), .C2(n20642), .A(n20598), .B(n20597), .ZN(
        P1_U3065) );
  AOI22_X1 U23538 ( .A1(n20982), .A2(n20612), .B1(n20981), .B2(n20611), .ZN(
        n20600) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20899), .ZN(n20599) );
  OAI211_X1 U23540 ( .C1(n9983), .C2(n20642), .A(n20600), .B(n20599), .ZN(
        P1_U3066) );
  AOI22_X1 U23541 ( .A1(n20987), .A2(n20612), .B1(n20986), .B2(n20611), .ZN(
        n20602) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20903), .ZN(n20601) );
  OAI211_X1 U23543 ( .C1(n20906), .C2(n20642), .A(n20602), .B(n20601), .ZN(
        P1_U3067) );
  AOI22_X1 U23544 ( .A1(n20993), .A2(n20612), .B1(n20992), .B2(n20611), .ZN(
        n20604) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20907), .ZN(n20603) );
  OAI211_X1 U23546 ( .C1(n20910), .C2(n20642), .A(n20604), .B(n20603), .ZN(
        P1_U3068) );
  AOI22_X1 U23547 ( .A1(n20999), .A2(n20612), .B1(n20998), .B2(n20611), .ZN(
        n20606) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20911), .ZN(n20605) );
  OAI211_X1 U23549 ( .C1(n9979), .C2(n20642), .A(n20606), .B(n20605), .ZN(
        P1_U3069) );
  AOI22_X1 U23550 ( .A1(n21004), .A2(n20612), .B1(n21003), .B2(n20611), .ZN(
        n20608) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20915), .ZN(n20607) );
  OAI211_X1 U23552 ( .C1(n20918), .C2(n20642), .A(n20608), .B(n20607), .ZN(
        P1_U3070) );
  AOI22_X1 U23553 ( .A1(n21010), .A2(n20612), .B1(n21009), .B2(n20611), .ZN(
        n20610) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n20919), .ZN(n20609) );
  OAI211_X1 U23555 ( .C1(n20922), .C2(n20642), .A(n20610), .B(n20609), .ZN(
        P1_U3071) );
  AOI22_X1 U23556 ( .A1(n21018), .A2(n20612), .B1(n21016), .B2(n20611), .ZN(
        n20616) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20614), .B1(
        n20613), .B2(n9976), .ZN(n20615) );
  OAI211_X1 U23558 ( .C1(n9981), .C2(n20642), .A(n20616), .B(n20615), .ZN(
        P1_U3072) );
  NOR2_X1 U23559 ( .A1(n20889), .A2(n20617), .ZN(n20637) );
  AOI21_X1 U23560 ( .B1(n20679), .B2(n20736), .A(n20637), .ZN(n20618) );
  OAI22_X1 U23561 ( .A1(n20618), .A2(n20967), .B1(n20617), .B2(n21028), .ZN(
        n20636) );
  AOI22_X1 U23562 ( .A1(n20969), .A2(n20637), .B1(n20968), .B2(n20636), .ZN(
        n20622) );
  INV_X1 U23563 ( .A(n20617), .ZN(n20620) );
  OAI211_X1 U23564 ( .C1(n20686), .C2(n21220), .A(n20842), .B(n20618), .ZN(
        n20619) );
  OAI211_X1 U23565 ( .C1(n20842), .C2(n20620), .A(n20974), .B(n20619), .ZN(
        n20639) );
  INV_X1 U23566 ( .A(n20642), .ZN(n20633) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20639), .B1(
        n20633), .B2(n20895), .ZN(n20621) );
  OAI211_X1 U23568 ( .C1(n20898), .C2(n20677), .A(n20622), .B(n20621), .ZN(
        P1_U3073) );
  AOI22_X1 U23569 ( .A1(n20982), .A2(n20637), .B1(n20981), .B2(n20636), .ZN(
        n20624) );
  INV_X1 U23570 ( .A(n20677), .ZN(n20638) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n9982), .ZN(n20623) );
  OAI211_X1 U23572 ( .C1(n20985), .C2(n20642), .A(n20624), .B(n20623), .ZN(
        P1_U3074) );
  AOI22_X1 U23573 ( .A1(n20987), .A2(n20637), .B1(n20986), .B2(n20636), .ZN(
        n20626) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20639), .B1(
        n20633), .B2(n20903), .ZN(n20625) );
  OAI211_X1 U23575 ( .C1(n20906), .C2(n20677), .A(n20626), .B(n20625), .ZN(
        P1_U3075) );
  AOI22_X1 U23576 ( .A1(n20993), .A2(n20637), .B1(n20992), .B2(n20636), .ZN(
        n20628) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20994), .ZN(n20627) );
  OAI211_X1 U23578 ( .C1(n20997), .C2(n20642), .A(n20628), .B(n20627), .ZN(
        P1_U3076) );
  AOI22_X1 U23579 ( .A1(n20999), .A2(n20637), .B1(n20998), .B2(n20636), .ZN(
        n20630) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n9978), .ZN(n20629) );
  OAI211_X1 U23581 ( .C1(n21002), .C2(n20642), .A(n20630), .B(n20629), .ZN(
        P1_U3077) );
  AOI22_X1 U23582 ( .A1(n21004), .A2(n20637), .B1(n21003), .B2(n20636), .ZN(
        n20632) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n21005), .ZN(n20631) );
  OAI211_X1 U23584 ( .C1(n21008), .C2(n20642), .A(n20632), .B(n20631), .ZN(
        P1_U3078) );
  AOI22_X1 U23585 ( .A1(n21010), .A2(n20637), .B1(n21009), .B2(n20636), .ZN(
        n20635) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20639), .B1(
        n20633), .B2(n20919), .ZN(n20634) );
  OAI211_X1 U23587 ( .C1(n20922), .C2(n20677), .A(n20635), .B(n20634), .ZN(
        P1_U3079) );
  AOI22_X1 U23588 ( .A1(n21018), .A2(n20637), .B1(n21016), .B2(n20636), .ZN(
        n20641) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n9980), .ZN(n20640) );
  OAI211_X1 U23590 ( .C1(n9977), .C2(n20642), .A(n20641), .B(n20640), .ZN(
        P1_U3080) );
  INV_X1 U23591 ( .A(n20685), .ZN(n20680) );
  OR2_X1 U23592 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20680), .ZN(
        n20671) );
  OAI22_X1 U23593 ( .A1(n20708), .A2(n20898), .B1(n20840), .B2(n20671), .ZN(
        n20643) );
  INV_X1 U23594 ( .A(n20643), .ZN(n20652) );
  NAND3_X1 U23595 ( .A1(n20708), .A2(n20677), .A3(n20842), .ZN(n20644) );
  NAND2_X1 U23596 ( .A1(n20644), .A2(n20843), .ZN(n20647) );
  NAND2_X1 U23597 ( .A1(n20679), .A2(n20936), .ZN(n20649) );
  AOI22_X1 U23598 ( .A1(n20647), .A2(n20649), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20671), .ZN(n20646) );
  NAND3_X1 U23599 ( .A1(n20940), .A2(n20646), .A3(n20645), .ZN(n20674) );
  INV_X1 U23600 ( .A(n20647), .ZN(n20650) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20674), .B1(
        n20968), .B2(n20673), .ZN(n20651) );
  OAI211_X1 U23602 ( .C1(n20980), .C2(n20677), .A(n20652), .B(n20651), .ZN(
        P1_U3081) );
  OAI22_X1 U23603 ( .A1(n20708), .A2(n9983), .B1(n20855), .B2(n20671), .ZN(
        n20653) );
  INV_X1 U23604 ( .A(n20653), .ZN(n20655) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20674), .B1(
        n20981), .B2(n20673), .ZN(n20654) );
  OAI211_X1 U23606 ( .C1(n20985), .C2(n20677), .A(n20655), .B(n20654), .ZN(
        P1_U3082) );
  OAI22_X1 U23607 ( .A1(n20677), .A2(n20991), .B1(n20859), .B2(n20671), .ZN(
        n20656) );
  INV_X1 U23608 ( .A(n20656), .ZN(n20658) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20674), .B1(
        n20986), .B2(n20673), .ZN(n20657) );
  OAI211_X1 U23610 ( .C1(n20906), .C2(n20708), .A(n20658), .B(n20657), .ZN(
        P1_U3083) );
  OAI22_X1 U23611 ( .A1(n20708), .A2(n20910), .B1(n20863), .B2(n20671), .ZN(
        n20659) );
  INV_X1 U23612 ( .A(n20659), .ZN(n20661) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20674), .B1(
        n20992), .B2(n20673), .ZN(n20660) );
  OAI211_X1 U23614 ( .C1(n20997), .C2(n20677), .A(n20661), .B(n20660), .ZN(
        P1_U3084) );
  OAI22_X1 U23615 ( .A1(n20708), .A2(n9979), .B1(n20867), .B2(n20671), .ZN(
        n20662) );
  INV_X1 U23616 ( .A(n20662), .ZN(n20664) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20674), .B1(
        n20998), .B2(n20673), .ZN(n20663) );
  OAI211_X1 U23618 ( .C1(n21002), .C2(n20677), .A(n20664), .B(n20663), .ZN(
        P1_U3085) );
  OAI22_X1 U23619 ( .A1(n20677), .A2(n21008), .B1(n20871), .B2(n20671), .ZN(
        n20665) );
  INV_X1 U23620 ( .A(n20665), .ZN(n20667) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20674), .B1(
        n21003), .B2(n20673), .ZN(n20666) );
  OAI211_X1 U23622 ( .C1(n20918), .C2(n20708), .A(n20667), .B(n20666), .ZN(
        P1_U3086) );
  OAI22_X1 U23623 ( .A1(n20708), .A2(n20922), .B1(n20875), .B2(n20671), .ZN(
        n20668) );
  INV_X1 U23624 ( .A(n20668), .ZN(n20670) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20674), .B1(
        n21009), .B2(n20673), .ZN(n20669) );
  OAI211_X1 U23626 ( .C1(n21014), .C2(n20677), .A(n20670), .B(n20669), .ZN(
        P1_U3087) );
  OAI22_X1 U23627 ( .A1(n20708), .A2(n9981), .B1(n20880), .B2(n20671), .ZN(
        n20672) );
  INV_X1 U23628 ( .A(n20672), .ZN(n20676) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20674), .B1(
        n21016), .B2(n20673), .ZN(n20675) );
  OAI211_X1 U23630 ( .C1(n9977), .C2(n20677), .A(n20676), .B(n20675), .ZN(
        P1_U3088) );
  INV_X1 U23631 ( .A(n20678), .ZN(n20704) );
  AOI21_X1 U23632 ( .B1(n20679), .B2(n20963), .A(n20704), .ZN(n20682) );
  OAI22_X1 U23633 ( .A1(n20682), .A2(n20967), .B1(n20680), .B2(n21028), .ZN(
        n20703) );
  AOI22_X1 U23634 ( .A1(n20969), .A2(n20704), .B1(n20968), .B2(n20703), .ZN(
        n20688) );
  INV_X1 U23635 ( .A(n20686), .ZN(n20681) );
  OAI21_X1 U23636 ( .B1(n20681), .B2(n20967), .A(n20808), .ZN(n20683) );
  NAND2_X1 U23637 ( .A1(n20683), .A2(n20682), .ZN(n20684) );
  OAI211_X1 U23638 ( .C1(n20685), .C2(n20842), .A(n20974), .B(n20684), .ZN(
        n20705) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20705), .B1(
        n20732), .B2(n20977), .ZN(n20687) );
  OAI211_X1 U23640 ( .C1(n20980), .C2(n20708), .A(n20688), .B(n20687), .ZN(
        P1_U3089) );
  AOI22_X1 U23641 ( .A1(n20982), .A2(n20704), .B1(n20981), .B2(n20703), .ZN(
        n20690) );
  INV_X1 U23642 ( .A(n20708), .ZN(n20697) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20705), .B1(
        n20697), .B2(n20899), .ZN(n20689) );
  OAI211_X1 U23644 ( .C1(n9983), .C2(n20700), .A(n20690), .B(n20689), .ZN(
        P1_U3090) );
  AOI22_X1 U23645 ( .A1(n20987), .A2(n20704), .B1(n20986), .B2(n20703), .ZN(
        n20692) );
  INV_X1 U23646 ( .A(n20906), .ZN(n20988) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20705), .B1(
        n20732), .B2(n20988), .ZN(n20691) );
  OAI211_X1 U23648 ( .C1(n20991), .C2(n20708), .A(n20692), .B(n20691), .ZN(
        P1_U3091) );
  AOI22_X1 U23649 ( .A1(n20993), .A2(n20704), .B1(n20992), .B2(n20703), .ZN(
        n20694) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20705), .B1(
        n20732), .B2(n20994), .ZN(n20693) );
  OAI211_X1 U23651 ( .C1(n20997), .C2(n20708), .A(n20694), .B(n20693), .ZN(
        P1_U3092) );
  AOI22_X1 U23652 ( .A1(n20999), .A2(n20704), .B1(n20998), .B2(n20703), .ZN(
        n20696) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20705), .B1(
        n20697), .B2(n20911), .ZN(n20695) );
  OAI211_X1 U23654 ( .C1(n9979), .C2(n20700), .A(n20696), .B(n20695), .ZN(
        P1_U3093) );
  AOI22_X1 U23655 ( .A1(n21004), .A2(n20704), .B1(n21003), .B2(n20703), .ZN(
        n20699) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20705), .B1(
        n20697), .B2(n20915), .ZN(n20698) );
  OAI211_X1 U23657 ( .C1(n20918), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P1_U3094) );
  AOI22_X1 U23658 ( .A1(n21010), .A2(n20704), .B1(n21009), .B2(n20703), .ZN(
        n20702) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20705), .B1(
        n20732), .B2(n21011), .ZN(n20701) );
  OAI211_X1 U23660 ( .C1(n21014), .C2(n20708), .A(n20702), .B(n20701), .ZN(
        P1_U3095) );
  AOI22_X1 U23661 ( .A1(n21018), .A2(n20704), .B1(n21016), .B2(n20703), .ZN(
        n20707) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20705), .B1(
        n20732), .B2(n9980), .ZN(n20706) );
  OAI211_X1 U23663 ( .C1(n9977), .C2(n20708), .A(n20707), .B(n20706), .ZN(
        P1_U3096) );
  INV_X1 U23664 ( .A(n20838), .ZN(n20709) );
  NAND3_X1 U23665 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20764), .A3(
        n20839), .ZN(n20737) );
  NOR2_X1 U23666 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20737), .ZN(
        n20731) );
  AND2_X1 U23667 ( .A1(n20710), .A2(n20845), .ZN(n20806) );
  AOI21_X1 U23668 ( .B1(n20806), .B2(n20932), .A(n20731), .ZN(n20713) );
  NAND2_X1 U23669 ( .A1(n20711), .A2(n20768), .ZN(n20850) );
  OAI22_X1 U23670 ( .A1(n20713), .A2(n20967), .B1(n20774), .B2(n20850), .ZN(
        n20730) );
  AOI22_X1 U23671 ( .A1(n20969), .A2(n20731), .B1(n20968), .B2(n20730), .ZN(
        n20717) );
  INV_X1 U23672 ( .A(n20762), .ZN(n20712) );
  OAI21_X1 U23673 ( .B1(n20712), .B2(n20732), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20714) );
  NAND2_X1 U23674 ( .A1(n20714), .A2(n20713), .ZN(n20715) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20895), .ZN(n20716) );
  OAI211_X1 U23676 ( .C1(n20898), .C2(n20762), .A(n20717), .B(n20716), .ZN(
        P1_U3097) );
  AOI22_X1 U23677 ( .A1(n20982), .A2(n20731), .B1(n20981), .B2(n20730), .ZN(
        n20719) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20899), .ZN(n20718) );
  OAI211_X1 U23679 ( .C1(n9983), .C2(n20762), .A(n20719), .B(n20718), .ZN(
        P1_U3098) );
  AOI22_X1 U23680 ( .A1(n20987), .A2(n20731), .B1(n20986), .B2(n20730), .ZN(
        n20721) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20903), .ZN(n20720) );
  OAI211_X1 U23682 ( .C1(n20906), .C2(n20762), .A(n20721), .B(n20720), .ZN(
        P1_U3099) );
  AOI22_X1 U23683 ( .A1(n20993), .A2(n20731), .B1(n20992), .B2(n20730), .ZN(
        n20723) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20907), .ZN(n20722) );
  OAI211_X1 U23685 ( .C1(n20910), .C2(n20762), .A(n20723), .B(n20722), .ZN(
        P1_U3100) );
  AOI22_X1 U23686 ( .A1(n20999), .A2(n20731), .B1(n20998), .B2(n20730), .ZN(
        n20725) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20911), .ZN(n20724) );
  OAI211_X1 U23688 ( .C1(n9979), .C2(n20762), .A(n20725), .B(n20724), .ZN(
        P1_U3101) );
  AOI22_X1 U23689 ( .A1(n21004), .A2(n20731), .B1(n21003), .B2(n20730), .ZN(
        n20727) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20915), .ZN(n20726) );
  OAI211_X1 U23691 ( .C1(n20918), .C2(n20762), .A(n20727), .B(n20726), .ZN(
        P1_U3102) );
  AOI22_X1 U23692 ( .A1(n21010), .A2(n20731), .B1(n21009), .B2(n20730), .ZN(
        n20729) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n20919), .ZN(n20728) );
  OAI211_X1 U23694 ( .C1(n20922), .C2(n20762), .A(n20729), .B(n20728), .ZN(
        P1_U3103) );
  AOI22_X1 U23695 ( .A1(n21018), .A2(n20731), .B1(n21016), .B2(n20730), .ZN(
        n20735) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20733), .B1(
        n20732), .B2(n9976), .ZN(n20734) );
  OAI211_X1 U23697 ( .C1(n9981), .C2(n20762), .A(n20735), .B(n20734), .ZN(
        P1_U3104) );
  NOR2_X1 U23698 ( .A1(n20889), .A2(n20737), .ZN(n20758) );
  AOI21_X1 U23699 ( .B1(n20806), .B2(n20736), .A(n20758), .ZN(n20738) );
  OAI22_X1 U23700 ( .A1(n20738), .A2(n20967), .B1(n20737), .B2(n21028), .ZN(
        n20757) );
  AOI22_X1 U23701 ( .A1(n20969), .A2(n20758), .B1(n20968), .B2(n20757), .ZN(
        n20744) );
  INV_X1 U23702 ( .A(n20737), .ZN(n20741) );
  INV_X1 U23703 ( .A(n20815), .ZN(n20739) );
  OAI211_X1 U23704 ( .C1(n20739), .C2(n21220), .A(n20842), .B(n20738), .ZN(
        n20740) );
  OAI211_X1 U23705 ( .C1(n20842), .C2(n20741), .A(n20974), .B(n20740), .ZN(
        n20759) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n20977), .ZN(n20743) );
  OAI211_X1 U23707 ( .C1(n20980), .C2(n20762), .A(n20744), .B(n20743), .ZN(
        P1_U3105) );
  AOI22_X1 U23708 ( .A1(n20982), .A2(n20758), .B1(n20981), .B2(n20757), .ZN(
        n20746) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n9982), .ZN(n20745) );
  OAI211_X1 U23710 ( .C1(n20985), .C2(n20762), .A(n20746), .B(n20745), .ZN(
        P1_U3106) );
  AOI22_X1 U23711 ( .A1(n20987), .A2(n20758), .B1(n20986), .B2(n20757), .ZN(
        n20748) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n20988), .ZN(n20747) );
  OAI211_X1 U23713 ( .C1(n20991), .C2(n20762), .A(n20748), .B(n20747), .ZN(
        P1_U3107) );
  AOI22_X1 U23714 ( .A1(n20993), .A2(n20758), .B1(n20992), .B2(n20757), .ZN(
        n20750) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n20994), .ZN(n20749) );
  OAI211_X1 U23716 ( .C1(n20997), .C2(n20762), .A(n20750), .B(n20749), .ZN(
        P1_U3108) );
  AOI22_X1 U23717 ( .A1(n20999), .A2(n20758), .B1(n20998), .B2(n20757), .ZN(
        n20752) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n9978), .ZN(n20751) );
  OAI211_X1 U23719 ( .C1(n21002), .C2(n20762), .A(n20752), .B(n20751), .ZN(
        P1_U3109) );
  AOI22_X1 U23720 ( .A1(n21004), .A2(n20758), .B1(n21003), .B2(n20757), .ZN(
        n20754) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n21005), .ZN(n20753) );
  OAI211_X1 U23722 ( .C1(n21008), .C2(n20762), .A(n20754), .B(n20753), .ZN(
        P1_U3110) );
  AOI22_X1 U23723 ( .A1(n21010), .A2(n20758), .B1(n21009), .B2(n20757), .ZN(
        n20756) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n21011), .ZN(n20755) );
  OAI211_X1 U23725 ( .C1(n21014), .C2(n20762), .A(n20756), .B(n20755), .ZN(
        P1_U3111) );
  AOI22_X1 U23726 ( .A1(n21018), .A2(n20758), .B1(n21016), .B2(n20757), .ZN(
        n20761) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20759), .B1(
        n20766), .B2(n9980), .ZN(n20760) );
  OAI211_X1 U23728 ( .C1(n9977), .C2(n20762), .A(n20761), .B(n20760), .ZN(
        P1_U3112) );
  INV_X1 U23729 ( .A(n20933), .ZN(n20763) );
  NAND3_X1 U23730 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20764), .ZN(n20807) );
  NOR2_X1 U23731 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20807), .ZN(
        n20769) );
  INV_X1 U23732 ( .A(n20769), .ZN(n20797) );
  OAI22_X1 U23733 ( .A1(n20798), .A2(n20980), .B1(n20797), .B2(n20840), .ZN(
        n20765) );
  INV_X1 U23734 ( .A(n20765), .ZN(n20778) );
  OAI21_X1 U23735 ( .B1(n20834), .B2(n20766), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20767) );
  NAND2_X1 U23736 ( .A1(n20767), .A2(n20842), .ZN(n20776) );
  AND2_X1 U23737 ( .A1(n20806), .A2(n20936), .ZN(n20773) );
  OR2_X1 U23738 ( .A1(n20768), .A2(n20804), .ZN(n20931) );
  NAND2_X1 U23739 ( .A1(n20931), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20939) );
  OAI21_X1 U23740 ( .B1(n20847), .B2(n20769), .A(n20939), .ZN(n20770) );
  INV_X1 U23741 ( .A(n20770), .ZN(n20772) );
  OAI211_X1 U23742 ( .C1(n20776), .C2(n20773), .A(n20772), .B(n20771), .ZN(
        n20801) );
  INV_X1 U23743 ( .A(n20773), .ZN(n20775) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20801), .B1(
        n20968), .B2(n20800), .ZN(n20777) );
  OAI211_X1 U23745 ( .C1(n20898), .C2(n20829), .A(n20778), .B(n20777), .ZN(
        P1_U3113) );
  OAI22_X1 U23746 ( .A1(n20829), .A2(n9983), .B1(n20797), .B2(n20855), .ZN(
        n20779) );
  INV_X1 U23747 ( .A(n20779), .ZN(n20781) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20801), .B1(
        n20981), .B2(n20800), .ZN(n20780) );
  OAI211_X1 U23749 ( .C1(n20985), .C2(n20798), .A(n20781), .B(n20780), .ZN(
        P1_U3114) );
  OAI22_X1 U23750 ( .A1(n20798), .A2(n20991), .B1(n20797), .B2(n20859), .ZN(
        n20782) );
  INV_X1 U23751 ( .A(n20782), .ZN(n20784) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20801), .B1(
        n20986), .B2(n20800), .ZN(n20783) );
  OAI211_X1 U23753 ( .C1(n20906), .C2(n20829), .A(n20784), .B(n20783), .ZN(
        P1_U3115) );
  OAI22_X1 U23754 ( .A1(n20798), .A2(n20997), .B1(n20797), .B2(n20863), .ZN(
        n20785) );
  INV_X1 U23755 ( .A(n20785), .ZN(n20787) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20801), .B1(
        n20992), .B2(n20800), .ZN(n20786) );
  OAI211_X1 U23757 ( .C1(n20910), .C2(n20829), .A(n20787), .B(n20786), .ZN(
        P1_U3116) );
  OAI22_X1 U23758 ( .A1(n20798), .A2(n21002), .B1(n20797), .B2(n20867), .ZN(
        n20788) );
  INV_X1 U23759 ( .A(n20788), .ZN(n20790) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20801), .B1(
        n20998), .B2(n20800), .ZN(n20789) );
  OAI211_X1 U23761 ( .C1(n9979), .C2(n20829), .A(n20790), .B(n20789), .ZN(
        P1_U3117) );
  OAI22_X1 U23762 ( .A1(n20798), .A2(n21008), .B1(n20797), .B2(n20871), .ZN(
        n20791) );
  INV_X1 U23763 ( .A(n20791), .ZN(n20793) );
  AOI22_X1 U23764 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20801), .B1(
        n21003), .B2(n20800), .ZN(n20792) );
  OAI211_X1 U23765 ( .C1(n20918), .C2(n20829), .A(n20793), .B(n20792), .ZN(
        P1_U3118) );
  OAI22_X1 U23766 ( .A1(n20798), .A2(n21014), .B1(n20797), .B2(n20875), .ZN(
        n20794) );
  INV_X1 U23767 ( .A(n20794), .ZN(n20796) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20801), .B1(
        n21009), .B2(n20800), .ZN(n20795) );
  OAI211_X1 U23769 ( .C1(n20922), .C2(n20829), .A(n20796), .B(n20795), .ZN(
        P1_U3119) );
  OAI22_X1 U23770 ( .A1(n20798), .A2(n9977), .B1(n20797), .B2(n20880), .ZN(
        n20799) );
  INV_X1 U23771 ( .A(n20799), .ZN(n20803) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20801), .B1(
        n21016), .B2(n20800), .ZN(n20802) );
  OAI211_X1 U23773 ( .C1(n9981), .C2(n20829), .A(n20803), .B(n20802), .ZN(
        P1_U3120) );
  NOR2_X1 U23774 ( .A1(n20805), .A2(n20804), .ZN(n20833) );
  AOI21_X1 U23775 ( .B1(n20806), .B2(n20963), .A(n20833), .ZN(n20809) );
  OAI22_X1 U23776 ( .A1(n20809), .A2(n20967), .B1(n20807), .B2(n21028), .ZN(
        n20832) );
  AOI22_X1 U23777 ( .A1(n20969), .A2(n20833), .B1(n20968), .B2(n20832), .ZN(
        n20817) );
  INV_X1 U23778 ( .A(n20807), .ZN(n20812) );
  OAI21_X1 U23779 ( .B1(n20815), .B2(n20967), .A(n20808), .ZN(n20810) );
  NAND2_X1 U23780 ( .A1(n20810), .A2(n20809), .ZN(n20811) );
  OAI211_X1 U23781 ( .C1(n20842), .C2(n20812), .A(n20974), .B(n20811), .ZN(
        n20835) );
  INV_X1 U23782 ( .A(n20813), .ZN(n20814) );
  INV_X1 U23783 ( .A(n20886), .ZN(n20826) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20835), .B1(
        n20826), .B2(n20977), .ZN(n20816) );
  OAI211_X1 U23785 ( .C1(n20980), .C2(n20829), .A(n20817), .B(n20816), .ZN(
        P1_U3121) );
  AOI22_X1 U23786 ( .A1(n20982), .A2(n20833), .B1(n20981), .B2(n20832), .ZN(
        n20819) );
  AOI22_X1 U23787 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20899), .ZN(n20818) );
  OAI211_X1 U23788 ( .C1(n9983), .C2(n20886), .A(n20819), .B(n20818), .ZN(
        P1_U3122) );
  AOI22_X1 U23789 ( .A1(n20987), .A2(n20833), .B1(n20986), .B2(n20832), .ZN(
        n20821) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20835), .B1(
        n20826), .B2(n20988), .ZN(n20820) );
  OAI211_X1 U23791 ( .C1(n20991), .C2(n20829), .A(n20821), .B(n20820), .ZN(
        P1_U3123) );
  AOI22_X1 U23792 ( .A1(n20993), .A2(n20833), .B1(n20992), .B2(n20832), .ZN(
        n20823) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20835), .B1(
        n20826), .B2(n20994), .ZN(n20822) );
  OAI211_X1 U23794 ( .C1(n20997), .C2(n20829), .A(n20823), .B(n20822), .ZN(
        P1_U3124) );
  AOI22_X1 U23795 ( .A1(n20999), .A2(n20833), .B1(n20998), .B2(n20832), .ZN(
        n20825) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20835), .B1(
        n20826), .B2(n9978), .ZN(n20824) );
  OAI211_X1 U23797 ( .C1(n21002), .C2(n20829), .A(n20825), .B(n20824), .ZN(
        P1_U3125) );
  AOI22_X1 U23798 ( .A1(n21004), .A2(n20833), .B1(n21003), .B2(n20832), .ZN(
        n20828) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20835), .B1(
        n20826), .B2(n21005), .ZN(n20827) );
  OAI211_X1 U23800 ( .C1(n21008), .C2(n20829), .A(n20828), .B(n20827), .ZN(
        P1_U3126) );
  AOI22_X1 U23801 ( .A1(n21010), .A2(n20833), .B1(n21009), .B2(n20832), .ZN(
        n20831) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20919), .ZN(n20830) );
  OAI211_X1 U23803 ( .C1(n20922), .C2(n20886), .A(n20831), .B(n20830), .ZN(
        P1_U3127) );
  AOI22_X1 U23804 ( .A1(n21018), .A2(n20833), .B1(n21016), .B2(n20832), .ZN(
        n20837) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n9976), .ZN(n20836) );
  OAI211_X1 U23806 ( .C1(n9981), .C2(n20886), .A(n20837), .B(n20836), .ZN(
        P1_U3128) );
  NAND3_X1 U23807 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20839), .ZN(n20892) );
  NOR2_X1 U23808 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20892), .ZN(
        n20848) );
  INV_X1 U23809 ( .A(n20848), .ZN(n20879) );
  OAI22_X1 U23810 ( .A1(n20894), .A2(n20898), .B1(n20840), .B2(n20879), .ZN(
        n20841) );
  INV_X1 U23811 ( .A(n20841), .ZN(n20854) );
  NAND3_X1 U23812 ( .A1(n20886), .A2(n20842), .A3(n20894), .ZN(n20844) );
  NAND2_X1 U23813 ( .A1(n20844), .A2(n20843), .ZN(n20849) );
  NOR2_X1 U23814 ( .A1(n20845), .A2(n10122), .ZN(n20937) );
  NAND2_X1 U23815 ( .A1(n20937), .A2(n20932), .ZN(n20851) );
  AOI22_X1 U23816 ( .A1(n20849), .A2(n20851), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20850), .ZN(n20846) );
  OAI211_X1 U23817 ( .C1(n20848), .C2(n20847), .A(n20940), .B(n20846), .ZN(
        n20883) );
  INV_X1 U23818 ( .A(n20849), .ZN(n20852) );
  OAI22_X1 U23819 ( .A1(n20852), .A2(n20851), .B1(n20850), .B2(n20930), .ZN(
        n20882) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20883), .B1(
        n20968), .B2(n20882), .ZN(n20853) );
  OAI211_X1 U23821 ( .C1(n20980), .C2(n20886), .A(n20854), .B(n20853), .ZN(
        P1_U3129) );
  OAI22_X1 U23822 ( .A1(n20894), .A2(n9983), .B1(n20855), .B2(n20879), .ZN(
        n20856) );
  INV_X1 U23823 ( .A(n20856), .ZN(n20858) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20883), .B1(
        n20981), .B2(n20882), .ZN(n20857) );
  OAI211_X1 U23825 ( .C1(n20985), .C2(n20886), .A(n20858), .B(n20857), .ZN(
        P1_U3130) );
  OAI22_X1 U23826 ( .A1(n20894), .A2(n20906), .B1(n20859), .B2(n20879), .ZN(
        n20860) );
  INV_X1 U23827 ( .A(n20860), .ZN(n20862) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20883), .B1(
        n20986), .B2(n20882), .ZN(n20861) );
  OAI211_X1 U23829 ( .C1(n20991), .C2(n20886), .A(n20862), .B(n20861), .ZN(
        P1_U3131) );
  OAI22_X1 U23830 ( .A1(n20894), .A2(n20910), .B1(n20863), .B2(n20879), .ZN(
        n20864) );
  INV_X1 U23831 ( .A(n20864), .ZN(n20866) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20883), .B1(
        n20992), .B2(n20882), .ZN(n20865) );
  OAI211_X1 U23833 ( .C1(n20997), .C2(n20886), .A(n20866), .B(n20865), .ZN(
        P1_U3132) );
  OAI22_X1 U23834 ( .A1(n20894), .A2(n9979), .B1(n20867), .B2(n20879), .ZN(
        n20868) );
  INV_X1 U23835 ( .A(n20868), .ZN(n20870) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20883), .B1(
        n20998), .B2(n20882), .ZN(n20869) );
  OAI211_X1 U23837 ( .C1(n21002), .C2(n20886), .A(n20870), .B(n20869), .ZN(
        P1_U3133) );
  OAI22_X1 U23838 ( .A1(n20894), .A2(n20918), .B1(n20871), .B2(n20879), .ZN(
        n20872) );
  INV_X1 U23839 ( .A(n20872), .ZN(n20874) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20883), .B1(
        n21003), .B2(n20882), .ZN(n20873) );
  OAI211_X1 U23841 ( .C1(n21008), .C2(n20886), .A(n20874), .B(n20873), .ZN(
        P1_U3134) );
  OAI22_X1 U23842 ( .A1(n20894), .A2(n20922), .B1(n20875), .B2(n20879), .ZN(
        n20876) );
  INV_X1 U23843 ( .A(n20876), .ZN(n20878) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20883), .B1(
        n21009), .B2(n20882), .ZN(n20877) );
  OAI211_X1 U23845 ( .C1(n21014), .C2(n20886), .A(n20878), .B(n20877), .ZN(
        P1_U3135) );
  OAI22_X1 U23846 ( .A1(n20894), .A2(n9981), .B1(n20880), .B2(n20879), .ZN(
        n20881) );
  INV_X1 U23847 ( .A(n20881), .ZN(n20885) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20883), .B1(
        n21016), .B2(n20882), .ZN(n20884) );
  OAI211_X1 U23849 ( .C1(n9977), .C2(n20886), .A(n20885), .B(n20884), .ZN(
        P1_U3136) );
  INV_X1 U23850 ( .A(n20934), .ZN(n20888) );
  NOR2_X1 U23851 ( .A1(n20889), .A2(n20892), .ZN(n20924) );
  INV_X1 U23852 ( .A(n20924), .ZN(n20891) );
  NAND2_X1 U23853 ( .A1(n20937), .A2(n20842), .ZN(n20964) );
  OAI222_X1 U23854 ( .A1(n20891), .A2(n20967), .B1(n21028), .B2(n20892), .C1(
        n20890), .C2(n20964), .ZN(n20923) );
  AOI22_X1 U23855 ( .A1(n20969), .A2(n20924), .B1(n20968), .B2(n20923), .ZN(
        n20897) );
  INV_X1 U23856 ( .A(n20892), .ZN(n20893) );
  OAI21_X1 U23857 ( .B1(n20893), .B2(n20970), .A(n20974), .ZN(n20926) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20895), .ZN(n20896) );
  OAI211_X1 U23859 ( .C1(n20898), .C2(n20962), .A(n20897), .B(n20896), .ZN(
        P1_U3137) );
  AOI22_X1 U23860 ( .A1(n20982), .A2(n20924), .B1(n20981), .B2(n20923), .ZN(
        n20901) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20899), .ZN(n20900) );
  OAI211_X1 U23862 ( .C1(n9983), .C2(n20962), .A(n20901), .B(n20900), .ZN(
        P1_U3138) );
  AOI22_X1 U23863 ( .A1(n20987), .A2(n20924), .B1(n20986), .B2(n20923), .ZN(
        n20905) );
  AOI22_X1 U23864 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20903), .ZN(n20904) );
  OAI211_X1 U23865 ( .C1(n20906), .C2(n20962), .A(n20905), .B(n20904), .ZN(
        P1_U3139) );
  AOI22_X1 U23866 ( .A1(n20993), .A2(n20924), .B1(n20992), .B2(n20923), .ZN(
        n20909) );
  AOI22_X1 U23867 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20907), .ZN(n20908) );
  OAI211_X1 U23868 ( .C1(n20910), .C2(n20962), .A(n20909), .B(n20908), .ZN(
        P1_U3140) );
  AOI22_X1 U23869 ( .A1(n20999), .A2(n20924), .B1(n20998), .B2(n20923), .ZN(
        n20913) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20911), .ZN(n20912) );
  OAI211_X1 U23871 ( .C1(n9979), .C2(n20962), .A(n20913), .B(n20912), .ZN(
        P1_U3141) );
  AOI22_X1 U23872 ( .A1(n21004), .A2(n20924), .B1(n21003), .B2(n20923), .ZN(
        n20917) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20915), .ZN(n20916) );
  OAI211_X1 U23874 ( .C1(n20918), .C2(n20962), .A(n20917), .B(n20916), .ZN(
        P1_U3142) );
  AOI22_X1 U23875 ( .A1(n21010), .A2(n20924), .B1(n21009), .B2(n20923), .ZN(
        n20921) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n20919), .ZN(n20920) );
  OAI211_X1 U23877 ( .C1(n20922), .C2(n20962), .A(n20921), .B(n20920), .ZN(
        P1_U3143) );
  AOI22_X1 U23878 ( .A1(n21018), .A2(n20924), .B1(n21016), .B2(n20923), .ZN(
        n20928) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20926), .B1(
        n20925), .B2(n9976), .ZN(n20927) );
  OAI211_X1 U23880 ( .C1(n9981), .C2(n20962), .A(n20928), .B(n20927), .ZN(
        P1_U3144) );
  NOR2_X1 U23881 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20971), .ZN(
        n20957) );
  OAI22_X1 U23882 ( .A1(n20964), .A2(n20932), .B1(n20931), .B2(n20930), .ZN(
        n20956) );
  AOI22_X1 U23883 ( .A1(n20969), .A2(n20957), .B1(n20968), .B2(n20956), .ZN(
        n20943) );
  AOI21_X1 U23884 ( .B1(n20962), .B2(n21023), .A(n21220), .ZN(n20935) );
  AOI21_X1 U23885 ( .B1(n20937), .B2(n20936), .A(n20935), .ZN(n20938) );
  NOR2_X1 U23886 ( .A1(n20938), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20941) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n20977), .ZN(n20942) );
  OAI211_X1 U23888 ( .C1(n20980), .C2(n20962), .A(n20943), .B(n20942), .ZN(
        P1_U3145) );
  AOI22_X1 U23889 ( .A1(n20982), .A2(n20957), .B1(n20981), .B2(n20956), .ZN(
        n20945) );
  AOI22_X1 U23890 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n9982), .ZN(n20944) );
  OAI211_X1 U23891 ( .C1(n20985), .C2(n20962), .A(n20945), .B(n20944), .ZN(
        P1_U3146) );
  AOI22_X1 U23892 ( .A1(n20987), .A2(n20957), .B1(n20986), .B2(n20956), .ZN(
        n20947) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n20988), .ZN(n20946) );
  OAI211_X1 U23894 ( .C1(n20991), .C2(n20962), .A(n20947), .B(n20946), .ZN(
        P1_U3147) );
  AOI22_X1 U23895 ( .A1(n20993), .A2(n20957), .B1(n20992), .B2(n20956), .ZN(
        n20949) );
  AOI22_X1 U23896 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n20994), .ZN(n20948) );
  OAI211_X1 U23897 ( .C1(n20997), .C2(n20962), .A(n20949), .B(n20948), .ZN(
        P1_U3148) );
  AOI22_X1 U23898 ( .A1(n20999), .A2(n20957), .B1(n20998), .B2(n20956), .ZN(
        n20951) );
  AOI22_X1 U23899 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n9978), .ZN(n20950) );
  OAI211_X1 U23900 ( .C1(n21002), .C2(n20962), .A(n20951), .B(n20950), .ZN(
        P1_U3149) );
  AOI22_X1 U23901 ( .A1(n21004), .A2(n20957), .B1(n21003), .B2(n20956), .ZN(
        n20953) );
  AOI22_X1 U23902 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n21005), .ZN(n20952) );
  OAI211_X1 U23903 ( .C1(n21008), .C2(n20962), .A(n20953), .B(n20952), .ZN(
        P1_U3150) );
  AOI22_X1 U23904 ( .A1(n21010), .A2(n20957), .B1(n21009), .B2(n20956), .ZN(
        n20955) );
  AOI22_X1 U23905 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n21011), .ZN(n20954) );
  OAI211_X1 U23906 ( .C1(n21014), .C2(n20962), .A(n20955), .B(n20954), .ZN(
        P1_U3151) );
  AOI22_X1 U23907 ( .A1(n21018), .A2(n20957), .B1(n21016), .B2(n20956), .ZN(
        n20961) );
  AOI22_X1 U23908 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20959), .B1(
        n20958), .B2(n9980), .ZN(n20960) );
  OAI211_X1 U23909 ( .C1(n9977), .C2(n20962), .A(n20961), .B(n20960), .ZN(
        P1_U3152) );
  INV_X1 U23910 ( .A(n20966), .ZN(n21017) );
  INV_X1 U23911 ( .A(n20963), .ZN(n20965) );
  OAI222_X1 U23912 ( .A1(n20967), .A2(n20966), .B1(n21028), .B2(n20971), .C1(
        n20965), .C2(n20964), .ZN(n21015) );
  AOI22_X1 U23913 ( .A1(n20969), .A2(n21017), .B1(n20968), .B2(n21015), .ZN(
        n20979) );
  INV_X1 U23914 ( .A(n20970), .ZN(n20973) );
  OAI21_X1 U23915 ( .B1(n20973), .B2(n20972), .A(n20971), .ZN(n20975) );
  NAND2_X1 U23916 ( .A1(n20975), .A2(n20974), .ZN(n21020) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n20977), .ZN(n20978) );
  OAI211_X1 U23918 ( .C1(n20980), .C2(n21023), .A(n20979), .B(n20978), .ZN(
        P1_U3153) );
  AOI22_X1 U23919 ( .A1(n20982), .A2(n21017), .B1(n20981), .B2(n21015), .ZN(
        n20984) );
  AOI22_X1 U23920 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n9982), .ZN(n20983) );
  OAI211_X1 U23921 ( .C1(n20985), .C2(n21023), .A(n20984), .B(n20983), .ZN(
        P1_U3154) );
  AOI22_X1 U23922 ( .A1(n20987), .A2(n21017), .B1(n20986), .B2(n21015), .ZN(
        n20990) );
  AOI22_X1 U23923 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n20988), .ZN(n20989) );
  OAI211_X1 U23924 ( .C1(n20991), .C2(n21023), .A(n20990), .B(n20989), .ZN(
        P1_U3155) );
  AOI22_X1 U23925 ( .A1(n20993), .A2(n21017), .B1(n20992), .B2(n21015), .ZN(
        n20996) );
  AOI22_X1 U23926 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n20994), .ZN(n20995) );
  OAI211_X1 U23927 ( .C1(n20997), .C2(n21023), .A(n20996), .B(n20995), .ZN(
        P1_U3156) );
  AOI22_X1 U23928 ( .A1(n20999), .A2(n21017), .B1(n20998), .B2(n21015), .ZN(
        n21001) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n9978), .ZN(n21000) );
  OAI211_X1 U23930 ( .C1(n21002), .C2(n21023), .A(n21001), .B(n21000), .ZN(
        P1_U3157) );
  AOI22_X1 U23931 ( .A1(n21004), .A2(n21017), .B1(n21003), .B2(n21015), .ZN(
        n21007) );
  AOI22_X1 U23932 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21005), .ZN(n21006) );
  OAI211_X1 U23933 ( .C1(n21008), .C2(n21023), .A(n21007), .B(n21006), .ZN(
        P1_U3158) );
  AOI22_X1 U23934 ( .A1(n21010), .A2(n21017), .B1(n21009), .B2(n21015), .ZN(
        n21013) );
  AOI22_X1 U23935 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21011), .ZN(n21012) );
  OAI211_X1 U23936 ( .C1(n21014), .C2(n21023), .A(n21013), .B(n21012), .ZN(
        P1_U3159) );
  AOI22_X1 U23937 ( .A1(n21018), .A2(n21017), .B1(n21016), .B2(n21015), .ZN(
        n21022) );
  AOI22_X1 U23938 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n9980), .ZN(n21021) );
  OAI211_X1 U23939 ( .C1(n9977), .C2(n21023), .A(n21022), .B(n21021), .ZN(
        P1_U3160) );
  NOR2_X1 U23940 ( .A1(n21026), .A2(n21025), .ZN(n21029) );
  OAI21_X1 U23941 ( .B1(n21029), .B2(n21028), .A(n21027), .ZN(P1_U3163) );
  AND2_X1 U23942 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21094), .ZN(
        P1_U3164) );
  AND2_X1 U23943 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21094), .ZN(
        P1_U3165) );
  AND2_X1 U23944 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21094), .ZN(
        P1_U3166) );
  AND2_X1 U23945 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21094), .ZN(
        P1_U3167) );
  AND2_X1 U23946 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21094), .ZN(
        P1_U3168) );
  AND2_X1 U23947 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21094), .ZN(
        P1_U3169) );
  AND2_X1 U23948 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21094), .ZN(
        P1_U3170) );
  AND2_X1 U23949 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21094), .ZN(
        P1_U3171) );
  AND2_X1 U23950 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21094), .ZN(
        P1_U3172) );
  AND2_X1 U23951 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21094), .ZN(
        P1_U3173) );
  AND2_X1 U23952 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21094), .ZN(
        P1_U3174) );
  AND2_X1 U23953 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21094), .ZN(
        P1_U3175) );
  AND2_X1 U23954 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21094), .ZN(
        P1_U3176) );
  AND2_X1 U23955 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21094), .ZN(
        P1_U3177) );
  AND2_X1 U23956 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21094), .ZN(
        P1_U3178) );
  AND2_X1 U23957 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21094), .ZN(
        P1_U3179) );
  AND2_X1 U23958 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21094), .ZN(
        P1_U3180) );
  AND2_X1 U23959 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21094), .ZN(
        P1_U3181) );
  AND2_X1 U23960 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21094), .ZN(
        P1_U3182) );
  AND2_X1 U23961 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21094), .ZN(
        P1_U3183) );
  AND2_X1 U23962 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21094), .ZN(
        P1_U3184) );
  AND2_X1 U23963 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21094), .ZN(
        P1_U3185) );
  AND2_X1 U23964 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21094), .ZN(P1_U3186) );
  AND2_X1 U23965 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21094), .ZN(P1_U3187) );
  AND2_X1 U23966 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21094), .ZN(P1_U3188) );
  AND2_X1 U23967 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21094), .ZN(P1_U3189) );
  AND2_X1 U23968 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21094), .ZN(P1_U3190) );
  AND2_X1 U23969 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21094), .ZN(P1_U3191) );
  AND2_X1 U23970 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21094), .ZN(P1_U3192) );
  AND2_X1 U23971 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21094), .ZN(P1_U3193) );
  NOR2_X1 U23972 ( .A1(NA), .A2(n21327), .ZN(n21035) );
  NOR2_X1 U23973 ( .A1(n21038), .A2(n21327), .ZN(n21032) );
  NOR2_X1 U23974 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21031) );
  OAI22_X1 U23975 ( .A1(n21035), .A2(n21032), .B1(n21031), .B2(n21329), .ZN(
        n21033) );
  NAND2_X1 U23976 ( .A1(n21115), .A2(n21033), .ZN(n21034) );
  OAI221_X1 U23977 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_0__SCAN_IN), .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21043), .A(n21034), .ZN(P1_U3194) );
  AOI21_X1 U23978 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21035), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n21042) );
  AOI221_X1 U23979 ( .B1(NA), .B2(n21036), .C1(n21110), .C2(n21036), .A(n21329), .ZN(n21037) );
  OAI211_X1 U23980 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21327), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n21037), .ZN(n21041) );
  OAI211_X1 U23981 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21039), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21038), .ZN(n21040) );
  OAI211_X1 U23982 ( .C1(n21043), .C2(n21042), .A(n21041), .B(n21040), .ZN(
        P1_U3196) );
  NAND2_X1 U23983 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21116), .ZN(n21087) );
  INV_X1 U23984 ( .A(n21087), .ZN(n21076) );
  NOR2_X1 U23985 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21115), .ZN(n21073) );
  AOI22_X1 U23986 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n21115), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21073), .ZN(n21044) );
  OAI21_X1 U23987 ( .B1(n12958), .B2(n21082), .A(n21044), .ZN(P1_U3197) );
  AOI22_X1 U23988 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21115), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n21073), .ZN(n21045) );
  OAI21_X1 U23989 ( .B1(n12979), .B2(n21082), .A(n21045), .ZN(P1_U3198) );
  INV_X1 U23990 ( .A(n21073), .ZN(n21084) );
  OAI222_X1 U23991 ( .A1(n21087), .A2(n13444), .B1(n21046), .B2(n21064), .C1(
        n21265), .C2(n21084), .ZN(P1_U3199) );
  INV_X1 U23992 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21047) );
  OAI222_X1 U23993 ( .A1(n21084), .A2(n21218), .B1(n21047), .B2(n21064), .C1(
        n21265), .C2(n21082), .ZN(P1_U3200) );
  AOI22_X1 U23994 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21115), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21073), .ZN(n21048) );
  OAI21_X1 U23995 ( .B1(n21218), .B2(n21082), .A(n21048), .ZN(P1_U3201) );
  AOI22_X1 U23996 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21115), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21073), .ZN(n21049) );
  OAI21_X1 U23997 ( .B1(n13697), .B2(n21082), .A(n21049), .ZN(P1_U3202) );
  AOI22_X1 U23998 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21115), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21076), .ZN(n21050) );
  OAI21_X1 U23999 ( .B1(n21052), .B2(n21084), .A(n21050), .ZN(P1_U3203) );
  INV_X1 U24000 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21051) );
  OAI222_X1 U24001 ( .A1(n21087), .A2(n21052), .B1(n21051), .B2(n21064), .C1(
        n21326), .C2(n21084), .ZN(P1_U3204) );
  INV_X1 U24002 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21053) );
  OAI222_X1 U24003 ( .A1(n21082), .A2(n21326), .B1(n21053), .B2(n21064), .C1(
        n21054), .C2(n21084), .ZN(P1_U3205) );
  INV_X1 U24004 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21055) );
  OAI222_X1 U24005 ( .A1(n21084), .A2(n21290), .B1(n21055), .B2(n21064), .C1(
        n21054), .C2(n21082), .ZN(P1_U3206) );
  INV_X1 U24006 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21056) );
  OAI222_X1 U24007 ( .A1(n21084), .A2(n21453), .B1(n21056), .B2(n21064), .C1(
        n21290), .C2(n21082), .ZN(P1_U3207) );
  INV_X1 U24008 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21057) );
  OAI222_X1 U24009 ( .A1(n21087), .A2(n21453), .B1(n21057), .B2(n21064), .C1(
        n21289), .C2(n21084), .ZN(P1_U3208) );
  INV_X1 U24010 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21058) );
  OAI222_X1 U24011 ( .A1(n21084), .A2(n21350), .B1(n21058), .B2(n21064), .C1(
        n21289), .C2(n21082), .ZN(P1_U3209) );
  INV_X1 U24012 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21059) );
  OAI222_X1 U24013 ( .A1(n21082), .A2(n21350), .B1(n21059), .B2(n21064), .C1(
        n21308), .C2(n21084), .ZN(P1_U3210) );
  INV_X1 U24014 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21060) );
  OAI222_X1 U24015 ( .A1(n21087), .A2(n21308), .B1(n21060), .B2(n21116), .C1(
        n21062), .C2(n21084), .ZN(P1_U3211) );
  INV_X1 U24016 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21061) );
  OAI222_X1 U24017 ( .A1(n21087), .A2(n21062), .B1(n21061), .B2(n21116), .C1(
        n21225), .C2(n21084), .ZN(P1_U3212) );
  INV_X1 U24018 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21063) );
  OAI222_X1 U24019 ( .A1(n21084), .A2(n21236), .B1(n21063), .B2(n21116), .C1(
        n21225), .C2(n21082), .ZN(P1_U3213) );
  INV_X1 U24020 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21065) );
  OAI222_X1 U24021 ( .A1(n21084), .A2(n21180), .B1(n21065), .B2(n21064), .C1(
        n21236), .C2(n21087), .ZN(P1_U3214) );
  INV_X1 U24022 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21066) );
  OAI222_X1 U24023 ( .A1(n21087), .A2(n21180), .B1(n21066), .B2(n21116), .C1(
        n21068), .C2(n21084), .ZN(P1_U3215) );
  INV_X1 U24024 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21067) );
  OAI222_X1 U24025 ( .A1(n21087), .A2(n21068), .B1(n21067), .B2(n21116), .C1(
        n21340), .C2(n21084), .ZN(P1_U3216) );
  INV_X1 U24026 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21069) );
  OAI222_X1 U24027 ( .A1(n21084), .A2(n21232), .B1(n21069), .B2(n21116), .C1(
        n21340), .C2(n21082), .ZN(P1_U3217) );
  INV_X1 U24028 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21070) );
  INV_X1 U24029 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21307) );
  OAI222_X1 U24030 ( .A1(n21087), .A2(n21232), .B1(n21070), .B2(n21116), .C1(
        n21307), .C2(n21084), .ZN(P1_U3218) );
  INV_X1 U24031 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21071) );
  OAI222_X1 U24032 ( .A1(n21087), .A2(n21307), .B1(n21071), .B2(n21116), .C1(
        n21447), .C2(n21084), .ZN(P1_U3219) );
  INV_X1 U24033 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21072) );
  OAI222_X1 U24034 ( .A1(n21087), .A2(n21447), .B1(n21072), .B2(n21116), .C1(
        n21075), .C2(n21084), .ZN(P1_U3220) );
  AOI22_X1 U24035 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21073), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21115), .ZN(n21074) );
  OAI21_X1 U24036 ( .B1(n21075), .B2(n21082), .A(n21074), .ZN(P1_U3221) );
  AOI22_X1 U24037 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21076), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21115), .ZN(n21077) );
  OAI21_X1 U24038 ( .B1(n21079), .B2(n21084), .A(n21077), .ZN(P1_U3222) );
  INV_X1 U24039 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21078) );
  OAI222_X1 U24040 ( .A1(n21087), .A2(n21079), .B1(n21078), .B2(n21116), .C1(
        n21081), .C2(n21084), .ZN(P1_U3223) );
  INV_X1 U24041 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21080) );
  OAI222_X1 U24042 ( .A1(n21087), .A2(n21081), .B1(n21080), .B2(n21116), .C1(
        n21353), .C2(n21084), .ZN(P1_U3224) );
  INV_X1 U24043 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21083) );
  OAI222_X1 U24044 ( .A1(n21084), .A2(n21086), .B1(n21083), .B2(n21116), .C1(
        n21353), .C2(n21082), .ZN(P1_U3225) );
  INV_X1 U24045 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21085) );
  OAI222_X1 U24046 ( .A1(n21087), .A2(n21086), .B1(n21085), .B2(n21116), .C1(
        n21197), .C2(n21084), .ZN(P1_U3226) );
  INV_X1 U24047 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U24048 ( .A1(n21116), .A2(n21276), .B1(n21088), .B2(n21115), .ZN(
        P1_U3458) );
  INV_X1 U24049 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21209) );
  INV_X1 U24050 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U24051 ( .A1(n21116), .A2(n21209), .B1(n21089), .B2(n21115), .ZN(
        P1_U3459) );
  INV_X1 U24052 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21090) );
  AOI22_X1 U24053 ( .A1(n21116), .A2(n21282), .B1(n21090), .B2(n21115), .ZN(
        P1_U3460) );
  INV_X1 U24054 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21101) );
  INV_X1 U24055 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21091) );
  AOI22_X1 U24056 ( .A1(n21116), .A2(n21101), .B1(n21091), .B2(n21115), .ZN(
        P1_U3461) );
  INV_X1 U24057 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21097) );
  INV_X1 U24058 ( .A(n21092), .ZN(n21093) );
  AOI21_X1 U24059 ( .B1(n21097), .B2(n21094), .A(n21093), .ZN(P1_U3464) );
  AOI21_X1 U24060 ( .B1(n21094), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21093), 
        .ZN(n21095) );
  INV_X1 U24061 ( .A(n21095), .ZN(P1_U3465) );
  NOR3_X1 U24062 ( .A1(n21097), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n21096) );
  AOI221_X1 U24063 ( .B1(n21098), .B2(n21097), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n21096), .ZN(n21099) );
  INV_X1 U24064 ( .A(n21103), .ZN(n21100) );
  AOI22_X1 U24065 ( .A1(n21103), .A2(n21099), .B1(n21209), .B2(n21100), .ZN(
        P1_U3481) );
  NOR2_X1 U24066 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21102) );
  AOI22_X1 U24067 ( .A1(n21103), .A2(n21102), .B1(n21101), .B2(n21100), .ZN(
        P1_U3482) );
  AOI22_X1 U24068 ( .A1(n21116), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21223), 
        .B2(n21115), .ZN(P1_U3483) );
  OAI21_X1 U24069 ( .B1(n21104), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21106) );
  OAI22_X1 U24070 ( .A1(n21107), .A2(n21106), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21105), .ZN(n21114) );
  AOI211_X1 U24071 ( .C1(n21111), .C2(n21110), .A(n21109), .B(n21108), .ZN(
        n21113) );
  NAND2_X1 U24072 ( .A1(n21113), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21112) );
  OAI21_X1 U24073 ( .B1(n21114), .B2(n21113), .A(n21112), .ZN(P1_U3485) );
  AOI22_X1 U24074 ( .A1(n21116), .A2(n21324), .B1(n21465), .B2(n21115), .ZN(
        P1_U3486) );
  XOR2_X1 U24075 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_g39), .Z(n21123) );
  AOI22_X1 U24076 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .ZN(n21117) );
  OAI221_X1 U24077 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(n21117), .ZN(n21122)
         );
  AOI22_X1 U24078 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .ZN(n21118) );
  OAI221_X1 U24079 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_EBX_REG_21__SCAN_IN), .C2(keyinput_g94), .A(n21118), .ZN(n21121) );
  AOI22_X1 U24080 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(DATAI_20_), .B2(
        keyinput_g12), .ZN(n21119) );
  OAI221_X1 U24081 ( .B1(DATAI_2_), .B2(keyinput_g30), .C1(DATAI_20_), .C2(
        keyinput_g12), .A(n21119), .ZN(n21120) );
  NOR4_X1 U24082 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21151) );
  AOI22_X1 U24083 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .ZN(n21124) );
  OAI221_X1 U24084 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        P1_FLUSH_REG_SCAN_IN), .C2(keyinput_g46), .A(n21124), .ZN(n21131) );
  AOI22_X1 U24085 ( .A1(NA), .A2(keyinput_g34), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(keyinput_g93), .ZN(n21125) );
  OAI221_X1 U24086 ( .B1(NA), .B2(keyinput_g34), .C1(P1_EBX_REG_22__SCAN_IN), 
        .C2(keyinput_g93), .A(n21125), .ZN(n21130) );
  AOI22_X1 U24087 ( .A1(READY2), .A2(keyinput_g37), .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_g76), .ZN(n21126) );
  OAI221_X1 U24088 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput_g76), .A(n21126), .ZN(n21129) );
  AOI22_X1 U24089 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_g104), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(keyinput_g99), .ZN(n21127) );
  OAI221_X1 U24090 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .C1(
        P1_EBX_REG_16__SCAN_IN), .C2(keyinput_g99), .A(n21127), .ZN(n21128) );
  NOR4_X1 U24091 ( .A1(n21131), .A2(n21130), .A3(n21129), .A4(n21128), .ZN(
        n21150) );
  AOI22_X1 U24092 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_g84), .ZN(n21132) );
  OAI221_X1 U24093 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_g84), .A(n21132), .ZN(n21139) );
  AOI22_X1 U24094 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_g87), .ZN(n21133) );
  OAI221_X1 U24095 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(P1_EBX_REG_28__SCAN_IN), .C2(keyinput_g87), .A(n21133), .ZN(n21138) );
  AOI22_X1 U24096 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_g53), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_g115), .ZN(n21134) );
  OAI221_X1 U24097 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_g53), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_g115), .A(n21134), .ZN(n21137) );
  AOI22_X1 U24098 ( .A1(DATAI_24_), .A2(keyinput_g8), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(keyinput_g67), .ZN(n21135) );
  OAI221_X1 U24099 ( .B1(DATAI_24_), .B2(keyinput_g8), .C1(
        P1_REIP_REG_16__SCAN_IN), .C2(keyinput_g67), .A(n21135), .ZN(n21136)
         );
  NOR4_X1 U24100 ( .A1(n21139), .A2(n21138), .A3(n21137), .A4(n21136), .ZN(
        n21149) );
  AOI22_X1 U24101 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_EBX_REG_9__SCAN_IN), .B2(keyinput_g106), .ZN(n21140) );
  OAI221_X1 U24102 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_EBX_REG_9__SCAN_IN), .C2(keyinput_g106), .A(n21140), .ZN(n21147) );
  AOI22_X1 U24103 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput_g92), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_g90), .ZN(n21141) );
  OAI221_X1 U24104 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_g92), .C1(
        P1_EBX_REG_25__SCAN_IN), .C2(keyinput_g90), .A(n21141), .ZN(n21146) );
  AOI22_X1 U24105 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(keyinput_g102), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(keyinput_g96), .ZN(n21142) );
  OAI221_X1 U24106 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(keyinput_g102), .C1(
        P1_EBX_REG_19__SCAN_IN), .C2(keyinput_g96), .A(n21142), .ZN(n21145) );
  AOI22_X1 U24107 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        READY1), .B2(keyinput_g36), .ZN(n21143) );
  OAI221_X1 U24108 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        READY1), .C2(keyinput_g36), .A(n21143), .ZN(n21144) );
  NOR4_X1 U24109 ( .A1(n21147), .A2(n21146), .A3(n21145), .A4(n21144), .ZN(
        n21148) );
  NAND4_X1 U24110 ( .A1(n21151), .A2(n21150), .A3(n21149), .A4(n21148), .ZN(
        n21302) );
  AOI22_X1 U24111 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_g86), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_g121), .ZN(n21152) );
  OAI221_X1 U24112 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_g121), .A(n21152), .ZN(n21159)
         );
  AOI22_X1 U24113 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(keyinput_g82), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n21153) );
  OAI221_X1 U24114 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(keyinput_g82), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n21153), .ZN(n21158)
         );
  AOI22_X1 U24115 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput_g120), .ZN(n21154) );
  OAI221_X1 U24116 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_g120), .A(n21154), .ZN(n21157)
         );
  AOI22_X1 U24117 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .ZN(n21155) );
  OAI221_X1 U24118 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(
        P1_EBX_REG_14__SCAN_IN), .C2(keyinput_g101), .A(n21155), .ZN(n21156)
         );
  NOR4_X1 U24119 ( .A1(n21159), .A2(n21158), .A3(n21157), .A4(n21156), .ZN(
        n21189) );
  AOI22_X1 U24120 ( .A1(DATAI_16_), .A2(keyinput_g16), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_g118), .ZN(n21160) );
  OAI221_X1 U24121 ( .B1(DATAI_16_), .B2(keyinput_g16), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_g118), .A(n21160), .ZN(n21167)
         );
  AOI22_X1 U24122 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21161) );
  OAI221_X1 U24123 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21161), .ZN(n21166)
         );
  AOI22_X1 U24124 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n21162) );
  OAI221_X1 U24125 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n21162), .ZN(n21165)
         );
  AOI22_X1 U24126 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_g58), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(keyinput_g107), .ZN(n21163) );
  OAI221_X1 U24127 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .C1(
        P1_EBX_REG_8__SCAN_IN), .C2(keyinput_g107), .A(n21163), .ZN(n21164) );
  NOR4_X1 U24128 ( .A1(n21167), .A2(n21166), .A3(n21165), .A4(n21164), .ZN(
        n21188) );
  AOI22_X1 U24129 ( .A1(DATAI_4_), .A2(keyinput_g28), .B1(DATAI_21_), .B2(
        keyinput_g11), .ZN(n21168) );
  OAI221_X1 U24130 ( .B1(DATAI_4_), .B2(keyinput_g28), .C1(DATAI_21_), .C2(
        keyinput_g11), .A(n21168), .ZN(n21175) );
  AOI22_X1 U24131 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(keyinput_g73), .ZN(n21169) );
  OAI221_X1 U24132 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(keyinput_g73), .A(n21169), .ZN(n21174)
         );
  AOI22_X1 U24133 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_g77), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_g117), .ZN(n21170) );
  OAI221_X1 U24134 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_g77), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_g117), .A(n21170), .ZN(n21173)
         );
  AOI22_X1 U24135 ( .A1(DATAI_31_), .A2(keyinput_g1), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput_g95), .ZN(n21171) );
  OAI221_X1 U24136 ( .B1(DATAI_31_), .B2(keyinput_g1), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput_g95), .A(n21171), .ZN(n21172) );
  NOR4_X1 U24137 ( .A1(n21175), .A2(n21174), .A3(n21173), .A4(n21172), .ZN(
        n21187) );
  AOI22_X1 U24138 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(DATAI_10_), .B2(
        keyinput_g22), .ZN(n21176) );
  OAI221_X1 U24139 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(DATAI_10_), .C2(
        keyinput_g22), .A(n21176), .ZN(n21185) );
  AOI22_X1 U24140 ( .A1(DATAI_18_), .A2(keyinput_g14), .B1(DATAI_23_), .B2(
        keyinput_g9), .ZN(n21177) );
  OAI221_X1 U24141 ( .B1(DATAI_18_), .B2(keyinput_g14), .C1(DATAI_23_), .C2(
        keyinput_g9), .A(n21177), .ZN(n21184) );
  AOI22_X1 U24142 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .ZN(n21178) );
  OAI221_X1 U24143 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        P1_EBX_REG_27__SCAN_IN), .C2(keyinput_g88), .A(n21178), .ZN(n21183) );
  INV_X1 U24144 ( .A(DATAI_0_), .ZN(n21181) );
  AOI22_X1 U24145 ( .A1(n21181), .A2(keyinput_g32), .B1(n21180), .B2(
        keyinput_g64), .ZN(n21179) );
  OAI221_X1 U24146 ( .B1(n21181), .B2(keyinput_g32), .C1(n21180), .C2(
        keyinput_g64), .A(n21179), .ZN(n21182) );
  NOR4_X1 U24147 ( .A1(n21185), .A2(n21184), .A3(n21183), .A4(n21182), .ZN(
        n21186) );
  NAND4_X1 U24148 ( .A1(n21189), .A2(n21188), .A3(n21187), .A4(n21186), .ZN(
        n21301) );
  AOI22_X1 U24149 ( .A1(n21192), .A2(keyinput_g85), .B1(n21191), .B2(
        keyinput_g112), .ZN(n21190) );
  OAI221_X1 U24150 ( .B1(n21192), .B2(keyinput_g85), .C1(n21191), .C2(
        keyinput_g112), .A(n21190), .ZN(n21201) );
  AOI22_X1 U24151 ( .A1(n21350), .A2(keyinput_g69), .B1(n21447), .B2(
        keyinput_g59), .ZN(n21193) );
  OAI221_X1 U24152 ( .B1(n21350), .B2(keyinput_g69), .C1(n21447), .C2(
        keyinput_g59), .A(n21193), .ZN(n21200) );
  AOI22_X1 U24153 ( .A1(n21195), .A2(keyinput_g21), .B1(n21482), .B2(
        keyinput_g103), .ZN(n21194) );
  OAI221_X1 U24154 ( .B1(n21195), .B2(keyinput_g21), .C1(n21482), .C2(
        keyinput_g103), .A(n21194), .ZN(n21199) );
  INV_X1 U24155 ( .A(DATAI_19_), .ZN(n21349) );
  AOI22_X1 U24156 ( .A1(n21349), .A2(keyinput_g13), .B1(n21197), .B2(
        keyinput_g52), .ZN(n21196) );
  OAI221_X1 U24157 ( .B1(n21349), .B2(keyinput_g13), .C1(n21197), .C2(
        keyinput_g52), .A(n21196), .ZN(n21198) );
  NOR4_X1 U24158 ( .A1(n21201), .A2(n21200), .A3(n21199), .A4(n21198), .ZN(
        n21246) );
  INV_X1 U24159 ( .A(DATAI_6_), .ZN(n21204) );
  AOI22_X1 U24160 ( .A1(n21204), .A2(keyinput_g26), .B1(n21203), .B2(
        keyinput_g25), .ZN(n21202) );
  OAI221_X1 U24161 ( .B1(n21204), .B2(keyinput_g26), .C1(n21203), .C2(
        keyinput_g25), .A(n21202), .ZN(n21216) );
  INV_X1 U24162 ( .A(BS16), .ZN(n21206) );
  AOI22_X1 U24163 ( .A1(n21206), .A2(keyinput_g35), .B1(n21313), .B2(
        keyinput_g100), .ZN(n21205) );
  OAI221_X1 U24164 ( .B1(n21206), .B2(keyinput_g35), .C1(n21313), .C2(
        keyinput_g100), .A(n21205), .ZN(n21215) );
  AOI22_X1 U24165 ( .A1(n21209), .A2(keyinput_g50), .B1(n21208), .B2(
        keyinput_g20), .ZN(n21207) );
  OAI221_X1 U24166 ( .B1(n21209), .B2(keyinput_g50), .C1(n21208), .C2(
        keyinput_g20), .A(n21207), .ZN(n21214) );
  AOI22_X1 U24167 ( .A1(n21212), .A2(keyinput_g6), .B1(n21211), .B2(
        keyinput_g2), .ZN(n21210) );
  OAI221_X1 U24168 ( .B1(n21212), .B2(keyinput_g6), .C1(n21211), .C2(
        keyinput_g2), .A(n21210), .ZN(n21213) );
  NOR4_X1 U24169 ( .A1(n21216), .A2(n21215), .A3(n21214), .A4(n21213), .ZN(
        n21245) );
  AOI22_X1 U24170 ( .A1(n12979), .A2(keyinput_g81), .B1(keyinput_g78), .B2(
        n21218), .ZN(n21217) );
  OAI221_X1 U24171 ( .B1(n12979), .B2(keyinput_g81), .C1(n21218), .C2(
        keyinput_g78), .A(n21217), .ZN(n21230) );
  AOI22_X1 U24172 ( .A1(n21221), .A2(keyinput_g38), .B1(n21220), .B2(
        keyinput_g44), .ZN(n21219) );
  OAI221_X1 U24173 ( .B1(n21221), .B2(keyinput_g38), .C1(n21220), .C2(
        keyinput_g44), .A(n21219), .ZN(n21229) );
  INV_X1 U24174 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21356) );
  AOI22_X1 U24175 ( .A1(n21223), .A2(keyinput_g47), .B1(n21356), .B2(
        keyinput_g116), .ZN(n21222) );
  OAI221_X1 U24176 ( .B1(n21223), .B2(keyinput_g47), .C1(n21356), .C2(
        keyinput_g116), .A(n21222), .ZN(n21228) );
  AOI22_X1 U24177 ( .A1(n21226), .A2(keyinput_g126), .B1(keyinput_g66), .B2(
        n21225), .ZN(n21224) );
  OAI221_X1 U24178 ( .B1(n21226), .B2(keyinput_g126), .C1(n21225), .C2(
        keyinput_g66), .A(n21224), .ZN(n21227) );
  NOR4_X1 U24179 ( .A1(n21230), .A2(n21229), .A3(n21228), .A4(n21227), .ZN(
        n21244) );
  AOI22_X1 U24180 ( .A1(n21233), .A2(keyinput_g113), .B1(keyinput_g61), .B2(
        n21232), .ZN(n21231) );
  OAI221_X1 U24181 ( .B1(n21233), .B2(keyinput_g113), .C1(n21232), .C2(
        keyinput_g61), .A(n21231), .ZN(n21242) );
  INV_X1 U24182 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21355) );
  AOI22_X1 U24183 ( .A1(n21450), .A2(keyinput_g110), .B1(keyinput_g40), .B2(
        n21355), .ZN(n21234) );
  OAI221_X1 U24184 ( .B1(n21450), .B2(keyinput_g110), .C1(n21355), .C2(
        keyinput_g40), .A(n21234), .ZN(n21241) );
  AOI22_X1 U24185 ( .A1(n21236), .A2(keyinput_g65), .B1(n21340), .B2(
        keyinput_g62), .ZN(n21235) );
  OAI221_X1 U24186 ( .B1(n21236), .B2(keyinput_g65), .C1(n21340), .C2(
        keyinput_g62), .A(n21235), .ZN(n21240) );
  AOI22_X1 U24187 ( .A1(n21238), .A2(keyinput_g124), .B1(keyinput_g122), .B2(
        n21466), .ZN(n21237) );
  OAI221_X1 U24188 ( .B1(n21238), .B2(keyinput_g124), .C1(n21466), .C2(
        keyinput_g122), .A(n21237), .ZN(n21239) );
  NOR4_X1 U24189 ( .A1(n21242), .A2(n21241), .A3(n21240), .A4(n21239), .ZN(
        n21243) );
  NAND4_X1 U24190 ( .A1(n21246), .A2(n21245), .A3(n21244), .A4(n21243), .ZN(
        n21300) );
  AOI22_X1 U24191 ( .A1(n12796), .A2(keyinput_g83), .B1(n21248), .B2(
        keyinput_g109), .ZN(n21247) );
  OAI221_X1 U24192 ( .B1(n12796), .B2(keyinput_g83), .C1(n21248), .C2(
        keyinput_g109), .A(n21247), .ZN(n21257) );
  INV_X1 U24193 ( .A(DATAI_1_), .ZN(n21449) );
  AOI22_X1 U24194 ( .A1(n21449), .A2(keyinput_g31), .B1(n13444), .B2(
        keyinput_g80), .ZN(n21249) );
  OAI221_X1 U24195 ( .B1(n21449), .B2(keyinput_g31), .C1(n13444), .C2(
        keyinput_g80), .A(n21249), .ZN(n21256) );
  AOI22_X1 U24196 ( .A1(n21326), .A2(keyinput_g74), .B1(n21459), .B2(
        keyinput_g119), .ZN(n21250) );
  OAI221_X1 U24197 ( .B1(n21326), .B2(keyinput_g74), .C1(n21459), .C2(
        keyinput_g119), .A(n21250), .ZN(n21255) );
  AOI22_X1 U24198 ( .A1(n21253), .A2(keyinput_g18), .B1(keyinput_g45), .B2(
        n21252), .ZN(n21251) );
  OAI221_X1 U24199 ( .B1(n21253), .B2(keyinput_g18), .C1(n21252), .C2(
        keyinput_g45), .A(n21251), .ZN(n21254) );
  NOR4_X1 U24200 ( .A1(n21257), .A2(n21256), .A3(n21255), .A4(n21254), .ZN(
        n21298) );
  AOI22_X1 U24201 ( .A1(n21260), .A2(keyinput_g89), .B1(keyinput_g111), .B2(
        n21259), .ZN(n21258) );
  OAI221_X1 U24202 ( .B1(n21260), .B2(keyinput_g89), .C1(n21259), .C2(
        keyinput_g111), .A(n21258), .ZN(n21269) );
  INV_X1 U24203 ( .A(DATAI_5_), .ZN(n21460) );
  AOI22_X1 U24204 ( .A1(n21327), .A2(keyinput_g43), .B1(n21460), .B2(
        keyinput_g27), .ZN(n21261) );
  OAI221_X1 U24205 ( .B1(n21327), .B2(keyinput_g43), .C1(n21460), .C2(
        keyinput_g27), .A(n21261), .ZN(n21268) );
  AOI22_X1 U24206 ( .A1(n21263), .A2(keyinput_g7), .B1(keyinput_g33), .B2(
        n21329), .ZN(n21262) );
  OAI221_X1 U24207 ( .B1(n21263), .B2(keyinput_g7), .C1(n21329), .C2(
        keyinput_g33), .A(n21262), .ZN(n21267) );
  AOI22_X1 U24208 ( .A1(n21358), .A2(keyinput_g19), .B1(n21265), .B2(
        keyinput_g79), .ZN(n21264) );
  OAI221_X1 U24209 ( .B1(n21358), .B2(keyinput_g19), .C1(n21265), .C2(
        keyinput_g79), .A(n21264), .ZN(n21266) );
  NOR4_X1 U24210 ( .A1(n21269), .A2(n21268), .A3(n21267), .A4(n21266), .ZN(
        n21297) );
  AOI22_X1 U24211 ( .A1(n21479), .A2(keyinput_g91), .B1(keyinput_g68), .B2(
        n21308), .ZN(n21270) );
  OAI221_X1 U24212 ( .B1(n21479), .B2(keyinput_g91), .C1(n21308), .C2(
        keyinput_g68), .A(n21270), .ZN(n21280) );
  AOI22_X1 U24213 ( .A1(n21272), .A2(keyinput_g114), .B1(n21478), .B2(
        keyinput_g123), .ZN(n21271) );
  OAI221_X1 U24214 ( .B1(n21272), .B2(keyinput_g114), .C1(n21478), .C2(
        keyinput_g123), .A(n21271), .ZN(n21279) );
  AOI22_X1 U24215 ( .A1(n21485), .A2(keyinput_g98), .B1(keyinput_g3), .B2(
        n21274), .ZN(n21273) );
  OAI221_X1 U24216 ( .B1(n21485), .B2(keyinput_g98), .C1(n21274), .C2(
        keyinput_g3), .A(n21273), .ZN(n21278) );
  AOI22_X1 U24217 ( .A1(n21453), .A2(keyinput_g71), .B1(keyinput_g51), .B2(
        n21276), .ZN(n21275) );
  OAI221_X1 U24218 ( .B1(n21453), .B2(keyinput_g71), .C1(n21276), .C2(
        keyinput_g51), .A(n21275), .ZN(n21277) );
  NOR4_X1 U24219 ( .A1(n21280), .A2(n21279), .A3(n21278), .A4(n21277), .ZN(
        n21296) );
  AOI22_X1 U24220 ( .A1(n21282), .A2(keyinput_g49), .B1(n21337), .B2(
        keyinput_g108), .ZN(n21281) );
  OAI221_X1 U24221 ( .B1(n21282), .B2(keyinput_g49), .C1(n21337), .C2(
        keyinput_g108), .A(n21281), .ZN(n21294) );
  INV_X1 U24222 ( .A(DATAI_8_), .ZN(n21320) );
  AOI22_X1 U24223 ( .A1(n21284), .A2(keyinput_g4), .B1(keyinput_g24), .B2(
        n21320), .ZN(n21283) );
  OAI221_X1 U24224 ( .B1(n21284), .B2(keyinput_g4), .C1(n21320), .C2(
        keyinput_g24), .A(n21283), .ZN(n21293) );
  AOI22_X1 U24225 ( .A1(n21287), .A2(keyinput_g5), .B1(n21286), .B2(
        keyinput_g97), .ZN(n21285) );
  OAI221_X1 U24226 ( .B1(n21287), .B2(keyinput_g5), .C1(n21286), .C2(
        keyinput_g97), .A(n21285), .ZN(n21292) );
  AOI22_X1 U24227 ( .A1(n21290), .A2(keyinput_g72), .B1(n21289), .B2(
        keyinput_g70), .ZN(n21288) );
  OAI221_X1 U24228 ( .B1(n21290), .B2(keyinput_g72), .C1(n21289), .C2(
        keyinput_g70), .A(n21288), .ZN(n21291) );
  NOR4_X1 U24229 ( .A1(n21294), .A2(n21293), .A3(n21292), .A4(n21291), .ZN(
        n21295) );
  NAND4_X1 U24230 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21299) );
  NOR4_X1 U24231 ( .A1(n21302), .A2(n21301), .A3(n21300), .A4(n21299), .ZN(
        n21506) );
  INV_X1 U24232 ( .A(keyinput_f105), .ZN(n21503) );
  INV_X1 U24233 ( .A(READY2), .ZN(n21304) );
  AOI22_X1 U24234 ( .A1(n21305), .A2(keyinput_f107), .B1(keyinput_f37), .B2(
        n21304), .ZN(n21303) );
  OAI221_X1 U24235 ( .B1(n21305), .B2(keyinput_f107), .C1(n21304), .C2(
        keyinput_f37), .A(n21303), .ZN(n21318) );
  AOI22_X1 U24236 ( .A1(n21308), .A2(keyinput_f68), .B1(n21307), .B2(
        keyinput_f60), .ZN(n21306) );
  OAI221_X1 U24237 ( .B1(n21308), .B2(keyinput_f68), .C1(n21307), .C2(
        keyinput_f60), .A(n21306), .ZN(n21317) );
  INV_X1 U24238 ( .A(keyinput_f48), .ZN(n21310) );
  AOI22_X1 U24239 ( .A1(n21311), .A2(keyinput_f46), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n21310), .ZN(n21309) );
  OAI221_X1 U24240 ( .B1(n21311), .B2(keyinput_f46), .C1(n21310), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21309), .ZN(n21316) );
  AOI22_X1 U24241 ( .A1(n21314), .A2(keyinput_f115), .B1(n21313), .B2(
        keyinput_f100), .ZN(n21312) );
  OAI221_X1 U24242 ( .B1(n21314), .B2(keyinput_f115), .C1(n21313), .C2(
        keyinput_f100), .A(n21312), .ZN(n21315) );
  NOR4_X1 U24243 ( .A1(n21318), .A2(n21317), .A3(n21316), .A4(n21315), .ZN(
        n21501) );
  INV_X1 U24244 ( .A(DATAI_16_), .ZN(n21321) );
  AOI22_X1 U24245 ( .A1(n21321), .A2(keyinput_f16), .B1(n21320), .B2(
        keyinput_f24), .ZN(n21319) );
  OAI221_X1 U24246 ( .B1(n21321), .B2(keyinput_f16), .C1(n21320), .C2(
        keyinput_f24), .A(n21319), .ZN(n21334) );
  AOI22_X1 U24247 ( .A1(n21324), .A2(keyinput_f0), .B1(n21323), .B2(
        keyinput_f127), .ZN(n21322) );
  OAI221_X1 U24248 ( .B1(n21324), .B2(keyinput_f0), .C1(n21323), .C2(
        keyinput_f127), .A(n21322), .ZN(n21333) );
  AOI22_X1 U24249 ( .A1(n21327), .A2(keyinput_f43), .B1(n21326), .B2(
        keyinput_f74), .ZN(n21325) );
  OAI221_X1 U24250 ( .B1(n21327), .B2(keyinput_f43), .C1(n21326), .C2(
        keyinput_f74), .A(n21325), .ZN(n21332) );
  INV_X1 U24251 ( .A(DATAI_17_), .ZN(n21330) );
  AOI22_X1 U24252 ( .A1(n21330), .A2(keyinput_f15), .B1(keyinput_f33), .B2(
        n21329), .ZN(n21328) );
  OAI221_X1 U24253 ( .B1(n21330), .B2(keyinput_f15), .C1(n21329), .C2(
        keyinput_f33), .A(n21328), .ZN(n21331) );
  NOR4_X1 U24254 ( .A1(n21334), .A2(n21333), .A3(n21332), .A4(n21331), .ZN(
        n21500) );
  AOI22_X1 U24255 ( .A1(n21337), .A2(keyinput_f108), .B1(n21336), .B2(
        keyinput_f92), .ZN(n21335) );
  OAI221_X1 U24256 ( .B1(n21337), .B2(keyinput_f108), .C1(n21336), .C2(
        keyinput_f92), .A(n21335), .ZN(n21366) );
  INV_X1 U24257 ( .A(DATAI_23_), .ZN(n21339) );
  AOI22_X1 U24258 ( .A1(n21340), .A2(keyinput_f62), .B1(keyinput_f9), .B2(
        n21339), .ZN(n21338) );
  OAI221_X1 U24259 ( .B1(n21340), .B2(keyinput_f62), .C1(n21339), .C2(
        keyinput_f9), .A(n21338), .ZN(n21365) );
  XOR2_X1 U24260 ( .A(READY1), .B(keyinput_f36), .Z(n21345) );
  INV_X1 U24261 ( .A(keyinput_f51), .ZN(n21342) );
  AOI22_X1 U24262 ( .A1(n21343), .A2(keyinput_f23), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n21342), .ZN(n21341) );
  OAI221_X1 U24263 ( .B1(n21343), .B2(keyinput_f23), .C1(n21342), .C2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A(n21341), .ZN(n21344) );
  AOI211_X1 U24264 ( .C1(n21347), .C2(keyinput_f42), .A(n21345), .B(n21344), 
        .ZN(n21346) );
  OAI21_X1 U24265 ( .B1(n21347), .B2(keyinput_f42), .A(n21346), .ZN(n21364) );
  OAI22_X1 U24266 ( .A1(n21350), .A2(keyinput_f69), .B1(n21349), .B2(
        keyinput_f13), .ZN(n21348) );
  AOI221_X1 U24267 ( .B1(n21350), .B2(keyinput_f69), .C1(keyinput_f13), .C2(
        n21349), .A(n21348), .ZN(n21362) );
  INV_X1 U24268 ( .A(DATAI_20_), .ZN(n21352) );
  OAI22_X1 U24269 ( .A1(n21353), .A2(keyinput_f54), .B1(n21352), .B2(
        keyinput_f12), .ZN(n21351) );
  AOI221_X1 U24270 ( .B1(n21353), .B2(keyinput_f54), .C1(keyinput_f12), .C2(
        n21352), .A(n21351), .ZN(n21361) );
  OAI22_X1 U24271 ( .A1(n21356), .A2(keyinput_f116), .B1(n21355), .B2(
        keyinput_f40), .ZN(n21354) );
  AOI221_X1 U24272 ( .B1(n21356), .B2(keyinput_f116), .C1(keyinput_f40), .C2(
        n21355), .A(n21354), .ZN(n21360) );
  OAI22_X1 U24273 ( .A1(n12958), .A2(keyinput_f82), .B1(n21358), .B2(
        keyinput_f19), .ZN(n21357) );
  AOI221_X1 U24274 ( .B1(n12958), .B2(keyinput_f82), .C1(keyinput_f19), .C2(
        n21358), .A(n21357), .ZN(n21359) );
  NAND4_X1 U24275 ( .A1(n21362), .A2(n21361), .A3(n21360), .A4(n21359), .ZN(
        n21363) );
  NOR4_X1 U24276 ( .A1(n21366), .A2(n21365), .A3(n21364), .A4(n21363), .ZN(
        n21499) );
  OAI22_X1 U24277 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_f96), .B1(
        P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .ZN(n21367) );
  AOI221_X1 U24278 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .C1(
        keyinput_f112), .C2(P1_EBX_REG_3__SCAN_IN), .A(n21367), .ZN(n21374) );
  OAI22_X1 U24279 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput_f126), .B1(
        keyinput_f78), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n21368) );
  AOI221_X1 U24280 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .C1(
        P1_REIP_REG_5__SCAN_IN), .C2(keyinput_f78), .A(n21368), .ZN(n21373) );
  OAI22_X1 U24281 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_f79), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(keyinput_f72), .ZN(n21369) );
  AOI221_X1 U24282 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_f79), .C1(
        keyinput_f72), .C2(P1_REIP_REG_11__SCAN_IN), .A(n21369), .ZN(n21372)
         );
  OAI22_X1 U24283 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_W_R_N_REG_SCAN_IN), .B2(keyinput_f47), .ZN(n21370) );
  AOI221_X1 U24284 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f47), .C2(P1_W_R_N_REG_SCAN_IN), .A(n21370), .ZN(n21371) );
  NAND4_X1 U24285 ( .A1(n21374), .A2(n21373), .A3(n21372), .A4(n21371), .ZN(
        n21497) );
  OAI22_X1 U24286 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_f125), .B1(
        DATAI_30_), .B2(keyinput_f2), .ZN(n21375) );
  AOI221_X1 U24287 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(keyinput_f125), .C1(
        keyinput_f2), .C2(DATAI_30_), .A(n21375), .ZN(n21400) );
  OAI22_X1 U24288 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_f80), .B1(
        DATAI_29_), .B2(keyinput_f3), .ZN(n21376) );
  AOI221_X1 U24289 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_f80), .C1(
        keyinput_f3), .C2(DATAI_29_), .A(n21376), .ZN(n21379) );
  OAI22_X1 U24290 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_f109), .B1(
        keyinput_f30), .B2(DATAI_2_), .ZN(n21377) );
  AOI221_X1 U24291 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_f109), .C1(
        DATAI_2_), .C2(keyinput_f30), .A(n21377), .ZN(n21378) );
  OAI211_X1 U24292 ( .C1(n12796), .C2(keyinput_f83), .A(n21379), .B(n21378), 
        .ZN(n21380) );
  AOI21_X1 U24293 ( .B1(n12796), .B2(keyinput_f83), .A(n21380), .ZN(n21399) );
  AOI22_X1 U24294 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput_f81), .B1(
        DATAI_31_), .B2(keyinput_f1), .ZN(n21381) );
  OAI221_X1 U24295 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_f81), .C1(
        DATAI_31_), .C2(keyinput_f1), .A(n21381), .ZN(n21388) );
  AOI22_X1 U24296 ( .A1(keyinput_f50), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        DATAI_0_), .B2(keyinput_f32), .ZN(n21382) );
  OAI221_X1 U24297 ( .B1(keyinput_f50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), 
        .C1(DATAI_0_), .C2(keyinput_f32), .A(n21382), .ZN(n21387) );
  AOI22_X1 U24298 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .ZN(n21383) );
  OAI221_X1 U24299 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(
        P1_EBX_REG_28__SCAN_IN), .C2(keyinput_f87), .A(n21383), .ZN(n21386) );
  AOI22_X1 U24300 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .ZN(n21384) );
  OAI221_X1 U24301 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_EBX_REG_14__SCAN_IN), .C2(keyinput_f101), .A(n21384), .ZN(n21385)
         );
  NOR4_X1 U24302 ( .A1(n21388), .A2(n21387), .A3(n21386), .A4(n21385), .ZN(
        n21398) );
  AOI22_X1 U24303 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_f56), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(keyinput_f97), .ZN(n21389) );
  OAI221_X1 U24304 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_f56), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_f97), .A(n21389), .ZN(n21396) );
  AOI22_X1 U24305 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(keyinput_f94), .ZN(n21390) );
  OAI221_X1 U24306 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_EBX_REG_21__SCAN_IN), .C2(keyinput_f94), .A(n21390), .ZN(n21395) );
  AOI22_X1 U24307 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .ZN(n21391) );
  OAI221_X1 U24308 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_f55), .A(n21391), .ZN(n21394)
         );
  AOI22_X1 U24309 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_f75), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21392) );
  OAI221_X1 U24310 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21392), .ZN(n21393)
         );
  NOR4_X1 U24311 ( .A1(n21396), .A2(n21395), .A3(n21394), .A4(n21393), .ZN(
        n21397) );
  NAND4_X1 U24312 ( .A1(n21400), .A2(n21399), .A3(n21398), .A4(n21397), .ZN(
        n21496) );
  AOI22_X1 U24313 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_f64), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_f121), .ZN(n21401) );
  OAI221_X1 U24314 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_f64), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_f121), .A(n21401), .ZN(n21408)
         );
  AOI22_X1 U24315 ( .A1(keyinput_f35), .A2(BS16), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(keyinput_f90), .ZN(n21402) );
  OAI221_X1 U24316 ( .B1(keyinput_f35), .B2(BS16), .C1(P1_EBX_REG_25__SCAN_IN), 
        .C2(keyinput_f90), .A(n21402), .ZN(n21407) );
  AOI22_X1 U24317 ( .A1(DATAI_6_), .A2(keyinput_f26), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .ZN(n21403) );
  OAI221_X1 U24318 ( .B1(DATAI_6_), .B2(keyinput_f26), .C1(
        P1_EBX_REG_4__SCAN_IN), .C2(keyinput_f111), .A(n21403), .ZN(n21406) );
  AOI22_X1 U24319 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .ZN(n21404) );
  OAI221_X1 U24320 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_f85), .A(n21404), .ZN(n21405) );
  NOR4_X1 U24321 ( .A1(n21408), .A2(n21407), .A3(n21406), .A4(n21405), .ZN(
        n21436) );
  AOI22_X1 U24322 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_f89), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n21409) );
  OAI221_X1 U24323 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n21409), .ZN(n21416)
         );
  AOI22_X1 U24324 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .ZN(n21410) );
  OAI221_X1 U24325 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        P1_EAX_REG_23__SCAN_IN), .C2(keyinput_f124), .A(n21410), .ZN(n21415)
         );
  AOI22_X1 U24326 ( .A1(DATAI_18_), .A2(keyinput_f14), .B1(
        P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .ZN(n21411) );
  OAI221_X1 U24327 ( .B1(DATAI_18_), .B2(keyinput_f14), .C1(
        P1_EBX_REG_20__SCAN_IN), .C2(keyinput_f95), .A(n21411), .ZN(n21414) );
  AOI22_X1 U24328 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .ZN(n21412) );
  OAI221_X1 U24329 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(
        P1_EBX_REG_1__SCAN_IN), .C2(keyinput_f114), .A(n21412), .ZN(n21413) );
  NOR4_X1 U24330 ( .A1(n21416), .A2(n21415), .A3(n21414), .A4(n21413), .ZN(
        n21435) );
  AOI22_X1 U24331 ( .A1(DATAI_11_), .A2(keyinput_f21), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .ZN(n21417) );
  OAI221_X1 U24332 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_f84), .A(n21417), .ZN(n21424) );
  AOI22_X1 U24333 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_f77), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .ZN(n21418) );
  OAI221_X1 U24334 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_f77), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21418), .ZN(n21423)
         );
  AOI22_X1 U24335 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(
        P1_EBX_REG_9__SCAN_IN), .B2(keyinput_f106), .ZN(n21419) );
  OAI221_X1 U24336 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(
        P1_EBX_REG_9__SCAN_IN), .C2(keyinput_f106), .A(n21419), .ZN(n21422) );
  AOI22_X1 U24337 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput_f73), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(keyinput_f99), .ZN(n21420) );
  OAI221_X1 U24338 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput_f73), .C1(
        P1_EBX_REG_16__SCAN_IN), .C2(keyinput_f99), .A(n21420), .ZN(n21421) );
  NOR4_X1 U24339 ( .A1(n21424), .A2(n21423), .A3(n21422), .A4(n21421), .ZN(
        n21434) );
  AOI22_X1 U24340 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_f38), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n21425) );
  OAI221_X1 U24341 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n21425), .ZN(n21432)
         );
  AOI22_X1 U24342 ( .A1(DATAI_10_), .A2(keyinput_f22), .B1(DATAI_14_), .B2(
        keyinput_f18), .ZN(n21426) );
  OAI221_X1 U24343 ( .B1(DATAI_10_), .B2(keyinput_f22), .C1(DATAI_14_), .C2(
        keyinput_f18), .A(n21426), .ZN(n21431) );
  AOI22_X1 U24344 ( .A1(keyinput_f49), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n21427) );
  OAI221_X1 U24345 ( .B1(keyinput_f49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), 
        .C1(P1_REIP_REG_25__SCAN_IN), .C2(keyinput_f58), .A(n21427), .ZN(
        n21430) );
  AOI22_X1 U24346 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(keyinput_f70), .ZN(n21428) );
  OAI221_X1 U24347 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(
        P1_REIP_REG_13__SCAN_IN), .C2(keyinput_f70), .A(n21428), .ZN(n21429)
         );
  NOR4_X1 U24348 ( .A1(n21432), .A2(n21431), .A3(n21430), .A4(n21429), .ZN(
        n21433) );
  NAND4_X1 U24349 ( .A1(n21436), .A2(n21435), .A3(n21434), .A4(n21433), .ZN(
        n21495) );
  AOI22_X1 U24350 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_f76), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .ZN(n21437) );
  OAI221_X1 U24351 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_f76), .C1(
        P1_EBX_REG_11__SCAN_IN), .C2(keyinput_f104), .A(n21437), .ZN(n21444)
         );
  AOI22_X1 U24352 ( .A1(DATAI_12_), .A2(keyinput_f20), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n21438) );
  OAI221_X1 U24353 ( .B1(DATAI_12_), .B2(keyinput_f20), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_f53), .A(n21438), .ZN(n21443)
         );
  AOI22_X1 U24354 ( .A1(keyinput_f34), .A2(NA), .B1(keyinput_f39), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n21439) );
  OAI221_X1 U24355 ( .B1(keyinput_f34), .B2(NA), .C1(keyinput_f39), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n21439), .ZN(n21442) );
  AOI22_X1 U24356 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_f67), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .ZN(n21440) );
  OAI221_X1 U24357 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_f102), .A(n21440), .ZN(n21441)
         );
  NOR4_X1 U24358 ( .A1(n21444), .A2(n21443), .A3(n21442), .A4(n21441), .ZN(
        n21493) );
  AOI22_X1 U24359 ( .A1(DATAI_27_), .A2(keyinput_f5), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(keyinput_f113), .ZN(n21445) );
  OAI221_X1 U24360 ( .B1(DATAI_27_), .B2(keyinput_f5), .C1(
        P1_EBX_REG_2__SCAN_IN), .C2(keyinput_f113), .A(n21445), .ZN(n21457) );
  AOI22_X1 U24361 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_f86), .B1(n21447), .B2(keyinput_f59), .ZN(n21446) );
  OAI221_X1 U24362 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_f86), .C1(
        n21447), .C2(keyinput_f59), .A(n21446), .ZN(n21456) );
  AOI22_X1 U24363 ( .A1(n21450), .A2(keyinput_f110), .B1(keyinput_f31), .B2(
        n21449), .ZN(n21448) );
  OAI221_X1 U24364 ( .B1(n21450), .B2(keyinput_f110), .C1(n21449), .C2(
        keyinput_f31), .A(n21448), .ZN(n21455) );
  INV_X1 U24365 ( .A(DATAI_3_), .ZN(n21452) );
  AOI22_X1 U24366 ( .A1(n21453), .A2(keyinput_f71), .B1(keyinput_f29), .B2(
        n21452), .ZN(n21451) );
  OAI221_X1 U24367 ( .B1(n21453), .B2(keyinput_f71), .C1(n21452), .C2(
        keyinput_f29), .A(n21451), .ZN(n21454) );
  NOR4_X1 U24368 ( .A1(n21457), .A2(n21456), .A3(n21455), .A4(n21454), .ZN(
        n21492) );
  AOI22_X1 U24369 ( .A1(n21460), .A2(keyinput_f27), .B1(n21459), .B2(
        keyinput_f119), .ZN(n21458) );
  OAI221_X1 U24370 ( .B1(n21460), .B2(keyinput_f27), .C1(n21459), .C2(
        keyinput_f119), .A(n21458), .ZN(n21473) );
  INV_X1 U24371 ( .A(DATAI_21_), .ZN(n21463) );
  INV_X1 U24372 ( .A(DATAI_22_), .ZN(n21462) );
  AOI22_X1 U24373 ( .A1(n21463), .A2(keyinput_f11), .B1(n21462), .B2(
        keyinput_f10), .ZN(n21461) );
  OAI221_X1 U24374 ( .B1(n21463), .B2(keyinput_f11), .C1(n21462), .C2(
        keyinput_f10), .A(n21461), .ZN(n21472) );
  AOI22_X1 U24375 ( .A1(n21466), .A2(keyinput_f122), .B1(keyinput_f41), .B2(
        n21465), .ZN(n21464) );
  OAI221_X1 U24376 ( .B1(n21466), .B2(keyinput_f122), .C1(n21465), .C2(
        keyinput_f41), .A(n21464), .ZN(n21471) );
  AOI22_X1 U24377 ( .A1(n21469), .A2(keyinput_f8), .B1(n21468), .B2(
        keyinput_f93), .ZN(n21467) );
  OAI221_X1 U24378 ( .B1(n21469), .B2(keyinput_f8), .C1(n21468), .C2(
        keyinput_f93), .A(n21467), .ZN(n21470) );
  NOR4_X1 U24379 ( .A1(n21473), .A2(n21472), .A3(n21471), .A4(n21470), .ZN(
        n21491) );
  INV_X1 U24380 ( .A(DATAI_4_), .ZN(n21476) );
  AOI22_X1 U24381 ( .A1(n21476), .A2(keyinput_f28), .B1(n21475), .B2(
        keyinput_f117), .ZN(n21474) );
  OAI221_X1 U24382 ( .B1(n21476), .B2(keyinput_f28), .C1(n21475), .C2(
        keyinput_f117), .A(n21474), .ZN(n21489) );
  AOI22_X1 U24383 ( .A1(n21479), .A2(keyinput_f91), .B1(n21478), .B2(
        keyinput_f123), .ZN(n21477) );
  OAI221_X1 U24384 ( .B1(n21479), .B2(keyinput_f91), .C1(n21478), .C2(
        keyinput_f123), .A(n21477), .ZN(n21488) );
  AOI22_X1 U24385 ( .A1(n21482), .A2(keyinput_f103), .B1(n21481), .B2(
        keyinput_f88), .ZN(n21480) );
  OAI221_X1 U24386 ( .B1(n21482), .B2(keyinput_f103), .C1(n21481), .C2(
        keyinput_f88), .A(n21480), .ZN(n21487) );
  AOI22_X1 U24387 ( .A1(n21485), .A2(keyinput_f98), .B1(n21484), .B2(
        keyinput_f120), .ZN(n21483) );
  OAI221_X1 U24388 ( .B1(n21485), .B2(keyinput_f98), .C1(n21484), .C2(
        keyinput_f120), .A(n21483), .ZN(n21486) );
  NOR4_X1 U24389 ( .A1(n21489), .A2(n21488), .A3(n21487), .A4(n21486), .ZN(
        n21490) );
  NAND4_X1 U24390 ( .A1(n21493), .A2(n21492), .A3(n21491), .A4(n21490), .ZN(
        n21494) );
  NOR4_X1 U24391 ( .A1(n21497), .A2(n21496), .A3(n21495), .A4(n21494), .ZN(
        n21498) );
  NAND4_X1 U24392 ( .A1(n21501), .A2(n21500), .A3(n21499), .A4(n21498), .ZN(
        n21502) );
  OAI221_X1 U24393 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(n21503), .C1(n21507), 
        .C2(keyinput_f105), .A(n21502), .ZN(n21504) );
  OAI21_X1 U24394 ( .B1(n21507), .B2(keyinput_g105), .A(n21504), .ZN(n21505)
         );
  AOI211_X1 U24395 ( .C1(n21507), .C2(keyinput_g105), .A(n21506), .B(n21505), 
        .ZN(n21509) );
  AOI22_X1 U24396 ( .A1(n16721), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16723), .ZN(n21508) );
  XNOR2_X1 U24397 ( .A(n21509), .B(n21508), .ZN(U355) );
  NOR2_X1 U11340 ( .A1(n10438), .A2(n10437), .ZN(n10576) );
  INV_X1 U11285 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13184) );
  INV_X2 U11589 ( .A(n13142), .ZN(n13155) );
  CLKBUF_X1 U11292 ( .A(n11494), .Z(n11439) );
  CLKBUF_X1 U11360 ( .A(n11444), .Z(n11461) );
  INV_X2 U11379 ( .A(n18083), .ZN(n18055) );
  XNOR2_X1 U12819 ( .A(n14249), .B(n14247), .ZN(n15235) );
  OR2_X1 U13177 ( .A1(n10618), .A2(n19564), .ZN(n21510) );
endmodule

