

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314;

  INV_X4 U4936 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  BUF_X2 U4937 ( .A(n6349), .Z(n4431) );
  INV_X1 U4938 ( .A(n5080), .ZN(n5427) );
  AOI22_X1 U4939 ( .A1(n10094), .A2(keyinput21), .B1(keyinput58), .B2(n10093), 
        .ZN(n10092) );
  OAI221_X1 U4940 ( .B1(n10094), .B2(keyinput21), .C1(n10093), .C2(keyinput58), 
        .A(n10092), .ZN(n10098) );
  NAND2_X1 U4941 ( .A1(n6864), .A2(n5046), .ZN(n5047) );
  INV_X1 U4942 ( .A(n7735), .ZN(n7726) );
  INV_X1 U4943 ( .A(n6925), .ZN(n5455) );
  INV_X1 U4944 ( .A(n6926), .ZN(n5663) );
  AND2_X1 U4945 ( .A1(n5160), .A2(n5159), .ZN(n9906) );
  INV_X1 U4946 ( .A(n6065), .ZN(n7713) );
  INV_X1 U4947 ( .A(n9051), .ZN(n8712) );
  NAND2_X1 U4948 ( .A1(n6148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6144) );
  AND2_X1 U4949 ( .A1(n5601), .A2(n5600), .ZN(n8306) );
  AOI211_X1 U4950 ( .C1(n9358), .C2(n9673), .A(n9357), .B(n9356), .ZN(n9421)
         );
  NAND4_X1 U4951 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n9868)
         );
  NAND3_X1 U4952 ( .A1(n4852), .A2(n4851), .A3(n4850), .ZN(n9472) );
  AND4_X1 U4953 ( .A1(n4555), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4430)
         );
  NOR2_X2 U4954 ( .A1(n9230), .A2(n6127), .ZN(n6128) );
  AOI21_X2 U4955 ( .B1(n8279), .B2(n9927), .A(n4512), .ZN(n4736) );
  AND2_X2 U4956 ( .A1(n6812), .A2(n5180), .ZN(n5183) );
  NAND2_X1 U4957 ( .A1(n6750), .A2(n5143), .ZN(n6872) );
  XNOR2_X2 U4958 ( .A(n5674), .B(n5673), .ZN(n5683) );
  INV_X1 U4959 ( .A(n7682), .ZN(n6003) );
  XNOR2_X2 U4960 ( .A(n5030), .B(n5029), .ZN(n7652) );
  NAND2_X4 U4961 ( .A1(n6360), .A2(n6352), .ZN(n6361) );
  INV_X2 U4962 ( .A(n6351), .ZN(n6352) );
  AND2_X4 U4963 ( .A1(n5048), .A2(n5047), .ZN(n5078) );
  XNOR2_X2 U4964 ( .A(n6144), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6156) );
  OR2_X2 U4965 ( .A1(n8328), .A2(n5526), .ZN(n4763) );
  XNOR2_X2 U4966 ( .A(n5042), .B(n5041), .ZN(n5660) );
  AOI21_X1 U4967 ( .B1(n7988), .B2(n4912), .A(n4473), .ZN(n4911) );
  AND2_X1 U4968 ( .A1(n4913), .A2(n7989), .ZN(n4912) );
  NOR2_X1 U4969 ( .A1(n8038), .A2(n8331), .ZN(n7992) );
  NAND2_X1 U4970 ( .A1(n4923), .A2(n4922), .ZN(n9939) );
  NAND2_X2 U4971 ( .A1(n7914), .A2(n7911), .ZN(n7843) );
  NAND2_X2 U4972 ( .A1(n7907), .A2(n7890), .ZN(n7838) );
  NAND4_X1 U4973 ( .A1(n5132), .A2(n5131), .A3(n5130), .A4(n5129), .ZN(n8196)
         );
  NAND4_X1 U4974 ( .A1(n5111), .A2(n5110), .A3(n5109), .A4(n5108), .ZN(n8197)
         );
  CLKBUF_X2 U4975 ( .A(n5146), .Z(n5404) );
  NAND2_X1 U4976 ( .A1(n5789), .A2(n5788), .ZN(n9074) );
  INV_X4 U4977 ( .A(n5835), .ZN(n6293) );
  AND2_X2 U4978 ( .A1(n9472), .A2(n5756), .ZN(n5804) );
  OAI21_X1 U4979 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8025) );
  AND2_X1 U4980 ( .A1(n4659), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U4981 ( .A1(n8309), .A2(n8308), .ZN(n8310) );
  OR2_X1 U4982 ( .A1(n8062), .A2(n9368), .ZN(n4659) );
  OR4_X1 U4983 ( .A1(n8687), .A2(n8693), .A3(n8694), .A4(n8792), .ZN(n8698) );
  NAND2_X1 U4984 ( .A1(n6096), .A2(n4450), .ZN(n8062) );
  INV_X1 U4985 ( .A(n8844), .ZN(n4685) );
  OAI21_X1 U4986 ( .B1(n8746), .B2(n4488), .A(n4445), .ZN(n8687) );
  AND2_X1 U4987 ( .A1(n7678), .A2(n7677), .ZN(n8844) );
  NAND2_X1 U4988 ( .A1(n8327), .A2(n4912), .ZN(n4909) );
  NAND2_X1 U4989 ( .A1(n9206), .A2(n6130), .ZN(n9207) );
  AND2_X1 U4990 ( .A1(n4911), .A2(n4495), .ZN(n4908) );
  AND2_X1 U4991 ( .A1(n9205), .A2(n9000), .ZN(n9221) );
  OAI21_X1 U4992 ( .B1(n7654), .B2(n7653), .A(n7657), .ZN(n7663) );
  AND2_X1 U4993 ( .A1(n9009), .A2(n8808), .ZN(n9182) );
  OR2_X1 U4994 ( .A1(n9227), .A2(n8801), .ZN(n9205) );
  AOI21_X1 U4995 ( .B1(n6128), .B2(n4635), .A(n4634), .ZN(n4633) );
  OR2_X1 U4996 ( .A1(n5652), .A2(n8077), .ZN(n7989) );
  AND2_X1 U4997 ( .A1(n8993), .A2(n9234), .ZN(n9248) );
  NAND2_X1 U4998 ( .A1(n5534), .A2(n5533), .ZN(n8038) );
  OAI21_X1 U4999 ( .B1(n8783), .B2(n8781), .A(n8780), .ZN(n8580) );
  NOR2_X1 U5000 ( .A1(n9379), .A2(n4681), .ZN(n4680) );
  XNOR2_X1 U5001 ( .A(n5532), .B(n5531), .ZN(n7614) );
  NAND2_X1 U5002 ( .A1(n5501), .A2(n5500), .ZN(n8507) );
  AND2_X1 U5003 ( .A1(n5483), .A2(n5482), .ZN(n8350) );
  NAND2_X1 U5004 ( .A1(n9939), .A2(n7933), .ZN(n7213) );
  NAND2_X1 U5005 ( .A1(n5543), .A2(n5542), .ZN(n8321) );
  OAI21_X1 U5006 ( .B1(n7125), .B2(n4623), .A(n4441), .ZN(n4628) );
  NAND2_X1 U5007 ( .A1(n6997), .A2(n5009), .ZN(n7125) );
  NAND2_X1 U5008 ( .A1(n7344), .A2(n7343), .ZN(n7342) );
  OR2_X1 U5009 ( .A1(n5413), .A2(n5412), .ZN(n5417) );
  NAND2_X1 U5010 ( .A1(n5366), .A2(n5365), .ZN(n8540) );
  NAND2_X1 U5011 ( .A1(n8750), .A2(n6789), .ZN(n6908) );
  NAND2_X1 U5012 ( .A1(n5911), .A2(n5910), .ZN(n7229) );
  XNOR2_X1 U5013 ( .A(n5299), .B(n5296), .ZN(n6419) );
  NAND2_X1 U5014 ( .A1(n5201), .A2(n5200), .ZN(n9917) );
  NAND2_X1 U5015 ( .A1(n4722), .A2(n4720), .ZN(n5265) );
  OR2_X1 U5016 ( .A1(n6937), .A2(n6952), .ZN(n6839) );
  INV_X1 U5017 ( .A(n6918), .ZN(n7111) );
  NAND2_X1 U5018 ( .A1(n4833), .A2(n5189), .ZN(n5213) );
  AOI21_X1 U5019 ( .B1(n6576), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6425), .ZN(
        n6427) );
  AND2_X1 U5020 ( .A1(n4819), .A2(n4818), .ZN(n7704) );
  NAND2_X2 U5021 ( .A1(n7068), .A2(n9621), .ZN(n9624) );
  INV_X1 U5022 ( .A(n6361), .ZN(n8635) );
  AND2_X1 U5023 ( .A1(n5034), .A2(n5033), .ZN(n5039) );
  NAND4_X2 U5024 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n8198)
         );
  AND3_X1 U5025 ( .A1(n5101), .A2(n5100), .A3(n5099), .ZN(n6561) );
  AND3_X1 U5026 ( .A1(n5122), .A2(n5121), .A3(n5120), .ZN(n9896) );
  MUX2_X1 U5027 ( .A(n6182), .B(n7837), .S(n8024), .Z(n6184) );
  CLKBUF_X1 U5028 ( .A(n5084), .Z(n6929) );
  XNOR2_X1 U5029 ( .A(n8820), .B(n9074), .ZN(n6438) );
  BUF_X2 U5030 ( .A(n5089), .Z(n5156) );
  NAND2_X1 U5031 ( .A1(n5032), .A2(n5035), .ZN(n5146) );
  INV_X2 U5032 ( .A(n6273), .ZN(n8257) );
  INV_X1 U5033 ( .A(n7665), .ZN(n5032) );
  AND3_X1 U5034 ( .A1(n5786), .A2(n5785), .A3(n5784), .ZN(n5789) );
  NAND3_X1 U5035 ( .A1(n5797), .A2(n5796), .A3(n5795), .ZN(n6723) );
  XNOR2_X1 U5036 ( .A(n5677), .B(n5676), .ZN(n8033) );
  NAND2_X1 U5037 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U5038 ( .A1(n8553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5027) );
  XNOR2_X1 U5039 ( .A(n6001), .B(n6000), .ZN(n6349) );
  OAI21_X1 U5040 ( .B1(n5680), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U5041 ( .A1(n5680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  OR2_X1 U5042 ( .A1(n5040), .A2(n5079), .ZN(n5042) );
  OR2_X1 U5043 ( .A1(n5028), .A2(n5079), .ZN(n5030) );
  INV_X1 U5044 ( .A(n5812), .ZN(n6065) );
  CLKBUF_X1 U5045 ( .A(n6138), .Z(n8054) );
  NAND2_X1 U5046 ( .A1(n5672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  CLKBUF_X1 U5047 ( .A(n5679), .Z(n5680) );
  XNOR2_X1 U5048 ( .A(n6152), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10044) );
  OR3_X1 U5049 ( .A1(n9467), .A2(n4853), .A3(n5745), .ZN(n4852) );
  NAND2_X1 U5050 ( .A1(n4969), .A2(n4497), .ZN(n5624) );
  AND3_X2 U5051 ( .A1(n5023), .A2(n5398), .A3(n4469), .ZN(n5620) );
  OAI21_X1 U5052 ( .B1(n5078), .B2(n4925), .A(n4924), .ZN(n5075) );
  CLKBUF_X1 U5053 ( .A(n5078), .Z(n7671) );
  AND2_X1 U5054 ( .A1(n5806), .A2(n4551), .ZN(n5729) );
  NAND2_X1 U5055 ( .A1(n5053), .A2(n5013), .ZN(n5097) );
  NOR2_X1 U5056 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5196) );
  INV_X1 U5057 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5195) );
  NOR2_X1 U5058 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5015) );
  INV_X1 U5059 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5300) );
  INV_X1 U5060 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5221) );
  INV_X1 U5061 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10016) );
  NOR2_X2 U5062 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6865) );
  AND2_X1 U5063 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6864) );
  OAI21_X2 U5064 ( .B1(n4559), .B2(n4560), .A(n4567), .ZN(n8744) );
  NOR2_X2 U5065 ( .A1(n5022), .A2(n5021), .ZN(n5398) );
  INV_X4 U5066 ( .A(n8630), .ZN(n4574) );
  OAI21_X2 U5067 ( .B1(n4738), .B2(n4518), .A(n4748), .ZN(n8380) );
  NAND2_X1 U5068 ( .A1(n6184), .A2(n6183), .ZN(n4432) );
  OAI21_X2 U5069 ( .B1(n5647), .B2(n4665), .A(n4663), .ZN(n7793) );
  NAND2_X2 U5070 ( .A1(n8378), .A2(n8381), .ZN(n5647) );
  OAI222_X1 U5071 ( .A1(n8562), .A2(n7650), .B1(P2_U3151), .B2(n5683), .C1(
        n7649), .C2(n8555), .ZN(P2_U3271) );
  AOI21_X1 U5072 ( .B1(n7963), .B2(n4468), .A(n4718), .ZN(n4717) );
  NAND2_X1 U5073 ( .A1(n7966), .A2(n7961), .ZN(n4718) );
  OAI21_X1 U5074 ( .B1(n4831), .B2(n4832), .A(n8002), .ZN(n4829) );
  AOI21_X1 U5075 ( .B1(n4845), .B2(n4846), .A(n5315), .ZN(n4843) );
  OR2_X1 U5076 ( .A1(n9523), .A2(n7568), .ZN(n7944) );
  OR2_X1 U5077 ( .A1(n8692), .A2(n8684), .ZN(n9012) );
  NOR2_X1 U5078 ( .A1(n6101), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U5079 ( .A1(n5212), .A2(n5214), .ZN(n4731) );
  INV_X1 U5080 ( .A(n5404), .ZN(n5613) );
  NOR2_X1 U5081 ( .A1(n5642), .A2(n7962), .ZN(n4926) );
  INV_X1 U5082 ( .A(n5804), .ZN(n6133) );
  INV_X4 U5083 ( .A(n5078), .ZN(n7676) );
  NAND2_X1 U5084 ( .A1(n7677), .A2(n7676), .ZN(n5843) );
  NAND2_X1 U5085 ( .A1(n8924), .A2(n9020), .ZN(n4612) );
  NAND2_X1 U5086 ( .A1(n8921), .A2(n4616), .ZN(n4613) );
  INV_X1 U5087 ( .A(n7124), .ZN(n4624) );
  NAND2_X1 U5088 ( .A1(n4588), .A2(n7100), .ZN(n8826) );
  OR2_X1 U5089 ( .A1(n7301), .A2(n7305), .ZN(n7302) );
  NAND2_X1 U5090 ( .A1(n6696), .A2(n9707), .ZN(n6699) );
  OR2_X1 U5091 ( .A1(n9697), .A2(n6686), .ZN(n6698) );
  AOI21_X1 U5092 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8234), .A(n9802), .ZN(
        n8206) );
  INV_X1 U5093 ( .A(n4745), .ZN(n4744) );
  OR2_X1 U5094 ( .A1(n9942), .A2(n8190), .ZN(n4773) );
  OR2_X1 U5095 ( .A1(n9942), .A2(n7458), .ZN(n7933) );
  INV_X1 U5096 ( .A(n9906), .ZN(n4734) );
  INV_X1 U5097 ( .A(n8531), .ZN(n5643) );
  NAND2_X1 U5098 ( .A1(n5026), .A2(n4465), .ZN(n5679) );
  INV_X1 U5099 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U5100 ( .A1(n4459), .A2(n4570), .ZN(n4569) );
  INV_X1 U5101 ( .A(n8614), .ZN(n4570) );
  OR2_X1 U5102 ( .A1(n7382), .A2(n7490), .ZN(n8952) );
  INV_X1 U5103 ( .A(n7601), .ZN(n6170) );
  NAND2_X1 U5104 ( .A1(n4515), .A2(n4514), .ZN(n7670) );
  INV_X1 U5105 ( .A(n7662), .ZN(n4514) );
  INV_X1 U5106 ( .A(n7663), .ZN(n4515) );
  AND2_X1 U5107 ( .A1(n5739), .A2(n6145), .ZN(n4594) );
  INV_X1 U5108 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5739) );
  AND2_X1 U5109 ( .A1(n10180), .A2(n5744), .ZN(n4880) );
  AND2_X1 U5110 ( .A1(n4592), .A2(n4591), .ZN(n6142) );
  NOR2_X1 U5111 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  NAND2_X1 U5112 ( .A1(n4838), .A2(n4836), .ZN(n5393) );
  AOI21_X1 U5113 ( .B1(n5357), .B2(n4839), .A(n4837), .ZN(n4836) );
  INV_X1 U5114 ( .A(n5373), .ZN(n4837) );
  INV_X1 U5115 ( .A(n5280), .ZN(n4848) );
  AND2_X1 U5116 ( .A1(n5239), .A2(n5218), .ZN(n5219) );
  NAND2_X1 U5117 ( .A1(n5214), .A2(n5194), .ZN(n5212) );
  OR2_X1 U5118 ( .A1(n4935), .A2(n7048), .ZN(n4934) );
  INV_X1 U5119 ( .A(n4939), .ZN(n4935) );
  OR2_X1 U5120 ( .A1(n5223), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5267) );
  INV_X1 U5121 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7475) );
  INV_X1 U5122 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4928) );
  NOR2_X1 U5123 ( .A1(n8250), .A2(n4901), .ZN(n8251) );
  NOR2_X1 U5124 ( .A1(n8262), .A2(n8199), .ZN(n4901) );
  NAND2_X1 U5125 ( .A1(n4753), .A2(n4750), .ZN(n8292) );
  INV_X1 U5126 ( .A(n4751), .ZN(n4750) );
  OAI21_X1 U5127 ( .B1(n4758), .B2(n4752), .A(n4756), .ZN(n4751) );
  INV_X1 U5128 ( .A(n4664), .ZN(n4663) );
  OAI21_X1 U5129 ( .B1(n4435), .B2(n4665), .A(n7970), .ZN(n4664) );
  INV_X1 U5130 ( .A(n7972), .ZN(n4665) );
  AND4_X1 U5131 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n8395)
         );
  AND2_X1 U5132 ( .A1(n4771), .A2(n4773), .ZN(n4770) );
  INV_X1 U5133 ( .A(n7851), .ZN(n4771) );
  OR2_X1 U5134 ( .A1(n7080), .A2(n5295), .ZN(n4772) );
  NAND2_X1 U5135 ( .A1(n6270), .A2(n6250), .ZN(n6212) );
  OR2_X1 U5136 ( .A1(n8523), .A2(n8393), .ZN(n7959) );
  AND4_X1 U5137 ( .A1(n5410), .A2(n5409), .A3(n5408), .A4(n5407), .ZN(n8382)
         );
  AOI21_X1 U5138 ( .B1(n4918), .B2(n4921), .A(n4916), .ZN(n4915) );
  INV_X1 U5139 ( .A(n7947), .ZN(n4921) );
  NOR2_X1 U5140 ( .A1(n5721), .A2(n5698), .ZN(n6209) );
  AOI21_X1 U5141 ( .B1(n4996), .B2(n8672), .A(n4466), .ZN(n4994) );
  NAND2_X1 U5142 ( .A1(n4978), .A2(n4980), .ZN(n4977) );
  INV_X1 U5143 ( .A(n8565), .ZN(n4978) );
  AND2_X1 U5144 ( .A1(n6049), .A2(n6048), .ZN(n8713) );
  AOI21_X1 U5145 ( .B1(n4633), .B2(n4636), .A(n4632), .ZN(n4631) );
  OR2_X1 U5146 ( .A1(n7541), .A2(n7491), .ZN(n8957) );
  NAND2_X1 U5147 ( .A1(n7256), .A2(n5931), .ZN(n7486) );
  OR2_X1 U5148 ( .A1(n4431), .A2(n6357), .ZN(n7135) );
  AOI21_X1 U5149 ( .B1(n4776), .B2(n4780), .A(n4474), .ZN(n4775) );
  NAND2_X1 U5150 ( .A1(n9450), .A2(n9057), .ZN(n6022) );
  NAND2_X1 U5151 ( .A1(n7503), .A2(n5946), .ZN(n5947) );
  OR2_X1 U5152 ( .A1(n7541), .A2(n9061), .ZN(n5946) );
  NAND2_X2 U5153 ( .A1(n6257), .A2(n6138), .ZN(n7677) );
  NAND4_X1 U5154 ( .A1(n4880), .A2(n4593), .A3(n6142), .A4(n4594), .ZN(n5753)
         );
  AND2_X1 U5155 ( .A1(n5738), .A2(n5747), .ZN(n4593) );
  NAND2_X1 U5156 ( .A1(n5580), .A2(n5579), .ZN(n8452) );
  NAND2_X1 U5157 ( .A1(n6084), .A2(n6083), .ZN(n8692) );
  OR2_X1 U5158 ( .A1(n7682), .A2(n8055), .ZN(n6083) );
  INV_X1 U5159 ( .A(n8684), .ZN(n9050) );
  NAND2_X1 U5160 ( .A1(n4438), .A2(n4480), .ZN(n4610) );
  NAND2_X1 U5161 ( .A1(n8922), .A2(n4616), .ZN(n4614) );
  NAND2_X1 U5162 ( .A1(n8925), .A2(n9020), .ZN(n4615) );
  NAND2_X1 U5163 ( .A1(n4438), .A2(n4812), .ZN(n4611) );
  AND2_X1 U5164 ( .A1(n4610), .A2(n8944), .ZN(n4609) );
  AOI21_X1 U5165 ( .B1(n4609), .B2(n4611), .A(n4607), .ZN(n4606) );
  NOR2_X1 U5166 ( .A1(n7963), .A2(n7962), .ZN(n4714) );
  NAND2_X1 U5167 ( .A1(n7961), .A2(n8397), .ZN(n4713) );
  NAND2_X1 U5168 ( .A1(n7967), .A2(n7959), .ZN(n4716) );
  AOI21_X1 U5169 ( .B1(n7975), .B2(n8007), .A(n7984), .ZN(n4709) );
  NAND2_X1 U5170 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  NOR2_X1 U5171 ( .A1(n7990), .A2(n8007), .ZN(n4702) );
  NAND2_X1 U5172 ( .A1(n4707), .A2(n7991), .ZN(n4703) );
  NAND2_X1 U5173 ( .A1(n4706), .A2(n4705), .ZN(n4704) );
  NOR2_X1 U5174 ( .A1(n7988), .A2(n8005), .ZN(n4705) );
  NAND2_X1 U5175 ( .A1(n4707), .A2(n7986), .ZN(n4706) );
  OR2_X1 U5176 ( .A1(n8009), .A2(n8008), .ZN(n4697) );
  INV_X1 U5177 ( .A(n4619), .ZN(n4618) );
  OAI21_X1 U5178 ( .B1(n4452), .B2(n4622), .A(n4620), .ZN(n4619) );
  INV_X1 U5179 ( .A(n7236), .ZN(n4622) );
  NOR2_X1 U5180 ( .A1(n4624), .A2(n7236), .ZN(n4623) );
  INV_X1 U5181 ( .A(n4682), .ZN(n4681) );
  INV_X1 U5182 ( .A(n8911), .ZN(n4862) );
  NOR2_X1 U5183 ( .A1(n4724), .A2(n5257), .ZN(n4723) );
  INV_X1 U5184 ( .A(n4726), .ZN(n4724) );
  NOR2_X1 U5185 ( .A1(n5170), .A2(n4907), .ZN(n4905) );
  INV_X1 U5186 ( .A(SI_5_), .ZN(n4907) );
  INV_X1 U5187 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5045) );
  NAND2_X1 U5188 ( .A1(n4952), .A2(n7569), .ZN(n4951) );
  INV_X1 U5189 ( .A(n7482), .ZN(n4952) );
  OR2_X1 U5190 ( .A1(n7482), .A2(n7568), .ZN(n4949) );
  OR2_X1 U5191 ( .A1(n4950), .A2(n4953), .ZN(n4947) );
  NOR2_X1 U5192 ( .A1(n8189), .A2(n4433), .ZN(n4950) );
  NAND2_X1 U5193 ( .A1(n4433), .A2(n8189), .ZN(n4948) );
  NOR2_X1 U5194 ( .A1(n5008), .A2(n7756), .ZN(n7757) );
  NOR2_X1 U5195 ( .A1(n7755), .A2(n8361), .ZN(n7756) );
  NAND2_X1 U5196 ( .A1(n7047), .A2(n7055), .ZN(n4939) );
  NAND2_X1 U5197 ( .A1(n8021), .A2(n4667), .ZN(n4666) );
  AND2_X1 U5198 ( .A1(n8481), .A2(n8273), .ZN(n8022) );
  NAND2_X1 U5199 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  OR2_X1 U5200 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  NAND2_X1 U5201 ( .A1(n7618), .A2(n7617), .ZN(n7620) );
  NOR2_X1 U5202 ( .A1(n9825), .A2(n10197), .ZN(n4519) );
  AOI21_X1 U5203 ( .B1(n4759), .B2(n4764), .A(n4757), .ZN(n4756) );
  INV_X1 U5204 ( .A(n8000), .ZN(n4757) );
  OR2_X1 U5205 ( .A1(n5367), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U5206 ( .A1(n9942), .A2(n7458), .ZN(n7932) );
  OR2_X1 U5207 ( .A1(n7050), .A2(n7305), .ZN(n7922) );
  AND2_X1 U5208 ( .A1(n7897), .A2(n6839), .ZN(n7920) );
  OR2_X1 U5209 ( .A1(n8197), .A2(n9896), .ZN(n7907) );
  NAND2_X1 U5210 ( .A1(n5685), .A2(n5682), .ZN(n6181) );
  INV_X1 U5211 ( .A(n7992), .ZN(n4913) );
  OR2_X1 U5212 ( .A1(n8496), .A2(n8307), .ZN(n7998) );
  AND2_X1 U5213 ( .A1(n5649), .A2(n8188), .ZN(n7976) );
  OR2_X1 U5214 ( .A1(n8513), .A2(n7796), .ZN(n7970) );
  AND2_X1 U5215 ( .A1(n8540), .A2(n8430), .ZN(n4749) );
  OR2_X1 U5216 ( .A1(n6243), .A2(n5697), .ZN(n5719) );
  INV_X1 U5217 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5041) );
  INV_X1 U5218 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4973) );
  OAI21_X1 U5219 ( .B1(n5006), .B2(n4572), .A(n4569), .ZN(n4568) );
  NOR2_X1 U5220 ( .A1(n4562), .A2(n4571), .ZN(n4561) );
  OR2_X1 U5221 ( .A1(n8616), .A2(n4572), .ZN(n4571) );
  INV_X1 U5222 ( .A(n4994), .ZN(n4562) );
  NAND2_X1 U5223 ( .A1(n4617), .A2(n4624), .ZN(n4625) );
  NAND2_X1 U5224 ( .A1(n7125), .A2(n7123), .ZN(n4617) );
  INV_X1 U5225 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5948) );
  INV_X1 U5226 ( .A(n9012), .ZN(n4855) );
  INV_X1 U5227 ( .A(n6128), .ZN(n4636) );
  AOI21_X1 U5228 ( .B1(n7584), .B2(n4870), .A(n4655), .ZN(n4654) );
  INV_X1 U5229 ( .A(n4868), .ZN(n4655) );
  AOI21_X1 U5230 ( .B1(n4870), .B2(n4873), .A(n4869), .ZN(n4868) );
  INV_X1 U5231 ( .A(n9336), .ZN(n4873) );
  AND2_X1 U5232 ( .A1(n9316), .A2(n9301), .ZN(n9283) );
  NOR2_X1 U5233 ( .A1(n4817), .A2(n4640), .ZN(n4814) );
  INV_X1 U5234 ( .A(n5907), .ZN(n4816) );
  NOR2_X1 U5235 ( .A1(n4812), .A2(n4808), .ZN(n4807) );
  INV_X1 U5236 ( .A(n5858), .ZN(n4811) );
  NAND2_X1 U5237 ( .A1(n6964), .A2(n6966), .ZN(n8923) );
  NOR2_X1 U5238 ( .A1(n6964), .A2(n9626), .ZN(n4678) );
  AND2_X1 U5239 ( .A1(n6114), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U5240 ( .A1(n4866), .A2(n8826), .ZN(n4865) );
  INV_X1 U5241 ( .A(n6112), .ZN(n4866) );
  INV_X1 U5242 ( .A(n8826), .ZN(n4867) );
  NAND2_X1 U5243 ( .A1(n9071), .A2(n7704), .ZN(n8911) );
  AOI21_X1 U5244 ( .B1(n9182), .B2(n4859), .A(n4858), .ZN(n4857) );
  INV_X1 U5245 ( .A(n8808), .ZN(n4858) );
  INV_X1 U5246 ( .A(n9182), .ZN(n4860) );
  NAND2_X1 U5247 ( .A1(n8726), .A2(n9060), .ZN(n4790) );
  OR2_X1 U5248 ( .A1(n7031), .A2(n7363), .ZN(n7263) );
  INV_X1 U5249 ( .A(n7704), .ZN(n6586) );
  NAND2_X1 U5250 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  AND2_X1 U5251 ( .A1(n6105), .A2(n9035), .ZN(n6409) );
  NAND2_X1 U5252 ( .A1(n6156), .A2(n6158), .ZN(n6171) );
  AOI21_X1 U5253 ( .B1(n5550), .B2(n5549), .A(n4511), .ZN(n5570) );
  AND2_X1 U5254 ( .A1(n6097), .A2(n10180), .ZN(n6143) );
  INV_X1 U5255 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5043) );
  AND2_X1 U5256 ( .A1(n5422), .A2(n5416), .ZN(n4849) );
  AND2_X1 U5257 ( .A1(n5394), .A2(n5379), .ZN(n5392) );
  OAI21_X1 U5258 ( .B1(n5265), .B2(n4844), .A(n4843), .ZN(n5319) );
  INV_X1 U5259 ( .A(n4845), .ZN(n4844) );
  INV_X1 U5260 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5955) );
  AOI21_X1 U5261 ( .B1(n4730), .B2(n4728), .A(n4727), .ZN(n4726) );
  INV_X1 U5262 ( .A(n5239), .ZN(n4727) );
  INV_X1 U5263 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4552) );
  NOR2_X1 U5264 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4553) );
  NAND2_X1 U5265 ( .A1(n5078), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U5266 ( .A1(n8158), .A2(n8307), .ZN(n4967) );
  NAND2_X1 U5267 ( .A1(n8157), .A2(n4968), .ZN(n4966) );
  OR2_X1 U5268 ( .A1(n8158), .A2(n8307), .ZN(n4968) );
  NAND2_X1 U5269 ( .A1(n7004), .A2(n6937), .ZN(n4940) );
  INV_X1 U5270 ( .A(n5519), .ZN(n5518) );
  NAND2_X1 U5271 ( .A1(n4958), .A2(n4961), .ZN(n4956) );
  INV_X1 U5272 ( .A(n6624), .ZN(n4958) );
  OR2_X1 U5273 ( .A1(n6189), .A2(n6604), .ZN(n4961) );
  NAND2_X1 U5274 ( .A1(n4929), .A2(n4931), .ZN(n7457) );
  INV_X1 U5275 ( .A(n4932), .ZN(n4931) );
  OAI21_X1 U5276 ( .B1(n4934), .B2(n4933), .A(n7302), .ZN(n4932) );
  OR3_X1 U5277 ( .A1(n7833), .A2(n5705), .A3(n8024), .ZN(n6194) );
  NAND2_X1 U5278 ( .A1(n4886), .A2(n9688), .ZN(n4885) );
  NAND2_X1 U5279 ( .A1(n6536), .A2(n6546), .ZN(n6539) );
  OAI21_X1 U5280 ( .B1(n6696), .B2(n9707), .A(n6699), .ZN(n9697) );
  AND2_X1 U5281 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  XNOR2_X1 U5282 ( .A(n7409), .B(n9715), .ZN(n7411) );
  OR2_X1 U5283 ( .A1(n9740), .A2(n9739), .ZN(n4882) );
  OAI21_X1 U5284 ( .B1(n9724), .B2(n9723), .A(n4506), .ZN(n9732) );
  NAND2_X1 U5285 ( .A1(n9732), .A2(n9731), .ZN(n9730) );
  XNOR2_X1 U5286 ( .A(n7620), .B(n7630), .ZN(n9770) );
  NAND2_X1 U5287 ( .A1(n4889), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5288 ( .A1(n8204), .A2(n4889), .ZN(n4887) );
  INV_X1 U5289 ( .A(n9803), .ZN(n4889) );
  NOR2_X1 U5290 ( .A1(n8293), .A2(n8394), .ZN(n8296) );
  OR2_X1 U5291 ( .A1(n5562), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U5292 ( .A1(n5465), .A2(n10135), .ZN(n5502) );
  INV_X1 U5293 ( .A(n5466), .ZN(n5465) );
  INV_X1 U5294 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U5295 ( .A1(n4772), .A2(n4773), .ZN(n7214) );
  NAND2_X1 U5296 ( .A1(n7040), .A2(n4700), .ZN(n4923) );
  NAND2_X1 U5297 ( .A1(n7933), .A2(n7932), .ZN(n7930) );
  OR2_X1 U5298 ( .A1(n5245), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5271) );
  AND4_X1 U5299 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n7476)
         );
  NAND2_X1 U5300 ( .A1(n4670), .A2(n4672), .ZN(n4669) );
  NAND2_X1 U5301 ( .A1(n4673), .A2(n7013), .ZN(n4670) );
  INV_X1 U5302 ( .A(n7843), .ZN(n4732) );
  AND2_X1 U5303 ( .A1(n5686), .A2(n6245), .ZN(n6649) );
  NAND2_X1 U5304 ( .A1(n8310), .A2(n4475), .ZN(n8288) );
  INV_X1 U5305 ( .A(n8291), .ZN(n5657) );
  XNOR2_X1 U5306 ( .A(n8448), .B(n8306), .ZN(n8291) );
  AND2_X1 U5307 ( .A1(n4495), .A2(n7998), .ZN(n8318) );
  NAND2_X1 U5308 ( .A1(n8501), .A2(n8077), .ZN(n4767) );
  OR2_X1 U5309 ( .A1(n7992), .A2(n4473), .ZN(n7995) );
  INV_X1 U5310 ( .A(n8321), .ZN(n8331) );
  NAND2_X1 U5311 ( .A1(n4927), .A2(n7979), .ZN(n8338) );
  NAND2_X1 U5312 ( .A1(n8369), .A2(n5460), .ZN(n8359) );
  OR2_X1 U5313 ( .A1(n5643), .A2(n8411), .ZN(n4748) );
  NAND2_X1 U5314 ( .A1(n4740), .A2(n4471), .ZN(n4518) );
  AND2_X1 U5315 ( .A1(n7959), .A2(n7966), .ZN(n8381) );
  NAND2_X1 U5316 ( .A1(n5646), .A2(n7964), .ZN(n8378) );
  AOI21_X1 U5317 ( .B1(n7835), .B2(n4746), .A(n4749), .ZN(n4745) );
  INV_X1 U5318 ( .A(n7856), .ZN(n4746) );
  NOR2_X1 U5319 ( .A1(n4749), .A2(n7855), .ZN(n4747) );
  INV_X1 U5320 ( .A(n7835), .ZN(n8419) );
  INV_X4 U5321 ( .A(n5156), .ZN(n7822) );
  OR2_X1 U5322 ( .A1(n7856), .A2(n7855), .ZN(n8429) );
  AOI21_X1 U5323 ( .B1(n4770), .B2(n5295), .A(n4442), .ZN(n4768) );
  AND2_X1 U5324 ( .A1(n6216), .A2(n8005), .ZN(n9866) );
  NAND2_X1 U5325 ( .A1(n4662), .A2(n7944), .ZN(n7326) );
  NAND2_X1 U5326 ( .A1(n7500), .A2(n7837), .ZN(n9919) );
  INV_X1 U5327 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5622) );
  INV_X1 U5328 ( .A(n5097), .ZN(n4894) );
  AND2_X1 U5329 ( .A1(n5079), .A2(n5013), .ZN(n4895) );
  OAI21_X1 U5330 ( .B1(n6908), .B2(n6798), .A(n6797), .ZN(n6799) );
  OR2_X1 U5331 ( .A1(n7281), .A2(n7282), .ZN(n4991) );
  NAND2_X1 U5332 ( .A1(n8565), .A2(n8566), .ZN(n4979) );
  AND2_X1 U5333 ( .A1(n4598), .A2(n4601), .ZN(n8717) );
  AOI21_X1 U5334 ( .B1(n6782), .B2(n6781), .A(n5002), .ZN(n8752) );
  AND3_X1 U5335 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n6426) );
  NAND2_X1 U5336 ( .A1(n4991), .A2(n7377), .ZN(n4989) );
  NAND2_X1 U5337 ( .A1(n4995), .A2(n4451), .ZN(n4566) );
  INV_X1 U5338 ( .A(n8731), .ZN(n4976) );
  NAND2_X1 U5339 ( .A1(n4602), .A2(n4508), .ZN(n4601) );
  INV_X1 U5340 ( .A(n4979), .ZN(n4602) );
  NOR2_X1 U5341 ( .A1(n4976), .A2(n4604), .ZN(n4599) );
  INV_X1 U5342 ( .A(n4974), .ZN(n4596) );
  AOI21_X1 U5343 ( .B1(n8731), .B2(n4975), .A(n4467), .ZN(n4974) );
  INV_X1 U5344 ( .A(n8720), .ZN(n4975) );
  AND2_X1 U5345 ( .A1(n10044), .A2(n8822), .ZN(n8900) );
  AND4_X1 U5346 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n7490)
         );
  AND4_X1 U5347 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n7276)
         );
  AND4_X1 U5348 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n7227)
         );
  AND4_X1 U5349 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n7127)
         );
  AND4_X1 U5350 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n6898)
         );
  NAND2_X1 U5351 ( .A1(n5823), .A2(n4589), .ZN(n4588) );
  NOR2_X1 U5352 ( .A1(n4457), .A2(n4590), .ZN(n4589) );
  NOR2_X1 U5353 ( .A1(n9472), .A2(n5756), .ZN(n5812) );
  INV_X1 U5354 ( .A(n9472), .ZN(n4558) );
  INV_X1 U5355 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5954) );
  INV_X1 U5356 ( .A(n4688), .ZN(n4687) );
  OR2_X1 U5357 ( .A1(n9167), .A2(n7719), .ZN(n4688) );
  AOI21_X1 U5358 ( .B1(n4779), .B2(n6072), .A(n4476), .ZN(n4778) );
  INV_X1 U5359 ( .A(n6061), .ZN(n4779) );
  NAND2_X1 U5360 ( .A1(n9207), .A2(n9003), .ZN(n9181) );
  INV_X1 U5361 ( .A(n8997), .ZN(n4634) );
  INV_X1 U5362 ( .A(n9248), .ZN(n4635) );
  OR2_X1 U5363 ( .A1(n9247), .A2(n4636), .ZN(n4630) );
  NAND2_X1 U5364 ( .A1(n9231), .A2(n6050), .ZN(n9219) );
  NAND2_X1 U5365 ( .A1(n9247), .A2(n9248), .ZN(n9246) );
  NOR2_X1 U5366 ( .A1(n9343), .A2(n9399), .ZN(n9316) );
  INV_X1 U5367 ( .A(n9450), .ZN(n9301) );
  NAND2_X1 U5368 ( .A1(n7584), .A2(n8969), .ZN(n9331) );
  NAND2_X1 U5369 ( .A1(n4645), .A2(n4643), .ZN(n7555) );
  AOI21_X1 U5370 ( .B1(n4646), .B2(n4648), .A(n4644), .ZN(n4643) );
  INV_X1 U5371 ( .A(n8870), .ZN(n4644) );
  OR2_X1 U5372 ( .A1(n4649), .A2(n6119), .ZN(n4648) );
  INV_X1 U5373 ( .A(n8832), .ZN(n4649) );
  NAND2_X1 U5374 ( .A1(n4647), .A2(n8832), .ZN(n4646) );
  INV_X1 U5375 ( .A(n4650), .ZN(n4647) );
  NAND2_X1 U5376 ( .A1(n4652), .A2(n8952), .ZN(n7487) );
  AND2_X1 U5377 ( .A1(n4651), .A2(n8952), .ZN(n4650) );
  OR2_X1 U5378 ( .A1(n7259), .A2(n6119), .ZN(n4652) );
  OAI21_X1 U5379 ( .B1(n7166), .B2(n8867), .A(n8951), .ZN(n7259) );
  NAND2_X1 U5380 ( .A1(n7033), .A2(n8929), .ZN(n7166) );
  AOI21_X1 U5381 ( .B1(n8850), .B2(n4640), .A(n4637), .ZN(n4638) );
  NAND2_X1 U5382 ( .A1(n4543), .A2(n8914), .ZN(n6825) );
  NAND2_X1 U5383 ( .A1(n7342), .A2(n5895), .ZN(n6978) );
  NAND2_X1 U5384 ( .A1(n6978), .A2(n8851), .ZN(n6977) );
  OR2_X1 U5385 ( .A1(n6964), .A2(n9068), .ZN(n5881) );
  NAND2_X1 U5386 ( .A1(n6584), .A2(n5845), .ZN(n6634) );
  NAND2_X1 U5387 ( .A1(n6634), .A2(n8855), .ZN(n6633) );
  NAND2_X1 U5388 ( .A1(n8823), .A2(n4878), .ZN(n4877) );
  INV_X1 U5389 ( .A(n9329), .ZN(n9314) );
  NAND2_X1 U5390 ( .A1(n6451), .A2(n8857), .ZN(n6450) );
  NAND2_X1 U5391 ( .A1(n8853), .A2(n6725), .ZN(n6441) );
  INV_X1 U5392 ( .A(n9342), .ZN(n9317) );
  AND2_X1 U5393 ( .A1(n4658), .A2(n4657), .ZN(n6141) );
  INV_X1 U5394 ( .A(n4793), .ZN(n9231) );
  OAI21_X1 U5395 ( .B1(n9278), .B2(n4797), .A(n4794), .ZN(n4793) );
  NAND2_X1 U5396 ( .A1(n4802), .A2(n6039), .ZN(n4797) );
  INV_X1 U5397 ( .A(n4795), .ZN(n4794) );
  NAND2_X1 U5398 ( .A1(n4802), .A2(n4806), .ZN(n4798) );
  OR2_X1 U5399 ( .A1(n4439), .A2(n9264), .ZN(n4801) );
  INV_X1 U5400 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6024) );
  NOR2_X1 U5401 ( .A1(n9399), .A2(n8785), .ZN(n6013) );
  NOR2_X1 U5402 ( .A1(n4792), .A2(n4789), .ZN(n4788) );
  INV_X1 U5403 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5404 ( .A1(n4786), .A2(n4790), .ZN(n4785) );
  INV_X1 U5405 ( .A(n8872), .ZN(n4786) );
  AOI21_X2 U5406 ( .B1(n7486), .B2(n5945), .A(n4453), .ZN(n7503) );
  AND2_X1 U5407 ( .A1(n8957), .A2(n8960), .ZN(n8870) );
  NAND2_X1 U5408 ( .A1(n7257), .A2(n7258), .ZN(n7256) );
  INV_X1 U5409 ( .A(n7677), .ZN(n6002) );
  XNOR2_X1 U5410 ( .A(n4588), .B(n7100), .ZN(n6510) );
  OR2_X1 U5411 ( .A1(n4689), .A2(n4492), .ZN(n6440) );
  AND2_X1 U5412 ( .A1(n6409), .A2(n6350), .ZN(n9411) );
  XNOR2_X1 U5413 ( .A(n7675), .B(n7674), .ZN(n8552) );
  XNOR2_X1 U5414 ( .A(n4556), .B(n5747), .ZN(n6138) );
  OR2_X1 U5415 ( .A1(n5746), .A2(n5745), .ZN(n4556) );
  NOR2_X1 U5416 ( .A1(n6099), .A2(n5751), .ZN(n5746) );
  NAND2_X1 U5417 ( .A1(n5743), .A2(n4880), .ZN(n5751) );
  XNOR2_X1 U5418 ( .A(n4557), .B(n5744), .ZN(n6257) );
  OR2_X1 U5419 ( .A1(n5742), .A2(n5745), .ZN(n4557) );
  NOR2_X1 U5420 ( .A1(n6099), .A2(n5741), .ZN(n5742) );
  OR2_X1 U5421 ( .A1(n5740), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5741) );
  INV_X1 U5422 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U5423 ( .B1(n6149), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U5424 ( .A(n6154), .B(n4592), .ZN(n9036) );
  XNOR2_X1 U5425 ( .A(n6100), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U5426 ( .A1(n6099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6100) );
  XNOR2_X1 U5427 ( .A(n6103), .B(n6102), .ZN(n8885) );
  INV_X1 U5428 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6102) );
  INV_X1 U5429 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5997) );
  INV_X1 U5430 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U5431 ( .A(n5393), .B(n5392), .ZN(n6878) );
  XNOR2_X1 U5432 ( .A(n4841), .B(n5374), .ZN(n6807) );
  OAI21_X1 U5433 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n4841) );
  NAND2_X1 U5434 ( .A1(n4842), .A2(n4845), .ZN(n5316) );
  NAND2_X1 U5435 ( .A1(n5281), .A2(n5280), .ZN(n5299) );
  OAI21_X1 U5436 ( .B1(n5213), .B2(n5212), .A(n4675), .ZN(n5220) );
  NAND2_X1 U5437 ( .A1(n4725), .A2(n4730), .ZN(n5240) );
  NOR2_X1 U5438 ( .A1(n5219), .A2(n4728), .ZN(n4675) );
  NOR2_X1 U5439 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4551) );
  NAND2_X1 U5440 ( .A1(n6560), .A2(n6559), .ZN(n6558) );
  AND4_X1 U5441 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n8169)
         );
  AND3_X1 U5442 ( .A1(n5438), .A2(n5437), .A3(n5436), .ZN(n8393) );
  NOR2_X1 U5443 ( .A1(n6944), .A2(n6945), .ZN(n6950) );
  NAND2_X1 U5444 ( .A1(n6213), .A2(n9863), .ZN(n8182) );
  NAND2_X1 U5445 ( .A1(n5589), .A2(n5588), .ZN(n8320) );
  INV_X1 U5446 ( .A(n8382), .ZN(n8411) );
  INV_X1 U5447 ( .A(n8169), .ZN(n8430) );
  OAI21_X1 U5448 ( .B1(n6543), .B2(n6310), .A(n4522), .ZN(n6315) );
  NAND2_X1 U5449 ( .A1(n6543), .A2(n6310), .ZN(n4522) );
  AND2_X1 U5450 ( .A1(n5224), .A2(n5267), .ZN(n9746) );
  XNOR2_X1 U5451 ( .A(n8251), .B(n4520), .ZN(n8270) );
  AOI21_X1 U5452 ( .B1(n8269), .B2(n9852), .A(n4539), .ZN(n4538) );
  INV_X1 U5453 ( .A(n8259), .ZN(n4520) );
  OAI21_X1 U5454 ( .B1(n4735), .B2(n9873), .A(n4736), .ZN(n8280) );
  INV_X1 U5455 ( .A(n5602), .ZN(n8448) );
  INV_X1 U5456 ( .A(n9863), .ZN(n8437) );
  AND2_X1 U5457 ( .A1(n8452), .A2(n9943), .ZN(n4517) );
  OAI22_X1 U5458 ( .A1(n6572), .A2(n6571), .B1(n6570), .B2(n6569), .ZN(n6782)
         );
  INV_X1 U5459 ( .A(n9443), .ZN(n9269) );
  INV_X1 U5460 ( .A(n7090), .ZN(n6469) );
  INV_X1 U5461 ( .A(n8570), .ZN(n9060) );
  INV_X1 U5462 ( .A(n6801), .ZN(n9070) );
  INV_X1 U5463 ( .A(n4431), .ZN(n9156) );
  NAND2_X1 U5464 ( .A1(n4875), .A2(n7718), .ZN(n9176) );
  NAND2_X1 U5465 ( .A1(n4876), .A2(n9329), .ZN(n4875) );
  XNOR2_X1 U5466 ( .A(n7712), .B(n7711), .ZN(n4876) );
  NAND2_X1 U5467 ( .A1(n9667), .A2(n6411), .ZN(n9621) );
  INV_X1 U5468 ( .A(n6410), .ZN(n6411) );
  NAND2_X1 U5469 ( .A1(n6095), .A2(n8881), .ZN(n6096) );
  AOI21_X1 U5470 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(n9674), .A(n4482), .ZN(
        n4825) );
  AOI21_X1 U5471 ( .B1(n6141), .B2(n9368), .A(n9674), .ZN(n4824) );
  INV_X1 U5472 ( .A(n6141), .ZN(n4822) );
  OR2_X1 U5473 ( .A1(n5753), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5752) );
  MUX2_X1 U5474 ( .A(n7939), .B(n7938), .S(n8007), .Z(n7940) );
  OAI21_X1 U5475 ( .B1(n4605), .B2(n4611), .A(n4610), .ZN(n8946) );
  OAI21_X1 U5476 ( .B1(n8918), .B2(n4608), .A(n4606), .ZN(n8950) );
  INV_X1 U5477 ( .A(n4609), .ZN(n4608) );
  OAI22_X1 U5478 ( .A1(n4715), .A2(n8005), .B1(n4712), .B2(n4711), .ZN(n7969)
         );
  NAND2_X1 U5479 ( .A1(n8381), .A2(n4472), .ZN(n4711) );
  NAND2_X1 U5480 ( .A1(n4583), .A2(n4462), .ZN(n4582) );
  NAND2_X1 U5481 ( .A1(n8940), .A2(n8939), .ZN(n4583) );
  NOR2_X1 U5482 ( .A1(n8943), .A2(n4616), .ZN(n4581) );
  OAI211_X1 U5483 ( .C1(n4585), .C2(n4584), .A(n8964), .B(n4580), .ZN(n8974)
         );
  NAND2_X1 U5484 ( .A1(n8963), .A2(n4616), .ZN(n4584) );
  NOR2_X1 U5485 ( .A1(n4443), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U5486 ( .A1(n4582), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U5487 ( .A1(n4710), .A2(n4709), .ZN(n4708) );
  NAND2_X1 U5488 ( .A1(n4704), .A2(n4701), .ZN(n7996) );
  INV_X1 U5489 ( .A(n7999), .ZN(n4831) );
  NAND2_X1 U5490 ( .A1(n4624), .A2(n4621), .ZN(n4620) );
  INV_X1 U5491 ( .A(n7123), .ZN(n4621) );
  INV_X1 U5492 ( .A(n9008), .ZN(n4578) );
  OAI21_X1 U5493 ( .B1(n8996), .B2(n8995), .A(n4486), .ZN(n4579) );
  NOR2_X1 U5494 ( .A1(n4760), .A2(n5654), .ZN(n4759) );
  INV_X1 U5495 ( .A(n4765), .ZN(n4760) );
  OAI21_X1 U5496 ( .B1(n4577), .B2(n4576), .A(n4575), .ZN(n9013) );
  NAND2_X1 U5497 ( .A1(n9010), .A2(n9020), .ZN(n4575) );
  OR2_X1 U5498 ( .A1(n9010), .A2(n9007), .ZN(n4576) );
  AOI21_X1 U5499 ( .B1(n4579), .B2(n4461), .A(n4578), .ZN(n4577) );
  AND2_X1 U5500 ( .A1(n8965), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U5501 ( .A1(n9336), .A2(n4872), .ZN(n4871) );
  INV_X1 U5502 ( .A(n8969), .ZN(n4872) );
  NOR2_X1 U5503 ( .A1(n9269), .A2(n9390), .ZN(n4682) );
  INV_X1 U5504 ( .A(n10044), .ZN(n6105) );
  NAND2_X1 U5505 ( .A1(n5610), .A2(n5609), .ZN(n7656) );
  OR2_X1 U5506 ( .A1(n5547), .A2(n5546), .ZN(n5551) );
  INV_X1 U5507 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5733) );
  NOR2_X1 U5508 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5734) );
  INV_X1 U5509 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5396) );
  NOR2_X1 U5510 ( .A1(n5374), .A2(n4840), .ZN(n4839) );
  INV_X1 U5511 ( .A(n5356), .ZN(n4840) );
  INV_X1 U5512 ( .A(SI_14_), .ZN(n5321) );
  INV_X1 U5513 ( .A(n7052), .ZN(n4933) );
  NOR2_X1 U5514 ( .A1(n4933), .A2(n4938), .ZN(n4930) );
  AND2_X1 U5515 ( .A1(n7831), .A2(n7867), .ZN(n4528) );
  AND2_X1 U5516 ( .A1(n8446), .A2(n8184), .ZN(n8006) );
  NAND2_X1 U5517 ( .A1(n8017), .A2(n8016), .ZN(n4693) );
  NAND2_X1 U5518 ( .A1(n4885), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U5519 ( .A1(n8239), .A2(n9794), .ZN(n8240) );
  AND2_X1 U5520 ( .A1(n9847), .A2(n4542), .ZN(n8223) );
  NAND2_X1 U5521 ( .A1(n9843), .A2(n8221), .ZN(n4542) );
  INV_X1 U5522 ( .A(n4759), .ZN(n4758) );
  NAND2_X1 U5523 ( .A1(n4761), .A2(n5526), .ZN(n4752) );
  NOR2_X1 U5524 ( .A1(n4758), .A2(n4762), .ZN(n4754) );
  INV_X1 U5525 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10241) );
  BUF_X1 U5526 ( .A(n5634), .Z(n7879) );
  AND2_X1 U5527 ( .A1(n7979), .A2(n7977), .ZN(n7861) );
  OR2_X1 U5528 ( .A1(n5643), .A2(n8382), .ZN(n7964) );
  INV_X1 U5529 ( .A(n7953), .ZN(n4916) );
  AOI21_X1 U5530 ( .B1(n7947), .B2(n4920), .A(n4919), .ZN(n4918) );
  INV_X1 U5531 ( .A(n7948), .ZN(n4920) );
  INV_X1 U5532 ( .A(n7952), .ZN(n4919) );
  XNOR2_X1 U5533 ( .A(n5684), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5699) );
  INV_X1 U5534 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5535 ( .A1(n6360), .A2(n6353), .ZN(n6424) );
  NAND2_X1 U5536 ( .A1(n4588), .A2(n6773), .ZN(n6784) );
  AOI22_X1 U5537 ( .A1(n8754), .A2(n6773), .B1(n8635), .B2(n4588), .ZN(n6787)
         );
  NAND2_X1 U5538 ( .A1(n4628), .A2(n4477), .ZN(n7531) );
  NAND2_X1 U5539 ( .A1(n4989), .A2(n7386), .ZN(n4987) );
  NAND2_X1 U5540 ( .A1(n5824), .A2(n5825), .ZN(n4590) );
  NOR2_X1 U5541 ( .A1(n4679), .A2(n7373), .ZN(n6982) );
  INV_X1 U5542 ( .A(n6106), .ZN(n4878) );
  OR2_X1 U5543 ( .A1(n7719), .A2(n7706), .ZN(n9016) );
  INV_X1 U5544 ( .A(n4778), .ZN(n4777) );
  AND2_X1 U5545 ( .A1(n9283), .A2(n4493), .ZN(n9238) );
  OAI21_X1 U5546 ( .B1(n4437), .B2(n4796), .A(n4454), .ZN(n4795) );
  INV_X1 U5547 ( .A(n6039), .ZN(n4796) );
  OR2_X1 U5548 ( .A1(n9432), .A2(n8713), .ZN(n8997) );
  NAND2_X1 U5549 ( .A1(n9283), .A2(n4680), .ZN(n9253) );
  NAND2_X1 U5550 ( .A1(n9283), .A2(n9290), .ZN(n9284) );
  NAND2_X1 U5551 ( .A1(n7506), .A2(n4478), .ZN(n9343) );
  AND2_X1 U5552 ( .A1(n7506), .A2(n7511), .ZN(n7561) );
  NAND2_X1 U5553 ( .A1(n6830), .A2(n4676), .ZN(n4679) );
  NOR2_X1 U5554 ( .A1(n7352), .A2(n4677), .ZN(n4676) );
  INV_X1 U5555 ( .A(n4678), .ZN(n4677) );
  NAND2_X1 U5556 ( .A1(n4544), .A2(n8909), .ZN(n6637) );
  OR2_X1 U5557 ( .A1(n6519), .A2(n8754), .ZN(n6587) );
  XNOR2_X1 U5558 ( .A(n7656), .B(n7655), .ZN(n7654) );
  AND2_X1 U5559 ( .A1(n5571), .A2(n5559), .ZN(n5569) );
  AND2_X1 U5560 ( .A1(n5545), .A2(n5514), .ZN(n5553) );
  INV_X1 U5561 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10169) );
  INV_X1 U5562 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10135) );
  AND2_X1 U5563 ( .A1(n5439), .A2(n5421), .ZN(n5422) );
  AOI21_X1 U5564 ( .B1(n5264), .B2(n4847), .A(n4444), .ZN(n4845) );
  AOI21_X1 U5565 ( .B1(n4721), .B2(n4726), .A(n4490), .ZN(n4720) );
  NAND2_X1 U5566 ( .A1(n5213), .A2(n4723), .ZN(n4722) );
  OR2_X1 U5567 ( .A1(n5265), .A2(n5264), .ZN(n5281) );
  NAND2_X1 U5568 ( .A1(n5213), .A2(n5214), .ZN(n4725) );
  OAI21_X1 U5569 ( .B1(n5155), .B2(n5170), .A(n5173), .ZN(n4835) );
  NAND2_X1 U5570 ( .A1(n5139), .A2(n5138), .ZN(n5154) );
  INV_X1 U5571 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5728) );
  NOR2_X1 U5572 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5806) );
  OAI21_X1 U5573 ( .B1(n7676), .B2(n5051), .A(n5800), .ZN(n5073) );
  NAND2_X1 U5574 ( .A1(n6865), .A2(n5045), .ZN(n5048) );
  INV_X1 U5575 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5046) );
  NAND2_X1 U5576 ( .A1(n4947), .A2(n4948), .ZN(n4946) );
  NAND2_X1 U5577 ( .A1(n4951), .A2(n4949), .ZN(n4944) );
  INV_X1 U5578 ( .A(n7480), .ZN(n4945) );
  AOI21_X1 U5579 ( .B1(n7730), .B2(n8179), .A(n8126), .ZN(n4942) );
  INV_X1 U5580 ( .A(n5386), .ZN(n5385) );
  NAND2_X1 U5581 ( .A1(n4957), .A2(n4955), .ZN(n6943) );
  NAND2_X1 U5582 ( .A1(n4960), .A2(n4956), .ZN(n4955) );
  NAND2_X1 U5583 ( .A1(n4943), .A2(n7725), .ZN(n8175) );
  INV_X1 U5584 ( .A(n8178), .ZN(n4943) );
  NAND2_X1 U5585 ( .A1(n5629), .A2(n8255), .ZN(n4699) );
  NOR2_X1 U5586 ( .A1(n8025), .A2(n8265), .ZN(n4668) );
  NAND2_X1 U5587 ( .A1(n4883), .A2(n6539), .ZN(n9679) );
  INV_X1 U5588 ( .A(n4884), .ZN(n4883) );
  NAND2_X1 U5589 ( .A1(n6688), .A2(n4540), .ZN(n9704) );
  OR2_X1 U5590 ( .A1(n6689), .A2(n6690), .ZN(n4540) );
  OR2_X1 U5591 ( .A1(n6711), .A2(n4525), .ZN(n6714) );
  NAND2_X1 U5592 ( .A1(n9704), .A2(n9703), .ZN(n9702) );
  INV_X1 U5593 ( .A(n6698), .ZN(n6700) );
  NOR2_X1 U5594 ( .A1(n7430), .A2(n4531), .ZN(n9724) );
  NOR2_X1 U5595 ( .A1(n4533), .A2(n4532), .ZN(n4531) );
  INV_X1 U5596 ( .A(n7432), .ZN(n4532) );
  INV_X1 U5597 ( .A(n7431), .ZN(n4533) );
  NAND2_X1 U5598 ( .A1(n4524), .A2(n4523), .ZN(n9736) );
  NAND2_X1 U5599 ( .A1(n9730), .A2(n7435), .ZN(n9750) );
  XNOR2_X1 U5600 ( .A(n7424), .B(n9746), .ZN(n9748) );
  XNOR2_X1 U5601 ( .A(n7413), .B(n9746), .ZN(n9755) );
  AND2_X1 U5602 ( .A1(n4882), .A2(n4881), .ZN(n7413) );
  NAND2_X1 U5603 ( .A1(n7428), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4881) );
  NOR2_X1 U5604 ( .A1(n9755), .A2(n5227), .ZN(n9754) );
  OR2_X1 U5605 ( .A1(n5267), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5283) );
  OAI21_X1 U5606 ( .B1(n9770), .B2(n4891), .A(n4890), .ZN(n9786) );
  NAND2_X1 U5607 ( .A1(n4892), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4891) );
  INV_X1 U5608 ( .A(n9787), .ZN(n4892) );
  NOR2_X1 U5609 ( .A1(n9770), .A2(n7043), .ZN(n9769) );
  NOR2_X1 U5610 ( .A1(n5283), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5301) );
  AOI21_X1 U5611 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7637), .A(n9786), .ZN(
        n8201) );
  XOR2_X1 U5612 ( .A(n8241), .B(n8240), .Z(n9811) );
  NOR2_X1 U5613 ( .A1(n8207), .A2(n9818), .ZN(n9836) );
  XNOR2_X1 U5614 ( .A(n8243), .B(n9843), .ZN(n9846) );
  NAND2_X1 U5615 ( .A1(n9846), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U5616 ( .A1(n9829), .A2(n8220), .ZN(n9848) );
  NAND2_X1 U5617 ( .A1(n9848), .A2(n9849), .ZN(n9847) );
  AND2_X1 U5618 ( .A1(n5198), .A2(n5197), .ZN(n5397) );
  OR2_X1 U5619 ( .A1(n9855), .A2(n8414), .ZN(n4903) );
  INV_X1 U5620 ( .A(n8268), .ZN(n4539) );
  OR2_X1 U5621 ( .A1(n8448), .A2(n8186), .ZN(n5603) );
  INV_X1 U5622 ( .A(n5670), .ZN(n4512) );
  OR2_X1 U5623 ( .A1(n5595), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8274) );
  AND2_X1 U5624 ( .A1(n5594), .A2(n5593), .ZN(n5602) );
  NAND2_X1 U5625 ( .A1(n8168), .A2(n8307), .ZN(n4765) );
  NAND2_X1 U5626 ( .A1(n4436), .A2(n4470), .ZN(n4764) );
  NAND2_X1 U5627 ( .A1(n5536), .A2(n5535), .ZN(n5562) );
  OR2_X1 U5628 ( .A1(n5502), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5503) );
  OR2_X1 U5629 ( .A1(n5503), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5519) );
  OR2_X1 U5630 ( .A1(n5452), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5466) );
  OR2_X1 U5631 ( .A1(n5405), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U5632 ( .A1(n5431), .A2(n10241), .ZN(n5452) );
  INV_X1 U5633 ( .A(n5432), .ZN(n5431) );
  NAND2_X1 U5634 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  INV_X1 U5635 ( .A(n8409), .ZN(n4743) );
  AOI21_X1 U5636 ( .B1(n4741), .B2(n4744), .A(n4489), .ZN(n4740) );
  NOR2_X1 U5637 ( .A1(n8409), .A2(n4747), .ZN(n4741) );
  NAND2_X1 U5638 ( .A1(n5346), .A2(n10147), .ZN(n5367) );
  INV_X1 U5639 ( .A(n5289), .ZN(n5288) );
  OR2_X1 U5640 ( .A1(n5271), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5289) );
  INV_X1 U5641 ( .A(n8190), .ZN(n7458) );
  INV_X1 U5642 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5229) );
  INV_X1 U5643 ( .A(n7849), .ZN(n5638) );
  OR2_X1 U5644 ( .A1(n5631), .A2(n7920), .ZN(n7015) );
  OR2_X1 U5645 ( .A1(n5203), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5231) );
  AND2_X1 U5646 ( .A1(n7897), .A2(n7896), .ZN(n7846) );
  OR2_X1 U5647 ( .A1(n5144), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U5648 ( .A1(n5637), .A2(n7907), .ZN(n6748) );
  AND2_X1 U5649 ( .A1(n6868), .A2(n7910), .ZN(n7842) );
  AND2_X1 U5650 ( .A1(n8024), .A2(n8255), .ZN(n6678) );
  NAND2_X1 U5651 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND2_X1 U5652 ( .A1(n8371), .A2(n8370), .ZN(n8369) );
  NAND2_X1 U5653 ( .A1(n6217), .A2(n8005), .ZN(n8394) );
  AND3_X1 U5654 ( .A1(n6655), .A2(n9919), .A3(n5659), .ZN(n9927) );
  OR2_X1 U5655 ( .A1(n5707), .A2(n6649), .ZN(n6215) );
  INV_X1 U5656 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U5657 ( .A1(n4973), .A2(n5043), .ZN(n4971) );
  INV_X1 U5658 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5676) );
  INV_X1 U5659 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5673) );
  INV_X1 U5660 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5024) );
  AND2_X1 U5661 ( .A1(n5023), .A2(n5398), .ZN(n4969) );
  OR2_X1 U5662 ( .A1(n5097), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U5663 ( .A1(n7125), .A2(n4452), .ZN(n7235) );
  INV_X1 U5664 ( .A(n4625), .ZN(n7234) );
  INV_X1 U5665 ( .A(n6466), .ZN(n8681) );
  OR2_X1 U5666 ( .A1(n5860), .A2(n5859), .ZN(n5873) );
  NOR2_X1 U5667 ( .A1(n4451), .A2(n4561), .ZN(n4560) );
  NOR2_X1 U5668 ( .A1(n8663), .A2(n4568), .ZN(n4567) );
  NOR2_X1 U5669 ( .A1(n8762), .A2(n4997), .ZN(n4996) );
  INV_X1 U5670 ( .A(n8590), .ZN(n4997) );
  NOR2_X1 U5671 ( .A1(n6017), .A2(n8764), .ZN(n6019) );
  OR2_X1 U5672 ( .A1(n6027), .A2(n8774), .ZN(n6033) );
  BUF_X1 U5673 ( .A(n6424), .Z(n8629) );
  NOR2_X1 U5674 ( .A1(n4626), .A2(n7234), .ZN(n7237) );
  INV_X1 U5675 ( .A(n4627), .ZN(n4626) );
  NAND2_X1 U5676 ( .A1(n7237), .A2(n7238), .ZN(n7283) );
  NAND2_X1 U5677 ( .A1(n8054), .A2(n8900), .ZN(n8798) );
  NAND2_X1 U5678 ( .A1(n6421), .A2(n4573), .ZN(n6423) );
  NAND2_X1 U5679 ( .A1(n4574), .A2(n6440), .ZN(n4573) );
  AND2_X1 U5680 ( .A1(n4983), .A2(n8639), .ZN(n4982) );
  NAND2_X1 U5681 ( .A1(n8710), .A2(n4984), .ZN(n4983) );
  INV_X1 U5682 ( .A(n8626), .ZN(n4984) );
  INV_X1 U5683 ( .A(n8710), .ZN(n4985) );
  INV_X1 U5684 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U5685 ( .A1(n6098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6152) );
  INV_X1 U5686 ( .A(n8847), .ZN(n9033) );
  AND4_X1 U5687 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n8799)
         );
  AND4_X1 U5688 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n6980)
         );
  AND4_X1 U5689 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n6966)
         );
  AND4_X1 U5690 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n6801)
         );
  OR2_X1 U5691 ( .A1(n6360), .A2(n6575), .ZN(n6261) );
  AOI21_X1 U5692 ( .B1(n4857), .B2(n4860), .A(n4855), .ZN(n4854) );
  INV_X1 U5693 ( .A(n8800), .ZN(n9042) );
  NAND2_X1 U5694 ( .A1(n4654), .A2(n4653), .ZN(n9298) );
  INV_X1 U5695 ( .A(n9294), .ZN(n4653) );
  INV_X1 U5696 ( .A(n4654), .ZN(n9295) );
  OR2_X1 U5697 ( .A1(n6007), .A2(n10167), .ZN(n6017) );
  NAND2_X1 U5698 ( .A1(n9331), .A2(n9336), .ZN(n9330) );
  NAND2_X1 U5699 ( .A1(n5976), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U5700 ( .A1(n7581), .A2(n6122), .ZN(n7584) );
  AND2_X1 U5701 ( .A1(n5963), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5976) );
  INV_X1 U5702 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5936) );
  INV_X1 U5703 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5771) );
  AOI21_X1 U5704 ( .B1(n8849), .B2(n4816), .A(n4485), .ZN(n4815) );
  NAND2_X1 U5705 ( .A1(n7165), .A2(n8867), .ZN(n7164) );
  NOR2_X1 U5706 ( .A1(n5887), .A2(n10200), .ZN(n5900) );
  AOI21_X1 U5707 ( .B1(n6826), .B2(n4811), .A(n4484), .ZN(n4810) );
  NAND2_X1 U5708 ( .A1(n6830), .A2(n4678), .ZN(n7345) );
  NAND2_X1 U5709 ( .A1(n6830), .A2(n6835), .ZN(n6891) );
  NOR2_X1 U5710 ( .A1(n6587), .A2(n6586), .ZN(n6635) );
  AND2_X1 U5711 ( .A1(n6635), .A2(n7111), .ZN(n6830) );
  NAND2_X1 U5712 ( .A1(n7100), .A2(n6516), .ZN(n5004) );
  NOR2_X1 U5713 ( .A1(n6452), .A2(n6469), .ZN(n6520) );
  OR2_X1 U5714 ( .A1(n6440), .A2(n7324), .ZN(n6452) );
  AND2_X1 U5715 ( .A1(n8058), .A2(n4660), .ZN(n4657) );
  NAND2_X1 U5716 ( .A1(n4661), .A2(n9329), .ZN(n4658) );
  OR2_X1 U5717 ( .A1(n8896), .A2(n7686), .ZN(n9352) );
  NAND2_X1 U5718 ( .A1(n6063), .A2(n6062), .ZN(n9362) );
  NAND2_X1 U5719 ( .A1(n6005), .A2(n6004), .ZN(n9399) );
  AND2_X1 U5720 ( .A1(n9310), .A2(n8970), .ZN(n9336) );
  INV_X1 U5721 ( .A(n4783), .ZN(n4782) );
  OAI21_X1 U5722 ( .B1(n4785), .B2(n4784), .A(n5983), .ZN(n4783) );
  NAND2_X1 U5723 ( .A1(n5974), .A2(n5973), .ZN(n8575) );
  NAND2_X1 U5724 ( .A1(n4641), .A2(n5880), .ZN(n6964) );
  NAND2_X1 U5725 ( .A1(n6255), .A2(n5855), .ZN(n4641) );
  NAND2_X1 U5726 ( .A1(n6511), .A2(n6510), .ZN(n6509) );
  XNOR2_X1 U5727 ( .A(n7654), .B(SI_29_), .ZN(n7681) );
  XNOR2_X1 U5728 ( .A(n5570), .B(n5569), .ZN(n7611) );
  XNOR2_X1 U5729 ( .A(n5527), .B(n5553), .ZN(n7599) );
  AND2_X1 U5730 ( .A1(n5548), .A2(n5496), .ZN(n5497) );
  OR2_X1 U5731 ( .A1(n5879), .A2(n5760), .ZN(n5778) );
  INV_X1 U5732 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U5733 ( .A1(n4719), .A2(n4726), .ZN(n5258) );
  OR2_X1 U5734 ( .A1(n5213), .A2(n4729), .ZN(n4719) );
  NOR2_X1 U5735 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4555) );
  NOR2_X1 U5736 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4554) );
  NOR2_X1 U5737 ( .A1(n8065), .A2(n4965), .ZN(n4964) );
  INV_X1 U5738 ( .A(n4967), .ZN(n4965) );
  NAND2_X1 U5739 ( .A1(n4954), .A2(n7766), .ZN(n8074) );
  NAND2_X1 U5740 ( .A1(n7005), .A2(n4940), .ZN(n7049) );
  INV_X1 U5741 ( .A(n9879), .ZN(n5059) );
  AND2_X1 U5742 ( .A1(n7804), .A2(n8093), .ZN(n8095) );
  NOR2_X1 U5743 ( .A1(n7480), .A2(n7482), .ZN(n7481) );
  INV_X1 U5744 ( .A(n4956), .ZN(n4959) );
  NAND2_X1 U5745 ( .A1(n6558), .A2(n4961), .ZN(n6623) );
  NAND2_X1 U5746 ( .A1(n4936), .A2(n4934), .ZN(n7053) );
  NAND2_X1 U5747 ( .A1(n7005), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U5748 ( .A1(n7053), .A2(n7052), .ZN(n7303) );
  NAND2_X1 U5749 ( .A1(n5304), .A2(n5303), .ZN(n9523) );
  OAI22_X1 U5750 ( .A1(n6595), .A2(n6594), .B1(n9867), .B2(n6187), .ZN(n6603)
         );
  AND2_X1 U5751 ( .A1(n6197), .A2(n6196), .ZN(n8160) );
  INV_X1 U5752 ( .A(n8032), .ZN(n4827) );
  AND2_X1 U5753 ( .A1(n6932), .A2(n6931), .ZN(n8273) );
  NAND2_X1 U5754 ( .A1(n5488), .A2(n5487), .ZN(n8361) );
  AND4_X1 U5755 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n7305)
         );
  NAND4_X1 U5756 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n8193)
         );
  NAND2_X1 U5757 ( .A1(n5454), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5150) );
  OR2_X1 U5758 ( .A1(n5084), .A2(n9878), .ZN(n5070) );
  OR2_X1 U5759 ( .A1(n6270), .A2(n6180), .ZN(n8225) );
  NAND2_X1 U5760 ( .A1(n6314), .A2(n6315), .ZN(n6545) );
  NAND2_X1 U5761 ( .A1(n4885), .A2(n6539), .ZN(n9681) );
  NOR2_X1 U5762 ( .A1(n9689), .A2(n4541), .ZN(n6533) );
  AND2_X1 U5763 ( .A1(n6531), .A2(n9688), .ZN(n4541) );
  NAND2_X1 U5764 ( .A1(n6533), .A2(n6532), .ZN(n6688) );
  XNOR2_X1 U5765 ( .A(n7411), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9719) );
  INV_X1 U5766 ( .A(n4882), .ZN(n9738) );
  OR2_X1 U5767 ( .A1(n7419), .A2(n7418), .ZN(n7618) );
  XNOR2_X1 U5768 ( .A(n8201), .B(n8202), .ZN(n7623) );
  NOR2_X1 U5769 ( .A1(n7623), .A2(n5306), .ZN(n8203) );
  AND2_X1 U5770 ( .A1(n5342), .A2(n5328), .ZN(n9793) );
  OAI21_X1 U5771 ( .B1(n9855), .B2(n4900), .A(n4898), .ZN(n8250) );
  NAND2_X1 U5772 ( .A1(n4899), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4900) );
  AND2_X1 U5773 ( .A1(n6279), .A2(n8257), .ZN(n9852) );
  NOR2_X1 U5774 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  NAND2_X1 U5775 ( .A1(n4772), .A2(n4770), .ZN(n7216) );
  AND2_X1 U5776 ( .A1(n5640), .A2(n7931), .ZN(n4922) );
  NAND2_X1 U5777 ( .A1(n4923), .A2(n7931), .ZN(n7084) );
  NAND2_X1 U5778 ( .A1(n5226), .A2(n5225), .ZN(n7050) );
  INV_X1 U5779 ( .A(n6677), .ZN(n8413) );
  INV_X1 U5780 ( .A(n8403), .ZN(n8438) );
  OR2_X1 U5781 ( .A1(n6212), .A2(n6211), .ZN(n9863) );
  OR2_X1 U5782 ( .A1(n6652), .A2(n9864), .ZN(n8403) );
  NAND2_X1 U5783 ( .A1(n7821), .A2(n7820), .ZN(n8481) );
  NAND2_X1 U5784 ( .A1(n8552), .A2(n7822), .ZN(n7821) );
  NAND2_X1 U5785 ( .A1(n7827), .A2(n7826), .ZN(n8485) );
  NAND2_X1 U5786 ( .A1(n8310), .A2(n5656), .ZN(n8290) );
  NAND2_X1 U5787 ( .A1(n4766), .A2(n4436), .ZN(n8319) );
  NAND2_X1 U5788 ( .A1(n4909), .A2(n4911), .ZN(n8317) );
  NAND2_X1 U5789 ( .A1(n4763), .A2(n4767), .ZN(n7776) );
  INV_X1 U5790 ( .A(n4910), .ZN(n7775) );
  AOI21_X1 U5791 ( .B1(n5651), .B2(n5650), .A(n7990), .ZN(n4910) );
  INV_X1 U5792 ( .A(n8327), .ZN(n5651) );
  NAND2_X1 U5793 ( .A1(n5464), .A2(n5463), .ZN(n8513) );
  NAND2_X1 U5794 ( .A1(n5647), .A2(n4435), .ZN(n8356) );
  NAND2_X1 U5795 ( .A1(n5451), .A2(n5450), .ZN(n8518) );
  NAND2_X1 U5796 ( .A1(n5647), .A2(n7959), .ZN(n8368) );
  NAND2_X1 U5797 ( .A1(n5430), .A2(n5429), .ZN(n8523) );
  AND2_X1 U5798 ( .A1(n5403), .A2(n5402), .ZN(n8531) );
  NAND2_X1 U5799 ( .A1(n5383), .A2(n5382), .ZN(n8534) );
  INV_X1 U5800 ( .A(n4739), .ZN(n8410) );
  AOI21_X1 U5801 ( .B1(n8428), .B2(n4747), .A(n4745), .ZN(n4739) );
  NAND2_X1 U5802 ( .A1(n5641), .A2(n7960), .ZN(n8408) );
  AOI21_X1 U5803 ( .B1(n8428), .B2(n7854), .A(n7856), .ZN(n8420) );
  NAND2_X1 U5804 ( .A1(n5345), .A2(n5344), .ZN(n8547) );
  INV_X1 U5805 ( .A(n8530), .ZN(n8546) );
  NAND2_X1 U5806 ( .A1(n4917), .A2(n7947), .ZN(n8427) );
  NAND2_X1 U5807 ( .A1(n7326), .A2(n7948), .ZN(n4917) );
  INV_X2 U5808 ( .A(n9944), .ZN(n9946) );
  AND2_X1 U5809 ( .A1(n6201), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6250) );
  INV_X1 U5810 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8554) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7502) );
  XNOR2_X1 U5812 ( .A(n5623), .B(n5622), .ZN(n7500) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7271) );
  INV_X1 U5814 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7180) );
  INV_X1 U5815 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6976) );
  INV_X1 U5816 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6921) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6810) );
  INV_X1 U5818 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6731) );
  INV_X1 U5819 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6663) );
  INV_X1 U5820 ( .A(n9793), .ZN(n8234) );
  INV_X1 U5821 ( .A(n9776), .ZN(n7637) );
  INV_X1 U5822 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6345) );
  INV_X1 U5823 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6307) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10244) );
  AND2_X1 U5825 ( .A1(n6228), .A2(P2_U3151), .ZN(n8560) );
  INV_X1 U5826 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6238) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6227) );
  INV_X1 U5828 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6226) );
  OR2_X1 U5829 ( .A1(n5053), .A2(n4897), .ZN(n4896) );
  NOR2_X1 U5830 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  NAND2_X1 U5831 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4897) );
  NAND2_X1 U5832 ( .A1(n5055), .A2(n5054), .ZN(n6291) );
  NAND2_X1 U5833 ( .A1(n6075), .A2(n6074), .ZN(n9188) );
  NAND2_X1 U5834 ( .A1(n5934), .A2(n5933), .ZN(n9410) );
  INV_X1 U5835 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U5836 ( .A1(n4565), .A2(n4564), .ZN(n8665) );
  AOI21_X1 U5837 ( .B1(n5006), .B2(n8616), .A(n4572), .ZN(n4564) );
  INV_X1 U5838 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10167) );
  OR2_X1 U5839 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  AND2_X1 U5840 ( .A1(n8650), .A2(n8649), .ZN(n8693) );
  NAND2_X1 U5841 ( .A1(n4990), .A2(n4991), .ZN(n7388) );
  AND2_X1 U5842 ( .A1(n4600), .A2(n4979), .ZN(n8719) );
  AOI22_X1 U5843 ( .A1(n9070), .A2(n8784), .B1(n9042), .B2(n4588), .ZN(n7699)
         );
  NAND2_X1 U5844 ( .A1(n8730), .A2(n8731), .ZN(n8729) );
  NAND2_X1 U5845 ( .A1(n8717), .A2(n8720), .ZN(n8730) );
  INV_X1 U5846 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U5847 ( .A1(n8674), .A2(n8590), .ZN(n8761) );
  NAND2_X1 U5848 ( .A1(n6413), .A2(n9040), .ZN(n8775) );
  NAND2_X1 U5849 ( .A1(n4990), .A2(n4988), .ZN(n4986) );
  INV_X1 U5850 ( .A(n4989), .ZN(n4988) );
  INV_X1 U5851 ( .A(n8775), .ZN(n8805) );
  NAND2_X1 U5852 ( .A1(n4597), .A2(n4595), .ZN(n8783) );
  NOR2_X1 U5853 ( .A1(n4483), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5854 ( .A1(n8709), .A2(n8710), .ZN(n8708) );
  INV_X1 U5855 ( .A(n8794), .ZN(n4548) );
  INV_X1 U5856 ( .A(n8795), .ZN(n4549) );
  OAI21_X1 U5857 ( .B1(n8746), .B2(n4985), .A(n4982), .ZN(n8796) );
  AND2_X1 U5858 ( .A1(n6413), .A2(n6405), .ZN(n8797) );
  NAND2_X1 U5859 ( .A1(n9362), .A2(n8790), .ZN(n4546) );
  INV_X1 U5860 ( .A(n8797), .ZN(n8792) );
  NAND2_X1 U5861 ( .A1(n6578), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8803) );
  NAND2_X1 U5862 ( .A1(n5765), .A2(n5764), .ZN(n7541) );
  INV_X1 U5863 ( .A(n8713), .ZN(n9053) );
  INV_X1 U5864 ( .A(n4588), .ZN(n6516) );
  AND2_X1 U5865 ( .A1(n5794), .A2(n5793), .ZN(n5797) );
  OAI21_X1 U5866 ( .B1(n7708), .B2(n4686), .A(n4684), .ZN(n5007) );
  NAND2_X1 U5867 ( .A1(n4687), .A2(n8844), .ZN(n4686) );
  OAI21_X1 U5868 ( .B1(n7708), .B2(n4688), .A(n4685), .ZN(n4684) );
  OR3_X1 U5869 ( .A1(n9164), .A2(n9163), .A3(n9317), .ZN(n9353) );
  NOR2_X1 U5870 ( .A1(n7708), .A2(n4688), .ZN(n9164) );
  AND2_X1 U5871 ( .A1(n4658), .A2(n4660), .ZN(n8056) );
  NAND2_X1 U5872 ( .A1(n9181), .A2(n9182), .ZN(n9180) );
  NAND2_X1 U5873 ( .A1(n9219), .A2(n6061), .ZN(n9197) );
  NAND2_X1 U5874 ( .A1(n4633), .A2(n4630), .ZN(n9215) );
  NAND2_X1 U5875 ( .A1(n6128), .A2(n9246), .ZN(n9232) );
  NAND2_X1 U5876 ( .A1(n4805), .A2(n4803), .ZN(n9263) );
  NAND2_X1 U5877 ( .A1(n9278), .A2(n4800), .ZN(n4805) );
  NAND2_X1 U5878 ( .A1(n4642), .A2(n4646), .ZN(n7504) );
  OR2_X1 U5879 ( .A1(n7259), .A2(n4648), .ZN(n4642) );
  NAND2_X1 U5880 ( .A1(n4652), .A2(n4650), .ZN(n7489) );
  NAND2_X1 U5881 ( .A1(n5783), .A2(n5782), .ZN(n7363) );
  NAND2_X1 U5882 ( .A1(n4639), .A2(n4638), .ZN(n7035) );
  NAND2_X1 U5883 ( .A1(n7030), .A2(n8849), .ZN(n7029) );
  NAND2_X1 U5884 ( .A1(n6977), .A2(n5907), .ZN(n7030) );
  NAND2_X1 U5885 ( .A1(n6824), .A2(n6826), .ZN(n6823) );
  NAND2_X1 U5886 ( .A1(n6633), .A2(n5858), .ZN(n6824) );
  INV_X1 U5887 ( .A(n9318), .ZN(n9629) );
  INV_X1 U5888 ( .A(n9324), .ZN(n9627) );
  NAND2_X1 U5889 ( .A1(n9624), .A2(n7073), .ZN(n9324) );
  NAND2_X1 U5890 ( .A1(n6113), .A2(n6112), .ZN(n6505) );
  NAND2_X1 U5891 ( .A1(n6441), .A2(n6106), .ZN(n6453) );
  NOR2_X2 U5892 ( .A1(n9321), .A2(n9156), .ZN(n9318) );
  INV_X1 U5893 ( .A(n8692), .ZN(n7705) );
  AND2_X1 U5894 ( .A1(n7691), .A2(n9352), .ZN(n9349) );
  NOR2_X1 U5895 ( .A1(n9176), .A2(n4456), .ZN(n7790) );
  AND2_X1 U5896 ( .A1(n7719), .A2(n9411), .ZN(n4874) );
  OAI21_X1 U5897 ( .B1(n9278), .B2(n4799), .A(n4437), .ZN(n9245) );
  AND2_X1 U5898 ( .A1(n6026), .A2(n6025), .ZN(n9443) );
  NAND2_X1 U5899 ( .A1(n6016), .A2(n6015), .ZN(n9450) );
  NAND2_X1 U5900 ( .A1(n4787), .A2(n4785), .ZN(n7580) );
  NAND2_X1 U5901 ( .A1(n5947), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5902 ( .A1(n5962), .A2(n5961), .ZN(n8726) );
  NAND2_X1 U5903 ( .A1(n5947), .A2(n4791), .ZN(n7554) );
  NAND2_X1 U5904 ( .A1(n5922), .A2(n5921), .ZN(n7382) );
  OR2_X1 U5905 ( .A1(n6237), .A2(n5843), .ZN(n4819) );
  AND2_X1 U5906 ( .A1(n5844), .A2(n4458), .ZN(n4818) );
  AND3_X1 U5907 ( .A1(n5822), .A2(n5821), .A3(n5820), .ZN(n7074) );
  AND3_X1 U5908 ( .A1(n5811), .A2(n5810), .A3(n5809), .ZN(n7090) );
  NOR2_X1 U5909 ( .A1(n9637), .A2(n9636), .ZN(n9664) );
  AND2_X1 U5910 ( .A1(n6360), .A2(n6155), .ZN(n9667) );
  NAND2_X1 U5911 ( .A1(n5745), .A2(n4853), .ZN(n4850) );
  INV_X1 U5912 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5754) );
  OAI21_X1 U5913 ( .B1(n6099), .B2(n5753), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5755) );
  CLKBUF_X1 U5914 ( .A(n6257), .Z(n7819) );
  OR2_X1 U5915 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  XNOR2_X1 U5916 ( .A(n6150), .B(n5738), .ZN(n7601) );
  INV_X1 U5917 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7313) );
  INV_X1 U5918 ( .A(n8822), .ZN(n9035) );
  INV_X1 U5919 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U5920 ( .A1(n5999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6001) );
  INV_X1 U5921 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6808) );
  INV_X1 U5922 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6747) );
  INV_X1 U5923 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5853) );
  INV_X1 U5924 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6236) );
  INV_X1 U5925 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6233) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U5927 ( .A1(n4535), .A2(n9851), .ZN(n4534) );
  XNOR2_X1 U5928 ( .A(n8263), .B(n8264), .ZN(n4535) );
  AOI21_X1 U5929 ( .B1(n7828), .B2(n5724), .A(n5723), .ZN(n5725) );
  OR2_X1 U5930 ( .A1(n8494), .A2(n8550), .ZN(n4516) );
  OAI21_X1 U5931 ( .B1(n4550), .B2(n4547), .A(n4545), .ZN(P1_U3240) );
  AND2_X1 U5932 ( .A1(n8806), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U5933 ( .A1(n8796), .A2(n8797), .ZN(n4550) );
  AOI21_X1 U5934 ( .B1(n8708), .B2(n4549), .A(n4548), .ZN(n4547) );
  OAI21_X1 U5935 ( .B1(n6516), .B2(n6670), .A(n4587), .ZN(P1_U3558) );
  NAND2_X1 U5936 ( .A1(n6670), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4587) );
  AOI21_X1 U5937 ( .B1(n4824), .B2(n4822), .A(n4821), .ZN(n4820) );
  INV_X1 U5938 ( .A(n4824), .ZN(n4823) );
  INV_X1 U5939 ( .A(n4825), .ZN(n4821) );
  INV_X1 U5940 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U5941 ( .A1(n5988), .A2(n5987), .ZN(n9459) );
  INV_X1 U5942 ( .A(n8945), .ZN(n4607) );
  NAND3_X2 U5943 ( .A1(n5039), .A2(n5038), .A3(n5037), .ZN(n9867) );
  AND2_X1 U5944 ( .A1(n7460), .A2(n8190), .ZN(n4433) );
  AND2_X1 U5945 ( .A1(n4566), .A2(n4569), .ZN(n4434) );
  AND2_X1 U5946 ( .A1(n7967), .A2(n7959), .ZN(n4435) );
  OR2_X1 U5947 ( .A1(n8114), .A2(n8331), .ZN(n4436) );
  AND2_X1 U5948 ( .A1(n4798), .A2(n4801), .ZN(n4437) );
  AND2_X1 U5949 ( .A1(n5652), .A2(n8077), .ZN(n7988) );
  AND2_X1 U5950 ( .A1(n4613), .A2(n4612), .ZN(n4438) );
  INV_X1 U5951 ( .A(n7828), .ZN(n8281) );
  NAND2_X1 U5952 ( .A1(n5612), .A2(n5611), .ZN(n7828) );
  AND2_X1 U5953 ( .A1(n9269), .A2(n9055), .ZN(n4439) );
  AND2_X1 U5954 ( .A1(n4992), .A2(n7238), .ZN(n4440) );
  AND3_X1 U5955 ( .A1(n7386), .A2(n4440), .A3(n4618), .ZN(n4441) );
  NAND2_X1 U5956 ( .A1(n7684), .A2(n7683), .ZN(n7719) );
  OR2_X1 U5957 ( .A1(n8540), .A2(n8169), .ZN(n7960) );
  INV_X1 U5958 ( .A(n8077), .ZN(n8341) );
  AND2_X1 U5959 ( .A1(n5525), .A2(n5524), .ZN(n8077) );
  AND2_X1 U5960 ( .A1(n9523), .A2(n8189), .ZN(n4442) );
  AND2_X1 U5961 ( .A1(n8961), .A2(n8960), .ZN(n4443) );
  AND2_X1 U5962 ( .A1(n5297), .A2(SI_12_), .ZN(n4444) );
  OR2_X1 U5963 ( .A1(n4982), .A2(n4449), .ZN(n4445) );
  INV_X1 U5964 ( .A(n8168), .ZN(n8496) );
  AND2_X1 U5965 ( .A1(n5561), .A2(n5560), .ZN(n8168) );
  INV_X1 U5966 ( .A(n7021), .ZN(n4673) );
  AND2_X1 U5967 ( .A1(n4455), .A2(n8739), .ZN(n4446) );
  XNOR2_X1 U5968 ( .A(n5044), .B(n5043), .ZN(n5661) );
  NAND2_X1 U5969 ( .A1(n7506), .A2(n4455), .ZN(n4447) );
  AND4_X1 U5970 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n7462)
         );
  NOR2_X1 U5971 ( .A1(n8850), .A2(n6825), .ZN(n4448) );
  INV_X1 U5972 ( .A(n8210), .ZN(n4899) );
  XNOR2_X1 U5973 ( .A(n5426), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8255) );
  INV_X1 U5975 ( .A(n5940), .ZN(n6044) );
  OR2_X1 U5976 ( .A1(n8656), .A2(n8655), .ZN(n4449) );
  NAND2_X1 U5977 ( .A1(n7677), .A2(n7671), .ZN(n5805) );
  OR2_X1 U5979 ( .A1(n6095), .A2(n8881), .ZN(n4450) );
  INV_X1 U5980 ( .A(n7929), .ZN(n4700) );
  NAND2_X1 U5981 ( .A1(n5729), .A2(n5728), .ZN(n5828) );
  AND2_X1 U5982 ( .A1(n4994), .A2(n4459), .ZN(n4451) );
  AND2_X1 U5983 ( .A1(n7123), .A2(n7124), .ZN(n4452) );
  XNOR2_X1 U5984 ( .A(n5755), .B(n5754), .ZN(n9474) );
  INV_X1 U5985 ( .A(n9715), .ZN(n7433) );
  NAND2_X1 U5986 ( .A1(n4763), .A2(n4761), .ZN(n4766) );
  INV_X1 U5987 ( .A(n5214), .ZN(n4728) );
  AND2_X1 U5988 ( .A1(n7530), .A2(n7529), .ZN(n4453) );
  INV_X1 U5989 ( .A(n9003), .ZN(n4859) );
  OR2_X1 U5990 ( .A1(n9379), .A2(n9054), .ZN(n4454) );
  AND2_X1 U5991 ( .A1(n7562), .A2(n7511), .ZN(n4455) );
  NAND2_X1 U5992 ( .A1(n6156), .A2(n6151), .ZN(n6360) );
  INV_X1 U5993 ( .A(n8971), .ZN(n4869) );
  INV_X1 U5994 ( .A(n9000), .ZN(n4632) );
  OR2_X1 U5995 ( .A1(n9169), .A2(n4874), .ZN(n4456) );
  INV_X1 U5996 ( .A(n7837), .ZN(n7833) );
  XNOR2_X1 U5997 ( .A(n5625), .B(n5025), .ZN(n7837) );
  NAND2_X1 U5998 ( .A1(n6041), .A2(n6040), .ZN(n9432) );
  INV_X1 U5999 ( .A(n9432), .ZN(n9242) );
  AND2_X1 U6000 ( .A1(n6293), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U6001 ( .A1(n5749), .A2(n5748), .ZN(n9390) );
  OR2_X1 U6002 ( .A1(n7677), .A2(n9099), .ZN(n4458) );
  AND2_X1 U6003 ( .A1(n8613), .A2(n8612), .ZN(n4459) );
  AND4_X1 U6004 ( .A1(n7868), .A2(n7867), .A3(n7866), .A4(n7865), .ZN(n4460)
         );
  AND3_X1 U6005 ( .A1(n8999), .A2(n9221), .A3(n6129), .ZN(n4461) );
  NAND2_X1 U6006 ( .A1(n4966), .A2(n4964), .ZN(n8063) );
  INV_X1 U6007 ( .A(n8937), .ZN(n4651) );
  AND2_X1 U6008 ( .A1(n8963), .A2(n8938), .ZN(n4462) );
  NAND2_X2 U6009 ( .A1(n9472), .A2(n9474), .ZN(n5835) );
  OR2_X1 U6010 ( .A1(n5080), .A2(n6329), .ZN(n4463) );
  INV_X1 U6011 ( .A(n7569), .ZN(n4953) );
  AND3_X1 U6012 ( .A1(n7834), .A2(n7833), .A3(n7832), .ZN(n4464) );
  AND3_X1 U6013 ( .A1(n5676), .A2(n5673), .A3(n5703), .ZN(n4465) );
  AND2_X1 U6014 ( .A1(n8595), .A2(n8594), .ZN(n4466) );
  AND2_X1 U6015 ( .A1(n8578), .A2(n8577), .ZN(n4467) );
  NAND2_X1 U6016 ( .A1(n6032), .A2(n6031), .ZN(n9379) );
  NAND2_X1 U6017 ( .A1(n4966), .A2(n4967), .ZN(n8064) );
  NAND2_X1 U6018 ( .A1(n4969), .A2(n5024), .ZN(n5626) );
  AND2_X1 U6019 ( .A1(n7964), .A2(n7958), .ZN(n4468) );
  AND2_X1 U6020 ( .A1(n4497), .A2(n5025), .ZN(n4469) );
  INV_X1 U6021 ( .A(n4806), .ZN(n4800) );
  OR2_X1 U6022 ( .A1(n8168), .A2(n8307), .ZN(n4470) );
  OR2_X1 U6023 ( .A1(n8531), .A2(n8382), .ZN(n4471) );
  AND2_X1 U6024 ( .A1(n7964), .A2(n8005), .ZN(n4472) );
  AND2_X1 U6025 ( .A1(n8038), .A2(n8331), .ZN(n4473) );
  AND2_X1 U6026 ( .A1(n6139), .A2(n8799), .ZN(n4474) );
  INV_X1 U6027 ( .A(n5982), .ZN(n4784) );
  AND2_X1 U6028 ( .A1(n5657), .A2(n5656), .ZN(n4475) );
  AND2_X1 U6029 ( .A1(n9362), .A2(n9051), .ZN(n4476) );
  AND2_X1 U6030 ( .A1(n4987), .A2(n7527), .ZN(n4477) );
  AND4_X1 U6031 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n6791)
         );
  AND2_X1 U6032 ( .A1(n4446), .A2(n9344), .ZN(n4478) );
  AND2_X1 U6033 ( .A1(n7983), .A2(n7985), .ZN(n4479) );
  AND2_X1 U6034 ( .A1(n4615), .A2(n4614), .ZN(n4480) );
  NAND3_X1 U6035 ( .A1(n8025), .A2(n8265), .A3(n8024), .ZN(n4481) );
  NOR2_X1 U6036 ( .A1(n7705), .A2(n9442), .ZN(n4482) );
  NOR2_X1 U6037 ( .A1(n4976), .A2(n4601), .ZN(n4483) );
  INV_X1 U6038 ( .A(n4792), .ZN(n4791) );
  NOR2_X1 U6039 ( .A1(n7511), .A2(n7491), .ZN(n4792) );
  NOR2_X1 U6040 ( .A1(n9626), .A2(n9069), .ZN(n4484) );
  INV_X1 U6041 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5049) );
  INV_X1 U6042 ( .A(n4804), .ZN(n4803) );
  NOR2_X1 U6043 ( .A1(n9290), .A2(n8814), .ZN(n4804) );
  INV_X1 U6044 ( .A(n7100), .ZN(n8754) );
  AND3_X1 U6045 ( .A1(n5832), .A2(n5831), .A3(n5830), .ZN(n7100) );
  INV_X1 U6046 ( .A(n4762), .ZN(n4761) );
  NAND2_X1 U6047 ( .A1(n4491), .A2(n4767), .ZN(n4762) );
  NOR2_X1 U6048 ( .A1(n7229), .A2(n9065), .ZN(n4485) );
  AND2_X1 U6049 ( .A1(n9233), .A2(n8994), .ZN(n4486) );
  NAND2_X1 U6050 ( .A1(n8039), .A2(n8103), .ZN(n8106) );
  NAND2_X1 U6051 ( .A1(n5417), .A2(n5416), .ZN(n4487) );
  INV_X1 U6052 ( .A(n4938), .ZN(n4937) );
  NAND2_X1 U6053 ( .A1(n4939), .A2(n4940), .ZN(n4938) );
  OR2_X1 U6054 ( .A1(n4449), .A2(n4985), .ZN(n4488) );
  INV_X1 U6055 ( .A(n4604), .ZN(n4603) );
  NAND2_X1 U6056 ( .A1(n4977), .A2(n4508), .ZN(n4604) );
  NOR2_X1 U6057 ( .A1(n8134), .A2(n8395), .ZN(n4489) );
  INV_X1 U6058 ( .A(n4802), .ZN(n4799) );
  NOR2_X1 U6059 ( .A1(n4439), .A2(n4804), .ZN(n4802) );
  AND2_X1 U6060 ( .A1(n5256), .A2(SI_10_), .ZN(n4490) );
  OR2_X1 U6061 ( .A1(n8038), .A2(n8321), .ZN(n4491) );
  OR2_X1 U6062 ( .A1(n8518), .A2(n8383), .ZN(n7967) );
  INV_X1 U6063 ( .A(n8501), .ZN(n5652) );
  AND2_X1 U6064 ( .A1(n5516), .A2(n5515), .ZN(n8501) );
  NAND2_X1 U6065 ( .A1(n6752), .A2(n6191), .ZN(n4960) );
  OR2_X1 U6066 ( .A1(n8481), .A2(n8273), .ZN(n8021) );
  AND2_X1 U6067 ( .A1(n9012), .A2(n8809), .ZN(n8881) );
  NOR2_X1 U6068 ( .A1(n7677), .A2(n6373), .ZN(n4492) );
  AND2_X1 U6069 ( .A1(n4680), .A2(n9242), .ZN(n4493) );
  NAND2_X1 U6070 ( .A1(n8106), .A2(n8041), .ZN(n8157) );
  AND2_X1 U6071 ( .A1(n4788), .A2(n5982), .ZN(n4494) );
  INV_X1 U6072 ( .A(n9167), .ZN(n9420) );
  NAND2_X1 U6073 ( .A1(n7680), .A2(n7679), .ZN(n9167) );
  NAND2_X1 U6074 ( .A1(n4563), .A2(n5006), .ZN(n8770) );
  INV_X1 U6075 ( .A(n4847), .ZN(n4846) );
  NOR2_X1 U6076 ( .A1(n5298), .A2(n4848), .ZN(n4847) );
  NOR2_X1 U6077 ( .A1(n4777), .A2(n9182), .ZN(n4776) );
  NAND2_X1 U6078 ( .A1(n8496), .A2(n8307), .ZN(n4495) );
  INV_X1 U6079 ( .A(n4730), .ZN(n4729) );
  AND2_X1 U6080 ( .A1(n4731), .A2(n5219), .ZN(n4730) );
  AND2_X1 U6081 ( .A1(n4903), .A2(n4902), .ZN(n4496) );
  AND2_X1 U6082 ( .A1(n8115), .A2(n8116), .ZN(n7730) );
  INV_X1 U6083 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5747) );
  INV_X1 U6084 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5013) );
  INV_X1 U6085 ( .A(n6072), .ZN(n4780) );
  AND2_X1 U6086 ( .A1(n5024), .A2(n4970), .ZN(n4497) );
  AND2_X2 U6087 ( .A1(n6422), .A2(n6361), .ZN(n8630) );
  NAND2_X1 U6088 ( .A1(n7235), .A2(n7236), .ZN(n4627) );
  AND2_X1 U6089 ( .A1(n8175), .A2(n7730), .ZN(n4498) );
  INV_X1 U6090 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4925) );
  INV_X1 U6091 ( .A(n8849), .ZN(n4817) );
  AND2_X1 U6092 ( .A1(n7506), .A2(n4446), .ZN(n4499) );
  NAND2_X1 U6093 ( .A1(n6349), .A2(n8885), .ZN(n6350) );
  INV_X1 U6094 ( .A(n8855), .ZN(n4808) );
  AOI21_X1 U6095 ( .B1(n7457), .B2(n7456), .A(n7455), .ZN(n7480) );
  INV_X1 U6096 ( .A(n8962), .ZN(n4586) );
  OR2_X1 U6097 ( .A1(n6139), .A2(n9387), .ZN(n4500) );
  INV_X1 U6098 ( .A(n8307), .ZN(n8187) );
  AND2_X1 U6099 ( .A1(n5568), .A2(n5567), .ZN(n8307) );
  INV_X1 U6100 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U6101 ( .A1(n5509), .A2(n5508), .ZN(n8188) );
  INV_X1 U6102 ( .A(n8188), .ZN(n8332) );
  NOR2_X1 U6103 ( .A1(n6118), .A2(n8850), .ZN(n4501) );
  AND2_X1 U6104 ( .A1(n4986), .A2(n7386), .ZN(n4502) );
  NOR2_X1 U6105 ( .A1(n9769), .A2(n7621), .ZN(n4503) );
  NOR2_X1 U6106 ( .A1(n8203), .A2(n8204), .ZN(n4504) );
  INV_X1 U6107 ( .A(n8383), .ZN(n8360) );
  AND3_X1 U6108 ( .A1(n5458), .A2(n5457), .A3(n5456), .ZN(n8383) );
  INV_X1 U6109 ( .A(n6937), .ZN(n8194) );
  AND4_X1 U6110 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n6937)
         );
  NAND2_X1 U6111 ( .A1(n9283), .A2(n4682), .ZN(n4683) );
  AND2_X1 U6112 ( .A1(n8674), .A2(n4996), .ZN(n4505) );
  OR2_X1 U6113 ( .A1(n7434), .A2(n7433), .ZN(n4506) );
  INV_X1 U6114 ( .A(n7568), .ZN(n8189) );
  AND4_X1 U6115 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n7568)
         );
  NOR2_X1 U6116 ( .A1(n7481), .A2(n4433), .ZN(n4507) );
  NAND2_X4 U6117 ( .A1(n6184), .A2(n6183), .ZN(n7735) );
  INV_X1 U6118 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4591) );
  INV_X1 U6119 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4592) );
  INV_X1 U6120 ( .A(n8007), .ZN(n8005) );
  NAND2_X1 U6121 ( .A1(n8030), .A2(n7833), .ZN(n8007) );
  INV_X1 U6122 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5327) );
  INV_X1 U6123 ( .A(n9825), .ZN(n8232) );
  OAI21_X1 U6124 ( .B1(n6673), .B2(n6185), .A(n7879), .ZN(n9862) );
  OR2_X1 U6125 ( .A1(n8573), .A2(n8572), .ZN(n4508) );
  XOR2_X1 U6126 ( .A(n8565), .B(n8566), .Z(n4509) );
  INV_X1 U6127 ( .A(n6273), .ZN(n8213) );
  INV_X1 U6128 ( .A(n5661), .ZN(n6273) );
  AND2_X1 U6129 ( .A1(n6558), .A2(n4959), .ZN(n4510) );
  NOR2_X1 U6130 ( .A1(n5555), .A2(n5554), .ZN(n4511) );
  NAND4_X2 U6131 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n8195)
         );
  INV_X1 U6132 ( .A(n8195), .ZN(n4733) );
  AND2_X1 U6133 ( .A1(n7069), .A2(n9414), .ZN(n9368) );
  NAND2_X1 U6134 ( .A1(n5628), .A2(n5624), .ZN(n8024) );
  INV_X1 U6135 ( .A(n8255), .ZN(n8265) );
  NAND2_X1 U6136 ( .A1(n4674), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U6137 ( .A1(n8418), .A2(n7957), .ZN(n5641) );
  NAND2_X1 U6138 ( .A1(n6886), .A2(n7924), .ZN(n7040) );
  NAND2_X1 U6139 ( .A1(n4828), .A2(n4699), .ZN(n4698) );
  INV_X1 U6140 ( .A(n4835), .ZN(n4834) );
  NAND3_X1 U6141 ( .A1(n4513), .A2(n4529), .A3(n4481), .ZN(n4530) );
  NAND2_X1 U6142 ( .A1(n4521), .A2(n4698), .ZN(n4513) );
  NAND3_X1 U6143 ( .A1(n7834), .A2(n8021), .A3(n4460), .ZN(n4526) );
  NAND2_X1 U6144 ( .A1(n5417), .A2(n4849), .ZN(n5440) );
  NAND2_X1 U6145 ( .A1(n4904), .A2(n4834), .ZN(n5187) );
  OAI21_X1 U6146 ( .B1(n5478), .B2(n5477), .A(n5476), .ZN(n5492) );
  NAND2_X1 U6147 ( .A1(n4631), .A2(n4629), .ZN(n9206) );
  NAND2_X1 U6148 ( .A1(n9360), .A2(n4500), .ZN(P1_U3549) );
  NAND2_X1 U6149 ( .A1(n5462), .A2(n5461), .ZN(n5478) );
  NAND2_X1 U6150 ( .A1(n5395), .A2(n5394), .ZN(n5413) );
  OAI21_X1 U6151 ( .B1(n5492), .B2(n5491), .A(n5490), .ZN(n5498) );
  INV_X1 U6152 ( .A(n4766), .ZN(n4755) );
  NAND2_X1 U6153 ( .A1(n9906), .A2(n8195), .ZN(n7914) );
  NAND2_X1 U6154 ( .A1(n8493), .A2(n4516), .ZN(P2_U3454) );
  NAND2_X1 U6155 ( .A1(n4769), .A2(n4768), .ZN(n7328) );
  NOR2_X1 U6156 ( .A1(n8451), .A2(n4517), .ZN(n8491) );
  NAND2_X1 U6157 ( .A1(n5151), .A2(SI_5_), .ZN(n4906) );
  NAND2_X1 U6158 ( .A1(n4732), .A2(n5181), .ZN(n6813) );
  NOR2_X2 U6159 ( .A1(n8428), .A2(n4742), .ZN(n4738) );
  AOI21_X1 U6160 ( .B1(n7411), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7410), .ZN(
        n9740) );
  NOR2_X1 U6161 ( .A1(n9834), .A2(n4519), .ZN(n8208) );
  INV_X1 U6162 ( .A(n4537), .ZN(n4536) );
  INV_X1 U6163 ( .A(n6536), .ZN(n4886) );
  XNOR2_X1 U6164 ( .A(n5213), .B(n5212), .ZN(n6255) );
  NAND2_X1 U6165 ( .A1(n8288), .A2(n5658), .ZN(n7831) );
  NAND2_X1 U6166 ( .A1(n7213), .A2(n7943), .ZN(n4662) );
  NAND2_X1 U6167 ( .A1(n5187), .A2(n5186), .ZN(n4833) );
  NAND2_X1 U6168 ( .A1(n4909), .A2(n4908), .ZN(n5653) );
  NAND2_X1 U6169 ( .A1(n4671), .A2(n4669), .ZN(n7017) );
  NAND2_X1 U6170 ( .A1(n7793), .A2(n7977), .ZN(n4927) );
  OR2_X2 U6171 ( .A1(n4828), .A2(n8265), .ZN(n4521) );
  NAND2_X1 U6172 ( .A1(n6585), .A2(n8856), .ZN(n6584) );
  INV_X1 U6173 ( .A(n9309), .ZN(n6014) );
  INV_X1 U6174 ( .A(n9293), .ZN(n6023) );
  NAND2_X1 U6175 ( .A1(n4658), .A2(n4656), .ZN(n6177) );
  NAND2_X1 U6176 ( .A1(n4430), .A2(n5737), .ZN(n6101) );
  OAI22_X1 U6177 ( .A1(n4925), .A2(n5805), .B1(n5843), .B2(n6229), .ZN(n4689)
         );
  INV_X1 U6178 ( .A(n7015), .ZN(n4674) );
  OAI21_X1 U6179 ( .B1(n4666), .B2(n4528), .A(n4464), .ZN(n4527) );
  NAND2_X1 U6180 ( .A1(n4527), .A2(n4526), .ZN(n8026) );
  NAND2_X1 U6181 ( .A1(n5498), .A2(n5497), .ZN(n5550) );
  NAND2_X1 U6182 ( .A1(n5319), .A2(n5318), .ZN(n5341) );
  NAND2_X1 U6183 ( .A1(n9736), .A2(n9735), .ZN(n9734) );
  NAND2_X1 U6184 ( .A1(n7423), .A2(n7433), .ZN(n4523) );
  NAND2_X1 U6185 ( .A1(n9716), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U6186 ( .A1(n4536), .A2(n4534), .ZN(P2_U3201) );
  OAI21_X1 U6187 ( .B1(n8270), .B2(n9856), .A(n4538), .ZN(n4537) );
  INV_X1 U6188 ( .A(n6714), .ZN(n6716) );
  AND2_X1 U6189 ( .A1(n6712), .A2(n9707), .ZN(n4525) );
  NOR2_X1 U6190 ( .A1(n4730), .A2(n5257), .ZN(n4721) );
  NAND2_X1 U6191 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  INV_X4 U6192 ( .A(n5078), .ZN(n6228) );
  NAND2_X1 U6193 ( .A1(n8019), .A2(n8020), .ZN(n4691) );
  NAND2_X1 U6194 ( .A1(n4668), .A2(n4828), .ZN(n4529) );
  INV_X1 U6195 ( .A(n7830), .ZN(n4667) );
  NAND2_X1 U6196 ( .A1(n5448), .A2(n5447), .ZN(n5462) );
  NAND2_X1 U6197 ( .A1(n8026), .A2(n5629), .ZN(n4828) );
  NAND3_X1 U6198 ( .A1(n7955), .A2(n8419), .A3(n7954), .ZN(n7956) );
  NAND2_X1 U6199 ( .A1(n4530), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U6200 ( .A1(n4830), .A2(n4829), .ZN(n8017) );
  NAND2_X1 U6201 ( .A1(n4692), .A2(n4691), .ZN(n4690) );
  NOR2_X1 U6202 ( .A1(n4714), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U6203 ( .A1(n7974), .A2(n8005), .ZN(n4710) );
  INV_X1 U6204 ( .A(n4695), .ZN(n4694) );
  INV_X1 U6205 ( .A(n4969), .ZN(n5425) );
  INV_X1 U6206 ( .A(n6637), .ZN(n4543) );
  NAND2_X1 U6207 ( .A1(n4861), .A2(n4863), .ZN(n4544) );
  INV_X1 U6208 ( .A(n5729), .ZN(n5826) );
  NAND2_X2 U6209 ( .A1(n4558), .A2(n5756), .ZN(n5940) );
  INV_X1 U6210 ( .A(n4995), .ZN(n4559) );
  NAND2_X1 U6211 ( .A1(n4995), .A2(n4994), .ZN(n8699) );
  OR2_X1 U6212 ( .A1(n8699), .A2(n8616), .ZN(n4563) );
  NAND2_X1 U6213 ( .A1(n8699), .A2(n5006), .ZN(n4565) );
  INV_X1 U6214 ( .A(n8772), .ZN(n4572) );
  INV_X2 U6215 ( .A(n6440), .ZN(n8820) );
  AND3_X1 U6216 ( .A1(n4594), .A2(n6142), .A3(n5738), .ZN(n5743) );
  NAND3_X1 U6217 ( .A1(n7535), .A2(n4599), .A3(n7545), .ZN(n4597) );
  NAND3_X1 U6218 ( .A1(n7535), .A2(n7545), .A3(n4603), .ZN(n4598) );
  NAND3_X1 U6219 ( .A1(n7535), .A2(n7545), .A3(n4977), .ZN(n4600) );
  INV_X1 U6220 ( .A(n8918), .ZN(n4605) );
  INV_X1 U6221 ( .A(n9020), .ZN(n4616) );
  NAND3_X1 U6222 ( .A1(n4625), .A2(n4440), .A3(n4627), .ZN(n4990) );
  NAND2_X1 U6223 ( .A1(n9247), .A2(n4633), .ZN(n4629) );
  INV_X1 U6224 ( .A(n8851), .ZN(n4640) );
  INV_X1 U6225 ( .A(n8928), .ZN(n4637) );
  NAND3_X1 U6226 ( .A1(n4640), .A2(n6825), .A3(n6118), .ZN(n4639) );
  NAND3_X1 U6227 ( .A1(n4639), .A2(n4638), .A3(n4817), .ZN(n7033) );
  AOI21_X1 U6228 ( .B1(n6118), .B2(n6825), .A(n8850), .ZN(n6979) );
  NAND2_X1 U6229 ( .A1(n7259), .A2(n4646), .ZN(n4645) );
  XNOR2_X1 U6230 ( .A(n7709), .B(n8881), .ZN(n4661) );
  INV_X1 U6231 ( .A(n8688), .ZN(n4660) );
  NAND3_X1 U6232 ( .A1(n6811), .A2(n7914), .A3(n4672), .ZN(n4671) );
  INV_X1 U6233 ( .A(n4679), .ZN(n6983) );
  INV_X1 U6234 ( .A(n4683), .ZN(n9268) );
  NOR2_X1 U6235 ( .A1(n7708), .A2(n7719), .ZN(n9162) );
  NOR2_X1 U6236 ( .A1(n4690), .A2(n8018), .ZN(n8023) );
  OAI21_X1 U6237 ( .B1(n8017), .B2(n4697), .A(n4696), .ZN(n4695) );
  INV_X1 U6238 ( .A(n8015), .ZN(n4696) );
  NAND3_X1 U6239 ( .A1(n7933), .A2(n7932), .A3(n4700), .ZN(n7935) );
  NAND2_X1 U6240 ( .A1(n7937), .A2(n7935), .ZN(n7936) );
  NAND2_X1 U6241 ( .A1(n4708), .A2(n4479), .ZN(n4707) );
  NOR2_X1 U6242 ( .A1(n4717), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U6243 ( .A1(n4734), .A2(n4733), .ZN(n7911) );
  XNOR2_X1 U6244 ( .A(n5619), .B(n7867), .ZN(n4735) );
  NOR2_X2 U6245 ( .A1(n8280), .A2(n5010), .ZN(n5727) );
  INV_X1 U6246 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6247 ( .A1(n4737), .A2(n4740), .ZN(n8391) );
  NAND2_X1 U6248 ( .A1(n8328), .A2(n4754), .ZN(n4753) );
  OAI21_X2 U6249 ( .B1(n4755), .B2(n4764), .A(n4765), .ZN(n8304) );
  NAND2_X1 U6250 ( .A1(n7080), .A2(n4770), .ZN(n4769) );
  NAND2_X1 U6251 ( .A1(n7328), .A2(n7853), .ZN(n7327) );
  OAI22_X2 U6252 ( .A1(n7794), .A2(n7861), .B1(n8361), .B2(n5489), .ZN(n8339)
         );
  AOI21_X2 U6253 ( .B1(n8359), .B2(n8358), .A(n5472), .ZN(n7794) );
  NAND2_X1 U6254 ( .A1(n6815), .A2(n5184), .ZN(n6842) );
  NOR2_X2 U6255 ( .A1(n8379), .A2(n5012), .ZN(n8371) );
  OAI21_X2 U6256 ( .B1(n6880), .B2(n5253), .A(n5252), .ZN(n7041) );
  OAI21_X1 U6257 ( .B1(n8298), .B2(n9873), .A(n8297), .ZN(n8447) );
  OR2_X1 U6258 ( .A1(n5146), .A2(n10212), .ZN(n5033) );
  NOR2_X4 U6259 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5053) );
  NAND2_X1 U6260 ( .A1(n5620), .A2(n5622), .ZN(n5671) );
  AOI21_X2 U6261 ( .B1(n6872), .B2(n5183), .A(n5182), .ZN(n6815) );
  OAI22_X2 U6262 ( .A1(n8339), .A2(n5510), .B1(n5649), .B2(n8332), .ZN(n8328)
         );
  NOR2_X2 U6263 ( .A1(n8380), .A2(n8381), .ZN(n8379) );
  NAND2_X1 U6264 ( .A1(n5028), .A2(n5029), .ZN(n8553) );
  NOR2_X1 U6265 ( .A1(n6813), .A2(n7916), .ZN(n5182) );
  NAND2_X1 U6266 ( .A1(n5060), .A2(n5059), .ZN(n5634) );
  NAND2_X2 U6267 ( .A1(n5179), .A2(n5178), .ZN(n6952) );
  NAND2_X1 U6268 ( .A1(n9186), .A2(n6139), .ZN(n6140) );
  NAND2_X1 U6269 ( .A1(n9219), .A2(n4776), .ZN(n4774) );
  NAND2_X1 U6270 ( .A1(n4774), .A2(n4775), .ZN(n6095) );
  OAI21_X1 U6271 ( .B1(n9219), .B2(n4780), .A(n4778), .ZN(n9179) );
  NAND2_X1 U6272 ( .A1(n5947), .A2(n4494), .ZN(n4781) );
  NAND2_X1 U6273 ( .A1(n4781), .A2(n4782), .ZN(n9335) );
  NOR2_X1 U6274 ( .A1(n9390), .A2(n9056), .ZN(n4806) );
  NAND2_X1 U6275 ( .A1(n6634), .A2(n4807), .ZN(n4809) );
  NAND2_X1 U6276 ( .A1(n4809), .A2(n4810), .ZN(n6890) );
  INV_X1 U6277 ( .A(n6826), .ZN(n4812) );
  NAND2_X1 U6278 ( .A1(n6978), .A2(n4814), .ZN(n4813) );
  NAND2_X1 U6279 ( .A1(n4813), .A2(n4815), .ZN(n7165) );
  OAI21_X1 U6280 ( .B1(n8062), .B2(n4823), .A(n4820), .ZN(P1_U3518) );
  NAND2_X1 U6281 ( .A1(n4826), .A2(n8031), .ZN(P2_U3296) );
  NAND3_X1 U6282 ( .A1(n7997), .A2(n8002), .A3(n8318), .ZN(n4830) );
  INV_X1 U6283 ( .A(n8308), .ZN(n4832) );
  NAND2_X1 U6284 ( .A1(n5358), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U6285 ( .A1(n5265), .A2(n4847), .ZN(n4842) );
  NAND2_X1 U6286 ( .A1(n5440), .A2(n5439), .ZN(n5448) );
  INV_X1 U6287 ( .A(n5448), .ZN(n5445) );
  NAND2_X1 U6288 ( .A1(n9467), .A2(n4853), .ZN(n4851) );
  INV_X1 U6289 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4853) );
  OAI21_X1 U6290 ( .B1(n9207), .B2(n4860), .A(n4857), .ZN(n7709) );
  NAND2_X1 U6291 ( .A1(n4856), .A2(n4854), .ZN(n7710) );
  NAND2_X1 U6292 ( .A1(n9207), .A2(n4857), .ZN(n4856) );
  AOI21_X1 U6293 ( .B1(n4864), .B2(n4867), .A(n4862), .ZN(n4861) );
  NAND2_X1 U6294 ( .A1(n6113), .A2(n4864), .ZN(n4863) );
  OAI21_X1 U6295 ( .B1(n6113), .B2(n4867), .A(n4864), .ZN(n8913) );
  NAND3_X1 U6296 ( .A1(n4879), .A2(n6111), .A3(n4877), .ZN(n6515) );
  NAND3_X1 U6297 ( .A1(n8853), .A2(n8823), .A3(n6725), .ZN(n4879) );
  INV_X1 U6298 ( .A(n6699), .ZN(n6702) );
  NAND2_X1 U6299 ( .A1(n4884), .A2(n6539), .ZN(n6537) );
  OAI21_X1 U6300 ( .B1(n7623), .B2(n4888), .A(n4887), .ZN(n9802) );
  NAND2_X1 U6301 ( .A1(n7621), .A2(n4892), .ZN(n4890) );
  NAND2_X2 U6302 ( .A1(n4896), .A2(n4893), .ZN(n6543) );
  INV_X1 U6303 ( .A(n8209), .ZN(n4902) );
  NAND2_X1 U6304 ( .A1(n8209), .A2(n4899), .ZN(n4898) );
  INV_X1 U6305 ( .A(n4903), .ZN(n9854) );
  NAND2_X1 U6306 ( .A1(n5151), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U6307 ( .A1(n4906), .A2(n5155), .ZN(n5171) );
  NAND2_X1 U6308 ( .A1(n7326), .A2(n4918), .ZN(n4914) );
  NAND2_X1 U6309 ( .A1(n4914), .A2(n4915), .ZN(n8418) );
  INV_X1 U6310 ( .A(n6884), .ZN(n5639) );
  NAND2_X1 U6311 ( .A1(n7017), .A2(n7922), .ZN(n6884) );
  XNOR2_X1 U6312 ( .A(n5075), .B(SI_1_), .ZN(n5072) );
  NAND2_X1 U6313 ( .A1(n5641), .A2(n4926), .ZN(n8398) );
  NAND2_X1 U6314 ( .A1(n8398), .A2(n5645), .ZN(n5646) );
  OAI21_X2 U6315 ( .B1(n8338), .B2(n7976), .A(n7978), .ZN(n8327) );
  NAND4_X1 U6316 ( .A1(n10016), .A2(n5300), .A3(n5221), .A4(n4928), .ZN(n5021)
         );
  NAND2_X1 U6317 ( .A1(n7005), .A2(n4930), .ZN(n4929) );
  NAND2_X1 U6318 ( .A1(n4941), .A2(n4942), .ZN(n7734) );
  NAND2_X1 U6319 ( .A1(n8178), .A2(n7730), .ZN(n4941) );
  AOI21_X2 U6320 ( .B1(n4945), .B2(n4944), .A(n4946), .ZN(n7572) );
  NAND3_X1 U6321 ( .A1(n4954), .A2(n7766), .A3(n8332), .ZN(n7767) );
  NAND2_X1 U6322 ( .A1(n7761), .A2(n7760), .ZN(n7766) );
  NAND2_X1 U6323 ( .A1(n7759), .A2(n7758), .ZN(n4954) );
  NAND3_X1 U6324 ( .A1(n6560), .A2(n6559), .A3(n4960), .ZN(n4957) );
  AND2_X1 U6325 ( .A1(n5063), .A2(n5062), .ZN(n4963) );
  INV_X1 U6326 ( .A(n6185), .ZN(n6186) );
  NAND3_X1 U6327 ( .A1(n4962), .A2(n5061), .A3(n5064), .ZN(n6185) );
  AND3_X1 U6328 ( .A1(n5063), .A2(n5062), .A3(n5633), .ZN(n4962) );
  NAND3_X1 U6329 ( .A1(n4963), .A2(n5061), .A3(n5064), .ZN(n5632) );
  INV_X1 U6330 ( .A(n5633), .ZN(n6654) );
  NOR2_X1 U6331 ( .A1(n5679), .A2(n4971), .ZN(n5040) );
  NOR2_X2 U6332 ( .A1(n5679), .A2(n4972), .ZN(n5028) );
  NAND3_X1 U6333 ( .A1(n5043), .A2(n4973), .A3(n5041), .ZN(n4972) );
  INV_X1 U6334 ( .A(n8783), .ZN(n8582) );
  NAND2_X1 U6335 ( .A1(n7535), .A2(n7545), .ZN(n4981) );
  INV_X1 U6336 ( .A(n8566), .ZN(n4980) );
  XNOR2_X1 U6337 ( .A(n4981), .B(n4509), .ZN(n7543) );
  NAND2_X1 U6338 ( .A1(n8746), .A2(n8626), .ZN(n8709) );
  INV_X1 U6339 ( .A(n7281), .ZN(n4992) );
  AND2_X1 U6340 ( .A1(n5729), .A2(n4993), .ZN(n5959) );
  AND2_X1 U6341 ( .A1(n5728), .A2(n5841), .ZN(n4993) );
  NAND2_X1 U6342 ( .A1(n8673), .A2(n4996), .ZN(n4995) );
  OR2_X1 U6343 ( .A1(n5455), .A2(n5165), .ZN(n5166) );
  NAND2_X1 U6344 ( .A1(n6576), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U6345 ( .A1(n6293), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5785) );
  INV_X1 U6346 ( .A(n9867), .ZN(n5060) );
  XNOR2_X1 U6347 ( .A(n7831), .B(n7867), .ZN(n8279) );
  INV_X1 U6348 ( .A(n5635), .ZN(n7839) );
  AOI21_X1 U6349 ( .B1(n7726), .B2(n6654), .A(n6186), .ZN(n6594) );
  NAND2_X1 U6350 ( .A1(n6652), .A2(n9863), .ZN(n9876) );
  INV_X1 U6351 ( .A(n9963), .ZN(n5726) );
  INV_X1 U6352 ( .A(n8471), .ZN(n5724) );
  INV_X2 U6353 ( .A(n9676), .ZN(n9678) );
  NAND2_X1 U6354 ( .A1(n6360), .A2(n6359), .ZN(n6422) );
  NAND2_X1 U6355 ( .A1(n6762), .A2(n7889), .ZN(n6734) );
  INV_X1 U6356 ( .A(n9186), .ZN(n9200) );
  INV_X1 U6357 ( .A(n9476), .ZN(n10046) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6073) );
  OR2_X1 U6359 ( .A1(n8281), .A2(n8530), .ZN(n4998) );
  AND2_X1 U6360 ( .A1(n6462), .A2(n6461), .ZN(n4999) );
  OR2_X1 U6361 ( .A1(n7705), .A2(n9387), .ZN(n5000) );
  OR2_X1 U6362 ( .A1(n6469), .A2(n9073), .ZN(n5001) );
  AND2_X1 U6363 ( .A1(n6780), .A2(n6779), .ZN(n5002) );
  OR2_X1 U6364 ( .A1(n6573), .A2(n9072), .ZN(n5003) );
  AND2_X1 U6365 ( .A1(n9301), .A2(n8591), .ZN(n5005) );
  AND2_X1 U6366 ( .A1(n8615), .A2(n8614), .ZN(n5006) );
  INV_X4 U6367 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U6368 ( .A(n9074), .ZN(n5802) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8036) );
  INV_X2 U6370 ( .A(n9674), .ZN(n9464) );
  INV_X1 U6371 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5025) );
  INV_X1 U6372 ( .A(n8518), .ZN(n5459) );
  NAND2_X1 U6373 ( .A1(n7809), .A2(n7754), .ZN(n5008) );
  AND2_X1 U6374 ( .A1(n6996), .A2(n6998), .ZN(n5009) );
  INV_X1 U6375 ( .A(n7352), .ZN(n5894) );
  AND2_X1 U6376 ( .A1(n8279), .A2(n9926), .ZN(n5010) );
  OR2_X1 U6377 ( .A1(n9428), .A2(n8801), .ZN(n5011) );
  AND2_X1 U6378 ( .A1(n8523), .A2(n8372), .ZN(n5012) );
  INV_X1 U6379 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5014) );
  INV_X1 U6380 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5017) );
  INV_X1 U6381 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5738) );
  OR2_X1 U6382 ( .A1(n8196), .A2(n6758), .ZN(n5142) );
  INV_X1 U6383 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5418) );
  INV_X1 U6384 ( .A(n7796), .ZN(n5471) );
  NAND2_X1 U6385 ( .A1(n6737), .A2(n5103), .ZN(n5123) );
  INV_X1 U6386 ( .A(n9188), .ZN(n6139) );
  INV_X1 U6387 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5744) );
  INV_X1 U6388 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10015) );
  INV_X1 U6389 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U6390 ( .A1(n8513), .A2(n5471), .ZN(n5472) );
  INV_X1 U6391 ( .A(n5347), .ZN(n5346) );
  NAND2_X1 U6392 ( .A1(n5459), .A2(n8383), .ZN(n5460) );
  NAND2_X1 U6393 ( .A1(n7570), .A2(n8431), .ZN(n5338) );
  NAND2_X1 U6394 ( .A1(n5080), .A2(n7671), .ZN(n5089) );
  INV_X1 U6395 ( .A(SI_22_), .ZN(n10199) );
  INV_X1 U6396 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5859) );
  INV_X1 U6397 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5872) );
  INV_X1 U6398 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5989) );
  NOR2_X1 U6399 ( .A1(n5914), .A2(n5771), .ZN(n5924) );
  OR2_X1 U6400 ( .A1(n7382), .A2(n9063), .ZN(n5931) );
  INV_X1 U6401 ( .A(SI_25_), .ZN(n10194) );
  INV_X1 U6402 ( .A(SI_20_), .ZN(n5441) );
  INV_X1 U6403 ( .A(SI_16_), .ZN(n10108) );
  INV_X1 U6404 ( .A(SI_11_), .ZN(n5260) );
  NOR2_X1 U6405 ( .A1(n8294), .A2(n8396), .ZN(n8295) );
  NAND2_X1 U6406 ( .A1(n5385), .A2(n5384), .ZN(n5405) );
  INV_X1 U6407 ( .A(n7327), .ZN(n7330) );
  OR2_X1 U6408 ( .A1(n8007), .A2(n6183), .ZN(n6655) );
  OR2_X1 U6409 ( .A1(n5873), .A2(n5872), .ZN(n5887) );
  NAND2_X1 U6410 ( .A1(n6786), .A2(n6788), .ZN(n6789) );
  NOR2_X1 U6411 ( .A1(n10093), .A2(n6053), .ZN(n6066) );
  NOR2_X1 U6412 ( .A1(n5939), .A2(n10272), .ZN(n5963) );
  INV_X1 U6413 ( .A(n9474), .ZN(n5756) );
  OR2_X1 U6414 ( .A1(n5990), .A2(n5989), .ZN(n6007) );
  OR2_X1 U6415 ( .A1(n5937), .A2(n5936), .ZN(n5939) );
  OR2_X1 U6416 ( .A1(n5912), .A2(n10169), .ZN(n5914) );
  OR2_X1 U6417 ( .A1(n6918), .A2(n9070), .ZN(n5858) );
  OR2_X1 U6418 ( .A1(n7373), .A2(n9066), .ZN(n5907) );
  NAND2_X1 U6419 ( .A1(n8820), .A2(n5802), .ZN(n5803) );
  AND2_X1 U6420 ( .A1(n5590), .A2(n5575), .ZN(n5576) );
  INV_X1 U6421 ( .A(SI_12_), .ZN(n5282) );
  AND2_X1 U6422 ( .A1(n7805), .A2(n7749), .ZN(n8093) );
  NAND2_X1 U6423 ( .A1(n5518), .A2(n5517), .ZN(n5537) );
  AND2_X1 U6424 ( .A1(n7803), .A2(n7746), .ZN(n8136) );
  XNOR2_X1 U6425 ( .A(n4432), .B(n9879), .ZN(n6187) );
  INV_X1 U6426 ( .A(n8320), .ZN(n8294) );
  INV_X1 U6427 ( .A(n5084), .ZN(n5454) );
  NAND2_X1 U6428 ( .A1(n5663), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5064) );
  NAND2_X2 U6429 ( .A1(n5660), .A2(n5661), .ZN(n5080) );
  INV_X1 U6430 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10147) );
  AND2_X1 U6431 ( .A1(n6272), .A2(n8559), .ZN(n6279) );
  XNOR2_X1 U6432 ( .A(n8292), .B(n8291), .ZN(n8298) );
  INV_X1 U6433 ( .A(n7861), .ZN(n7984) );
  INV_X1 U6434 ( .A(n7930), .ZN(n5640) );
  OR2_X1 U6435 ( .A1(n6645), .A2(n5687), .ZN(n5721) );
  INV_X1 U6436 ( .A(n8192), .ZN(n7449) );
  INV_X1 U6437 ( .A(n9866), .ZN(n8396) );
  INV_X1 U6438 ( .A(n8394), .ZN(n9869) );
  AND2_X1 U6439 ( .A1(n5705), .A2(n5630), .ZN(n9873) );
  NOR2_X1 U6440 ( .A1(n6463), .A2(n4999), .ZN(n6572) );
  INV_X1 U6441 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7698) );
  OR3_X1 U6442 ( .A1(n6577), .A2(n6576), .A3(n6575), .ZN(n6578) );
  NAND2_X1 U6443 ( .A1(n6773), .A2(n7324), .ZN(n6354) );
  NOR2_X1 U6444 ( .A1(n7067), .A2(n9665), .ZN(n6413) );
  AND3_X1 U6445 ( .A1(n6296), .A2(n6295), .A3(n6294), .ZN(n8896) );
  NOR2_X1 U6446 ( .A1(n6033), .A2(n10052), .ZN(n6042) );
  INV_X1 U6447 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10200) );
  INV_X1 U6448 ( .A(n8054), .ZN(n6371) );
  NAND2_X1 U6449 ( .A1(n6371), .A2(n8900), .ZN(n8800) );
  OR2_X1 U6450 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  INV_X1 U6451 ( .A(n8798), .ZN(n8784) );
  NOR2_X1 U6452 ( .A1(n9459), .A2(n9058), .ZN(n5996) );
  INV_X1 U6453 ( .A(n9061), .ZN(n7491) );
  INV_X1 U6454 ( .A(n9626), .ZN(n6835) );
  AND2_X1 U6455 ( .A1(n9667), .A2(n6407), .ZN(n7065) );
  INV_X1 U6456 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6000) );
  INV_X1 U6457 ( .A(n8170), .ZN(n8141) );
  INV_X1 U6458 ( .A(n8143), .ZN(n8172) );
  INV_X1 U6459 ( .A(n9884), .ZN(n6608) );
  INV_X1 U6460 ( .A(n8174), .ZN(n8164) );
  INV_X1 U6461 ( .A(n7500), .ZN(n8030) );
  AND3_X1 U6462 ( .A1(n5470), .A2(n5469), .A3(n5468), .ZN(n7796) );
  NAND2_X1 U6463 ( .A1(n5702), .A2(n5701), .ZN(n6270) );
  INV_X1 U6464 ( .A(n9692), .ZN(n9851) );
  INV_X1 U6465 ( .A(n9713), .ZN(n9842) );
  INV_X1 U6466 ( .A(n9876), .ZN(n6677) );
  AND2_X1 U6467 ( .A1(n5650), .A2(n7989), .ZN(n8329) );
  AND2_X1 U6468 ( .A1(n7944), .A2(n7943), .ZN(n7851) );
  INV_X1 U6469 ( .A(n9873), .ZN(n8433) );
  NOR2_X1 U6470 ( .A1(n9963), .A2(n10209), .ZN(n5723) );
  AND2_X1 U6471 ( .A1(n5721), .A2(n5720), .ZN(n6651) );
  AND2_X1 U6472 ( .A1(n7958), .A2(n8397), .ZN(n8409) );
  INV_X1 U6473 ( .A(n9919), .ZN(n9943) );
  OR2_X1 U6474 ( .A1(n9927), .A2(n9926), .ZN(n9938) );
  AND2_X1 U6475 ( .A1(n7500), .A2(n6678), .ZN(n9926) );
  XNOR2_X1 U6476 ( .A(n5704), .B(n5703), .ZN(n6201) );
  NAND2_X1 U6477 ( .A1(n6412), .A2(n9621), .ZN(n8790) );
  AND4_X1 U6478 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n8684)
         );
  AND2_X1 U6479 ( .A1(n6060), .A2(n6059), .ZN(n8801) );
  AND4_X1 U6480 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n8570)
         );
  AND2_X1 U6481 ( .A1(n6409), .A2(n8885), .ZN(n9342) );
  NAND2_X1 U6482 ( .A1(n6132), .A2(n6131), .ZN(n9329) );
  INV_X1 U6483 ( .A(n9328), .ZN(n9338) );
  NAND2_X1 U6484 ( .A1(n9676), .A2(n6090), .ZN(n6172) );
  INV_X1 U6485 ( .A(n9387), .ZN(n9405) );
  INV_X1 U6486 ( .A(n9368), .ZN(n9673) );
  INV_X1 U6487 ( .A(n6171), .ZN(n9636) );
  OAI22_X1 U6488 ( .A1(n6171), .A2(P1_D_REG_0__SCAN_IN), .B1(n6156), .B2(n6170), .ZN(n7064) );
  OR2_X1 U6489 ( .A1(n5778), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5919) );
  AND2_X1 U6490 ( .A1(n7671), .A2(P1_U3086), .ZN(n10045) );
  AND2_X1 U6491 ( .A1(n6208), .A2(n6207), .ZN(n8174) );
  INV_X1 U6492 ( .A(n8160), .ZN(n8177) );
  INV_X1 U6493 ( .A(n8306), .ZN(n8186) );
  INV_X1 U6494 ( .A(n7462), .ZN(n8431) );
  OR2_X1 U6495 ( .A1(P2_U3150), .A2(n6271), .ZN(n9713) );
  OR2_X1 U6496 ( .A1(n6334), .A2(n8257), .ZN(n9856) );
  NAND2_X1 U6497 ( .A1(n8413), .A2(n6733), .ZN(n8441) );
  INV_X1 U6498 ( .A(n8485), .ZN(n8446) );
  NAND2_X1 U6499 ( .A1(n9963), .A2(n9943), .ZN(n8471) );
  NAND2_X1 U6500 ( .A1(n9963), .A2(n9938), .ZN(n8479) );
  AND2_X2 U6501 ( .A1(n5722), .A2(n6651), .ZN(n9963) );
  OR2_X1 U6502 ( .A1(n9944), .A2(n9919), .ZN(n8530) );
  OR2_X1 U6503 ( .A1(n9944), .A2(n9932), .ZN(n8550) );
  AND3_X1 U6504 ( .A1(n9931), .A2(n9930), .A3(n9929), .ZN(n9960) );
  AND2_X1 U6505 ( .A1(n5711), .A2(n5710), .ZN(n9944) );
  INV_X1 U6506 ( .A(n6265), .ZN(n6266) );
  NAND2_X1 U6507 ( .A1(n6244), .A2(n6243), .ZN(n6265) );
  INV_X1 U6508 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10258) );
  INV_X1 U6509 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6302) );
  INV_X1 U6510 ( .A(n9379), .ZN(n9259) );
  INV_X1 U6511 ( .A(n8575), .ZN(n8739) );
  INV_X1 U6512 ( .A(n8790), .ZN(n8807) );
  AND4_X1 U6513 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n7706)
         );
  OAI21_X1 U6514 ( .B1(n9255), .B2(n5940), .A(n6038), .ZN(n9054) );
  INV_X1 U6515 ( .A(n6966), .ZN(n9068) );
  INV_X1 U6516 ( .A(n9518), .ZN(n9620) );
  AND2_X1 U6517 ( .A1(n9334), .A2(n9333), .ZN(n9403) );
  NAND2_X1 U6518 ( .A1(n9624), .A2(n7070), .ZN(n9328) );
  NAND2_X1 U6519 ( .A1(n9678), .A2(n9411), .ZN(n9387) );
  NAND2_X1 U6520 ( .A1(n9678), .A2(n9673), .ZN(n9407) );
  OR2_X1 U6521 ( .A1(n6176), .A2(n7064), .ZN(n9676) );
  NAND2_X1 U6522 ( .A1(n9464), .A2(n9411), .ZN(n9442) );
  NAND2_X1 U6523 ( .A1(n9464), .A2(n9673), .ZN(n9462) );
  OR2_X1 U6524 ( .A1(n6176), .A2(n6175), .ZN(n9674) );
  CLKBUF_X1 U6525 ( .A(n9664), .Z(n9655) );
  INV_X1 U6526 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10213) );
  NAND2_X1 U6527 ( .A1(n6148), .A2(n6147), .ZN(n7616) );
  INV_X1 U6528 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7177) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6304) );
  INV_X2 U6530 ( .A(n8225), .ZN(P2_U3893) );
  OAI21_X1 U6531 ( .B1(n5727), .B2(n5726), .A(n5725), .ZN(P2_U3488) );
  INV_X1 U6532 ( .A(n6670), .ZN(P1_U3973) );
  NAND4_X1 U6533 ( .A1(n5196), .A2(n5015), .A3(n5014), .A4(n5195), .ZN(n5016)
         );
  NOR2_X1 U6534 ( .A1(n5097), .A2(n5016), .ZN(n5023) );
  NAND2_X1 U6535 ( .A1(n5327), .A2(n5017), .ZN(n5362) );
  INV_X1 U6536 ( .A(n5362), .ZN(n5020) );
  NOR2_X1 U6537 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5019) );
  NOR2_X1 U6538 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5018) );
  NAND3_X1 U6539 ( .A1(n5020), .A2(n5019), .A3(n5018), .ZN(n5022) );
  INV_X1 U6540 ( .A(n5671), .ZN(n5026) );
  XNOR2_X2 U6541 ( .A(n5027), .B(n8554), .ZN(n7665) );
  NAND2_X2 U6542 ( .A1(n5032), .A2(n7652), .ZN(n5084) );
  INV_X1 U6543 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5031) );
  OR2_X1 U6544 ( .A1(n5084), .A2(n5031), .ZN(n5034) );
  INV_X1 U6545 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10212) );
  INV_X1 U6546 ( .A(n7652), .ZN(n5035) );
  NAND2_X4 U6547 ( .A1(n5035), .A2(n7665), .ZN(n6926) );
  INV_X1 U6548 ( .A(n6926), .ZN(n5036) );
  NAND2_X1 U6549 ( .A1(n5036), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5038) );
  AND2_X4 U6550 ( .A1(n7665), .A2(n7652), .ZN(n6925) );
  NAND2_X1 U6551 ( .A1(n6925), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6552 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5051) );
  AND2_X1 U6553 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6554 ( .A1(n7676), .A2(n5050), .ZN(n5800) );
  XNOR2_X1 U6555 ( .A(n5073), .B(n5072), .ZN(n5790) );
  OR2_X1 U6556 ( .A1(n5089), .A2(n5790), .ZN(n5056) );
  NAND2_X1 U6557 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5052) );
  MUX2_X1 U6558 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5052), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5055) );
  INV_X1 U6559 ( .A(n5053), .ZN(n5054) );
  INV_X1 U6560 ( .A(n6291), .ZN(n6329) );
  AND2_X1 U6561 ( .A1(n5056), .A2(n4463), .ZN(n5058) );
  NAND2_X4 U6562 ( .A1(n5080), .A2(n7676), .ZN(n7825) );
  OR2_X1 U6563 ( .A1(n7825), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5057) );
  NAND2_X2 U6564 ( .A1(n5058), .A2(n5057), .ZN(n9879) );
  NAND2_X1 U6565 ( .A1(n9867), .A2(n9879), .ZN(n7881) );
  NAND2_X2 U6566 ( .A1(n5634), .A2(n7881), .ZN(n6673) );
  INV_X1 U6567 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6653) );
  OR2_X1 U6568 ( .A1(n5146), .A2(n6653), .ZN(n5063) );
  OR2_X1 U6569 ( .A1(n5084), .A2(n10253), .ZN(n5062) );
  NAND2_X1 U6570 ( .A1(n6925), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6571 ( .A1(n7671), .A2(SI_0_), .ZN(n5065) );
  XNOR2_X1 U6572 ( .A(n5065), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8564) );
  MUX2_X1 U6573 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8564), .S(n5080), .Z(n5633) );
  NAND2_X1 U6574 ( .A1(n5632), .A2(n5633), .ZN(n6672) );
  NAND2_X1 U6575 ( .A1(n6673), .A2(n6672), .ZN(n5067) );
  OR2_X1 U6576 ( .A1(n9867), .A2(n5059), .ZN(n5066) );
  NAND2_X1 U6577 ( .A1(n5067), .A2(n5066), .ZN(n9865) );
  NAND2_X1 U6578 ( .A1(n6925), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5071) );
  INV_X1 U6579 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9878) );
  INV_X1 U6580 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6310) );
  OR2_X1 U6581 ( .A1(n6926), .A2(n6310), .ZN(n5069) );
  INV_X1 U6582 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6321) );
  OR2_X1 U6583 ( .A1(n5146), .A2(n6321), .ZN(n5068) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6225) );
  OR2_X1 U6585 ( .A1(n7825), .A2(n6225), .ZN(n5083) );
  INV_X1 U6586 ( .A(n5072), .ZN(n5074) );
  NAND2_X1 U6587 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  NAND2_X1 U6588 ( .A1(n5075), .A2(SI_1_), .ZN(n5076) );
  NAND2_X1 U6589 ( .A1(n5077), .A2(n5076), .ZN(n5091) );
  INV_X1 U6590 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6235) );
  MUX2_X1 U6591 ( .A(n6235), .B(n6225), .S(n5078), .Z(n5092) );
  XNOR2_X1 U6592 ( .A(n5092), .B(SI_2_), .ZN(n5090) );
  XNOR2_X1 U6593 ( .A(n5091), .B(n5090), .ZN(n6234) );
  OR2_X1 U6594 ( .A1(n5089), .A2(n6234), .ZN(n5082) );
  OR2_X1 U6595 ( .A1(n5080), .A2(n6543), .ZN(n5081) );
  XNOR2_X1 U6597 ( .A(n8198), .B(n9884), .ZN(n5635) );
  NAND2_X1 U6598 ( .A1(n9865), .A2(n5635), .ZN(n6736) );
  OR2_X1 U6599 ( .A1(n8198), .A2(n6608), .ZN(n6735) );
  NAND2_X1 U6600 ( .A1(n6925), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5088) );
  INV_X1 U6601 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6767) );
  OR2_X1 U6602 ( .A1(n5084), .A2(n6767), .ZN(n5087) );
  OR2_X1 U6603 ( .A1(n6926), .A2(n9950), .ZN(n5086) );
  OR2_X1 U6604 ( .A1(n5146), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6605 ( .A1(n7825), .A2(n6226), .ZN(n5101) );
  NAND2_X1 U6606 ( .A1(n5091), .A2(n5090), .ZN(n5095) );
  INV_X1 U6607 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6608 ( .A1(n5093), .A2(SI_2_), .ZN(n5094) );
  NAND2_X1 U6609 ( .A1(n5095), .A2(n5094), .ZN(n5113) );
  MUX2_X1 U6610 ( .A(n6226), .B(n6231), .S(n7676), .Z(n5114) );
  XNOR2_X1 U6611 ( .A(n5114), .B(SI_3_), .ZN(n5112) );
  XNOR2_X1 U6612 ( .A(n5113), .B(n5112), .ZN(n6230) );
  OR2_X1 U6613 ( .A1(n5156), .A2(n6230), .ZN(n5100) );
  NAND2_X1 U6614 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5096) );
  MUX2_X1 U6615 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5096), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5098) );
  NAND2_X1 U6616 ( .A1(n5098), .A2(n5133), .ZN(n6546) );
  OR2_X1 U6617 ( .A1(n5080), .A2(n6546), .ZN(n5099) );
  INV_X1 U6618 ( .A(n6561), .ZN(n9889) );
  OR2_X1 U6619 ( .A1(n9868), .A2(n9889), .ZN(n6737) );
  AND2_X1 U6620 ( .A1(n6735), .A2(n6737), .ZN(n5102) );
  NAND2_X1 U6621 ( .A1(n6736), .A2(n5102), .ZN(n5124) );
  OR2_X2 U6622 ( .A1(n9868), .A2(n6561), .ZN(n7889) );
  NAND2_X1 U6623 ( .A1(n9868), .A2(n6561), .ZN(n7904) );
  NAND2_X1 U6624 ( .A1(n7889), .A2(n7904), .ZN(n6764) );
  INV_X1 U6625 ( .A(n6764), .ZN(n5103) );
  NAND2_X1 U6626 ( .A1(n5454), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5111) );
  INV_X1 U6627 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6542) );
  OR2_X1 U6628 ( .A1(n6926), .A2(n6542), .ZN(n5110) );
  INV_X1 U6629 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5105) );
  INV_X1 U6630 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6631 ( .A1(n5105), .A2(n5104), .ZN(n5127) );
  NAND2_X1 U6632 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5106) );
  AND2_X1 U6633 ( .A1(n5127), .A2(n5106), .ZN(n6629) );
  OR2_X1 U6634 ( .A1(n5404), .A2(n6629), .ZN(n5109) );
  INV_X1 U6635 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5107) );
  OR2_X1 U6636 ( .A1(n5455), .A2(n5107), .ZN(n5108) );
  NAND2_X1 U6637 ( .A1(n5113), .A2(n5112), .ZN(n5117) );
  INV_X1 U6638 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6639 ( .A1(n5115), .A2(SI_3_), .ZN(n5116) );
  NAND2_X1 U6640 ( .A1(n5117), .A2(n5116), .ZN(n5135) );
  MUX2_X1 U6641 ( .A(n6227), .B(n6233), .S(n6228), .Z(n5136) );
  XNOR2_X1 U6642 ( .A(n5136), .B(SI_4_), .ZN(n5134) );
  XNOR2_X1 U6643 ( .A(n5135), .B(n5134), .ZN(n6232) );
  OR2_X1 U6644 ( .A1(n5156), .A2(n6232), .ZN(n5122) );
  OR2_X1 U6645 ( .A1(n7825), .A2(n6227), .ZN(n5121) );
  NAND2_X1 U6646 ( .A1(n5133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5119) );
  INV_X1 U6647 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5118) );
  XNOR2_X1 U6648 ( .A(n5119), .B(n5118), .ZN(n6707) );
  OR2_X1 U6649 ( .A1(n5080), .A2(n6707), .ZN(n5120) );
  NAND2_X1 U6650 ( .A1(n8197), .A2(n9896), .ZN(n7890) );
  NAND3_X1 U6651 ( .A1(n5124), .A2(n5123), .A3(n7838), .ZN(n6750) );
  INV_X1 U6652 ( .A(n9896), .ZN(n6743) );
  OR2_X1 U6653 ( .A1(n8197), .A2(n6743), .ZN(n6749) );
  NAND2_X1 U6654 ( .A1(n6925), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5132) );
  INV_X1 U6655 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6685) );
  OR2_X1 U6656 ( .A1(n6926), .A2(n6685), .ZN(n5131) );
  INV_X1 U6657 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6686) );
  OR2_X1 U6658 ( .A1(n6929), .A2(n6686), .ZN(n5130) );
  INV_X1 U6659 ( .A(n5127), .ZN(n5126) );
  INV_X1 U6660 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6661 ( .A1(n5126), .A2(n5125), .ZN(n5144) );
  NAND2_X1 U6662 ( .A1(n5127), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5128) );
  AND2_X1 U6663 ( .A1(n5144), .A2(n5128), .ZN(n6756) );
  OR2_X1 U6664 ( .A1(n5404), .A2(n6756), .ZN(n5129) );
  NOR2_X1 U6665 ( .A1(n5133), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6666 ( .A1(n5198), .A2(n5079), .ZN(n5157) );
  XNOR2_X1 U6667 ( .A(n5157), .B(n5195), .ZN(n9707) );
  NAND2_X1 U6668 ( .A1(n5135), .A2(n5134), .ZN(n5139) );
  INV_X1 U6669 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6670 ( .A1(n5137), .A2(SI_4_), .ZN(n5138) );
  MUX2_X1 U6671 ( .A(n6238), .B(n6236), .S(n7676), .Z(n5152) );
  XNOR2_X2 U6672 ( .A(n5154), .B(n5152), .ZN(n5151) );
  XNOR2_X1 U6673 ( .A(n5151), .B(SI_5_), .ZN(n6237) );
  OR2_X1 U6674 ( .A1(n6237), .A2(n5156), .ZN(n5141) );
  OR2_X1 U6675 ( .A1(n7825), .A2(n6238), .ZN(n5140) );
  OAI211_X1 U6676 ( .C1(n5080), .C2(n9707), .A(n5141), .B(n5140), .ZN(n6758)
         );
  AND2_X1 U6677 ( .A1(n6749), .A2(n5142), .ZN(n5143) );
  NAND2_X1 U6678 ( .A1(n8196), .A2(n6758), .ZN(n6871) );
  INV_X1 U6679 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6684) );
  OR2_X1 U6680 ( .A1(n6926), .A2(n6684), .ZN(n5149) );
  NAND2_X1 U6681 ( .A1(n5144), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5145) );
  AND2_X1 U6682 ( .A1(n5163), .A2(n5145), .ZN(n6940) );
  OR2_X1 U6683 ( .A1(n5404), .A2(n6940), .ZN(n5148) );
  NAND2_X1 U6684 ( .A1(n6925), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5147) );
  INV_X1 U6685 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6686 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6228), .Z(n5172) );
  XNOR2_X1 U6688 ( .A(n5172), .B(SI_6_), .ZN(n5170) );
  XNOR2_X1 U6689 ( .A(n5171), .B(n5170), .ZN(n6239) );
  NAND2_X1 U6690 ( .A1(n6239), .A2(n7822), .ZN(n5160) );
  INV_X2 U6691 ( .A(n7825), .ZN(n5428) );
  NAND2_X1 U6692 ( .A1(n5157), .A2(n5195), .ZN(n5158) );
  NAND2_X1 U6693 ( .A1(n5158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5175) );
  XNOR2_X1 U6694 ( .A(n5175), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7432) );
  AOI22_X1 U6695 ( .A1(n5428), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5427), .B2(
        n7432), .ZN(n5159) );
  INV_X1 U6696 ( .A(n9906), .ZN(n6948) );
  NAND2_X1 U6697 ( .A1(n8195), .A2(n6948), .ZN(n5181) );
  AND2_X1 U6698 ( .A1(n6871), .A2(n5181), .ZN(n6812) );
  NAND2_X1 U6699 ( .A1(n5663), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5169) );
  INV_X1 U6700 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6818) );
  OR2_X1 U6701 ( .A1(n5084), .A2(n6818), .ZN(n5168) );
  INV_X1 U6702 ( .A(n5163), .ZN(n5162) );
  INV_X1 U6703 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6704 ( .A1(n5162), .A2(n5161), .ZN(n5203) );
  NAND2_X1 U6705 ( .A1(n5163), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5164) );
  AND2_X1 U6706 ( .A1(n5203), .A2(n5164), .ZN(n6819) );
  OR2_X1 U6707 ( .A1(n5404), .A2(n6819), .ZN(n5167) );
  INV_X1 U6708 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6709 ( .A1(n5172), .A2(SI_6_), .ZN(n5173) );
  MUX2_X1 U6710 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6228), .Z(n5188) );
  XNOR2_X1 U6711 ( .A(n5188), .B(SI_7_), .ZN(n5185) );
  XNOR2_X1 U6712 ( .A(n5187), .B(n5185), .ZN(n6251) );
  NAND2_X1 U6713 ( .A1(n6251), .A2(n7822), .ZN(n5179) );
  INV_X1 U6714 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6715 ( .A1(n5175), .A2(n5174), .ZN(n5176) );
  NAND2_X1 U6716 ( .A1(n5176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5177) );
  XNOR2_X1 U6717 ( .A(n5177), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U6718 ( .A1(n5428), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5427), .B2(
        n9715), .ZN(n5178) );
  NAND2_X1 U6719 ( .A1(n6937), .A2(n6952), .ZN(n7894) );
  AND2_X2 U6720 ( .A1(n6839), .A2(n7894), .ZN(n7916) );
  INV_X1 U6721 ( .A(n7916), .ZN(n5180) );
  OR2_X1 U6722 ( .A1(n6952), .A2(n8194), .ZN(n5184) );
  INV_X1 U6723 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6724 ( .A1(n5188), .A2(SI_7_), .ZN(n5189) );
  INV_X1 U6725 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5190) );
  MUX2_X1 U6726 ( .A(n10244), .B(n5190), .S(n6228), .Z(n5192) );
  INV_X1 U6727 ( .A(SI_8_), .ZN(n5191) );
  NAND2_X1 U6728 ( .A1(n5192), .A2(n5191), .ZN(n5214) );
  INV_X1 U6729 ( .A(n5192), .ZN(n5193) );
  NAND2_X1 U6730 ( .A1(n5193), .A2(SI_8_), .ZN(n5194) );
  NAND2_X1 U6731 ( .A1(n6255), .A2(n7822), .ZN(n5201) );
  AND2_X1 U6732 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  OR2_X1 U6733 ( .A1(n5397), .A2(n5079), .ZN(n5199) );
  XNOR2_X1 U6734 ( .A(n5199), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U6735 ( .A1(n5428), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5427), .B2(
        n9729), .ZN(n5200) );
  NAND2_X1 U6736 ( .A1(n6925), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5208) );
  INV_X1 U6737 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6738 ( .A1(n6926), .A2(n5202), .ZN(n5207) );
  INV_X1 U6739 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7412) );
  OR2_X1 U6740 ( .A1(n5084), .A2(n7412), .ZN(n5206) );
  NAND2_X1 U6741 ( .A1(n5203), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5204) );
  AND2_X1 U6742 ( .A1(n5231), .A2(n5204), .ZN(n7009) );
  OR2_X1 U6743 ( .A1(n5404), .A2(n7009), .ZN(n5205) );
  NAND2_X1 U6744 ( .A1(n9917), .A2(n8193), .ZN(n5209) );
  NAND2_X1 U6745 ( .A1(n6842), .A2(n5209), .ZN(n5211) );
  OR2_X1 U6746 ( .A1(n9917), .A2(n8193), .ZN(n5210) );
  NAND2_X1 U6747 ( .A1(n5211), .A2(n5210), .ZN(n7020) );
  MUX2_X1 U6748 ( .A(n6302), .B(n6304), .S(n6228), .Z(n5216) );
  INV_X1 U6749 ( .A(SI_9_), .ZN(n5215) );
  NAND2_X1 U6750 ( .A1(n5216), .A2(n5215), .ZN(n5239) );
  INV_X1 U6751 ( .A(n5216), .ZN(n5217) );
  NAND2_X1 U6752 ( .A1(n5217), .A2(SI_9_), .ZN(n5218) );
  NAND2_X1 U6753 ( .A1(n5240), .A2(n5220), .ZN(n6301) );
  NAND2_X1 U6754 ( .A1(n6301), .A2(n7822), .ZN(n5226) );
  NAND2_X1 U6755 ( .A1(n5397), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6756 ( .A1(n5223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5222) );
  MUX2_X1 U6757 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5222), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5224) );
  AOI22_X1 U6758 ( .A1(n5428), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5427), .B2(
        n9746), .ZN(n5225) );
  NAND2_X1 U6759 ( .A1(n6925), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5236) );
  INV_X1 U6760 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5227) );
  OR2_X1 U6761 ( .A1(n5084), .A2(n5227), .ZN(n5235) );
  INV_X1 U6762 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5228) );
  OR2_X1 U6763 ( .A1(n6926), .A2(n5228), .ZN(n5234) );
  INV_X1 U6764 ( .A(n5231), .ZN(n5230) );
  NAND2_X1 U6765 ( .A1(n5230), .A2(n5229), .ZN(n5245) );
  NAND2_X1 U6766 ( .A1(n5231), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5232) );
  AND2_X1 U6767 ( .A1(n5245), .A2(n5232), .ZN(n7054) );
  OR2_X1 U6768 ( .A1(n5404), .A2(n7054), .ZN(n5233) );
  NAND2_X1 U6769 ( .A1(n7050), .A2(n7305), .ZN(n7901) );
  NAND2_X1 U6770 ( .A1(n7922), .A2(n7901), .ZN(n7021) );
  NAND2_X1 U6771 ( .A1(n7020), .A2(n7021), .ZN(n5238) );
  INV_X1 U6772 ( .A(n7305), .ZN(n7051) );
  OR2_X1 U6773 ( .A1(n7050), .A2(n7051), .ZN(n5237) );
  NAND2_X1 U6774 ( .A1(n5238), .A2(n5237), .ZN(n6880) );
  INV_X1 U6775 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5241) );
  MUX2_X1 U6776 ( .A(n6307), .B(n5241), .S(n7676), .Z(n5255) );
  XNOR2_X1 U6777 ( .A(n5255), .B(SI_10_), .ZN(n5254) );
  XNOR2_X1 U6778 ( .A(n5258), .B(n5254), .ZN(n6305) );
  NAND2_X1 U6779 ( .A1(n6305), .A2(n7822), .ZN(n5244) );
  NAND2_X1 U6780 ( .A1(n5267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5242) );
  XNOR2_X1 U6781 ( .A(n5242), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7438) );
  AOI22_X1 U6782 ( .A1(n5428), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5427), .B2(
        n7438), .ZN(n5243) );
  NAND2_X1 U6783 ( .A1(n5244), .A2(n5243), .ZN(n9925) );
  NAND2_X1 U6784 ( .A1(n5663), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5251) );
  INV_X1 U6785 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7415) );
  OR2_X1 U6786 ( .A1(n5084), .A2(n7415), .ZN(n5250) );
  NAND2_X1 U6787 ( .A1(n5245), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5246) );
  AND2_X1 U6788 ( .A1(n5271), .A2(n5246), .ZN(n7308) );
  OR2_X1 U6789 ( .A1(n5404), .A2(n7308), .ZN(n5249) );
  INV_X1 U6790 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5247) );
  OR2_X1 U6791 ( .A1(n5455), .A2(n5247), .ZN(n5248) );
  NAND4_X1 U6792 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n8192)
         );
  NOR2_X1 U6793 ( .A1(n9925), .A2(n8192), .ZN(n5253) );
  NAND2_X1 U6794 ( .A1(n9925), .A2(n8192), .ZN(n5252) );
  INV_X1 U6795 ( .A(n5254), .ZN(n5257) );
  INV_X1 U6796 ( .A(n5255), .ZN(n5256) );
  INV_X1 U6797 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5259) );
  MUX2_X1 U6798 ( .A(n6345), .B(n5259), .S(n6228), .Z(n5261) );
  NAND2_X1 U6799 ( .A1(n5261), .A2(n5260), .ZN(n5280) );
  INV_X1 U6800 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6801 ( .A1(n5262), .A2(SI_11_), .ZN(n5263) );
  NAND2_X1 U6802 ( .A1(n5280), .A2(n5263), .ZN(n5264) );
  NAND2_X1 U6803 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6804 ( .A1(n5281), .A2(n5266), .ZN(n6342) );
  NAND2_X1 U6805 ( .A1(n6342), .A2(n7822), .ZN(n5270) );
  NAND2_X1 U6806 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6807 ( .A(n5268), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9761) );
  AOI22_X1 U6808 ( .A1(n5428), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5427), .B2(
        n9761), .ZN(n5269) );
  NAND2_X1 U6809 ( .A1(n5270), .A2(n5269), .ZN(n9936) );
  NAND2_X1 U6810 ( .A1(n6925), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5277) );
  INV_X1 U6811 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7043) );
  OR2_X1 U6812 ( .A1(n5084), .A2(n7043), .ZN(n5276) );
  NAND2_X1 U6813 ( .A1(n5271), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5272) );
  AND2_X1 U6814 ( .A1(n5289), .A2(n5272), .ZN(n7402) );
  OR2_X1 U6815 ( .A1(n5404), .A2(n7402), .ZN(n5275) );
  INV_X1 U6816 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5273) );
  OR2_X1 U6817 ( .A1(n6926), .A2(n5273), .ZN(n5274) );
  XNOR2_X1 U6818 ( .A(n9936), .B(n7476), .ZN(n7929) );
  NAND2_X1 U6819 ( .A1(n7041), .A2(n7929), .ZN(n5279) );
  INV_X1 U6820 ( .A(n7476), .ZN(n8191) );
  NAND2_X1 U6821 ( .A1(n9936), .A2(n8191), .ZN(n5278) );
  NAND2_X1 U6822 ( .A1(n5279), .A2(n5278), .ZN(n7080) );
  MUX2_X1 U6823 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7676), .Z(n5297) );
  XNOR2_X1 U6824 ( .A(n5297), .B(n5282), .ZN(n5296) );
  NAND2_X1 U6825 ( .A1(n6419), .A2(n7822), .ZN(n5286) );
  OR2_X1 U6826 ( .A1(n5301), .A2(n5079), .ZN(n5284) );
  XNOR2_X1 U6827 ( .A(n5284), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U6828 ( .A1(n5428), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5427), .B2(
        n9776), .ZN(n5285) );
  NAND2_X1 U6829 ( .A1(n5286), .A2(n5285), .ZN(n9942) );
  NAND2_X1 U6830 ( .A1(n6925), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5294) );
  INV_X1 U6831 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5287) );
  OR2_X1 U6832 ( .A1(n6926), .A2(n5287), .ZN(n5293) );
  INV_X1 U6833 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7082) );
  OR2_X1 U6834 ( .A1(n6929), .A2(n7082), .ZN(n5292) );
  NAND2_X1 U6835 ( .A1(n5288), .A2(n7475), .ZN(n5309) );
  NAND2_X1 U6836 ( .A1(n5289), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5290) );
  AND2_X1 U6837 ( .A1(n5309), .A2(n5290), .ZN(n7479) );
  OR2_X1 U6838 ( .A1(n5404), .A2(n7479), .ZN(n5291) );
  NAND4_X1 U6839 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n8190)
         );
  AND2_X1 U6840 ( .A1(n9942), .A2(n8190), .ZN(n5295) );
  INV_X1 U6841 ( .A(n5296), .ZN(n5298) );
  MUX2_X1 U6842 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6228), .Z(n5317) );
  XNOR2_X1 U6843 ( .A(n5317), .B(SI_13_), .ZN(n5315) );
  XNOR2_X1 U6844 ( .A(n5316), .B(n5315), .ZN(n6582) );
  NAND2_X1 U6845 ( .A1(n6582), .A2(n7822), .ZN(n5304) );
  NAND2_X1 U6846 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NAND2_X1 U6847 ( .A1(n5302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U6848 ( .A(n5325), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8202) );
  AOI22_X1 U6849 ( .A1(n5428), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5427), .B2(
        n8202), .ZN(n5303) );
  NAND2_X1 U6850 ( .A1(n6925), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5314) );
  INV_X1 U6851 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6852 ( .A1(n6926), .A2(n5305), .ZN(n5313) );
  INV_X1 U6853 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5306) );
  OR2_X1 U6854 ( .A1(n6929), .A2(n5306), .ZN(n5312) );
  INV_X1 U6855 ( .A(n5309), .ZN(n5308) );
  NAND2_X1 U6856 ( .A1(n5308), .A2(n5307), .ZN(n5331) );
  NAND2_X1 U6857 ( .A1(n5309), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5310) );
  AND2_X1 U6858 ( .A1(n5331), .A2(n5310), .ZN(n7465) );
  OR2_X1 U6859 ( .A1(n5404), .A2(n7465), .ZN(n5311) );
  NAND2_X1 U6860 ( .A1(n9523), .A2(n7568), .ZN(n7943) );
  NAND2_X1 U6861 ( .A1(n5317), .A2(SI_13_), .ZN(n5318) );
  INV_X1 U6862 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5320) );
  MUX2_X1 U6863 ( .A(n6663), .B(n5320), .S(n6228), .Z(n5322) );
  NAND2_X1 U6864 ( .A1(n5322), .A2(n5321), .ZN(n5339) );
  INV_X1 U6865 ( .A(n5322), .ZN(n5323) );
  NAND2_X1 U6866 ( .A1(n5323), .A2(SI_14_), .ZN(n5324) );
  NAND2_X1 U6867 ( .A1(n5339), .A2(n5324), .ZN(n5340) );
  XNOR2_X1 U6868 ( .A(n5341), .B(n5340), .ZN(n6611) );
  NAND2_X1 U6869 ( .A1(n6611), .A2(n7822), .ZN(n5330) );
  NAND2_X1 U6870 ( .A1(n5325), .A2(n10015), .ZN(n5326) );
  NAND2_X1 U6871 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6872 ( .A1(n5364), .A2(n5327), .ZN(n5342) );
  OR2_X1 U6873 ( .A1(n5364), .A2(n5327), .ZN(n5328) );
  AOI22_X1 U6874 ( .A1(n5428), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5427), .B2(
        n9793), .ZN(n5329) );
  NAND2_X1 U6875 ( .A1(n5330), .A2(n5329), .ZN(n7570) );
  NAND2_X1 U6876 ( .A1(n6925), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5337) );
  OR2_X2 U6877 ( .A1(n5331), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6878 ( .A1(n5331), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5332) );
  AND2_X1 U6879 ( .A1(n5347), .A2(n5332), .ZN(n7334) );
  OR2_X1 U6880 ( .A1(n5404), .A2(n7334), .ZN(n5336) );
  INV_X1 U6881 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6882 ( .A1(n6929), .A2(n5333), .ZN(n5335) );
  INV_X1 U6883 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8233) );
  OR2_X1 U6884 ( .A1(n6926), .A2(n8233), .ZN(n5334) );
  OR2_X1 U6885 ( .A1(n7570), .A2(n7462), .ZN(n7947) );
  NAND2_X1 U6886 ( .A1(n7570), .A2(n7462), .ZN(n7948) );
  NAND2_X1 U6887 ( .A1(n7947), .A2(n7948), .ZN(n7853) );
  AND2_X2 U6888 ( .A1(n7327), .A2(n5338), .ZN(n8428) );
  OAI21_X2 U6889 ( .B1(n5341), .B2(n5340), .A(n5339), .ZN(n5358) );
  MUX2_X1 U6890 ( .A(n6731), .B(n6747), .S(n6228), .Z(n5354) );
  XNOR2_X1 U6891 ( .A(n5354), .B(SI_15_), .ZN(n5353) );
  XNOR2_X1 U6892 ( .A(n5358), .B(n5353), .ZN(n6730) );
  NAND2_X1 U6893 ( .A1(n6730), .A2(n7822), .ZN(n5345) );
  NAND2_X1 U6894 ( .A1(n5342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5343) );
  XNOR2_X1 U6895 ( .A(n5343), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9809) );
  AOI22_X1 U6896 ( .A1(n5428), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9809), .B2(
        n5427), .ZN(n5344) );
  NAND2_X1 U6897 ( .A1(n6925), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5352) );
  INV_X1 U6898 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8476) );
  OR2_X1 U6899 ( .A1(n6926), .A2(n8476), .ZN(n5351) );
  INV_X1 U6900 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8434) );
  OR2_X1 U6901 ( .A1(n5084), .A2(n8434), .ZN(n5350) );
  NAND2_X1 U6902 ( .A1(n5347), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5348) );
  AND2_X1 U6903 ( .A1(n5367), .A2(n5348), .ZN(n8435) );
  OR2_X1 U6904 ( .A1(n5404), .A2(n8435), .ZN(n5349) );
  NAND4_X1 U6905 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n8422)
         );
  NAND2_X1 U6906 ( .A1(n8547), .A2(n8422), .ZN(n7854) );
  NOR2_X1 U6907 ( .A1(n8547), .A2(n8422), .ZN(n7856) );
  INV_X1 U6908 ( .A(n5353), .ZN(n5357) );
  INV_X1 U6909 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6910 ( .A1(n5355), .A2(SI_15_), .ZN(n5356) );
  MUX2_X1 U6911 ( .A(n6810), .B(n6808), .S(n6228), .Z(n5359) );
  NAND2_X1 U6912 ( .A1(n5359), .A2(n10108), .ZN(n5373) );
  INV_X1 U6913 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6914 ( .A1(n5360), .A2(SI_16_), .ZN(n5361) );
  NAND2_X1 U6915 ( .A1(n5373), .A2(n5361), .ZN(n5374) );
  NAND2_X1 U6916 ( .A1(n6807), .A2(n7822), .ZN(n5366) );
  NAND2_X1 U6917 ( .A1(n5362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6918 ( .A1(n5364), .A2(n5363), .ZN(n5380) );
  XNOR2_X1 U6919 ( .A(n5380), .B(n10016), .ZN(n9825) );
  AOI22_X1 U6920 ( .A1(n5428), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9825), .B2(
        n5427), .ZN(n5365) );
  NAND2_X1 U6921 ( .A1(n6925), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5372) );
  INV_X1 U6922 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10197) );
  OR2_X1 U6923 ( .A1(n5084), .A2(n10197), .ZN(n5371) );
  NAND2_X1 U6924 ( .A1(n5367), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5368) );
  AND2_X1 U6925 ( .A1(n5386), .A2(n5368), .ZN(n8118) );
  OR2_X1 U6926 ( .A1(n5404), .A2(n8118), .ZN(n5370) );
  INV_X1 U6927 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10255) );
  OR2_X1 U6928 ( .A1(n6926), .A2(n10255), .ZN(n5369) );
  NAND2_X1 U6929 ( .A1(n8540), .A2(n8169), .ZN(n7957) );
  NAND2_X1 U6930 ( .A1(n7960), .A2(n7957), .ZN(n7835) );
  MUX2_X1 U6931 ( .A(n6921), .B(n5375), .S(n6228), .Z(n5377) );
  INV_X1 U6932 ( .A(SI_17_), .ZN(n5376) );
  NAND2_X1 U6933 ( .A1(n5377), .A2(n5376), .ZN(n5394) );
  INV_X1 U6934 ( .A(n5377), .ZN(n5378) );
  NAND2_X1 U6935 ( .A1(n5378), .A2(SI_17_), .ZN(n5379) );
  NAND2_X1 U6936 ( .A1(n6878), .A2(n7822), .ZN(n5383) );
  OAI21_X1 U6937 ( .B1(n5380), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5381) );
  XNOR2_X1 U6938 ( .A(n5381), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U6939 ( .A1(n9843), .A2(n5427), .B1(n5428), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6940 ( .A1(n6925), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5391) );
  INV_X1 U6941 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10123) );
  OR2_X1 U6942 ( .A1(n6926), .A2(n10123), .ZN(n5390) );
  INV_X1 U6943 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8414) );
  OR2_X1 U6944 ( .A1(n6929), .A2(n8414), .ZN(n5389) );
  INV_X1 U6945 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6946 ( .A1(n5386), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5387) );
  AND2_X1 U6947 ( .A1(n5405), .A2(n5387), .ZN(n8129) );
  OR2_X1 U6948 ( .A1(n5404), .A2(n8129), .ZN(n5388) );
  OR2_X1 U6949 ( .A1(n8534), .A2(n8395), .ZN(n7958) );
  NAND2_X1 U6950 ( .A1(n8534), .A2(n8395), .ZN(n8397) );
  INV_X1 U6951 ( .A(n8534), .ZN(n8134) );
  NAND2_X1 U6952 ( .A1(n5393), .A2(n5392), .ZN(n5395) );
  MUX2_X1 U6953 ( .A(n6976), .B(n5396), .S(n6228), .Z(n5414) );
  XNOR2_X1 U6954 ( .A(n5414), .B(SI_18_), .ZN(n5411) );
  XNOR2_X1 U6955 ( .A(n5413), .B(n5411), .ZN(n6923) );
  NAND2_X1 U6956 ( .A1(n6923), .A2(n7822), .ZN(n5403) );
  INV_X1 U6957 ( .A(n5397), .ZN(n5400) );
  INV_X1 U6958 ( .A(n5398), .ZN(n5399) );
  OAI21_X1 U6959 ( .B1(n5400), .B2(n5399), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5401) );
  XNOR2_X1 U6960 ( .A(n5401), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8262) );
  AOI22_X1 U6961 ( .A1(n5428), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5427), .B2(
        n8262), .ZN(n5402) );
  NAND2_X1 U6962 ( .A1(n5405), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6963 ( .A1(n5432), .A2(n5406), .ZN(n8401) );
  NAND2_X1 U6964 ( .A1(n5613), .A2(n8401), .ZN(n5410) );
  INV_X1 U6965 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10165) );
  OR2_X1 U6966 ( .A1(n6926), .A2(n10165), .ZN(n5409) );
  INV_X1 U6967 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8199) );
  OR2_X1 U6968 ( .A1(n6929), .A2(n8199), .ZN(n5408) );
  INV_X1 U6969 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8528) );
  OR2_X1 U6970 ( .A1(n5455), .A2(n8528), .ZN(n5407) );
  INV_X1 U6971 ( .A(n5411), .ZN(n5412) );
  INV_X1 U6972 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6973 ( .A1(n5415), .A2(SI_18_), .ZN(n5416) );
  MUX2_X1 U6974 ( .A(n5418), .B(n10110), .S(n6228), .Z(n5419) );
  INV_X1 U6975 ( .A(SI_19_), .ZN(n10227) );
  NAND2_X1 U6976 ( .A1(n5419), .A2(n10227), .ZN(n5439) );
  INV_X1 U6977 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U6978 ( .A1(n5420), .A2(SI_19_), .ZN(n5421) );
  INV_X1 U6979 ( .A(n5422), .ZN(n5423) );
  NAND2_X1 U6980 ( .A1(n4487), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U6981 ( .A1(n5440), .A2(n5424), .ZN(n7061) );
  NAND2_X1 U6982 ( .A1(n7061), .A2(n7822), .ZN(n5430) );
  NAND2_X1 U6983 ( .A1(n5425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5426) );
  AOI22_X1 U6984 ( .A1(n5428), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8255), .B2(
        n5427), .ZN(n5429) );
  NAND2_X1 U6985 ( .A1(n5432), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6986 ( .A1(n5452), .A2(n5433), .ZN(n8387) );
  NAND2_X1 U6987 ( .A1(n8387), .A2(n5613), .ZN(n5438) );
  INV_X1 U6988 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8465) );
  OR2_X1 U6989 ( .A1(n6926), .A2(n8465), .ZN(n5435) );
  INV_X1 U6990 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8386) );
  OR2_X1 U6991 ( .A1(n5084), .A2(n8386), .ZN(n5434) );
  AND2_X1 U6992 ( .A1(n5435), .A2(n5434), .ZN(n5437) );
  INV_X1 U6993 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10170) );
  OR2_X1 U6994 ( .A1(n5455), .A2(n10170), .ZN(n5436) );
  NAND2_X1 U6995 ( .A1(n8523), .A2(n8393), .ZN(n7966) );
  INV_X1 U6996 ( .A(n8393), .ZN(n8372) );
  MUX2_X1 U6997 ( .A(n7180), .B(n7177), .S(n6228), .Z(n5442) );
  NAND2_X1 U6998 ( .A1(n5442), .A2(n5441), .ZN(n5461) );
  INV_X1 U6999 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U7000 ( .A1(n5443), .A2(SI_20_), .ZN(n5444) );
  NAND2_X1 U7001 ( .A1(n5461), .A2(n5444), .ZN(n5446) );
  NAND2_X1 U7002 ( .A1(n5445), .A2(n5446), .ZN(n5449) );
  INV_X1 U7003 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U7004 ( .A1(n5449), .A2(n5462), .ZN(n7178) );
  NAND2_X1 U7005 ( .A1(n7178), .A2(n7822), .ZN(n5451) );
  OR2_X1 U7006 ( .A1(n7825), .A2(n7180), .ZN(n5450) );
  NAND2_X1 U7007 ( .A1(n5452), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U7008 ( .A1(n5466), .A2(n5453), .ZN(n8375) );
  NAND2_X1 U7009 ( .A1(n8375), .A2(n5613), .ZN(n5458) );
  AOI22_X1 U7010 ( .A1(n5454), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n5663), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5457) );
  INV_X1 U7011 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10127) );
  OR2_X1 U7012 ( .A1(n5455), .A2(n10127), .ZN(n5456) );
  NAND2_X1 U7013 ( .A1(n8518), .A2(n8383), .ZN(n8355) );
  NAND2_X1 U7014 ( .A1(n7967), .A2(n8355), .ZN(n8370) );
  MUX2_X1 U7015 ( .A(n7271), .B(n7313), .S(n7676), .Z(n5474) );
  XNOR2_X1 U7016 ( .A(n5474), .B(SI_21_), .ZN(n5473) );
  XNOR2_X1 U7017 ( .A(n5478), .B(n5473), .ZN(n7270) );
  NAND2_X1 U7018 ( .A1(n7270), .A2(n7822), .ZN(n5464) );
  OR2_X1 U7019 ( .A1(n7825), .A2(n7271), .ZN(n5463) );
  NAND2_X1 U7020 ( .A1(n5466), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7021 ( .A1(n5502), .A2(n5467), .ZN(n8364) );
  NAND2_X1 U7022 ( .A1(n8364), .A2(n5613), .ZN(n5470) );
  AOI22_X1 U7023 ( .A1(n6925), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5454), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5469) );
  INV_X1 U7024 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10178) );
  OR2_X1 U7025 ( .A1(n6926), .A2(n10178), .ZN(n5468) );
  NAND2_X1 U7026 ( .A1(n8513), .A2(n7796), .ZN(n5648) );
  NAND2_X1 U7027 ( .A1(n7970), .A2(n5648), .ZN(n8358) );
  INV_X1 U7028 ( .A(n8513), .ZN(n8101) );
  INV_X1 U7029 ( .A(n5473), .ZN(n5477) );
  INV_X1 U7030 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U7031 ( .A1(n5475), .A2(SI_21_), .ZN(n5476) );
  MUX2_X1 U7032 ( .A(n7502), .B(n6024), .S(n6228), .Z(n5479) );
  NAND2_X1 U7033 ( .A1(n5479), .A2(n10199), .ZN(n5490) );
  INV_X1 U7034 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U7035 ( .A1(n5480), .A2(SI_22_), .ZN(n5481) );
  NAND2_X1 U7036 ( .A1(n5490), .A2(n5481), .ZN(n5491) );
  XNOR2_X1 U7037 ( .A(n5492), .B(n5491), .ZN(n10047) );
  NAND2_X1 U7038 ( .A1(n10047), .A2(n7822), .ZN(n5483) );
  OR2_X1 U7039 ( .A1(n7825), .A2(n7502), .ZN(n5482) );
  XNOR2_X1 U7040 ( .A(n5502), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U7041 ( .A1(n8348), .A2(n5613), .ZN(n5488) );
  INV_X1 U7042 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U7043 ( .A1(n5454), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7044 ( .A1(n5663), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5484) );
  OAI211_X1 U7045 ( .C1(n7797), .C2(n5455), .A(n5485), .B(n5484), .ZN(n5486)
         );
  INV_X1 U7046 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U7047 ( .A1(n8350), .A2(n8361), .ZN(n7979) );
  INV_X1 U7048 ( .A(n8350), .ZN(n5489) );
  INV_X1 U7049 ( .A(n8361), .ZN(n7750) );
  NAND2_X1 U7050 ( .A1(n5489), .A2(n7750), .ZN(n7977) );
  INV_X1 U7051 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7526) );
  MUX2_X1 U7052 ( .A(n10258), .B(n7526), .S(n6228), .Z(n5494) );
  INV_X1 U7053 ( .A(SI_23_), .ZN(n5493) );
  NAND2_X1 U7054 ( .A1(n5494), .A2(n5493), .ZN(n5548) );
  INV_X1 U7055 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U7056 ( .A1(n5495), .A2(SI_23_), .ZN(n5496) );
  OR2_X1 U7057 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U7058 ( .A1(n5550), .A2(n5499), .ZN(n7524) );
  NAND2_X1 U7059 ( .A1(n7524), .A2(n7822), .ZN(n5501) );
  OR2_X1 U7060 ( .A1(n7825), .A2(n10258), .ZN(n5500) );
  NAND2_X1 U7061 ( .A1(n5503), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7062 ( .A1(n5519), .A2(n5504), .ZN(n8344) );
  NAND2_X1 U7063 ( .A1(n8344), .A2(n5613), .ZN(n5509) );
  INV_X1 U7064 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10065) );
  NAND2_X1 U7065 ( .A1(n6925), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7066 ( .A1(n5454), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5505) );
  OAI211_X1 U7067 ( .C1(n6926), .C2(n10065), .A(n5506), .B(n5505), .ZN(n5507)
         );
  INV_X1 U7068 ( .A(n5507), .ZN(n5508) );
  NOR2_X1 U7069 ( .A1(n8507), .A2(n8188), .ZN(n5510) );
  INV_X1 U7070 ( .A(n8507), .ZN(n5649) );
  NAND2_X1 U7071 ( .A1(n5550), .A2(n5548), .ZN(n5527) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7649) );
  INV_X1 U7073 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U7074 ( .A(n7649), .B(n7600), .S(n6228), .Z(n5512) );
  INV_X1 U7075 ( .A(SI_24_), .ZN(n5511) );
  NAND2_X1 U7076 ( .A1(n5512), .A2(n5511), .ZN(n5545) );
  INV_X1 U7077 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U7078 ( .A1(n5513), .A2(SI_24_), .ZN(n5514) );
  NAND2_X1 U7079 ( .A1(n7599), .A2(n7822), .ZN(n5516) );
  OR2_X1 U7080 ( .A1(n7825), .A2(n7649), .ZN(n5515) );
  INV_X1 U7081 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7082 ( .A1(n5519), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7083 ( .A1(n5537), .A2(n5520), .ZN(n8333) );
  NAND2_X1 U7084 ( .A1(n8333), .A2(n5613), .ZN(n5525) );
  INV_X1 U7085 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U7086 ( .A1(n5663), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7087 ( .A1(n5454), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5521) );
  OAI211_X1 U7088 ( .C1(n10269), .C2(n5455), .A(n5522), .B(n5521), .ZN(n5523)
         );
  INV_X1 U7089 ( .A(n5523), .ZN(n5524) );
  NOR2_X1 U7090 ( .A1(n8501), .A2(n8077), .ZN(n5526) );
  NAND2_X1 U7091 ( .A1(n5527), .A2(n5553), .ZN(n5528) );
  NAND2_X1 U7092 ( .A1(n5528), .A2(n5545), .ZN(n5532) );
  INV_X1 U7093 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10247) );
  INV_X1 U7094 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7615) );
  MUX2_X1 U7095 ( .A(n10247), .B(n7615), .S(n6228), .Z(n5529) );
  NAND2_X1 U7096 ( .A1(n5529), .A2(n10194), .ZN(n5544) );
  INV_X1 U7097 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7098 ( .A1(n5530), .A2(SI_25_), .ZN(n5552) );
  AND2_X1 U7099 ( .A1(n5544), .A2(n5552), .ZN(n5531) );
  NAND2_X1 U7100 ( .A1(n7614), .A2(n7822), .ZN(n5534) );
  OR2_X1 U7101 ( .A1(n7825), .A2(n10247), .ZN(n5533) );
  INV_X1 U7102 ( .A(n5537), .ZN(n5536) );
  INV_X1 U7103 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7104 ( .A1(n5537), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7105 ( .A1(n5562), .A2(n5538), .ZN(n8111) );
  NAND2_X1 U7106 ( .A1(n8111), .A2(n5613), .ZN(n5543) );
  INV_X1 U7107 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U7108 ( .A1(n6925), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7109 ( .A1(n5454), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U7110 ( .C1(n6926), .C2(n10089), .A(n5540), .B(n5539), .ZN(n5541)
         );
  INV_X1 U7111 ( .A(n5541), .ZN(n5542) );
  INV_X1 U7112 ( .A(n8038), .ZN(n8114) );
  INV_X1 U7113 ( .A(n5552), .ZN(n5547) );
  AND2_X1 U7114 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  AND2_X1 U7115 ( .A1(n5548), .A2(n5551), .ZN(n5549) );
  INV_X1 U7116 ( .A(n5551), .ZN(n5555) );
  AND2_X1 U7117 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7666) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7612) );
  MUX2_X1 U7120 ( .A(n7666), .B(n7612), .S(n7676), .Z(n5557) );
  INV_X1 U7121 ( .A(SI_26_), .ZN(n5556) );
  NAND2_X1 U7122 ( .A1(n5557), .A2(n5556), .ZN(n5571) );
  INV_X1 U7123 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U7124 ( .A1(n5558), .A2(SI_26_), .ZN(n5559) );
  NAND2_X1 U7125 ( .A1(n7611), .A2(n7822), .ZN(n5561) );
  OR2_X1 U7126 ( .A1(n7825), .A2(n7666), .ZN(n5560) );
  NAND2_X1 U7127 ( .A1(n5562), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7128 ( .A1(n5583), .A2(n5563), .ZN(n8324) );
  NAND2_X1 U7129 ( .A1(n8324), .A2(n5613), .ZN(n5568) );
  INV_X1 U7130 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U7131 ( .A1(n5454), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5565) );
  INV_X1 U7132 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10266) );
  OR2_X1 U7133 ( .A1(n6926), .A2(n10266), .ZN(n5564) );
  OAI211_X1 U7134 ( .C1(n10243), .C2(n5455), .A(n5565), .B(n5564), .ZN(n5566)
         );
  INV_X1 U7135 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7136 ( .A1(n5570), .A2(n5569), .ZN(n5572) );
  NAND2_X1 U7137 ( .A1(n5572), .A2(n5571), .ZN(n5577) );
  MUX2_X1 U7138 ( .A(n8036), .B(n6073), .S(n6228), .Z(n5573) );
  INV_X1 U7139 ( .A(SI_27_), .ZN(n10207) );
  NAND2_X1 U7140 ( .A1(n5573), .A2(n10207), .ZN(n5590) );
  INV_X1 U7141 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7142 ( .A1(n5574), .A2(SI_27_), .ZN(n5575) );
  NAND2_X1 U7143 ( .A1(n5577), .A2(n5576), .ZN(n5591) );
  OR2_X1 U7144 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  NAND2_X1 U7145 ( .A1(n5591), .A2(n5578), .ZN(n7818) );
  NAND2_X1 U7146 ( .A1(n7818), .A2(n7822), .ZN(n5580) );
  OR2_X1 U7147 ( .A1(n7825), .A2(n8036), .ZN(n5579) );
  INV_X1 U7148 ( .A(n5583), .ZN(n5582) );
  INV_X1 U7149 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7150 ( .A1(n5582), .A2(n5581), .ZN(n5595) );
  NAND2_X1 U7151 ( .A1(n5583), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7152 ( .A1(n5595), .A2(n5584), .ZN(n8312) );
  NAND2_X1 U7153 ( .A1(n8312), .A2(n5613), .ZN(n5589) );
  INV_X1 U7154 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U7155 ( .A1(n6925), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7156 ( .A1(n5454), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7157 ( .C1(n6926), .C2(n10067), .A(n5586), .B(n5585), .ZN(n5587)
         );
  INV_X1 U7158 ( .A(n5587), .ZN(n5588) );
  NOR2_X1 U7159 ( .A1(n8452), .A2(n8320), .ZN(n5654) );
  NAND2_X1 U7160 ( .A1(n8452), .A2(n8320), .ZN(n8000) );
  NAND2_X1 U7161 ( .A1(n5591), .A2(n5590), .ZN(n5606) );
  MUX2_X1 U7162 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7676), .Z(n5607) );
  INV_X1 U7163 ( .A(SI_28_), .ZN(n10182) );
  XNOR2_X1 U7164 ( .A(n5607), .B(n10182), .ZN(n5605) );
  XNOR2_X1 U7165 ( .A(n5606), .B(n5605), .ZN(n8053) );
  NAND2_X1 U7166 ( .A1(n8053), .A2(n7822), .ZN(n5594) );
  INV_X1 U7167 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5592) );
  OR2_X1 U7168 ( .A1(n7825), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U7169 ( .A1(n5595), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7170 ( .A1(n8274), .A2(n5596), .ZN(n8048) );
  NAND2_X1 U7171 ( .A1(n8048), .A2(n5613), .ZN(n5601) );
  INV_X1 U7172 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U7173 ( .A1(n5663), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7174 ( .A1(n5454), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5597) );
  OAI211_X1 U7175 ( .C1(n10237), .C2(n5455), .A(n5598), .B(n5597), .ZN(n5599)
         );
  INV_X1 U7176 ( .A(n5599), .ZN(n5600) );
  NOR2_X1 U7177 ( .A1(n5602), .A2(n8306), .ZN(n5604) );
  OAI21_X1 U7178 ( .B1(n8292), .B2(n5604), .A(n5603), .ZN(n5619) );
  NAND2_X1 U7179 ( .A1(n5606), .A2(n5605), .ZN(n5610) );
  INV_X1 U7180 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7181 ( .A1(n5608), .A2(n10182), .ZN(n5609) );
  INV_X1 U7182 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7651) );
  INV_X1 U7183 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9477) );
  MUX2_X1 U7184 ( .A(n7651), .B(n9477), .S(n6228), .Z(n7655) );
  NAND2_X1 U7185 ( .A1(n7681), .A2(n7822), .ZN(n5612) );
  OR2_X1 U7186 ( .A1(n7825), .A2(n7651), .ZN(n5611) );
  INV_X1 U7187 ( .A(n8274), .ZN(n5614) );
  NAND2_X1 U7188 ( .A1(n5614), .A2(n5613), .ZN(n6932) );
  INV_X1 U7189 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U7190 ( .A1(n5454), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5616) );
  INV_X1 U7191 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10209) );
  OR2_X1 U7192 ( .A1(n6926), .A2(n10209), .ZN(n5615) );
  OAI211_X1 U7193 ( .C1(n5455), .C2(n10091), .A(n5616), .B(n5615), .ZN(n5617)
         );
  INV_X1 U7194 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7195 ( .A1(n6932), .A2(n5618), .ZN(n8185) );
  XNOR2_X1 U7196 ( .A(n7828), .B(n8185), .ZN(n7867) );
  INV_X1 U7197 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7198 ( .A1(n5621), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7199 ( .A1(n8030), .A2(n8255), .ZN(n5705) );
  NAND2_X1 U7200 ( .A1(n5624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7201 ( .A1(n5626), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5627) );
  MUX2_X1 U7202 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5627), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5628) );
  INV_X1 U7203 ( .A(n8024), .ZN(n5629) );
  NAND2_X1 U7204 ( .A1(n7833), .A2(n5629), .ZN(n5630) );
  INV_X1 U7205 ( .A(n8193), .ZN(n7055) );
  NAND2_X1 U7206 ( .A1(n9917), .A2(n7055), .ZN(n7896) );
  INV_X1 U7207 ( .A(n7896), .ZN(n5631) );
  OR2_X1 U7208 ( .A1(n9917), .A2(n7055), .ZN(n7897) );
  AND2_X1 U7209 ( .A1(n7916), .A2(n7896), .ZN(n7013) );
  NAND2_X1 U7210 ( .A1(n9862), .A2(n7839), .ZN(n5636) );
  OR2_X1 U7211 ( .A1(n8198), .A2(n9884), .ZN(n7874) );
  NAND2_X1 U7212 ( .A1(n5636), .A2(n7874), .ZN(n6763) );
  NAND2_X1 U7213 ( .A1(n6763), .A2(n5103), .ZN(n6762) );
  INV_X1 U7214 ( .A(n7838), .ZN(n7905) );
  NAND2_X1 U7215 ( .A1(n6734), .A2(n7905), .ZN(n5637) );
  INV_X1 U7216 ( .A(n6758), .ZN(n9899) );
  OR2_X1 U7217 ( .A1(n8196), .A2(n9899), .ZN(n6868) );
  NAND2_X1 U7218 ( .A1(n8196), .A2(n9899), .ZN(n7910) );
  NAND2_X1 U7219 ( .A1(n6748), .A2(n7842), .ZN(n6869) );
  AND2_X1 U7220 ( .A1(n7911), .A2(n6868), .ZN(n7908) );
  NAND2_X1 U7221 ( .A1(n6869), .A2(n7908), .ZN(n6811) );
  OR2_X1 U7222 ( .A1(n9925), .A2(n7449), .ZN(n7923) );
  NAND2_X1 U7223 ( .A1(n9925), .A2(n7449), .ZN(n7924) );
  NAND2_X1 U7224 ( .A1(n7923), .A2(n7924), .ZN(n7849) );
  NAND2_X1 U7225 ( .A1(n5639), .A2(n5638), .ZN(n6886) );
  NAND2_X1 U7226 ( .A1(n9936), .A2(n7476), .ZN(n7931) );
  INV_X1 U7227 ( .A(n8422), .ZN(n8120) );
  NAND2_X1 U7228 ( .A1(n8547), .A2(n8120), .ZN(n7952) );
  OR2_X1 U7229 ( .A1(n8547), .A2(n8120), .ZN(n7953) );
  INV_X1 U7230 ( .A(n7958), .ZN(n5642) );
  NAND2_X1 U7231 ( .A1(n5643), .A2(n8382), .ZN(n7961) );
  NAND2_X1 U7232 ( .A1(n7964), .A2(n7961), .ZN(n8390) );
  INV_X1 U7233 ( .A(n8397), .ZN(n5644) );
  NOR2_X1 U7234 ( .A1(n8390), .A2(n5644), .ZN(n5645) );
  AND2_X1 U7235 ( .A1(n5648), .A2(n8355), .ZN(n7972) );
  NAND2_X1 U7236 ( .A1(n8507), .A2(n8332), .ZN(n7978) );
  INV_X1 U7237 ( .A(n7988), .ZN(n5650) );
  NAND2_X1 U7238 ( .A1(n5653), .A2(n7998), .ZN(n8309) );
  INV_X1 U7239 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7240 ( .A1(n5655), .A2(n8000), .ZN(n8308) );
  OR2_X1 U7241 ( .A1(n8452), .A2(n8294), .ZN(n5656) );
  NAND2_X1 U7242 ( .A1(n8448), .A2(n8306), .ZN(n5658) );
  NAND2_X1 U7243 ( .A1(n8024), .A2(n8265), .ZN(n6183) );
  NAND2_X1 U7244 ( .A1(n8030), .A2(n8265), .ZN(n5715) );
  NAND2_X1 U7245 ( .A1(n5715), .A2(n6183), .ZN(n5659) );
  INV_X1 U7246 ( .A(n5660), .ZN(n8027) );
  NAND2_X1 U7247 ( .A1(n8027), .A2(n6273), .ZN(n5662) );
  NAND2_X1 U7248 ( .A1(n5080), .A2(n5662), .ZN(n6217) );
  INV_X1 U7249 ( .A(n6217), .ZN(n6216) );
  INV_X1 U7250 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7251 ( .A1(n5663), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7252 ( .A1(n5454), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5664) );
  OAI211_X1 U7253 ( .C1(n5666), .C2(n5455), .A(n5665), .B(n5664), .ZN(n5667)
         );
  INV_X1 U7254 ( .A(n5667), .ZN(n5668) );
  NAND2_X1 U7255 ( .A1(n6932), .A2(n5668), .ZN(n8184) );
  AND2_X1 U7256 ( .A1(n5080), .A2(P2_B_REG_SCAN_IN), .ZN(n5669) );
  NOR2_X1 U7257 ( .A1(n8394), .A2(n5669), .ZN(n8271) );
  AOI22_X1 U7258 ( .A1(n9866), .A2(n8186), .B1(n8184), .B2(n8271), .ZN(n5670)
         );
  NAND2_X1 U7259 ( .A1(n5671), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7260 ( .A1(n5704), .A2(n5703), .ZN(n5672) );
  XNOR2_X1 U7261 ( .A(n5683), .B(P2_B_REG_SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7262 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U7263 ( .A1(n5678), .A2(n8033), .ZN(n5685) );
  INV_X1 U7264 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5681) );
  AND2_X1 U7265 ( .A1(n5681), .A2(n5699), .ZN(n5682) );
  XOR2_X1 U7266 ( .A(n5684), .B(P2_IR_REG_26__SCAN_IN), .Z(n7667) );
  NAND2_X1 U7267 ( .A1(n5683), .A2(n7667), .ZN(n6248) );
  NAND2_X1 U7268 ( .A1(n6181), .A2(n6248), .ZN(n6645) );
  NAND2_X1 U7269 ( .A1(n5685), .A2(n5699), .ZN(n6243) );
  OR2_X1 U7270 ( .A1(n6243), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7271 ( .A1(n8033), .A2(n7667), .ZN(n6245) );
  INV_X1 U7272 ( .A(n6649), .ZN(n5687) );
  NOR2_X1 U7273 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n10018) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5690) );
  NOR4_X1 U7275 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5689) );
  NOR4_X1 U7276 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5688) );
  AND4_X1 U7277 ( .A1(n10018), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n5696)
         );
  NOR4_X1 U7278 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5694) );
  NOR4_X1 U7279 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7280 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7281 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5691) );
  AND4_X1 U7282 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n5695)
         );
  AND2_X1 U7283 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  INV_X1 U7284 ( .A(n5719), .ZN(n5698) );
  INV_X1 U7285 ( .A(n8033), .ZN(n5702) );
  INV_X1 U7286 ( .A(n5683), .ZN(n5700) );
  OR2_X1 U7287 ( .A1(n6212), .A2(n6655), .ZN(n6214) );
  OAI21_X1 U7288 ( .B1(n6212), .B2(n6194), .A(n6214), .ZN(n5706) );
  NAND2_X1 U7289 ( .A1(n6209), .A2(n5706), .ZN(n5711) );
  NAND2_X1 U7290 ( .A1(n6645), .A2(n5719), .ZN(n5707) );
  INV_X1 U7291 ( .A(n6215), .ZN(n5709) );
  INV_X1 U7292 ( .A(n6212), .ZN(n6244) );
  AND2_X1 U7293 ( .A1(n8007), .A2(n9919), .ZN(n6192) );
  NAND2_X1 U7294 ( .A1(n6192), .A2(n6194), .ZN(n5708) );
  OR2_X1 U7295 ( .A1(n9919), .A2(n6678), .ZN(n9864) );
  NAND2_X1 U7296 ( .A1(n5708), .A2(n9864), .ZN(n6199) );
  NAND3_X1 U7297 ( .A1(n5709), .A2(n6244), .A3(n6199), .ZN(n5710) );
  NAND2_X1 U7298 ( .A1(n5727), .A2(n9946), .ZN(n5713) );
  OR2_X1 U7299 ( .A1(n9946), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7300 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  NAND2_X1 U7301 ( .A1(n5714), .A2(n4998), .ZN(P2_U3456) );
  AND2_X1 U7302 ( .A1(n9926), .A2(n7837), .ZN(n6210) );
  NOR2_X1 U7303 ( .A1(n6645), .A2(n6210), .ZN(n5717) );
  OR2_X1 U7304 ( .A1(n5715), .A2(n8024), .ZN(n5716) );
  AND2_X1 U7305 ( .A1(n5716), .A2(n8007), .ZN(n6646) );
  MUX2_X1 U7306 ( .A(n6649), .B(n5717), .S(n6646), .Z(n5722) );
  AND2_X1 U7307 ( .A1(n8005), .A2(n6183), .ZN(n6202) );
  NOR2_X1 U7308 ( .A1(n6212), .A2(n6202), .ZN(n5718) );
  AND2_X1 U7309 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NOR2_X2 U7310 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5951) );
  NOR2_X1 U7311 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5732) );
  NOR2_X1 U7312 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5731) );
  NOR2_X1 U7313 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5730) );
  NAND4_X1 U7314 ( .A1(n5951), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5736)
         );
  NAND4_X1 U7315 ( .A1(n5734), .A2(n5733), .A3(n5948), .A4(n5955), .ZN(n5735)
         );
  INV_X1 U7316 ( .A(n6097), .ZN(n6099) );
  INV_X1 U7317 ( .A(n5743), .ZN(n5740) );
  INV_X1 U7318 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5745) );
  INV_X2 U7319 ( .A(n5843), .ZN(n5855) );
  NAND2_X1 U7320 ( .A1(n7270), .A2(n5855), .ZN(n5749) );
  OR2_X1 U7321 ( .A1(n7682), .A2(n7313), .ZN(n5748) );
  INV_X1 U7322 ( .A(n9390), .ZN(n9290) );
  NAND2_X1 U7323 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5833) );
  NOR2_X1 U7324 ( .A1(n5833), .A2(n7698), .ZN(n5846) );
  NAND2_X1 U7325 ( .A1(n5846), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7326 ( .A1(n5900), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7327 ( .A1(n5924), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7328 ( .A1(n6019), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7329 ( .A1(n6019), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7330 ( .A1(n6027), .A2(n5750), .ZN(n9286) );
  NOR2_X2 U7331 ( .A1(n6099), .A2(n5752), .ZN(n9467) );
  AOI22_X1 U7332 ( .A1(n5804), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n7713), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7333 ( .A1(n6293), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5757) );
  OAI211_X1 U7334 ( .C1(n9286), .C2(n5940), .A(n5758), .B(n5757), .ZN(n9056)
         );
  INV_X1 U7335 ( .A(n9056), .ZN(n8814) );
  NAND2_X1 U7336 ( .A1(n6730), .A2(n5855), .ZN(n5765) );
  NAND2_X1 U7337 ( .A1(n4430), .A2(n5948), .ZN(n5879) );
  INV_X1 U7338 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5759) );
  NAND4_X1 U7339 ( .A1(n5949), .A2(n5759), .A3(n5955), .A4(n5954), .ZN(n5760)
         );
  OAI21_X1 U7340 ( .B1(n5919), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5932) );
  INV_X1 U7341 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7342 ( .A1(n5932), .A2(n5761), .ZN(n5762) );
  NAND2_X1 U7343 ( .A1(n5762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5763) );
  XNOR2_X1 U7344 ( .A(n5763), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9587) );
  AOI22_X1 U7345 ( .A1(n6003), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6002), .B2(
        n9587), .ZN(n5764) );
  INV_X1 U7346 ( .A(n7541), .ZN(n7511) );
  INV_X1 U7347 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9579) );
  OR2_X1 U7348 ( .A1(n6133), .A2(n9579), .ZN(n5770) );
  AND2_X1 U7349 ( .A1(n5939), .A2(n10272), .ZN(n5766) );
  OR2_X1 U7350 ( .A1(n5766), .A2(n5963), .ZN(n7537) );
  OR2_X1 U7351 ( .A1(n5940), .A2(n7537), .ZN(n5769) );
  NAND2_X1 U7352 ( .A1(n7713), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7353 ( .A1(n6293), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5767) );
  NAND4_X1 U7354 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n9061)
         );
  NAND2_X1 U7355 ( .A1(n6293), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5777) );
  INV_X1 U7356 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7181) );
  OR2_X1 U7357 ( .A1(n6133), .A2(n7181), .ZN(n5776) );
  INV_X1 U7358 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7359) );
  OR2_X1 U7359 ( .A1(n6065), .A2(n7359), .ZN(n5775) );
  INV_X1 U7360 ( .A(n5924), .ZN(n5773) );
  NAND2_X1 U7361 ( .A1(n5914), .A2(n5771), .ZN(n5772) );
  NAND2_X1 U7362 ( .A1(n5773), .A2(n5772), .ZN(n7358) );
  OR2_X1 U7363 ( .A1(n5940), .A2(n7358), .ZN(n5774) );
  INV_X1 U7364 ( .A(n7276), .ZN(n9064) );
  NAND2_X1 U7365 ( .A1(n6419), .A2(n5855), .ZN(n5783) );
  NAND2_X1 U7366 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  MUX2_X1 U7367 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5779), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5780) );
  NAND2_X1 U7368 ( .A1(n5780), .A2(n5919), .ZN(n7195) );
  INV_X1 U7369 ( .A(n7195), .ZN(n5781) );
  AOI22_X1 U7370 ( .A1(n6003), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6002), .B2(
        n5781), .ZN(n5782) );
  NAND2_X1 U7371 ( .A1(n5812), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7372 ( .A1(n5804), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5784) );
  INV_X1 U7373 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5787) );
  OR2_X1 U7374 ( .A1(n5940), .A2(n5787), .ZN(n5788) );
  INV_X1 U7375 ( .A(n5790), .ZN(n6229) );
  INV_X1 U7376 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7377 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5791) );
  XNOR2_X1 U7378 ( .A(n5792), .B(n5791), .ZN(n6373) );
  NAND2_X1 U7379 ( .A1(n5812), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7380 ( .A1(n5804), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7381 ( .A1(n6293), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5796) );
  INV_X1 U7382 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7314) );
  OR2_X1 U7383 ( .A1(n5940), .A2(n7314), .ZN(n5795) );
  INV_X1 U7384 ( .A(SI_0_), .ZN(n5799) );
  INV_X1 U7385 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5798) );
  OAI21_X1 U7386 ( .B1(n7671), .B2(n5799), .A(n5798), .ZN(n5801) );
  AND2_X1 U7387 ( .A1(n5800), .A2(n5801), .ZN(n9479) );
  MUX2_X1 U7388 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9479), .S(n7677), .Z(n7324) );
  NAND2_X1 U7389 ( .A1(n6723), .A2(n7324), .ZN(n6437) );
  NAND2_X1 U7390 ( .A1(n6436), .A2(n5803), .ZN(n6451) );
  NAND2_X1 U7391 ( .A1(n5812), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6110) );
  INV_X1 U7392 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6473) );
  OR2_X1 U7393 ( .A1(n5940), .A2(n6473), .ZN(n6109) );
  NAND2_X1 U7394 ( .A1(n6293), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7395 ( .A1(n5804), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6107) );
  NAND4_X1 U7396 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n9073)
         );
  OR2_X1 U7397 ( .A1(n5843), .A2(n6234), .ZN(n5811) );
  OR2_X1 U7398 ( .A1(n5805), .A2(n6235), .ZN(n5810) );
  OR2_X1 U7399 ( .A1(n5806), .A2(n5745), .ZN(n5808) );
  INV_X1 U7400 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7401 ( .A1(n5808), .A2(n5807), .ZN(n5817) );
  OAI21_X1 U7402 ( .B1(n5808), .B2(n5807), .A(n5817), .ZN(n6372) );
  OR2_X1 U7403 ( .A1(n7677), .A2(n6372), .ZN(n5809) );
  XNOR2_X1 U7404 ( .A(n9073), .B(n7090), .ZN(n8857) );
  NAND2_X1 U7405 ( .A1(n6450), .A2(n5001), .ZN(n6522) );
  NAND2_X1 U7406 ( .A1(n5812), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5816) );
  OR2_X1 U7407 ( .A1(n5940), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7408 ( .A1(n5804), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7409 ( .A1(n6293), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5813) );
  NAND4_X1 U7410 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n9072)
         );
  OR2_X1 U7411 ( .A1(n5843), .A2(n6230), .ZN(n5822) );
  OR2_X1 U7412 ( .A1(n5805), .A2(n6231), .ZN(n5821) );
  NAND2_X1 U7413 ( .A1(n5817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5819) );
  INV_X1 U7414 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U7415 ( .A(n5819), .B(n5818), .ZN(n6393) );
  OR2_X1 U7416 ( .A1(n7677), .A2(n6393), .ZN(n5820) );
  XNOR2_X1 U7417 ( .A(n9072), .B(n7074), .ZN(n8858) );
  NAND2_X1 U7418 ( .A1(n6522), .A2(n8858), .ZN(n6521) );
  INV_X1 U7419 ( .A(n7074), .ZN(n6573) );
  NAND2_X1 U7420 ( .A1(n6521), .A2(n5003), .ZN(n6511) );
  NAND2_X1 U7421 ( .A1(n5804), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5825) );
  OAI21_X1 U7422 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5833), .ZN(n8755) );
  OR2_X1 U7423 ( .A1(n5940), .A2(n8755), .ZN(n5824) );
  NAND2_X1 U7424 ( .A1(n7713), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5823) );
  OR2_X1 U7425 ( .A1(n5843), .A2(n6232), .ZN(n5832) );
  OR2_X1 U7426 ( .A1(n7682), .A2(n6233), .ZN(n5831) );
  NAND2_X1 U7427 ( .A1(n5826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5827) );
  MUX2_X1 U7428 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5827), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5829) );
  NAND2_X1 U7429 ( .A1(n5829), .A2(n5828), .ZN(n6389) );
  OR2_X1 U7430 ( .A1(n7677), .A2(n6389), .ZN(n5830) );
  NAND2_X1 U7431 ( .A1(n6509), .A2(n5004), .ZN(n6585) );
  NAND2_X1 U7432 ( .A1(n5804), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5840) );
  INV_X1 U7433 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6479) );
  OR2_X1 U7434 ( .A1(n6065), .A2(n6479), .ZN(n5839) );
  AND2_X1 U7435 ( .A1(n5833), .A2(n7698), .ZN(n5834) );
  OR2_X1 U7436 ( .A1(n5834), .A2(n5846), .ZN(n7249) );
  OR2_X1 U7437 ( .A1(n5940), .A2(n7249), .ZN(n5838) );
  INV_X1 U7438 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5836) );
  OR2_X1 U7439 ( .A1(n5835), .A2(n5836), .ZN(n5837) );
  NAND2_X1 U7440 ( .A1(n5828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5842) );
  INV_X1 U7441 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7442 ( .A(n5842), .B(n5841), .ZN(n9099) );
  OR2_X1 U7443 ( .A1(n7682), .A2(n6236), .ZN(n5844) );
  NAND2_X1 U7444 ( .A1(n6791), .A2(n6586), .ZN(n8909) );
  INV_X1 U7445 ( .A(n6791), .ZN(n9071) );
  NAND2_X1 U7446 ( .A1(n8909), .A2(n8911), .ZN(n8856) );
  NAND2_X1 U7447 ( .A1(n6791), .A2(n7704), .ZN(n5845) );
  NAND2_X1 U7448 ( .A1(n5804), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5852) );
  INV_X1 U7449 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7109) );
  OR2_X1 U7450 ( .A1(n6065), .A2(n7109), .ZN(n5851) );
  OR2_X1 U7451 ( .A1(n5846), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7452 ( .A1(n5860), .A2(n5847), .ZN(n7110) );
  OR2_X1 U7453 ( .A1(n5940), .A2(n7110), .ZN(n5850) );
  INV_X1 U7454 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5848) );
  OR2_X1 U7455 ( .A1(n5835), .A2(n5848), .ZN(n5849) );
  OR2_X1 U7456 ( .A1(n5959), .A2(n5745), .ZN(n5854) );
  XNOR2_X1 U7457 ( .A(n5854), .B(n5853), .ZN(n9113) );
  NAND2_X1 U7458 ( .A1(n6239), .A2(n5855), .ZN(n5857) );
  INV_X1 U7459 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6242) );
  OR2_X1 U7460 ( .A1(n7682), .A2(n6242), .ZN(n5856) );
  OAI211_X1 U7461 ( .C1(n7677), .C2(n9113), .A(n5857), .B(n5856), .ZN(n6918)
         );
  NAND2_X1 U7462 ( .A1(n6801), .A2(n6918), .ZN(n8914) );
  NAND2_X1 U7463 ( .A1(n9070), .A2(n7111), .ZN(n8910) );
  NAND2_X1 U7464 ( .A1(n8914), .A2(n8910), .ZN(n8855) );
  NAND2_X1 U7465 ( .A1(n6293), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7466 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U7467 ( .A1(n5873), .A2(n5861), .ZN(n9622) );
  OR2_X1 U7468 ( .A1(n5940), .A2(n9622), .ZN(n5865) );
  INV_X1 U7469 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9623) );
  OR2_X1 U7470 ( .A1(n6065), .A2(n9623), .ZN(n5864) );
  INV_X1 U7471 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5862) );
  OR2_X1 U7472 ( .A1(n6133), .A2(n5862), .ZN(n5863) );
  NAND2_X1 U7473 ( .A1(n6251), .A2(n5855), .ZN(n5869) );
  OR2_X1 U7474 ( .A1(n4430), .A2(n5745), .ZN(n5867) );
  XNOR2_X1 U7475 ( .A(n5867), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9498) );
  AOI22_X1 U7476 ( .A1(n6003), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6002), .B2(
        n9498), .ZN(n5868) );
  NAND2_X1 U7477 ( .A1(n5869), .A2(n5868), .ZN(n9626) );
  NAND2_X1 U7478 ( .A1(n6898), .A2(n9626), .ZN(n6893) );
  INV_X1 U7479 ( .A(n6898), .ZN(n9069) );
  NAND2_X1 U7480 ( .A1(n6835), .A2(n9069), .ZN(n6116) );
  NAND2_X1 U7481 ( .A1(n6893), .A2(n6116), .ZN(n6826) );
  NAND2_X1 U7482 ( .A1(n6293), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5878) );
  INV_X1 U7483 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7484 ( .A1(n6065), .A2(n5870), .ZN(n5877) );
  INV_X1 U7485 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5871) );
  OR2_X1 U7486 ( .A1(n6133), .A2(n5871), .ZN(n5876) );
  NAND2_X1 U7487 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  NAND2_X1 U7488 ( .A1(n5887), .A2(n5874), .ZN(n7146) );
  OR2_X1 U7489 ( .A1(n5940), .A2(n7146), .ZN(n5875) );
  NAND2_X1 U7490 ( .A1(n5879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U7491 ( .A(n5897), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9512) );
  AOI22_X1 U7492 ( .A1(n6003), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6002), .B2(
        n9512), .ZN(n5880) );
  OR2_X1 U7493 ( .A1(n6966), .A2(n6964), .ZN(n8920) );
  NAND2_X1 U7494 ( .A1(n8920), .A2(n8923), .ZN(n6896) );
  NAND2_X1 U7495 ( .A1(n6890), .A2(n6896), .ZN(n6889) );
  NAND2_X1 U7496 ( .A1(n6889), .A2(n5881), .ZN(n7344) );
  NAND2_X1 U7497 ( .A1(n6301), .A2(n5855), .ZN(n5885) );
  NAND2_X1 U7498 ( .A1(n5897), .A2(n5954), .ZN(n5882) );
  NAND2_X1 U7499 ( .A1(n5882), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7500 ( .A(n5883), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9136) );
  AOI22_X1 U7501 ( .A1(n6003), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6002), .B2(
        n9136), .ZN(n5884) );
  NAND2_X1 U7502 ( .A1(n5885), .A2(n5884), .ZN(n7352) );
  NAND2_X1 U7503 ( .A1(n6293), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5893) );
  INV_X1 U7504 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7505 ( .A1(n6133), .A2(n5886), .ZN(n5892) );
  INV_X1 U7506 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7350) );
  OR2_X1 U7507 ( .A1(n6065), .A2(n7350), .ZN(n5891) );
  INV_X1 U7508 ( .A(n5900), .ZN(n5889) );
  NAND2_X1 U7509 ( .A1(n5887), .A2(n10200), .ZN(n5888) );
  NAND2_X1 U7510 ( .A1(n5889), .A2(n5888), .ZN(n7349) );
  OR2_X1 U7511 ( .A1(n5940), .A2(n7349), .ZN(n5890) );
  OR2_X1 U7512 ( .A1(n7352), .A2(n6980), .ZN(n8926) );
  NAND2_X1 U7513 ( .A1(n7352), .A2(n6980), .ZN(n8944) );
  NAND2_X1 U7514 ( .A1(n8926), .A2(n8944), .ZN(n7343) );
  INV_X1 U7515 ( .A(n6980), .ZN(n9067) );
  NAND2_X1 U7516 ( .A1(n5894), .A2(n6980), .ZN(n5895) );
  NAND2_X1 U7517 ( .A1(n6305), .A2(n5855), .ZN(n5899) );
  OAI21_X1 U7518 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7519 ( .A1(n5897), .A2(n5896), .ZN(n5908) );
  XNOR2_X1 U7520 ( .A(n5908), .B(n5949), .ZN(n9488) );
  AOI22_X1 U7521 ( .A1(n6003), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6002), .B2(
        n9488), .ZN(n5898) );
  NAND2_X1 U7522 ( .A1(n5899), .A2(n5898), .ZN(n7373) );
  NAND2_X1 U7523 ( .A1(n5804), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5906) );
  INV_X1 U7524 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7369) );
  OR2_X1 U7525 ( .A1(n6065), .A2(n7369), .ZN(n5905) );
  OR2_X1 U7526 ( .A1(n5900), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7527 ( .A1(n5912), .A2(n5901), .ZN(n7368) );
  OR2_X1 U7528 ( .A1(n5940), .A2(n7368), .ZN(n5904) );
  INV_X1 U7529 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5902) );
  OR2_X1 U7530 ( .A1(n5835), .A2(n5902), .ZN(n5903) );
  OR2_X1 U7531 ( .A1(n7373), .A2(n7127), .ZN(n8945) );
  NAND2_X1 U7532 ( .A1(n7373), .A2(n7127), .ZN(n8928) );
  NAND2_X1 U7533 ( .A1(n8945), .A2(n8928), .ZN(n8851) );
  INV_X1 U7534 ( .A(n7127), .ZN(n9066) );
  NAND2_X1 U7535 ( .A1(n6342), .A2(n5855), .ZN(n5911) );
  OAI21_X1 U7536 ( .B1(n5908), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7537 ( .A(n5909), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9531) );
  AOI22_X1 U7538 ( .A1(n6003), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6002), .B2(
        n9531), .ZN(n5910) );
  NAND2_X1 U7539 ( .A1(n6293), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5918) );
  INV_X1 U7540 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7157) );
  OR2_X1 U7541 ( .A1(n6065), .A2(n7157), .ZN(n5917) );
  INV_X1 U7542 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6497) );
  OR2_X1 U7543 ( .A1(n6133), .A2(n6497), .ZN(n5916) );
  NAND2_X1 U7544 ( .A1(n5912), .A2(n10169), .ZN(n5913) );
  NAND2_X1 U7545 ( .A1(n5914), .A2(n5913), .ZN(n7240) );
  OR2_X1 U7546 ( .A1(n5940), .A2(n7240), .ZN(n5915) );
  OR2_X1 U7547 ( .A1(n7229), .A2(n7227), .ZN(n8929) );
  NAND2_X1 U7548 ( .A1(n7229), .A2(n7227), .ZN(n8931) );
  NAND2_X1 U7549 ( .A1(n8929), .A2(n8931), .ZN(n8849) );
  INV_X1 U7550 ( .A(n7227), .ZN(n9065) );
  OR2_X1 U7551 ( .A1(n7363), .A2(n7276), .ZN(n8933) );
  NAND2_X1 U7552 ( .A1(n7363), .A2(n7276), .ZN(n8951) );
  NAND2_X1 U7553 ( .A1(n8933), .A2(n8951), .ZN(n8867) );
  OAI21_X1 U7554 ( .B1(n9064), .B2(n7363), .A(n7164), .ZN(n7257) );
  NAND2_X1 U7555 ( .A1(n6582), .A2(n5855), .ZN(n5922) );
  NAND2_X1 U7556 ( .A1(n5919), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7557 ( .A(n5920), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U7558 ( .A1(n6003), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6002), .B2(
        n9553), .ZN(n5921) );
  NAND2_X1 U7559 ( .A1(n5804), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5930) );
  INV_X1 U7560 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5923) );
  OR2_X1 U7561 ( .A1(n6065), .A2(n5923), .ZN(n5929) );
  OR2_X1 U7562 ( .A1(n5924), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7563 ( .A1(n5937), .A2(n5925), .ZN(n7264) );
  OR2_X1 U7564 ( .A1(n5940), .A2(n7264), .ZN(n5928) );
  INV_X1 U7565 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7566 ( .A1(n5835), .A2(n5926), .ZN(n5927) );
  NAND2_X1 U7567 ( .A1(n7382), .A2(n7490), .ZN(n8955) );
  NAND2_X1 U7568 ( .A1(n8952), .A2(n8955), .ZN(n7258) );
  INV_X1 U7569 ( .A(n7490), .ZN(n9063) );
  NAND2_X1 U7570 ( .A1(n6611), .A2(n5855), .ZN(n5934) );
  XNOR2_X1 U7571 ( .A(n5932), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9566) );
  AOI22_X1 U7572 ( .A1(n6003), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6002), .B2(
        n9566), .ZN(n5933) );
  INV_X1 U7573 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7495) );
  OR2_X1 U7574 ( .A1(n6065), .A2(n7495), .ZN(n5944) );
  INV_X1 U7575 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7576 ( .A1(n6133), .A2(n5935), .ZN(n5943) );
  NAND2_X1 U7577 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7578 ( .A1(n5939), .A2(n5938), .ZN(n7550) );
  OR2_X1 U7579 ( .A1(n5940), .A2(n7550), .ZN(n5942) );
  NAND2_X1 U7580 ( .A1(n6293), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5941) );
  NAND4_X1 U7581 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n9062)
         );
  NAND2_X1 U7582 ( .A1(n9410), .A2(n9062), .ZN(n5945) );
  INV_X1 U7583 ( .A(n9410), .ZN(n7530) );
  INV_X1 U7584 ( .A(n9062), .ZN(n7529) );
  NAND2_X1 U7585 ( .A1(n6807), .A2(n5855), .ZN(n5962) );
  NOR2_X1 U7586 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5950) );
  NAND4_X1 U7587 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n5957)
         );
  INV_X1 U7588 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5953) );
  INV_X1 U7589 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5952) );
  NAND4_X1 U7590 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n5956)
         );
  NOR2_X1 U7591 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U7592 ( .A1(n5959), .A2(n5958), .ZN(n5969) );
  NAND2_X1 U7593 ( .A1(n5969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5960) );
  XNOR2_X1 U7594 ( .A(n5960), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U7595 ( .A1(n6003), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6002), .B2(
        n9599), .ZN(n5961) );
  NAND2_X1 U7596 ( .A1(n7713), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5968) );
  INV_X1 U7597 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10076) );
  OR2_X1 U7598 ( .A1(n5835), .A2(n10076), .ZN(n5967) );
  NOR2_X1 U7599 ( .A1(n5963), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5964) );
  OR2_X1 U7600 ( .A1(n5976), .A2(n5964), .ZN(n8724) );
  OR2_X1 U7601 ( .A1(n5940), .A2(n8724), .ZN(n5966) );
  INV_X1 U7602 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7189) );
  OR2_X1 U7603 ( .A1(n6133), .A2(n7189), .ZN(n5965) );
  OR2_X1 U7604 ( .A1(n8726), .A2(n8570), .ZN(n8962) );
  NAND2_X1 U7605 ( .A1(n8726), .A2(n8570), .ZN(n8963) );
  NAND2_X1 U7606 ( .A1(n8962), .A2(n8963), .ZN(n8872) );
  NAND2_X1 U7607 ( .A1(n6878), .A2(n5855), .ZN(n5974) );
  INV_X1 U7608 ( .A(n5969), .ZN(n5971) );
  INV_X1 U7609 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7610 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7611 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7612 ( .A(n5985), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9147) );
  AOI22_X1 U7613 ( .A1(n6003), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6002), .B2(
        n9147), .ZN(n5973) );
  INV_X1 U7614 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7615 ( .A1(n6065), .A2(n5975), .ZN(n5981) );
  OR2_X1 U7616 ( .A1(n5976), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7617 ( .A1(n5990), .A2(n5977), .ZN(n7589) );
  OR2_X1 U7618 ( .A1(n5940), .A2(n7589), .ZN(n5980) );
  INV_X1 U7619 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10077) );
  OR2_X1 U7620 ( .A1(n6133), .A2(n10077), .ZN(n5979) );
  NAND2_X1 U7621 ( .A1(n6293), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7622 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n9059)
         );
  NAND2_X1 U7623 ( .A1(n8575), .A2(n9059), .ZN(n5982) );
  INV_X1 U7624 ( .A(n9059), .ZN(n6121) );
  NAND2_X1 U7625 ( .A1(n8739), .A2(n6121), .ZN(n5983) );
  NAND2_X1 U7626 ( .A1(n6923), .A2(n5855), .ZN(n5988) );
  NAND2_X1 U7627 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7628 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7629 ( .A(n5998), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9613) );
  AOI22_X1 U7630 ( .A1(n6003), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6002), .B2(
        n9613), .ZN(n5987) );
  NAND2_X1 U7631 ( .A1(n7713), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7632 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  NAND2_X1 U7633 ( .A1(n6007), .A2(n5991), .ZN(n9340) );
  OR2_X1 U7634 ( .A1(n5940), .A2(n9340), .ZN(n5994) );
  NAND2_X1 U7635 ( .A1(n5804), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7636 ( .A1(n6293), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5992) );
  NAND4_X1 U7637 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9058)
         );
  INV_X1 U7638 ( .A(n9459), .ZN(n9344) );
  INV_X1 U7639 ( .A(n9058), .ZN(n6123) );
  OAI22_X2 U7640 ( .A1(n9335), .A2(n5996), .B1(n9344), .B2(n6123), .ZN(n9309)
         );
  NAND2_X1 U7641 ( .A1(n7061), .A2(n5855), .ZN(n6005) );
  NAND2_X1 U7642 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  AOI22_X1 U7643 ( .A1(n6003), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6002), .B2(
        n9156), .ZN(n6004) );
  NAND2_X1 U7644 ( .A1(n5804), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6012) );
  INV_X1 U7645 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7646 ( .A1(n6065), .A2(n6006), .ZN(n6011) );
  NAND2_X1 U7647 ( .A1(n6007), .A2(n10167), .ZN(n6008) );
  AND2_X1 U7648 ( .A1(n6017), .A2(n6008), .ZN(n9320) );
  NAND2_X1 U7649 ( .A1(n6044), .A2(n9320), .ZN(n6010) );
  NAND2_X1 U7650 ( .A1(n6293), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6009) );
  NAND4_X1 U7651 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8785)
         );
  INV_X1 U7652 ( .A(n9399), .ZN(n9325) );
  INV_X1 U7653 ( .A(n8785), .ZN(n6124) );
  OAI22_X2 U7654 ( .A1(n6014), .A2(n6013), .B1(n9325), .B2(n6124), .ZN(n9293)
         );
  NAND2_X1 U7655 ( .A1(n7178), .A2(n5855), .ZN(n6016) );
  OR2_X1 U7656 ( .A1(n7682), .A2(n7177), .ZN(n6015) );
  INV_X1 U7657 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10126) );
  AND2_X1 U7658 ( .A1(n6017), .A2(n8764), .ZN(n6018) );
  NOR2_X1 U7659 ( .A1(n6019), .A2(n6018), .ZN(n9302) );
  NAND2_X1 U7660 ( .A1(n9302), .A2(n6044), .ZN(n6021) );
  AOI22_X1 U7661 ( .A1(n7713), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n6293), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6020) );
  OAI211_X1 U7662 ( .C1(n6133), .C2(n10126), .A(n6021), .B(n6020), .ZN(n9057)
         );
  INV_X1 U7663 ( .A(n9057), .ZN(n8591) );
  AOI21_X2 U7664 ( .B1(n6023), .B2(n6022), .A(n5005), .ZN(n9278) );
  NAND2_X1 U7665 ( .A1(n10047), .A2(n5855), .ZN(n6026) );
  OR2_X1 U7666 ( .A1(n7682), .A2(n6024), .ZN(n6025) );
  INV_X1 U7667 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U7668 ( .A1(n6027), .A2(n8774), .ZN(n6028) );
  NAND2_X1 U7669 ( .A1(n6033), .A2(n6028), .ZN(n9270) );
  AOI22_X1 U7670 ( .A1(n5804), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n7713), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7671 ( .A1(n6293), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6029) );
  OAI211_X1 U7672 ( .C1(n9270), .C2(n5940), .A(n6030), .B(n6029), .ZN(n9055)
         );
  NAND2_X1 U7673 ( .A1(n9443), .A2(n9055), .ZN(n8810) );
  INV_X1 U7674 ( .A(n9055), .ZN(n8668) );
  NAND2_X1 U7675 ( .A1(n9269), .A2(n8668), .ZN(n8815) );
  NAND2_X1 U7676 ( .A1(n8810), .A2(n8815), .ZN(n9264) );
  NAND2_X1 U7677 ( .A1(n7524), .A2(n5855), .ZN(n6032) );
  OR2_X1 U7678 ( .A1(n7682), .A2(n7526), .ZN(n6031) );
  AND2_X1 U7679 ( .A1(n6033), .A2(n10052), .ZN(n6034) );
  OR2_X1 U7680 ( .A1(n6034), .A2(n6042), .ZN(n9255) );
  INV_X1 U7681 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U7682 ( .A1(n6293), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7683 ( .A1(n7713), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7684 ( .C1(n6133), .C2(n9380), .A(n6036), .B(n6035), .ZN(n6037)
         );
  INV_X1 U7685 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7686 ( .A1(n9379), .A2(n9054), .ZN(n6039) );
  NAND2_X1 U7687 ( .A1(n7599), .A2(n5855), .ZN(n6041) );
  OR2_X1 U7688 ( .A1(n7682), .A2(n7600), .ZN(n6040) );
  NAND2_X1 U7689 ( .A1(n6042), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6053) );
  OR2_X1 U7690 ( .A1(n6042), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6043) );
  AND2_X1 U7691 ( .A1(n6053), .A2(n6043), .ZN(n9239) );
  NAND2_X1 U7692 ( .A1(n9239), .A2(n6044), .ZN(n6049) );
  INV_X1 U7693 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U7694 ( .A1(n6293), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7695 ( .A1(n7713), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6045) );
  OAI211_X1 U7696 ( .C1(n6133), .C2(n9374), .A(n6046), .B(n6045), .ZN(n6047)
         );
  INV_X1 U7697 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7698 ( .A1(n9242), .A2(n8713), .ZN(n6050) );
  NAND2_X1 U7699 ( .A1(n9432), .A2(n9053), .ZN(n9218) );
  NAND2_X1 U7700 ( .A1(n7614), .A2(n5855), .ZN(n6052) );
  OR2_X1 U7701 ( .A1(n7682), .A2(n7615), .ZN(n6051) );
  AND2_X2 U7702 ( .A1(n6052), .A2(n6051), .ZN(n9428) );
  INV_X1 U7703 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U7704 ( .A1(n6053), .A2(n10093), .ZN(n6055) );
  INV_X1 U7705 ( .A(n6066), .ZN(n6054) );
  NAND2_X1 U7706 ( .A1(n6055), .A2(n6054), .ZN(n9223) );
  OR2_X1 U7707 ( .A1(n9223), .A2(n5940), .ZN(n6060) );
  INV_X1 U7708 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U7709 ( .A1(n6293), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7710 ( .A1(n5804), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6056) );
  OAI211_X1 U7711 ( .C1(n6065), .C2(n9222), .A(n6057), .B(n6056), .ZN(n6058)
         );
  INV_X1 U7712 ( .A(n6058), .ZN(n6059) );
  AND2_X1 U7713 ( .A1(n9218), .A2(n5011), .ZN(n6061) );
  NAND2_X1 U7714 ( .A1(n9428), .A2(n8801), .ZN(n9196) );
  NAND2_X1 U7715 ( .A1(n7611), .A2(n5855), .ZN(n6063) );
  OR2_X1 U7716 ( .A1(n7682), .A2(n7612), .ZN(n6062) );
  INV_X1 U7717 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7718 ( .A1(n6065), .A2(n6064), .ZN(n6070) );
  NAND2_X1 U7719 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6066), .ZN(n6077) );
  OAI21_X1 U7720 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6066), .A(n6077), .ZN(
        n9201) );
  OR2_X1 U7721 ( .A1(n5940), .A2(n9201), .ZN(n6069) );
  NAND2_X1 U7722 ( .A1(n6293), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7723 ( .A1(n5804), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6067) );
  NAND4_X1 U7724 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n9051)
         );
  OR2_X1 U7725 ( .A1(n9362), .A2(n9051), .ZN(n6071) );
  AND2_X1 U7726 ( .A1(n9196), .A2(n6071), .ZN(n6072) );
  NAND2_X1 U7727 ( .A1(n7818), .A2(n5855), .ZN(n6075) );
  OR2_X1 U7728 ( .A1(n7682), .A2(n6073), .ZN(n6074) );
  NAND2_X1 U7729 ( .A1(n7713), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6082) );
  INV_X1 U7730 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9422) );
  OR2_X1 U7731 ( .A1(n5835), .A2(n9422), .ZN(n6081) );
  INV_X1 U7732 ( .A(n6077), .ZN(n6076) );
  NAND2_X1 U7733 ( .A1(n6076), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6088) );
  INV_X1 U7734 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U7735 ( .A1(n6077), .A2(n8658), .ZN(n6078) );
  NAND2_X1 U7736 ( .A1(n6088), .A2(n6078), .ZN(n9189) );
  OR2_X1 U7737 ( .A1(n5940), .A2(n9189), .ZN(n6080) );
  INV_X1 U7738 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9359) );
  OR2_X1 U7739 ( .A1(n6133), .A2(n9359), .ZN(n6079) );
  OR2_X1 U7740 ( .A1(n9188), .A2(n8799), .ZN(n9009) );
  NAND2_X1 U7741 ( .A1(n9188), .A2(n8799), .ZN(n8808) );
  NAND2_X1 U7742 ( .A1(n8053), .A2(n5855), .ZN(n6084) );
  INV_X1 U7743 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U7744 ( .A1(n7713), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6094) );
  INV_X1 U7745 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7746 ( .A1(n5835), .A2(n6085), .ZN(n6093) );
  INV_X1 U7747 ( .A(n6088), .ZN(n6086) );
  NAND2_X1 U7748 ( .A1(n6086), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9170) );
  INV_X1 U7749 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7750 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  NAND2_X1 U7751 ( .A1(n9170), .A2(n6089), .ZN(n8690) );
  OR2_X1 U7752 ( .A1(n5940), .A2(n8690), .ZN(n6092) );
  INV_X1 U7753 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6090) );
  OR2_X1 U7754 ( .A1(n6133), .A2(n6090), .ZN(n6091) );
  NAND2_X1 U7755 ( .A1(n8692), .A2(n8684), .ZN(n8809) );
  INV_X1 U7756 ( .A(n6143), .ZN(n6098) );
  INV_X1 U7757 ( .A(n8900), .ZN(n7316) );
  INV_X1 U7758 ( .A(n6409), .ZN(n7317) );
  NAND2_X1 U7759 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7760 ( .A1(n4431), .A2(n10044), .ZN(n6358) );
  NAND2_X1 U7761 ( .A1(n6350), .A2(n6358), .ZN(n6104) );
  NAND3_X1 U7762 ( .A1(n7316), .A2(n7317), .A3(n6104), .ZN(n7069) );
  AND2_X1 U7763 ( .A1(n9156), .A2(n6105), .ZN(n9020) );
  NAND2_X1 U7764 ( .A1(n9020), .A2(n8885), .ZN(n9414) );
  INV_X1 U7765 ( .A(n6438), .ZN(n8853) );
  INV_X1 U7766 ( .A(n7324), .ZN(n6727) );
  NOR2_X1 U7767 ( .A1(n6723), .A2(n6727), .ZN(n6725) );
  NAND2_X1 U7768 ( .A1(n5802), .A2(n6440), .ZN(n6106) );
  NAND2_X1 U7769 ( .A1(n9073), .A2(n7090), .ZN(n8823) );
  AND4_X1 U7770 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6517)
         );
  NAND2_X1 U7771 ( .A1(n6517), .A2(n6469), .ZN(n6111) );
  NAND2_X1 U7772 ( .A1(n9072), .A2(n7074), .ZN(n8824) );
  NAND2_X1 U7773 ( .A1(n6515), .A2(n8824), .ZN(n6113) );
  INV_X1 U7774 ( .A(n9072), .ZN(n6568) );
  NAND2_X1 U7775 ( .A1(n6568), .A2(n6573), .ZN(n6112) );
  NAND2_X1 U7776 ( .A1(n6516), .A2(n8754), .ZN(n6114) );
  NAND2_X1 U7777 ( .A1(n8923), .A2(n6893), .ZN(n8919) );
  AND2_X1 U7778 ( .A1(n8919), .A2(n8920), .ZN(n7337) );
  NAND2_X1 U7779 ( .A1(n7337), .A2(n8926), .ZN(n6115) );
  NAND2_X1 U7780 ( .A1(n6115), .A2(n8944), .ZN(n8850) );
  AND2_X1 U7781 ( .A1(n8920), .A2(n6116), .ZN(n8925) );
  NAND2_X1 U7782 ( .A1(n8925), .A2(n8926), .ZN(n8862) );
  INV_X1 U7783 ( .A(n8910), .ZN(n6117) );
  NOR2_X1 U7784 ( .A1(n8862), .A2(n6117), .ZN(n6118) );
  INV_X1 U7785 ( .A(n8955), .ZN(n6119) );
  OR2_X1 U7786 ( .A1(n9410), .A2(n7529), .ZN(n8958) );
  NAND2_X1 U7787 ( .A1(n9410), .A2(n7529), .ZN(n8832) );
  NAND2_X1 U7788 ( .A1(n8958), .A2(n8832), .ZN(n8937) );
  NAND2_X1 U7789 ( .A1(n7541), .A2(n7491), .ZN(n8960) );
  INV_X1 U7790 ( .A(n8957), .ZN(n8941) );
  NOR2_X1 U7791 ( .A1(n8872), .A2(n8941), .ZN(n6120) );
  NAND2_X1 U7792 ( .A1(n7555), .A2(n6120), .ZN(n7581) );
  OR2_X1 U7793 ( .A1(n8575), .A2(n6121), .ZN(n8969) );
  NAND2_X1 U7794 ( .A1(n8575), .A2(n6121), .ZN(n8819) );
  NAND2_X1 U7795 ( .A1(n8969), .A2(n8819), .ZN(n7582) );
  INV_X1 U7796 ( .A(n8963), .ZN(n8835) );
  NOR2_X1 U7797 ( .A1(n7582), .A2(n8835), .ZN(n6122) );
  OR2_X1 U7798 ( .A1(n9459), .A2(n6123), .ZN(n9310) );
  NAND2_X1 U7799 ( .A1(n9459), .A2(n6123), .ZN(n8970) );
  OR2_X1 U7800 ( .A1(n9399), .A2(n6124), .ZN(n8977) );
  AND2_X1 U7801 ( .A1(n8977), .A2(n9310), .ZN(n8965) );
  NAND2_X1 U7802 ( .A1(n9399), .A2(n6124), .ZN(n8971) );
  OR2_X1 U7803 ( .A1(n9450), .A2(n8591), .ZN(n8978) );
  NAND2_X1 U7804 ( .A1(n9450), .A2(n8591), .ZN(n8966) );
  NAND2_X1 U7805 ( .A1(n8978), .A2(n8966), .ZN(n9294) );
  NAND2_X1 U7806 ( .A1(n9298), .A2(n8978), .ZN(n9280) );
  XNOR2_X1 U7807 ( .A(n9390), .B(n8814), .ZN(n9277) );
  NAND2_X1 U7808 ( .A1(n9390), .A2(n8814), .ZN(n8987) );
  OAI21_X1 U7809 ( .B1(n9280), .B2(n9277), .A(n8987), .ZN(n9265) );
  INV_X1 U7810 ( .A(n9264), .ZN(n9262) );
  NAND2_X1 U7811 ( .A1(n9265), .A2(n9262), .ZN(n6125) );
  NAND2_X1 U7812 ( .A1(n6125), .A2(n8815), .ZN(n9247) );
  NAND2_X1 U7813 ( .A1(n9259), .A2(n9054), .ZN(n8993) );
  INV_X1 U7814 ( .A(n9054), .ZN(n6126) );
  NAND2_X1 U7815 ( .A1(n9379), .A2(n6126), .ZN(n9234) );
  NAND2_X1 U7816 ( .A1(n9432), .A2(n8713), .ZN(n8998) );
  NAND2_X1 U7817 ( .A1(n8997), .A2(n8998), .ZN(n9230) );
  INV_X1 U7818 ( .A(n9234), .ZN(n6127) );
  INV_X1 U7819 ( .A(n9428), .ZN(n9227) );
  NAND2_X1 U7820 ( .A1(n9227), .A2(n8801), .ZN(n9000) );
  OR2_X1 U7821 ( .A1(n9362), .A2(n8712), .ZN(n9002) );
  NAND2_X1 U7822 ( .A1(n9362), .A2(n8712), .ZN(n9003) );
  NAND2_X1 U7823 ( .A1(n9002), .A2(n9003), .ZN(n9199) );
  INV_X1 U7824 ( .A(n9199), .ZN(n6129) );
  AND2_X1 U7825 ( .A1(n9205), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U7826 ( .A1(n9156), .A2(n10044), .ZN(n6132) );
  INV_X1 U7827 ( .A(n8885), .ZN(n8907) );
  NAND2_X1 U7828 ( .A1(n8822), .A2(n8907), .ZN(n6131) );
  NAND2_X1 U7829 ( .A1(n7713), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6137) );
  INV_X1 U7830 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7791) );
  OR2_X1 U7831 ( .A1(n6133), .A2(n7791), .ZN(n6136) );
  OR2_X1 U7832 ( .A1(n5940), .A2(n9170), .ZN(n6135) );
  INV_X1 U7833 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7720) );
  OR2_X1 U7834 ( .A1(n5835), .A2(n7720), .ZN(n6134) );
  OAI22_X1 U7835 ( .A1(n7706), .A2(n8798), .B1(n8799), .B2(n8800), .ZN(n8688)
         );
  NAND2_X1 U7836 ( .A1(n6520), .A2(n7074), .ZN(n6519) );
  INV_X1 U7837 ( .A(n7373), .ZN(n7128) );
  INV_X1 U7838 ( .A(n7229), .ZN(n7246) );
  NAND2_X1 U7839 ( .A1(n6982), .A2(n7246), .ZN(n7031) );
  OR2_X1 U7840 ( .A1(n7263), .A2(n7382), .ZN(n7494) );
  NOR2_X2 U7841 ( .A1(n7494), .A2(n9410), .ZN(n7506) );
  INV_X1 U7842 ( .A(n8726), .ZN(n7562) );
  NAND2_X1 U7843 ( .A1(n9428), .A2(n9238), .ZN(n9224) );
  NOR2_X2 U7844 ( .A1(n9224), .A2(n9362), .ZN(n9186) );
  INV_X1 U7845 ( .A(n6140), .ZN(n9187) );
  OR2_X2 U7846 ( .A1(n8692), .A2(n6140), .ZN(n7708) );
  OAI211_X1 U7847 ( .C1(n7705), .C2(n9187), .A(n9342), .B(n7708), .ZN(n8058)
         );
  NAND2_X1 U7848 ( .A1(n6143), .A2(n6142), .ZN(n6149) );
  NAND2_X1 U7849 ( .A1(n6146), .A2(n6145), .ZN(n6148) );
  NAND2_X1 U7850 ( .A1(n6149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U7851 ( .A1(n7616), .A2(n7601), .ZN(n6151) );
  NAND2_X1 U7852 ( .A1(n6152), .A2(n4591), .ZN(n6153) );
  NAND2_X1 U7853 ( .A1(n6153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6154) );
  AND2_X1 U7854 ( .A1(n9036), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7855 ( .A1(n8900), .A2(n6350), .ZN(n6407) );
  NAND2_X1 U7856 ( .A1(n7616), .A2(P1_B_REG_SCAN_IN), .ZN(n6157) );
  MUX2_X1 U7857 ( .A(n6157), .B(P1_B_REG_SCAN_IN), .S(n6170), .Z(n6158) );
  INV_X1 U7858 ( .A(n7616), .ZN(n6159) );
  OAI22_X1 U7859 ( .A1(n6171), .A2(P1_D_REG_1__SCAN_IN), .B1(n6156), .B2(n6159), .ZN(n6403) );
  NOR4_X1 U7860 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6163) );
  NOR4_X1 U7861 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6162) );
  NOR4_X1 U7862 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6161) );
  NOR4_X1 U7863 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6160) );
  NAND4_X1 U7864 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n6169)
         );
  NOR2_X1 U7865 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .ZN(
        n6167) );
  NOR4_X1 U7866 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6166) );
  NOR4_X1 U7867 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6165) );
  NOR4_X1 U7868 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7869 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n6168)
         );
  OAI21_X1 U7870 ( .B1(n6169), .B2(n6168), .A(n9636), .ZN(n6404) );
  NAND2_X1 U7871 ( .A1(n9342), .A2(n9156), .ZN(n6410) );
  NAND4_X1 U7872 ( .A1(n7065), .A2(n6403), .A3(n6404), .A4(n6410), .ZN(n6176)
         );
  OR2_X1 U7873 ( .A1(n6177), .A2(n9676), .ZN(n6173) );
  NAND2_X1 U7874 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  NAND2_X1 U7875 ( .A1(n6174), .A2(n5000), .ZN(P1_U3550) );
  INV_X1 U7876 ( .A(n7064), .ZN(n6175) );
  INV_X1 U7877 ( .A(n9036), .ZN(n6575) );
  OR2_X2 U7878 ( .A1(n6261), .A2(P1_U3086), .ZN(n6670) );
  NAND2_X1 U7879 ( .A1(n6270), .A2(n8007), .ZN(n6178) );
  NAND2_X1 U7880 ( .A1(n6178), .A2(n6201), .ZN(n6272) );
  NAND2_X1 U7881 ( .A1(n6272), .A2(n5080), .ZN(n6179) );
  NAND2_X1 U7882 ( .A1(n6179), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7883 ( .A(n6250), .ZN(n6180) );
  NAND3_X1 U7884 ( .A1(n6181), .A2(n7837), .A3(n6248), .ZN(n6182) );
  XNOR2_X1 U7885 ( .A(n7735), .B(n9899), .ZN(n6941) );
  XNOR2_X1 U7886 ( .A(n6941), .B(n8196), .ZN(n6942) );
  INV_X1 U7887 ( .A(n8197), .ZN(n6752) );
  XNOR2_X1 U7888 ( .A(n7735), .B(n9896), .ZN(n6190) );
  INV_X1 U7889 ( .A(n6190), .ZN(n6191) );
  INV_X1 U7890 ( .A(n9868), .ZN(n6604) );
  XNOR2_X1 U7891 ( .A(n7735), .B(n9889), .ZN(n6189) );
  XNOR2_X1 U7892 ( .A(n6187), .B(n9867), .ZN(n6595) );
  XNOR2_X1 U7893 ( .A(n7735), .B(n6608), .ZN(n6188) );
  XNOR2_X1 U7894 ( .A(n6188), .B(n8198), .ZN(n6602) );
  INV_X1 U7895 ( .A(n8198), .ZN(n6596) );
  AOI22_X1 U7896 ( .A1(n6603), .A2(n6602), .B1(n6596), .B2(n6188), .ZN(n6560)
         );
  XNOR2_X1 U7897 ( .A(n6189), .B(n9868), .ZN(n6559) );
  XNOR2_X1 U7898 ( .A(n6190), .B(n8197), .ZN(n6624) );
  XOR2_X1 U7899 ( .A(n6942), .B(n6943), .Z(n6198) );
  NAND2_X1 U7900 ( .A1(n6209), .A2(n6192), .ZN(n6193) );
  NAND2_X1 U7901 ( .A1(n6193), .A2(n6194), .ZN(n6197) );
  INV_X1 U7902 ( .A(n6194), .ZN(n6195) );
  NAND2_X1 U7903 ( .A1(n6215), .A2(n6195), .ZN(n6203) );
  AND2_X1 U7904 ( .A1(n6203), .A2(n6244), .ZN(n6196) );
  NOR2_X1 U7905 ( .A1(n6198), .A2(n8177), .ZN(n6223) );
  INV_X1 U7906 ( .A(n6199), .ZN(n6200) );
  OR2_X1 U7907 ( .A1(n6209), .A2(n6200), .ZN(n6205) );
  INV_X1 U7908 ( .A(n6201), .ZN(n7522) );
  NOR2_X1 U7909 ( .A1(n6202), .A2(n7522), .ZN(n6204) );
  NAND4_X1 U7910 ( .A1(n6205), .A2(n6204), .A3(n6270), .A4(n6203), .ZN(n6206)
         );
  NAND2_X1 U7911 ( .A1(n6206), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6208) );
  INV_X1 U7912 ( .A(n6214), .ZN(n8028) );
  NAND2_X1 U7913 ( .A1(n6215), .A2(n8028), .ZN(n6207) );
  NOR2_X1 U7914 ( .A1(n8174), .A2(n6756), .ZN(n6222) );
  NAND3_X1 U7915 ( .A1(n6209), .A2(n6244), .A3(n9943), .ZN(n6213) );
  INV_X1 U7916 ( .A(n6210), .ZN(n6211) );
  AND2_X1 U7917 ( .A1(n8182), .A2(n6758), .ZN(n6221) );
  NOR2_X1 U7918 ( .A1(n6215), .A2(n6214), .ZN(n6218) );
  NAND2_X1 U7919 ( .A1(n6218), .A2(n6216), .ZN(n8143) );
  NAND2_X1 U7920 ( .A1(n6218), .A2(n6217), .ZN(n8170) );
  OR2_X1 U7921 ( .A1(n8170), .A2(n4733), .ZN(n6219) );
  NAND2_X1 U7922 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9705) );
  OAI211_X1 U7923 ( .C1(n8143), .C2(n6752), .A(n6219), .B(n9705), .ZN(n6220)
         );
  OR4_X1 U7924 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(P2_U3167)
         );
  XNOR2_X1 U7925 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X2 U7926 ( .A(n8560), .ZN(n8555) );
  AND2_X1 U7927 ( .A1(n7671), .A2(P2_U3151), .ZN(n7521) );
  INV_X2 U7928 ( .A(n7521), .ZN(n8562) );
  OAI222_X1 U7929 ( .A1(n8555), .A2(n5049), .B1(n8562), .B2(n6229), .C1(
        P2_U3151), .C2(n6291), .ZN(P2_U3294) );
  OAI222_X1 U7930 ( .A1(n8555), .A2(n6225), .B1(n8562), .B2(n6234), .C1(
        P2_U3151), .C2(n6543), .ZN(P2_U3293) );
  OAI222_X1 U7931 ( .A1(n8555), .A2(n6226), .B1(n8562), .B2(n6230), .C1(
        P2_U3151), .C2(n6546), .ZN(P2_U3292) );
  OAI222_X1 U7932 ( .A1(n8555), .A2(n6227), .B1(n8562), .B2(n6232), .C1(
        P2_U3151), .C2(n6707), .ZN(P2_U3291) );
  INV_X1 U7933 ( .A(n10045), .ZN(n9478) );
  NAND2_X2 U7934 ( .A1(n6228), .A2(P1_U3086), .ZN(n9476) );
  OAI222_X1 U7935 ( .A1(n9478), .A2(n4925), .B1(n9476), .B2(n6229), .C1(
        P1_U3086), .C2(n6373), .ZN(P1_U3354) );
  OAI222_X1 U7936 ( .A1(n9478), .A2(n6231), .B1(n9476), .B2(n6230), .C1(
        P1_U3086), .C2(n6393), .ZN(P1_U3352) );
  OAI222_X1 U7937 ( .A1(n9478), .A2(n6233), .B1(n9476), .B2(n6232), .C1(
        P1_U3086), .C2(n6389), .ZN(P1_U3351) );
  OAI222_X1 U7938 ( .A1(n9478), .A2(n6235), .B1(n9476), .B2(n6234), .C1(
        P1_U3086), .C2(n6372), .ZN(P1_U3353) );
  OAI222_X1 U7939 ( .A1(n9478), .A2(n6236), .B1(n9476), .B2(n6237), .C1(
        P1_U3086), .C2(n9099), .ZN(P1_U3350) );
  OAI222_X1 U7940 ( .A1(n8555), .A2(n6238), .B1(n8562), .B2(n6237), .C1(
        P2_U3151), .C2(n9707), .ZN(P2_U3290) );
  INV_X1 U7941 ( .A(n6239), .ZN(n6241) );
  AOI22_X1 U7942 ( .A1(n7432), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8560), .ZN(n6240) );
  OAI21_X1 U7943 ( .B1(n6241), .B2(n8562), .A(n6240), .ZN(P2_U3289) );
  OAI222_X1 U7944 ( .A1(n9478), .A2(n6242), .B1(n9476), .B2(n6241), .C1(
        P1_U3086), .C2(n9113), .ZN(P1_U3349) );
  INV_X1 U7945 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6247) );
  INV_X1 U7946 ( .A(n6245), .ZN(n6246) );
  AOI22_X1 U7947 ( .A1(n6265), .A2(n6247), .B1(n6250), .B2(n6246), .ZN(
        P2_U3377) );
  INV_X1 U7948 ( .A(n6248), .ZN(n6249) );
  AOI22_X1 U7949 ( .A1(n6265), .A2(n5681), .B1(n6250), .B2(n6249), .ZN(
        P2_U3376) );
  INV_X1 U7950 ( .A(n6251), .ZN(n6253) );
  AOI22_X1 U7951 ( .A1(n9498), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10045), .ZN(n6252) );
  OAI21_X1 U7952 ( .B1(n6253), .B2(n9476), .A(n6252), .ZN(P1_U3348) );
  AND2_X1 U7953 ( .A1(n6265), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7954 ( .A1(n6265), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7955 ( .A1(n6265), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7956 ( .A1(n6265), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7957 ( .A1(n6265), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7958 ( .A1(n6265), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7959 ( .A1(n6265), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7960 ( .A1(n6265), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7961 ( .A1(n6265), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7962 ( .A1(n6265), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7963 ( .A1(n6265), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7964 ( .A1(n6265), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7965 ( .A1(n6265), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U7966 ( .A1(n6265), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7967 ( .A1(n6265), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7968 ( .A1(n6265), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7969 ( .A1(n6265), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7970 ( .A1(n6265), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7971 ( .A1(n6265), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7972 ( .A1(n6265), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7973 ( .A1(n6265), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  INV_X1 U7974 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6254) );
  OAI222_X1 U7975 ( .A1(n8555), .A2(n6254), .B1(n8562), .B2(n6253), .C1(
        P2_U3151), .C2(n7433), .ZN(P2_U3288) );
  INV_X1 U7976 ( .A(n6255), .ZN(n6267) );
  AOI22_X1 U7977 ( .A1(n9512), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10045), .ZN(n6256) );
  OAI21_X1 U7978 ( .B1(n6267), .B2(n9476), .A(n6256), .ZN(P1_U3347) );
  INV_X1 U7979 ( .A(n7819), .ZN(n9041) );
  INV_X1 U7980 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7315) );
  AOI21_X1 U7981 ( .B1(n9041), .B2(n7315), .A(n8054), .ZN(n6365) );
  OAI21_X1 U7982 ( .B1(n9041), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6365), .ZN(
        n6258) );
  XOR2_X1 U7983 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6258), .Z(n6264) );
  NAND2_X1 U7984 ( .A1(n8900), .A2(n9036), .ZN(n6259) );
  NAND2_X1 U7985 ( .A1(n7677), .A2(n6259), .ZN(n6262) );
  INV_X1 U7986 ( .A(n6261), .ZN(n6260) );
  OR3_X1 U7987 ( .A1(n6262), .A2(n6260), .A3(P1_U3086), .ZN(n6375) );
  AND3_X1 U7988 ( .A1(n6262), .A2(P1_STATE_REG_SCAN_IN), .A3(n6261), .ZN(n9518) );
  AOI22_X1 U7989 ( .A1(n9518), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6263) );
  OAI21_X1 U7990 ( .B1(n6264), .B2(n6375), .A(n6263), .ZN(P1_U3243) );
  INV_X1 U7991 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U7992 ( .A1(n6266), .A2(n10267), .ZN(P2_U3244) );
  INV_X1 U7993 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U7994 ( .A1(n6266), .A2(n10150), .ZN(P2_U3243) );
  INV_X1 U7995 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U7996 ( .A1(n6266), .A2(n10113), .ZN(P2_U3237) );
  INV_X1 U7997 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10088) );
  NOR2_X1 U7998 ( .A1(n6266), .A2(n10088), .ZN(P2_U3254) );
  INV_X1 U7999 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U8000 ( .A1(n6266), .A2(n10238), .ZN(P2_U3241) );
  INV_X1 U8001 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10121) );
  NOR2_X1 U8002 ( .A1(n6266), .A2(n10121), .ZN(P2_U3258) );
  INV_X1 U8003 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U8004 ( .A1(n6266), .A2(n10096), .ZN(P2_U3262) );
  INV_X1 U8005 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U8006 ( .A1(n6266), .A2(n10210), .ZN(P2_U3252) );
  INV_X1 U8007 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U8008 ( .A1(n6266), .A2(n10120), .ZN(P2_U3253) );
  INV_X1 U8009 ( .A(n9729), .ZN(n7428) );
  OAI222_X1 U8010 ( .A1(n8555), .A2(n10244), .B1(n8562), .B2(n6267), .C1(
        P2_U3151), .C2(n7428), .ZN(P2_U3287) );
  NOR2_X1 U8011 ( .A1(n9518), .A2(P1_U3973), .ZN(P1_U3085) );
  AND2_X1 U8012 ( .A1(n6272), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6268) );
  MUX2_X1 U8013 ( .A(P2_U3893), .B(n6268), .S(n5660), .Z(n6269) );
  NAND2_X1 U8014 ( .A1(n6269), .A2(n5080), .ZN(n9708) );
  INV_X1 U8015 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10246) );
  NOR2_X1 U8016 ( .A1(n6270), .A2(n7522), .ZN(n6271) );
  NOR2_X1 U8017 ( .A1(n5660), .A2(P2_U3151), .ZN(n8559) );
  NAND2_X1 U8018 ( .A1(n5053), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U8019 ( .A1(n6291), .A2(n6312), .ZN(n6277) );
  INV_X1 U8020 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U8021 ( .A1(n6274), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6275) );
  OR2_X1 U8022 ( .A1(n6275), .A2(n5053), .ZN(n6276) );
  NAND2_X1 U8023 ( .A1(n6277), .A2(n6276), .ZN(n6311) );
  XNOR2_X1 U8024 ( .A(n6311), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6278) );
  AOI22_X1 U8025 ( .A1(n9852), .A2(n6278), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n6285) );
  INV_X1 U8026 ( .A(n6279), .ZN(n6334) );
  INV_X1 U8027 ( .A(n9856), .ZN(n9718) );
  NOR2_X1 U8028 ( .A1(n10253), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U8029 ( .A1(n5053), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6316) );
  OAI21_X1 U8030 ( .B1(n6291), .B2(n6280), .A(n6316), .ZN(n6281) );
  OR2_X1 U8031 ( .A1(n6281), .A2(n5031), .ZN(n6317) );
  NAND2_X1 U8032 ( .A1(n6281), .A2(n5031), .ZN(n6282) );
  NAND2_X1 U8033 ( .A1(n6317), .A2(n6282), .ZN(n6283) );
  NAND2_X1 U8034 ( .A1(n9718), .A2(n6283), .ZN(n6284) );
  OAI211_X1 U8035 ( .C1(n10246), .C2(n9713), .A(n6285), .B(n6284), .ZN(n6286)
         );
  INV_X1 U8036 ( .A(n6286), .ZN(n6290) );
  MUX2_X1 U8037 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8213), .Z(n6326) );
  XNOR2_X1 U8038 ( .A(n6326), .B(n6329), .ZN(n6288) );
  INV_X1 U8039 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10253) );
  INV_X1 U8040 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6287) );
  MUX2_X1 U8041 ( .A(n10253), .B(n6287), .S(n8257), .Z(n6336) );
  NAND2_X1 U8042 ( .A1(n6336), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8043 ( .A1(n6288), .A2(n6335), .ZN(n6327) );
  NAND2_X1 U8044 ( .A1(P2_U3893), .A2(n5660), .ZN(n9692) );
  OAI211_X1 U8045 ( .C1(n6288), .C2(n6335), .A(n6327), .B(n9851), .ZN(n6289)
         );
  OAI211_X1 U8046 ( .C1(n9708), .C2(n6291), .A(n6290), .B(n6289), .ZN(P2_U3183) );
  MUX2_X1 U8047 ( .A(n6304), .B(n7305), .S(P2_U3893), .Z(n6292) );
  INV_X1 U8048 ( .A(n6292), .ZN(P2_U3500) );
  INV_X1 U8049 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U8050 ( .A1(n5804), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U8051 ( .A1(n7713), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U8052 ( .A1(n6293), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6294) );
  INV_X1 U8053 ( .A(n8896), .ZN(n9021) );
  NAND2_X1 U8054 ( .A1(n9021), .A2(P1_U3973), .ZN(n6297) );
  OAI21_X1 U8055 ( .B1(P1_U3973), .B2(n6298), .A(n6297), .ZN(P1_U3585) );
  INV_X1 U8056 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U8057 ( .A1(n6723), .A2(P1_U3973), .ZN(n6299) );
  OAI21_X1 U8058 ( .B1(P1_U3973), .B2(n6300), .A(n6299), .ZN(P1_U3554) );
  INV_X1 U8059 ( .A(n6301), .ZN(n6303) );
  INV_X1 U8060 ( .A(n9746), .ZN(n7436) );
  OAI222_X1 U8061 ( .A1(n8555), .A2(n6302), .B1(n8562), .B2(n6303), .C1(
        P2_U3151), .C2(n7436), .ZN(P2_U3286) );
  INV_X1 U8062 ( .A(n9136), .ZN(n6486) );
  OAI222_X1 U8063 ( .A1(n9478), .A2(n6304), .B1(n9476), .B2(n6303), .C1(
        P1_U3086), .C2(n6486), .ZN(P1_U3346) );
  INV_X1 U8064 ( .A(n6305), .ZN(n6308) );
  AOI22_X1 U8065 ( .A1(n9488), .A2(P1_STATE_REG_SCAN_IN), .B1(n10045), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U8066 ( .B1(n6308), .B2(n9476), .A(n6306), .ZN(P1_U3345) );
  INV_X1 U8067 ( .A(n7438), .ZN(n7632) );
  OAI222_X1 U8068 ( .A1(n8562), .A2(n6308), .B1(n7632), .B2(P2_U3151), .C1(
        n6307), .C2(n8555), .ZN(P2_U3285) );
  NAND2_X1 U8069 ( .A1(n8785), .A2(P1_U3973), .ZN(n6309) );
  OAI21_X1 U8070 ( .B1(n5418), .B2(P1_U3973), .A(n6309), .ZN(P1_U3573) );
  NAND2_X1 U8071 ( .A1(n6311), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U8072 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  OAI21_X1 U8073 ( .B1(n6315), .B2(n6314), .A(n6545), .ZN(n6325) );
  XNOR2_X1 U8074 ( .A(n6543), .B(n9878), .ZN(n6319) );
  NAND2_X1 U8075 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  NAND2_X1 U8076 ( .A1(n6319), .A2(n6318), .ZN(n6535) );
  OAI21_X1 U8077 ( .B1(n6319), .B2(n6318), .A(n6535), .ZN(n6320) );
  INV_X1 U8078 ( .A(n6320), .ZN(n6322) );
  OAI22_X1 U8079 ( .A1(n9856), .A2(n6322), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6321), .ZN(n6324) );
  INV_X1 U8080 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U8081 ( .A1(n9713), .A2(n10114), .ZN(n6323) );
  AOI211_X1 U8082 ( .C1(n9852), .C2(n6325), .A(n6324), .B(n6323), .ZN(n6333)
         );
  INV_X1 U8083 ( .A(n6326), .ZN(n6328) );
  OAI21_X1 U8084 ( .B1(n6329), .B2(n6328), .A(n6327), .ZN(n6331) );
  MUX2_X1 U8085 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8257), .Z(n6526) );
  XOR2_X1 U8086 ( .A(n6543), .B(n6526), .Z(n6330) );
  NAND2_X1 U8087 ( .A1(n6331), .A2(n6330), .ZN(n6527) );
  OAI211_X1 U8088 ( .C1(n6331), .C2(n6330), .A(n6527), .B(n9851), .ZN(n6332)
         );
  OAI211_X1 U8089 ( .C1(n9708), .C2(n6543), .A(n6333), .B(n6332), .ZN(P2_U3184) );
  INV_X1 U8090 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6341) );
  INV_X1 U8091 ( .A(n9708), .ZN(n9844) );
  NAND2_X1 U8092 ( .A1(n9844), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U8093 ( .A1(n6334), .A2(n9692), .ZN(n6338) );
  OAI21_X1 U8094 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6336), .A(n6335), .ZN(n6337) );
  AOI22_X1 U8095 ( .A1(n6338), .A2(n6337), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6339) );
  OAI211_X1 U8096 ( .C1(n9713), .C2(n6341), .A(n6340), .B(n6339), .ZN(P2_U3182) );
  INV_X1 U8097 ( .A(n6342), .ZN(n6344) );
  AOI22_X1 U8098 ( .A1(n9531), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10045), .ZN(n6343) );
  OAI21_X1 U8099 ( .B1(n6344), .B2(n9476), .A(n6343), .ZN(P1_U3344) );
  INV_X1 U8100 ( .A(n9761), .ZN(n7630) );
  OAI222_X1 U8101 ( .A1(n8555), .A2(n6345), .B1(n8562), .B2(n6344), .C1(
        P2_U3151), .C2(n7630), .ZN(P2_U3284) );
  INV_X1 U8102 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8103 ( .A1(n5632), .A2(n6654), .ZN(n7880) );
  NAND2_X1 U8104 ( .A1(n6185), .A2(n7880), .ZN(n6656) );
  OAI21_X1 U8105 ( .B1(n9938), .B2(n8433), .A(n6656), .ZN(n6346) );
  NAND2_X1 U8106 ( .A1(n9867), .A2(n9869), .ZN(n6657) );
  OAI211_X1 U8107 ( .C1(n9919), .C2(n6654), .A(n6346), .B(n6657), .ZN(n8480)
         );
  NAND2_X1 U8108 ( .A1(n8480), .A2(n9946), .ZN(n6347) );
  OAI21_X1 U8109 ( .B1(n6348), .B2(n9946), .A(n6347), .ZN(P2_U3390) );
  AND2_X1 U8110 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9076) );
  INV_X1 U8111 ( .A(n6360), .ZN(n6576) );
  NAND2_X1 U8112 ( .A1(n8822), .A2(n8885), .ZN(n6357) );
  OAI21_X1 U8113 ( .B1(n6350), .B2(n10044), .A(n7135), .ZN(n6351) );
  NAND2_X1 U8114 ( .A1(n6723), .A2(n8635), .ZN(n6355) );
  INV_X1 U8115 ( .A(n6357), .ZN(n6353) );
  INV_X2 U8116 ( .A(n6424), .ZN(n6773) );
  AND2_X1 U8117 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U8118 ( .A1(n6723), .A2(n6773), .ZN(n6362) );
  OAI21_X1 U8119 ( .B1(n8630), .B2(n6727), .A(n6362), .ZN(n6425) );
  XNOR2_X1 U8120 ( .A(n6426), .B(n6427), .ZN(n6416) );
  MUX2_X1 U8121 ( .A(n9076), .B(n6416), .S(n7819), .Z(n6363) );
  NAND2_X1 U8122 ( .A1(n6363), .A2(n6371), .ZN(n6364) );
  OAI211_X1 U8123 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6365), .A(n6364), .B(
        P1_U3973), .ZN(n6402) );
  XNOR2_X1 U8124 ( .A(n6372), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6370) );
  XNOR2_X1 U8125 ( .A(n6373), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U8126 ( .A1(n9077), .A2(n9076), .ZN(n9075) );
  INV_X1 U8127 ( .A(n6373), .ZN(n9078) );
  NAND2_X1 U8128 ( .A1(n9078), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8129 ( .A1(n9075), .A2(n6366), .ZN(n6369) );
  INV_X1 U8130 ( .A(n6375), .ZN(n6368) );
  NOR2_X1 U8131 ( .A1(n8054), .A2(n7819), .ZN(n6367) );
  NAND2_X1 U8132 ( .A1(n6368), .A2(n6367), .ZN(n9581) );
  INV_X1 U8133 ( .A(n9581), .ZN(n9605) );
  NAND2_X1 U8134 ( .A1(n6370), .A2(n6369), .ZN(n6385) );
  OAI211_X1 U8135 ( .C1(n6370), .C2(n6369), .A(n9605), .B(n6385), .ZN(n6381)
         );
  AOI22_X1 U8136 ( .A1(n9518), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6380) );
  NOR2_X2 U8137 ( .A1(n6375), .A2(n6371), .ZN(n9612) );
  INV_X1 U8138 ( .A(n6372), .ZN(n6390) );
  NAND2_X1 U8139 ( .A1(n9612), .A2(n6390), .ZN(n6379) );
  XNOR2_X1 U8140 ( .A(n6372), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6377) );
  XNOR2_X1 U8141 ( .A(n6373), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9081) );
  AND2_X1 U8142 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9080) );
  NAND2_X1 U8143 ( .A1(n9081), .A2(n9080), .ZN(n9079) );
  NAND2_X1 U8144 ( .A1(n9078), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8145 ( .A1(n9079), .A2(n6374), .ZN(n6376) );
  NOR2_X2 U8146 ( .A1(n6375), .A2(n9041), .ZN(n9597) );
  NAND2_X1 U8147 ( .A1(n6377), .A2(n6376), .ZN(n6392) );
  OAI211_X1 U8148 ( .C1(n6377), .C2(n6376), .A(n9597), .B(n6392), .ZN(n6378)
         );
  AND4_X1 U8149 ( .A1(n6381), .A2(n6380), .A3(n6379), .A4(n6378), .ZN(n6382)
         );
  NAND2_X1 U8150 ( .A1(n6402), .A2(n6382), .ZN(P1_U3245) );
  INV_X1 U8151 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6383) );
  MUX2_X1 U8152 ( .A(n6383), .B(P1_REG2_REG_4__SCAN_IN), .S(n6389), .Z(n6388)
         );
  INV_X1 U8153 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10152) );
  MUX2_X1 U8154 ( .A(n10152), .B(P1_REG2_REG_3__SCAN_IN), .S(n6393), .Z(n9095)
         );
  NAND2_X1 U8155 ( .A1(n6390), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8156 ( .A1(n6385), .A2(n6384), .ZN(n9094) );
  NAND2_X1 U8157 ( .A1(n9095), .A2(n9094), .ZN(n9093) );
  INV_X1 U8158 ( .A(n6393), .ZN(n9089) );
  NAND2_X1 U8159 ( .A1(n9089), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8160 ( .A1(n9093), .A2(n6386), .ZN(n6387) );
  NAND2_X1 U8161 ( .A1(n6387), .A2(n6388), .ZN(n6478) );
  OAI211_X1 U8162 ( .C1(n6388), .C2(n6387), .A(n9605), .B(n6478), .ZN(n6400)
         );
  AND2_X1 U8163 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8753) );
  AOI21_X1 U8164 ( .B1(n9518), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n8753), .ZN(
        n6399) );
  INV_X1 U8165 ( .A(n6389), .ZN(n6487) );
  NAND2_X1 U8166 ( .A1(n9612), .A2(n6487), .ZN(n6398) );
  INV_X1 U8167 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6512) );
  MUX2_X1 U8168 ( .A(n6512), .B(P1_REG1_REG_4__SCAN_IN), .S(n6389), .Z(n6396)
         );
  NAND2_X1 U8169 ( .A1(n6390), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U8170 ( .A1(n6392), .A2(n6391), .ZN(n9091) );
  XNOR2_X1 U8171 ( .A(n6393), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U8172 ( .A1(n9091), .A2(n9092), .ZN(n9090) );
  NAND2_X1 U8173 ( .A1(n9089), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8174 ( .A1(n9090), .A2(n6394), .ZN(n6395) );
  NAND2_X1 U8175 ( .A1(n6395), .A2(n6396), .ZN(n6489) );
  OAI211_X1 U8176 ( .C1(n6396), .C2(n6395), .A(n9597), .B(n6489), .ZN(n6397)
         );
  AND4_X1 U8177 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6401)
         );
  NAND2_X1 U8178 ( .A1(n6402), .A2(n6401), .ZN(P1_U3247) );
  INV_X1 U8179 ( .A(n6403), .ZN(n9466) );
  NAND2_X1 U8180 ( .A1(n9466), .A2(n6404), .ZN(n7067) );
  INV_X1 U8181 ( .A(n9667), .ZN(n9637) );
  OR2_X1 U8182 ( .A1(n7064), .A2(n9637), .ZN(n9665) );
  NOR2_X1 U8183 ( .A1(n9411), .A2(n8900), .ZN(n6405) );
  OR2_X1 U8184 ( .A1(n8885), .A2(P1_U3086), .ZN(n9034) );
  INV_X1 U8185 ( .A(n9034), .ZN(n6406) );
  INV_X1 U8186 ( .A(n9411), .ZN(n9669) );
  OAI22_X1 U8187 ( .A1(n7067), .A2(n7064), .B1(n6406), .B2(n9669), .ZN(n6408)
         );
  NAND2_X1 U8188 ( .A1(n6408), .A2(n6407), .ZN(n6577) );
  NOR2_X1 U8189 ( .A1(n6577), .A2(n9637), .ZN(n6474) );
  INV_X1 U8190 ( .A(n6474), .ZN(n6431) );
  AND2_X1 U8191 ( .A1(n6409), .A2(n8907), .ZN(n7073) );
  NAND2_X1 U8192 ( .A1(n6413), .A2(n7073), .ZN(n6412) );
  INV_X1 U8193 ( .A(n6350), .ZN(n9040) );
  NAND2_X1 U8194 ( .A1(n9074), .A2(n8784), .ZN(n7319) );
  OAI22_X1 U8195 ( .A1(n8807), .A2(n6727), .B1(n8775), .B2(n7319), .ZN(n6414)
         );
  AOI21_X1 U8196 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6431), .A(n6414), .ZN(
        n6415) );
  OAI21_X1 U8197 ( .B1(n6416), .B2(n8792), .A(n6415), .ZN(P1_U3232) );
  NOR2_X1 U8198 ( .A1(n8164), .A2(P2_U3151), .ZN(n6605) );
  INV_X1 U8199 ( .A(n8182), .ZN(n8167) );
  OAI22_X1 U8200 ( .A1(n8167), .A2(n6654), .B1(n5060), .B2(n8170), .ZN(n6417)
         );
  AOI21_X1 U8201 ( .B1(n8160), .B2(n6656), .A(n6417), .ZN(n6418) );
  OAI21_X1 U8202 ( .B1(n6605), .B2(n6653), .A(n6418), .ZN(P2_U3172) );
  INV_X1 U8203 ( .A(n6419), .ZN(n6434) );
  INV_X1 U8204 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6420) );
  OAI222_X1 U8205 ( .A1(n8562), .A2(n6434), .B1(n7637), .B2(P2_U3151), .C1(
        n6420), .C2(n8555), .ZN(P2_U3283) );
  NAND2_X1 U8206 ( .A1(n9074), .A2(n6773), .ZN(n6421) );
  XNOR2_X1 U8207 ( .A(n6423), .B(n6466), .ZN(n6459) );
  OAI22_X1 U8208 ( .A1(n5802), .A2(n6361), .B1(n8820), .B2(n8629), .ZN(n6460)
         );
  XNOR2_X1 U8209 ( .A(n6459), .B(n6460), .ZN(n6429) );
  OAI22_X1 U8210 ( .A1(n6427), .A2(n6426), .B1(n6466), .B2(n6425), .ZN(n6428)
         );
  NOR2_X1 U8211 ( .A1(n6429), .A2(n6428), .ZN(n6463) );
  AOI21_X1 U8212 ( .B1(n6429), .B2(n6428), .A(n6463), .ZN(n6433) );
  AOI22_X1 U8213 ( .A1(n8784), .A2(n9073), .B1(n6723), .B2(n9042), .ZN(n6444)
         );
  OAI22_X1 U8214 ( .A1(n6444), .A2(n8775), .B1(n8807), .B2(n8820), .ZN(n6430)
         );
  AOI21_X1 U8215 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6431), .A(n6430), .ZN(
        n6432) );
  OAI21_X1 U8216 ( .B1(n6433), .B2(n8792), .A(n6432), .ZN(P1_U3222) );
  INV_X1 U8217 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6435) );
  OAI222_X1 U8218 ( .A1(n9478), .A2(n6435), .B1(n9476), .B2(n6434), .C1(n7195), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8219 ( .A(n9414), .ZN(n6446) );
  OAI21_X1 U8220 ( .B1(n6438), .B2(n6437), .A(n6436), .ZN(n6445) );
  INV_X1 U8221 ( .A(n6452), .ZN(n6439) );
  AOI211_X1 U8222 ( .C1(n7324), .C2(n6440), .A(n9317), .B(n6439), .ZN(n7139)
         );
  INV_X1 U8223 ( .A(n6445), .ZN(n7143) );
  OAI21_X1 U8224 ( .B1(n8853), .B2(n6725), .A(n6441), .ZN(n6442) );
  NAND2_X1 U8225 ( .A1(n6442), .A2(n9329), .ZN(n6443) );
  OAI211_X1 U8226 ( .C1(n7143), .C2(n7069), .A(n6444), .B(n6443), .ZN(n7136)
         );
  AOI211_X1 U8227 ( .C1(n6446), .C2(n6445), .A(n7139), .B(n7136), .ZN(n6618)
         );
  INV_X1 U8228 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6447) );
  OAI22_X1 U8229 ( .A1(n9387), .A2(n8820), .B1(n9678), .B2(n6447), .ZN(n6448)
         );
  INV_X1 U8230 ( .A(n6448), .ZN(n6449) );
  OAI21_X1 U8231 ( .B1(n6618), .B2(n9676), .A(n6449), .ZN(P1_U3523) );
  OAI21_X1 U8232 ( .B1(n6451), .B2(n8857), .A(n6450), .ZN(n7093) );
  AOI211_X1 U8233 ( .C1(n6469), .C2(n6452), .A(n9317), .B(n6520), .ZN(n7092)
         );
  XNOR2_X1 U8234 ( .A(n8857), .B(n6453), .ZN(n6455) );
  OAI22_X1 U8235 ( .A1(n5802), .A2(n8800), .B1(n6568), .B2(n8798), .ZN(n6470)
         );
  INV_X1 U8236 ( .A(n6470), .ZN(n6454) );
  OAI21_X1 U8237 ( .B1(n6455), .B2(n9314), .A(n6454), .ZN(n7088) );
  AOI211_X1 U8238 ( .C1(n9673), .C2(n7093), .A(n7092), .B(n7088), .ZN(n6622)
         );
  INV_X1 U8239 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6456) );
  OAI22_X1 U8240 ( .A1(n9387), .A2(n7090), .B1(n9678), .B2(n6456), .ZN(n6457)
         );
  INV_X1 U8241 ( .A(n6457), .ZN(n6458) );
  OAI21_X1 U8242 ( .B1(n6622), .B2(n9676), .A(n6458), .ZN(P1_U3524) );
  INV_X1 U8243 ( .A(n6459), .ZN(n6462) );
  INV_X1 U8244 ( .A(n6460), .ZN(n6461) );
  NAND2_X1 U8245 ( .A1(n9073), .A2(n6773), .ZN(n6465) );
  OR2_X1 U8246 ( .A1(n7090), .A2(n8630), .ZN(n6464) );
  NAND2_X1 U8247 ( .A1(n6465), .A2(n6464), .ZN(n6467) );
  XNOR2_X1 U8248 ( .A(n6467), .B(n6466), .ZN(n6570) );
  OAI22_X1 U8249 ( .A1(n6517), .A2(n6361), .B1(n7090), .B2(n8629), .ZN(n6569)
         );
  XNOR2_X1 U8250 ( .A(n6570), .B(n6569), .ZN(n6571) );
  XNOR2_X1 U8251 ( .A(n6572), .B(n6571), .ZN(n6468) );
  NAND2_X1 U8252 ( .A1(n6468), .A2(n8797), .ZN(n6472) );
  AOI22_X1 U8253 ( .A1(n6470), .A2(n8805), .B1(n6469), .B2(n8790), .ZN(n6471)
         );
  OAI211_X1 U8254 ( .C1(n6474), .C2(n6473), .A(n6472), .B(n6471), .ZN(P1_U3237) );
  INV_X1 U8255 ( .A(n9612), .ZN(n6504) );
  XNOR2_X1 U8256 ( .A(n7195), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U8257 ( .A1(n9488), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6475) );
  OAI21_X1 U8258 ( .B1(n9488), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6475), .ZN(
        n9484) );
  NOR2_X1 U8259 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9136), .ZN(n6476) );
  AOI21_X1 U8260 ( .B1(n9136), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6476), .ZN(
        n9134) );
  NAND2_X1 U8261 ( .A1(n6487), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8262 ( .A1(n6478), .A2(n6477), .ZN(n9108) );
  MUX2_X1 U8263 ( .A(n6479), .B(P1_REG2_REG_5__SCAN_IN), .S(n9099), .Z(n9109)
         );
  NAND2_X1 U8264 ( .A1(n9108), .A2(n9109), .ZN(n9107) );
  OR2_X1 U8265 ( .A1(n9099), .A2(n6479), .ZN(n6480) );
  NAND2_X1 U8266 ( .A1(n9107), .A2(n6480), .ZN(n9122) );
  MUX2_X1 U8267 ( .A(n7109), .B(P1_REG2_REG_6__SCAN_IN), .S(n9113), .Z(n9123)
         );
  NAND2_X1 U8268 ( .A1(n9122), .A2(n9123), .ZN(n9121) );
  OR2_X1 U8269 ( .A1(n9113), .A2(n7109), .ZN(n6481) );
  NAND2_X1 U8270 ( .A1(n9121), .A2(n6481), .ZN(n9493) );
  XNOR2_X1 U8271 ( .A(n9498), .B(n9623), .ZN(n9494) );
  NAND2_X1 U8272 ( .A1(n9493), .A2(n9494), .ZN(n9492) );
  INV_X1 U8273 ( .A(n9492), .ZN(n6482) );
  AOI21_X1 U8274 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9498), .A(n6482), .ZN(
        n9510) );
  NAND2_X1 U8275 ( .A1(n9512), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6483) );
  OAI21_X1 U8276 ( .B1(n9512), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6483), .ZN(
        n9509) );
  NOR2_X1 U8277 ( .A1(n9510), .A2(n9509), .ZN(n9508) );
  AOI21_X1 U8278 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9512), .A(n9508), .ZN(
        n9133) );
  NAND2_X1 U8279 ( .A1(n9134), .A2(n9133), .ZN(n9132) );
  OAI21_X1 U8280 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9136), .A(n9132), .ZN(
        n9485) );
  NOR2_X1 U8281 ( .A1(n9484), .A2(n9485), .ZN(n9483) );
  AOI21_X1 U8282 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9488), .A(n9483), .ZN(
        n9526) );
  NAND2_X1 U8283 ( .A1(n9531), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6484) );
  OAI21_X1 U8284 ( .B1(n9531), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6484), .ZN(
        n9527) );
  NOR2_X1 U8285 ( .A1(n9526), .A2(n9527), .ZN(n9528) );
  AOI21_X1 U8286 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9531), .A(n9528), .ZN(
        n7193) );
  XNOR2_X1 U8287 ( .A(n7194), .B(n7193), .ZN(n6501) );
  INV_X1 U8288 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6485) );
  MUX2_X1 U8289 ( .A(n6485), .B(P1_REG1_REG_10__SCAN_IN), .S(n9488), .Z(n9481)
         );
  AOI22_X1 U8290 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9136), .B1(n6486), .B2(
        n5886), .ZN(n9129) );
  NAND2_X1 U8291 ( .A1(n6487), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8292 ( .A1(n6489), .A2(n6488), .ZN(n9105) );
  XNOR2_X1 U8293 ( .A(n9099), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U8294 ( .A1(n9105), .A2(n9106), .ZN(n9104) );
  INV_X1 U8295 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6490) );
  OR2_X1 U8296 ( .A1(n9099), .A2(n6490), .ZN(n6491) );
  NAND2_X1 U8297 ( .A1(n9104), .A2(n6491), .ZN(n9119) );
  XNOR2_X1 U8298 ( .A(n9113), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U8299 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  INV_X1 U8300 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6492) );
  OR2_X1 U8301 ( .A1(n9113), .A2(n6492), .ZN(n6493) );
  NAND2_X1 U8302 ( .A1(n9118), .A2(n6493), .ZN(n9496) );
  MUX2_X1 U8303 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n5862), .S(n9498), .Z(n9497)
         );
  NAND2_X1 U8304 ( .A1(n9496), .A2(n9497), .ZN(n9495) );
  NAND2_X1 U8305 ( .A1(n9498), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8306 ( .A1(n9495), .A2(n6494), .ZN(n9506) );
  OR2_X1 U8307 ( .A1(n9512), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U8308 ( .A1(n9512), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6495) );
  AND2_X1 U8309 ( .A1(n6496), .A2(n6495), .ZN(n9507) );
  AND2_X1 U8310 ( .A1(n9506), .A2(n9507), .ZN(n9515) );
  AOI21_X1 U8311 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9512), .A(n9515), .ZN(
        n9128) );
  NAND2_X1 U8312 ( .A1(n9129), .A2(n9128), .ZN(n9127) );
  OAI21_X1 U8313 ( .B1(n9136), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9127), .ZN(
        n9482) );
  NOR2_X1 U8314 ( .A1(n9481), .A2(n9482), .ZN(n9480) );
  AOI21_X1 U8315 ( .B1(n9488), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9480), .ZN(
        n9533) );
  MUX2_X1 U8316 ( .A(n6497), .B(P1_REG1_REG_11__SCAN_IN), .S(n9531), .Z(n9534)
         );
  NOR2_X1 U8317 ( .A1(n9533), .A2(n9534), .ZN(n9532) );
  AOI21_X1 U8318 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9531), .A(n9532), .ZN(
        n6499) );
  MUX2_X1 U8319 ( .A(n7181), .B(P1_REG1_REG_12__SCAN_IN), .S(n7195), .Z(n6498)
         );
  NAND2_X1 U8320 ( .A1(n6498), .A2(n6499), .ZN(n7183) );
  OAI21_X1 U8321 ( .B1(n6499), .B2(n6498), .A(n7183), .ZN(n6500) );
  AOI22_X1 U8322 ( .A1(n9605), .A2(n6501), .B1(n9597), .B2(n6500), .ZN(n6503)
         );
  AND2_X1 U8323 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7286) );
  AOI21_X1 U8324 ( .B1(n9518), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7286), .ZN(
        n6502) );
  OAI211_X1 U8325 ( .C1(n7195), .C2(n6504), .A(n6503), .B(n6502), .ZN(P1_U3255) );
  INV_X1 U8326 ( .A(n6510), .ZN(n8852) );
  XNOR2_X1 U8327 ( .A(n6505), .B(n8852), .ZN(n6507) );
  NAND2_X1 U8328 ( .A1(n9072), .A2(n9042), .ZN(n6506) );
  OAI21_X1 U8329 ( .B1(n6791), .B2(n8798), .A(n6506), .ZN(n8756) );
  AOI21_X1 U8330 ( .B1(n6507), .B2(n9329), .A(n8756), .ZN(n7098) );
  AOI21_X1 U8331 ( .B1(n6519), .B2(n8754), .A(n9317), .ZN(n6508) );
  NAND2_X1 U8332 ( .A1(n6508), .A2(n6587), .ZN(n7099) );
  AND2_X1 U8333 ( .A1(n7098), .A2(n7099), .ZN(n6666) );
  OAI21_X1 U8334 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(n7097) );
  INV_X1 U8335 ( .A(n9407), .ZN(n7293) );
  OAI22_X1 U8336 ( .A1(n9387), .A2(n7100), .B1(n9678), .B2(n6512), .ZN(n6513)
         );
  AOI21_X1 U8337 ( .B1(n7097), .B2(n7293), .A(n6513), .ZN(n6514) );
  OAI21_X1 U8338 ( .B1(n6666), .B2(n9676), .A(n6514), .ZN(P1_U3526) );
  XOR2_X1 U8339 ( .A(n8858), .B(n6515), .Z(n6518) );
  OAI22_X1 U8340 ( .A1(n6517), .A2(n8800), .B1(n6516), .B2(n8798), .ZN(n6574)
         );
  AOI21_X1 U8341 ( .B1(n6518), .B2(n9329), .A(n6574), .ZN(n7071) );
  OAI211_X1 U8342 ( .C1(n6520), .C2(n7074), .A(n6519), .B(n9342), .ZN(n7072)
         );
  AND2_X1 U8343 ( .A1(n7071), .A2(n7072), .ZN(n6669) );
  OAI21_X1 U8344 ( .B1(n6522), .B2(n8858), .A(n6521), .ZN(n7063) );
  INV_X1 U8345 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6523) );
  OAI22_X1 U8346 ( .A1(n9387), .A2(n7074), .B1(n9678), .B2(n6523), .ZN(n6524)
         );
  AOI21_X1 U8347 ( .B1(n7063), .B2(n7293), .A(n6524), .ZN(n6525) );
  OAI21_X1 U8348 ( .B1(n6669), .B2(n9676), .A(n6525), .ZN(P1_U3525) );
  INV_X1 U8349 ( .A(n6546), .ZN(n9688) );
  MUX2_X1 U8350 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8257), .Z(n6530) );
  INV_X1 U8351 ( .A(n6530), .ZN(n6531) );
  INV_X1 U8352 ( .A(n6543), .ZN(n6529) );
  INV_X1 U8353 ( .A(n6526), .ZN(n6528) );
  OAI21_X1 U8354 ( .B1(n6529), .B2(n6528), .A(n6527), .ZN(n9690) );
  XNOR2_X1 U8355 ( .A(n6530), .B(n6546), .ZN(n9691) );
  NOR2_X1 U8356 ( .A1(n9690), .A2(n9691), .ZN(n9689) );
  MUX2_X1 U8357 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8257), .Z(n6687) );
  XOR2_X1 U8358 ( .A(n6707), .B(n6687), .Z(n6532) );
  OAI211_X1 U8359 ( .C1(n6533), .C2(n6532), .A(n6688), .B(n9851), .ZN(n6557)
         );
  NAND2_X1 U8360 ( .A1(n6543), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8361 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  INV_X1 U8362 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6741) );
  XNOR2_X1 U8363 ( .A(n6707), .B(n6741), .ZN(n6538) );
  NAND2_X1 U8364 ( .A1(n6537), .A2(n6538), .ZN(n6695) );
  INV_X1 U8365 ( .A(n6538), .ZN(n6540) );
  NAND3_X1 U8366 ( .A1(n9679), .A2(n6540), .A3(n6539), .ZN(n6541) );
  AND2_X1 U8367 ( .A1(n6695), .A2(n6541), .ZN(n6554) );
  MUX2_X1 U8368 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6542), .S(n6707), .Z(n6551)
         );
  NAND2_X1 U8369 ( .A1(n6543), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8370 ( .A1(n6545), .A2(n6544), .ZN(n6547) );
  XNOR2_X1 U8371 ( .A(n6547), .B(n9688), .ZN(n9682) );
  NAND2_X1 U8372 ( .A1(n9682), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8373 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  NAND2_X1 U8374 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NAND2_X1 U8375 ( .A1(n6550), .A2(n6551), .ZN(n6709) );
  OAI21_X1 U8376 ( .B1(n6551), .B2(n6550), .A(n6709), .ZN(n6552) );
  NAND2_X1 U8377 ( .A1(n9852), .A2(n6552), .ZN(n6553) );
  NAND2_X1 U8378 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6625) );
  OAI211_X1 U8379 ( .C1(n6554), .C2(n9856), .A(n6553), .B(n6625), .ZN(n6555)
         );
  AOI21_X1 U8380 ( .B1(n9842), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6555), .ZN(
        n6556) );
  OAI211_X1 U8381 ( .C1(n9708), .C2(n6707), .A(n6557), .B(n6556), .ZN(P2_U3186) );
  OAI211_X1 U8382 ( .C1(n6560), .C2(n6559), .A(n6558), .B(n8160), .ZN(n6564)
         );
  NOR2_X1 U8383 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5105), .ZN(n9683) );
  OAI22_X1 U8384 ( .A1(n8167), .A2(n6561), .B1(n6752), .B2(n8170), .ZN(n6562)
         );
  AOI211_X1 U8385 ( .C1(n8172), .C2(n8198), .A(n9683), .B(n6562), .ZN(n6563)
         );
  OAI211_X1 U8386 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8174), .A(n6564), .B(
        n6563), .ZN(P2_U3158) );
  NAND2_X1 U8387 ( .A1(n9072), .A2(n6773), .ZN(n6566) );
  OR2_X1 U8388 ( .A1(n7074), .A2(n8630), .ZN(n6565) );
  NAND2_X1 U8389 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  XNOR2_X1 U8390 ( .A(n6567), .B(n6466), .ZN(n6777) );
  OAI22_X1 U8391 ( .A1(n6568), .A2(n6361), .B1(n7074), .B2(n8629), .ZN(n6778)
         );
  XOR2_X1 U8392 ( .A(n6777), .B(n6778), .Z(n6781) );
  XOR2_X1 U8393 ( .A(n6781), .B(n6782), .Z(n6581) );
  AOI22_X1 U8394 ( .A1(n6574), .A2(n8805), .B1(n6573), .B2(n8790), .ZN(n6580)
         );
  MUX2_X1 U8395 ( .A(n8803), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6579) );
  OAI211_X1 U8396 ( .C1(n6581), .C2(n8792), .A(n6580), .B(n6579), .ZN(P1_U3218) );
  INV_X1 U8397 ( .A(n6582), .ZN(n6593) );
  AOI22_X1 U8398 ( .A1(n9553), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10045), .ZN(n6583) );
  OAI21_X1 U8399 ( .B1(n6593), .B2(n9476), .A(n6583), .ZN(P1_U3342) );
  OAI21_X1 U8400 ( .B1(n6585), .B2(n8856), .A(n6584), .ZN(n7253) );
  NAND2_X1 U8401 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  NAND2_X1 U8402 ( .A1(n6588), .A2(n9342), .ZN(n6589) );
  NOR2_X1 U8403 ( .A1(n6635), .A2(n6589), .ZN(n7248) );
  XNOR2_X1 U8404 ( .A(n8913), .B(n8856), .ZN(n6590) );
  OAI21_X1 U8405 ( .B1(n6590), .B2(n9314), .A(n7699), .ZN(n7247) );
  AOI211_X1 U8406 ( .C1(n9673), .C2(n7253), .A(n7248), .B(n7247), .ZN(n6615)
         );
  OAI22_X1 U8407 ( .A1(n9387), .A2(n7704), .B1(n9678), .B2(n6490), .ZN(n6591)
         );
  INV_X1 U8408 ( .A(n6591), .ZN(n6592) );
  OAI21_X1 U8409 ( .B1(n6615), .B2(n9676), .A(n6592), .ZN(P1_U3527) );
  INV_X1 U8410 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10257) );
  INV_X1 U8411 ( .A(n8202), .ZN(n8236) );
  OAI222_X1 U8412 ( .A1(n8555), .A2(n10257), .B1(n8562), .B2(n6593), .C1(
        P2_U3151), .C2(n8236), .ZN(P2_U3282) );
  XOR2_X1 U8413 ( .A(n6595), .B(n6594), .Z(n6601) );
  INV_X1 U8414 ( .A(n5632), .ZN(n6597) );
  OAI22_X1 U8415 ( .A1(n6597), .A2(n8143), .B1(n8170), .B2(n6596), .ZN(n6599)
         );
  NOR2_X1 U8416 ( .A1(n6605), .A2(n10212), .ZN(n6598) );
  AOI211_X1 U8417 ( .C1(n5059), .C2(n8182), .A(n6599), .B(n6598), .ZN(n6600)
         );
  OAI21_X1 U8418 ( .B1(n8177), .B2(n6601), .A(n6600), .ZN(P2_U3162) );
  XOR2_X1 U8419 ( .A(n6603), .B(n6602), .Z(n6610) );
  OAI22_X1 U8420 ( .A1(n6604), .A2(n8170), .B1(n8143), .B2(n5060), .ZN(n6607)
         );
  NOR2_X1 U8421 ( .A1(n6605), .A2(n6321), .ZN(n6606) );
  AOI211_X1 U8422 ( .C1(n6608), .C2(n8182), .A(n6607), .B(n6606), .ZN(n6609)
         );
  OAI21_X1 U8423 ( .B1(n6610), .B2(n8177), .A(n6609), .ZN(P2_U3177) );
  INV_X1 U8424 ( .A(n6611), .ZN(n6662) );
  AOI22_X1 U8425 ( .A1(n9566), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10045), .ZN(n6612) );
  OAI21_X1 U8426 ( .B1(n6662), .B2(n9476), .A(n6612), .ZN(P1_U3341) );
  OAI22_X1 U8427 ( .A1(n9442), .A2(n7704), .B1(n9464), .B2(n5836), .ZN(n6613)
         );
  INV_X1 U8428 ( .A(n6613), .ZN(n6614) );
  OAI21_X1 U8429 ( .B1(n6615), .B2(n9674), .A(n6614), .ZN(P1_U3468) );
  INV_X1 U8430 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10124) );
  OAI22_X1 U8431 ( .A1(n9442), .A2(n8820), .B1(n9464), .B2(n10124), .ZN(n6616)
         );
  INV_X1 U8432 ( .A(n6616), .ZN(n6617) );
  OAI21_X1 U8433 ( .B1(n6618), .B2(n9674), .A(n6617), .ZN(P1_U3456) );
  INV_X1 U8434 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6619) );
  OAI22_X1 U8435 ( .A1(n9442), .A2(n7090), .B1(n9464), .B2(n6619), .ZN(n6620)
         );
  INV_X1 U8436 ( .A(n6620), .ZN(n6621) );
  OAI21_X1 U8437 ( .B1(n6622), .B2(n9674), .A(n6621), .ZN(P1_U3459) );
  AOI21_X1 U8438 ( .B1(n6624), .B2(n6623), .A(n4510), .ZN(n6632) );
  INV_X1 U8439 ( .A(n6625), .ZN(n6628) );
  INV_X1 U8440 ( .A(n8196), .ZN(n6626) );
  OAI22_X1 U8441 ( .A1(n8167), .A2(n9896), .B1(n6626), .B2(n8170), .ZN(n6627)
         );
  AOI211_X1 U8442 ( .C1(n8172), .C2(n9868), .A(n6628), .B(n6627), .ZN(n6631)
         );
  INV_X1 U8443 ( .A(n6629), .ZN(n6742) );
  NAND2_X1 U8444 ( .A1(n8164), .A2(n6742), .ZN(n6630) );
  OAI211_X1 U8445 ( .C1(n6632), .C2(n8177), .A(n6631), .B(n6630), .ZN(P2_U3170) );
  OAI21_X1 U8446 ( .B1(n6634), .B2(n8855), .A(n6633), .ZN(n7106) );
  OAI21_X1 U8447 ( .B1(n6635), .B2(n7111), .A(n9342), .ZN(n6636) );
  NOR2_X1 U8448 ( .A1(n6636), .A2(n6830), .ZN(n7113) );
  XNOR2_X1 U8449 ( .A(n6637), .B(n8855), .ZN(n6639) );
  OAI22_X1 U8450 ( .A1(n6898), .A2(n8798), .B1(n6791), .B2(n8800), .ZN(n6915)
         );
  INV_X1 U8451 ( .A(n6915), .ZN(n6638) );
  OAI21_X1 U8452 ( .B1(n6639), .B2(n9314), .A(n6638), .ZN(n7107) );
  AOI211_X1 U8453 ( .C1(n9673), .C2(n7106), .A(n7113), .B(n7107), .ZN(n6644)
         );
  OAI22_X1 U8454 ( .A1(n9442), .A2(n7111), .B1(n9464), .B2(n5848), .ZN(n6640)
         );
  INV_X1 U8455 ( .A(n6640), .ZN(n6641) );
  OAI21_X1 U8456 ( .B1(n6644), .B2(n9674), .A(n6641), .ZN(P1_U3471) );
  OAI22_X1 U8457 ( .A1(n9387), .A2(n7111), .B1(n9678), .B2(n6492), .ZN(n6642)
         );
  INV_X1 U8458 ( .A(n6642), .ZN(n6643) );
  OAI21_X1 U8459 ( .B1(n6644), .B2(n9676), .A(n6643), .ZN(P1_U3528) );
  INV_X1 U8460 ( .A(n6645), .ZN(n6648) );
  INV_X1 U8461 ( .A(n6646), .ZN(n6647) );
  MUX2_X1 U8462 ( .A(n6649), .B(n6648), .S(n6647), .Z(n6650) );
  OAI22_X1 U8463 ( .A1(n8403), .A2(n6654), .B1(n6653), .B2(n9863), .ZN(n6660)
         );
  NAND3_X1 U8464 ( .A1(n6656), .A2(n6655), .A3(n9919), .ZN(n6658) );
  AOI21_X1 U8465 ( .B1(n6658), .B2(n6657), .A(n6677), .ZN(n6659) );
  AOI211_X1 U8466 ( .C1(n6677), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6660), .B(
        n6659), .ZN(n6661) );
  INV_X1 U8467 ( .A(n6661), .ZN(P2_U3233) );
  OAI222_X1 U8468 ( .A1(n8555), .A2(n6663), .B1(n8562), .B2(n6662), .C1(
        P2_U3151), .C2(n8234), .ZN(P2_U3281) );
  INV_X1 U8469 ( .A(n9462), .ZN(n7296) );
  INV_X1 U8470 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10206) );
  OAI22_X1 U8471 ( .A1(n9442), .A2(n7100), .B1(n9464), .B2(n10206), .ZN(n6664)
         );
  AOI21_X1 U8472 ( .B1(n7097), .B2(n7296), .A(n6664), .ZN(n6665) );
  OAI21_X1 U8473 ( .B1(n6666), .B2(n9674), .A(n6665), .ZN(P1_U3465) );
  INV_X1 U8474 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10062) );
  OAI22_X1 U8475 ( .A1(n9442), .A2(n7074), .B1(n9464), .B2(n10062), .ZN(n6667)
         );
  AOI21_X1 U8476 ( .B1(n7063), .B2(n7296), .A(n6667), .ZN(n6668) );
  OAI21_X1 U8477 ( .B1(n6669), .B2(n9674), .A(n6668), .ZN(P1_U3462) );
  NAND2_X1 U8478 ( .A1(n6670), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6671) );
  OAI21_X1 U8479 ( .B1(n7706), .B2(n6670), .A(n6671), .ZN(P1_U3583) );
  INV_X1 U8480 ( .A(n6673), .ZN(n7836) );
  XNOR2_X1 U8481 ( .A(n7836), .B(n6672), .ZN(n6676) );
  AOI22_X1 U8482 ( .A1(n9866), .A2(n5632), .B1(n8198), .B2(n9869), .ZN(n6675)
         );
  XNOR2_X1 U8483 ( .A(n6185), .B(n6673), .ZN(n9882) );
  NAND2_X1 U8484 ( .A1(n9882), .A2(n9927), .ZN(n6674) );
  OAI211_X1 U8485 ( .C1(n6676), .C2(n9873), .A(n6675), .B(n6674), .ZN(n9880)
         );
  INV_X1 U8486 ( .A(n9880), .ZN(n6683) );
  AND2_X1 U8487 ( .A1(n7833), .A2(n6678), .ZN(n9875) );
  NAND2_X1 U8488 ( .A1(n8413), .A2(n9875), .ZN(n8286) );
  INV_X1 U8489 ( .A(n8286), .ZN(n6681) );
  AOI22_X1 U8490 ( .A1(n8438), .A2(n5059), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8437), .ZN(n6679) );
  OAI21_X1 U8491 ( .B1(n5031), .B2(n8413), .A(n6679), .ZN(n6680) );
  AOI21_X1 U8492 ( .B1(n6681), .B2(n9882), .A(n6680), .ZN(n6682) );
  OAI21_X1 U8493 ( .B1(n6683), .B2(n6677), .A(n6682), .ZN(P2_U3232) );
  INV_X1 U8494 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7406) );
  MUX2_X1 U8495 ( .A(n7406), .B(n6684), .S(n8257), .Z(n7431) );
  XNOR2_X1 U8496 ( .A(n7431), .B(n7432), .ZN(n6693) );
  INV_X1 U8497 ( .A(n9707), .ZN(n6710) );
  MUX2_X1 U8498 ( .A(n6686), .B(n6685), .S(n8257), .Z(n6691) );
  INV_X1 U8499 ( .A(n6707), .ZN(n6690) );
  INV_X1 U8500 ( .A(n6687), .ZN(n6689) );
  XNOR2_X1 U8501 ( .A(n6691), .B(n9707), .ZN(n9703) );
  OAI21_X1 U8502 ( .B1(n6710), .B2(n6691), .A(n9702), .ZN(n6692) );
  NOR2_X1 U8503 ( .A1(n6692), .A2(n6693), .ZN(n7430) );
  AOI21_X1 U8504 ( .B1(n6693), .B2(n6692), .A(n7430), .ZN(n6722) );
  INV_X1 U8505 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U8506 ( .A1(n6707), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6694) );
  MUX2_X1 U8507 ( .A(n7406), .B(P2_REG2_REG_6__SCAN_IN), .S(n7432), .Z(n6701)
         );
  INV_X1 U8508 ( .A(n6701), .ZN(n6697) );
  AOI21_X1 U8509 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(n7408) );
  NOR3_X1 U8510 ( .A1(n6702), .A2(n6701), .A3(n6700), .ZN(n6703) );
  OAI21_X1 U8511 ( .B1(n7408), .B2(n6703), .A(n9718), .ZN(n6705) );
  INV_X1 U8512 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10190) );
  NOR2_X1 U8513 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10190), .ZN(n6936) );
  INV_X1 U8514 ( .A(n6936), .ZN(n6704) );
  OAI211_X1 U8515 ( .C1(n6706), .C2(n9713), .A(n6705), .B(n6704), .ZN(n6720)
         );
  NAND2_X1 U8516 ( .A1(n6707), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8517 ( .A1(n6709), .A2(n6708), .ZN(n6712) );
  XNOR2_X1 U8518 ( .A(n6712), .B(n6710), .ZN(n9699) );
  NAND2_X1 U8519 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n9699), .ZN(n9698) );
  INV_X1 U8520 ( .A(n9698), .ZN(n6711) );
  MUX2_X1 U8521 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6684), .S(n7432), .Z(n6715)
         );
  INV_X1 U8522 ( .A(n6715), .ZN(n6713) );
  NAND2_X1 U8523 ( .A1(n6714), .A2(n6713), .ZN(n7422) );
  NAND2_X1 U8524 ( .A1(n6716), .A2(n6715), .ZN(n6718) );
  INV_X1 U8525 ( .A(n9852), .ZN(n6717) );
  AOI21_X1 U8526 ( .B1(n7422), .B2(n6718), .A(n6717), .ZN(n6719) );
  AOI211_X1 U8527 ( .C1(n9844), .C2(n7432), .A(n6720), .B(n6719), .ZN(n6721)
         );
  OAI21_X1 U8528 ( .B1(n6722), .B2(n9692), .A(n6721), .ZN(P2_U3188) );
  INV_X1 U8529 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U8530 ( .A1(n6723), .A2(n6727), .ZN(n8825) );
  INV_X1 U8531 ( .A(n8825), .ZN(n6724) );
  NOR2_X1 U8532 ( .A1(n6725), .A2(n6724), .ZN(n8854) );
  INV_X1 U8533 ( .A(n8854), .ZN(n7318) );
  OAI21_X1 U8534 ( .B1(n9329), .B2(n9673), .A(n7318), .ZN(n6726) );
  OAI211_X1 U8535 ( .C1(n6727), .C2(n7317), .A(n6726), .B(n7319), .ZN(n9416)
         );
  NAND2_X1 U8536 ( .A1(n9416), .A2(n9464), .ZN(n6728) );
  OAI21_X1 U8537 ( .B1(n9464), .B2(n6729), .A(n6728), .ZN(P1_U3453) );
  INV_X1 U8538 ( .A(n6730), .ZN(n6746) );
  INV_X1 U8539 ( .A(n9809), .ZN(n8241) );
  OAI222_X1 U8540 ( .A1(n8562), .A2(n6746), .B1(n8241), .B2(P2_U3151), .C1(
        n6731), .C2(n8555), .ZN(P2_U3280) );
  INV_X1 U8541 ( .A(n8799), .ZN(n8644) );
  NAND2_X1 U8542 ( .A1(n8644), .A2(P1_U3973), .ZN(n6732) );
  OAI21_X1 U8543 ( .B1(P1_U3973), .B2(n8036), .A(n6732), .ZN(P1_U3581) );
  OR2_X1 U8544 ( .A1(n9927), .A2(n9875), .ZN(n6733) );
  XNOR2_X1 U8545 ( .A(n6734), .B(n7838), .ZN(n9894) );
  NAND2_X1 U8546 ( .A1(n6736), .A2(n6735), .ZN(n6765) );
  NAND2_X1 U8547 ( .A1(n6765), .A2(n6764), .ZN(n6738) );
  NAND2_X1 U8548 ( .A1(n6738), .A2(n6737), .ZN(n6739) );
  XNOR2_X1 U8549 ( .A(n6739), .B(n7838), .ZN(n6740) );
  AOI222_X1 U8550 ( .A1(n8433), .A2(n6740), .B1(n9868), .B2(n9866), .C1(n8196), 
        .C2(n9869), .ZN(n9895) );
  MUX2_X1 U8551 ( .A(n6741), .B(n9895), .S(n9876), .Z(n6745) );
  AOI22_X1 U8552 ( .A1(n8438), .A2(n6743), .B1(n8437), .B2(n6742), .ZN(n6744)
         );
  OAI211_X1 U8553 ( .C1(n8441), .C2(n9894), .A(n6745), .B(n6744), .ZN(P2_U3229) );
  INV_X1 U8554 ( .A(n9587), .ZN(n7199) );
  OAI222_X1 U8555 ( .A1(n9478), .A2(n6747), .B1(n9476), .B2(n6746), .C1(n7199), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  OAI21_X1 U8556 ( .B1(n6748), .B2(n7842), .A(n6869), .ZN(n9902) );
  INV_X1 U8557 ( .A(n9902), .ZN(n6761) );
  NAND2_X1 U8558 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  XNOR2_X1 U8559 ( .A(n6751), .B(n7842), .ZN(n6755) );
  OAI22_X1 U8560 ( .A1(n4733), .A2(n8394), .B1(n6752), .B2(n8396), .ZN(n6753)
         );
  AOI21_X1 U8561 ( .B1(n9902), .B2(n9927), .A(n6753), .ZN(n6754) );
  OAI21_X1 U8562 ( .B1(n9873), .B2(n6755), .A(n6754), .ZN(n9900) );
  NAND2_X1 U8563 ( .A1(n9900), .A2(n9876), .ZN(n6760) );
  OAI22_X1 U8564 ( .A1(n8413), .A2(n6686), .B1(n6756), .B2(n9863), .ZN(n6757)
         );
  AOI21_X1 U8565 ( .B1(n8438), .B2(n6758), .A(n6757), .ZN(n6759) );
  OAI211_X1 U8566 ( .C1(n6761), .C2(n8286), .A(n6760), .B(n6759), .ZN(P2_U3228) );
  OAI21_X1 U8567 ( .B1(n6763), .B2(n5103), .A(n6762), .ZN(n9890) );
  INV_X1 U8568 ( .A(n9890), .ZN(n6770) );
  XNOR2_X1 U8569 ( .A(n6765), .B(n6764), .ZN(n6766) );
  AOI222_X1 U8570 ( .A1(n8433), .A2(n6766), .B1(n8198), .B2(n9866), .C1(n8197), 
        .C2(n9869), .ZN(n9892) );
  MUX2_X1 U8571 ( .A(n6767), .B(n9892), .S(n9876), .Z(n6769) );
  AOI22_X1 U8572 ( .A1(n8438), .A2(n9889), .B1(n5105), .B2(n8437), .ZN(n6768)
         );
  OAI211_X1 U8573 ( .C1(n6770), .C2(n8441), .A(n6769), .B(n6768), .ZN(P2_U3230) );
  NAND2_X1 U8574 ( .A1(n9626), .A2(n4574), .ZN(n6771) );
  OAI21_X1 U8575 ( .B1(n6898), .B2(n8629), .A(n6771), .ZN(n6772) );
  XNOR2_X1 U8576 ( .A(n6772), .B(n6466), .ZN(n6776) );
  NAND2_X1 U8577 ( .A1(n9626), .A2(n6773), .ZN(n6774) );
  OAI21_X1 U8578 ( .B1(n6898), .B2(n6361), .A(n6774), .ZN(n6775) );
  NOR2_X1 U8579 ( .A1(n6776), .A2(n6775), .ZN(n6961) );
  AOI21_X1 U8580 ( .B1(n6776), .B2(n6775), .A(n6961), .ZN(n6800) );
  INV_X1 U8581 ( .A(n6777), .ZN(n6780) );
  INV_X1 U8582 ( .A(n6778), .ZN(n6779) );
  OR2_X1 U8583 ( .A1(n7100), .A2(n8630), .ZN(n6783) );
  NAND2_X1 U8584 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  XNOR2_X1 U8585 ( .A(n6785), .B(n6466), .ZN(n6786) );
  XNOR2_X1 U8586 ( .A(n6786), .B(n6787), .ZN(n8751) );
  NAND2_X1 U8587 ( .A1(n8752), .A2(n8751), .ZN(n8750) );
  INV_X1 U8588 ( .A(n6787), .ZN(n6788) );
  OAI22_X1 U8589 ( .A1(n6791), .A2(n8629), .B1(n7704), .B2(n8630), .ZN(n6790)
         );
  XNOR2_X1 U8590 ( .A(n6790), .B(n6422), .ZN(n6909) );
  INV_X1 U8591 ( .A(n6909), .ZN(n6907) );
  OAI22_X1 U8592 ( .A1(n6791), .A2(n6361), .B1(n7704), .B2(n8629), .ZN(n6793)
         );
  INV_X1 U8593 ( .A(n6793), .ZN(n7696) );
  OAI22_X1 U8594 ( .A1(n6801), .A2(n8629), .B1(n7111), .B2(n8630), .ZN(n6792)
         );
  XNOR2_X1 U8595 ( .A(n6792), .B(n8681), .ZN(n6796) );
  INV_X1 U8596 ( .A(n6796), .ZN(n6912) );
  OAI22_X1 U8597 ( .A1(n6801), .A2(n6361), .B1(n7111), .B2(n8629), .ZN(n6911)
         );
  NAND2_X1 U8598 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  OAI21_X1 U8599 ( .B1(n6907), .B2(n7696), .A(n6910), .ZN(n6798) );
  OAI21_X1 U8600 ( .B1(n6909), .B2(n6793), .A(n6911), .ZN(n6795) );
  NOR3_X1 U8601 ( .A1(n6909), .A2(n6793), .A3(n6911), .ZN(n6794) );
  AOI21_X1 U8602 ( .B1(n6796), .B2(n6795), .A(n6794), .ZN(n6797) );
  NAND2_X1 U8603 ( .A1(n6799), .A2(n6800), .ZN(n6963) );
  OAI21_X1 U8604 ( .B1(n6800), .B2(n6799), .A(n6963), .ZN(n6805) );
  NOR2_X1 U8605 ( .A1(n8807), .A2(n6835), .ZN(n6804) );
  OAI22_X1 U8606 ( .A1(n6966), .A2(n8798), .B1(n6801), .B2(n8800), .ZN(n6829)
         );
  NAND2_X1 U8607 ( .A1(n6829), .A2(n8805), .ZN(n6802) );
  NAND2_X1 U8608 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9503) );
  OAI211_X1 U8609 ( .C1(n8803), .C2(n9622), .A(n6802), .B(n9503), .ZN(n6803)
         );
  AOI211_X1 U8610 ( .C1(n6805), .C2(n8797), .A(n6804), .B(n6803), .ZN(n6806)
         );
  INV_X1 U8611 ( .A(n6806), .ZN(P1_U3213) );
  INV_X1 U8612 ( .A(n6807), .ZN(n6809) );
  INV_X1 U8613 ( .A(n9599), .ZN(n7190) );
  OAI222_X1 U8614 ( .A1(n9478), .A2(n6808), .B1(n9476), .B2(n6809), .C1(
        P1_U3086), .C2(n7190), .ZN(P1_U3339) );
  OAI222_X1 U8615 ( .A1(n8555), .A2(n6810), .B1(n8562), .B2(n6809), .C1(
        P2_U3151), .C2(n8232), .ZN(P2_U3279) );
  NAND2_X1 U8616 ( .A1(n6811), .A2(n7914), .ZN(n7014) );
  NAND2_X1 U8617 ( .A1(n7014), .A2(n7916), .ZN(n6840) );
  OAI21_X1 U8618 ( .B1(n7014), .B2(n7916), .A(n6840), .ZN(n9911) );
  NAND2_X1 U8619 ( .A1(n6872), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8620 ( .A1(n6814), .A2(n6813), .ZN(n6816) );
  OAI21_X1 U8621 ( .B1(n6816), .B2(n5180), .A(n6815), .ZN(n6817) );
  AOI222_X1 U8622 ( .A1(n8433), .A2(n6817), .B1(n8193), .B2(n9869), .C1(n8195), 
        .C2(n9866), .ZN(n9909) );
  MUX2_X1 U8623 ( .A(n6818), .B(n9909), .S(n8413), .Z(n6821) );
  INV_X1 U8624 ( .A(n6819), .ZN(n6958) );
  AOI22_X1 U8625 ( .A1(n8438), .A2(n6952), .B1(n8437), .B2(n6958), .ZN(n6820)
         );
  OAI211_X1 U8626 ( .C1(n8441), .C2(n9911), .A(n6821), .B(n6820), .ZN(P2_U3226) );
  NAND2_X1 U8627 ( .A1(n8320), .A2(P2_U3893), .ZN(n6822) );
  OAI21_X1 U8628 ( .B1(P2_U3893), .B2(n6073), .A(n6822), .ZN(P2_U3518) );
  OAI21_X1 U8629 ( .B1(n6824), .B2(n6826), .A(n6823), .ZN(n9633) );
  INV_X1 U8630 ( .A(n9633), .ZN(n6831) );
  INV_X1 U8631 ( .A(n7069), .ZN(n7493) );
  NAND2_X1 U8632 ( .A1(n6825), .A2(n8910), .ZN(n8916) );
  XNOR2_X1 U8633 ( .A(n8916), .B(n4812), .ZN(n6827) );
  NOR2_X1 U8634 ( .A1(n6827), .A2(n9314), .ZN(n6828) );
  AOI211_X1 U8635 ( .C1(n9633), .C2(n7493), .A(n6829), .B(n6828), .ZN(n9635)
         );
  OAI211_X1 U8636 ( .C1(n6830), .C2(n6835), .A(n9342), .B(n6891), .ZN(n9630)
         );
  OAI211_X1 U8637 ( .C1(n6831), .C2(n9414), .A(n9635), .B(n9630), .ZN(n6837)
         );
  OAI22_X1 U8638 ( .A1(n9387), .A2(n6835), .B1(n9678), .B2(n5862), .ZN(n6832)
         );
  AOI21_X1 U8639 ( .B1(n6837), .B2(n9678), .A(n6832), .ZN(n6833) );
  INV_X1 U8640 ( .A(n6833), .ZN(P1_U3529) );
  INV_X1 U8641 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6834) );
  OAI22_X1 U8642 ( .A1(n9442), .A2(n6835), .B1(n9464), .B2(n6834), .ZN(n6836)
         );
  AOI21_X1 U8643 ( .B1(n6837), .B2(n9464), .A(n6836), .ZN(n6838) );
  INV_X1 U8644 ( .A(n6838), .ZN(P1_U3474) );
  NAND2_X1 U8645 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  XNOR2_X1 U8646 ( .A(n6841), .B(n7846), .ZN(n9914) );
  XNOR2_X1 U8647 ( .A(n6842), .B(n7846), .ZN(n6843) );
  OAI222_X1 U8648 ( .A1(n8394), .A2(n7305), .B1(n8396), .B2(n6937), .C1(n9873), 
        .C2(n6843), .ZN(n9915) );
  NAND2_X1 U8649 ( .A1(n9915), .A2(n9876), .ZN(n6846) );
  OAI22_X1 U8650 ( .A1(n8413), .A2(n7412), .B1(n7009), .B2(n9863), .ZN(n6844)
         );
  AOI21_X1 U8651 ( .B1(n8438), .B2(n9917), .A(n6844), .ZN(n6845) );
  OAI211_X1 U8652 ( .C1(n9914), .C2(n8441), .A(n6846), .B(n6845), .ZN(P2_U3225) );
  INV_X1 U8653 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9969) );
  NOR2_X1 U8654 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6847) );
  AOI21_X1 U8655 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6847), .ZN(n9975) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10068) );
  INV_X1 U8657 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U8658 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10068), .B2(n10050), .ZN(n9978) );
  NOR2_X1 U8659 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6848) );
  AOI21_X1 U8660 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6848), .ZN(n9981) );
  NOR2_X1 U8661 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6849) );
  AOI21_X1 U8662 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6849), .ZN(n9984) );
  NOR2_X1 U8663 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6850) );
  AOI21_X1 U8664 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6850), .ZN(n9987) );
  NOR2_X1 U8665 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6851) );
  AOI21_X1 U8666 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6851), .ZN(n9990) );
  NOR2_X1 U8667 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6852) );
  AOI21_X1 U8668 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6852), .ZN(n9993) );
  NOR2_X1 U8669 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6853) );
  AOI21_X1 U8670 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6853), .ZN(n9996) );
  NOR2_X1 U8671 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6854) );
  AOI21_X1 U8672 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6854), .ZN(n10299) );
  NOR2_X1 U8673 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6855) );
  AOI21_X1 U8674 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6855), .ZN(n10305) );
  NOR2_X1 U8675 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6856) );
  AOI21_X1 U8676 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6856), .ZN(n10302) );
  NOR2_X1 U8677 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6857) );
  AOI21_X1 U8678 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6857), .ZN(n10293) );
  NOR2_X1 U8679 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6858) );
  AOI21_X1 U8680 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6858), .ZN(n10296) );
  AND2_X1 U8681 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6859) );
  NOR2_X1 U8682 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6859), .ZN(n9965) );
  INV_X1 U8683 ( .A(n9965), .ZN(n9966) );
  NAND3_X1 U8684 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U8685 ( .A1(n10246), .A2(n9967), .ZN(n9964) );
  NAND2_X1 U8686 ( .A1(n9966), .A2(n9964), .ZN(n10308) );
  NAND2_X1 U8687 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6860) );
  OAI21_X1 U8688 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n6860), .ZN(n10307) );
  NOR2_X1 U8689 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  AOI21_X1 U8690 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10306), .ZN(n10311) );
  NAND2_X1 U8691 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6861) );
  OAI21_X1 U8692 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6861), .ZN(n10310) );
  NOR2_X1 U8693 ( .A1(n10311), .A2(n10310), .ZN(n10309) );
  AOI21_X1 U8694 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10309), .ZN(n10314) );
  NOR2_X1 U8695 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6862) );
  AOI21_X1 U8696 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6862), .ZN(n10313) );
  NAND2_X1 U8697 ( .A1(n10314), .A2(n10313), .ZN(n10312) );
  OAI21_X1 U8698 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10312), .ZN(n10295) );
  NAND2_X1 U8699 ( .A1(n10296), .A2(n10295), .ZN(n10294) );
  OAI21_X1 U8700 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10294), .ZN(n10292) );
  NAND2_X1 U8701 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  OAI21_X1 U8702 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10291), .ZN(n10301) );
  NAND2_X1 U8703 ( .A1(n10302), .A2(n10301), .ZN(n10300) );
  OAI21_X1 U8704 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10300), .ZN(n10304) );
  NAND2_X1 U8705 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  OAI21_X1 U8706 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10303), .ZN(n10298) );
  NAND2_X1 U8707 ( .A1(n10299), .A2(n10298), .ZN(n10297) );
  OAI21_X1 U8708 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10297), .ZN(n9995) );
  NAND2_X1 U8709 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OAI21_X1 U8710 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9994), .ZN(n9992) );
  NAND2_X1 U8711 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  OAI21_X1 U8712 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9991), .ZN(n9989) );
  NAND2_X1 U8713 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  OAI21_X1 U8714 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9988), .ZN(n9986) );
  NAND2_X1 U8715 ( .A1(n9987), .A2(n9986), .ZN(n9985) );
  OAI21_X1 U8716 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9985), .ZN(n9983) );
  NAND2_X1 U8717 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  OAI21_X1 U8718 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9982), .ZN(n9980) );
  NAND2_X1 U8719 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  OAI21_X1 U8720 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9979), .ZN(n9977) );
  NAND2_X1 U8721 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  OAI21_X1 U8722 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9976), .ZN(n9974) );
  NAND2_X1 U8723 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  OAI21_X1 U8724 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9973), .ZN(n9970) );
  NAND2_X1 U8725 ( .A1(n9969), .A2(n9970), .ZN(n6863) );
  NOR2_X1 U8726 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  AOI21_X1 U8727 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6863), .A(n9968), .ZN(
        n6867) );
  NOR2_X1 U8728 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  XNOR2_X1 U8729 ( .A(n6867), .B(n6866), .ZN(ADD_1068_U4) );
  NAND2_X1 U8730 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  XNOR2_X1 U8731 ( .A(n7843), .B(n6870), .ZN(n9904) );
  NAND2_X1 U8732 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  XOR2_X1 U8733 ( .A(n7843), .B(n6873), .Z(n6874) );
  AOI222_X1 U8734 ( .A1(n8433), .A2(n6874), .B1(n8194), .B2(n9869), .C1(n8196), 
        .C2(n9866), .ZN(n9905) );
  MUX2_X1 U8735 ( .A(n7406), .B(n9905), .S(n9876), .Z(n6877) );
  INV_X1 U8736 ( .A(n6940), .ZN(n6875) );
  AOI22_X1 U8737 ( .A1(n8438), .A2(n6948), .B1(n8437), .B2(n6875), .ZN(n6876)
         );
  OAI211_X1 U8738 ( .C1(n8441), .C2(n9904), .A(n6877), .B(n6876), .ZN(P2_U3227) );
  INV_X1 U8739 ( .A(n6878), .ZN(n6922) );
  AOI22_X1 U8740 ( .A1(n9147), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10045), .ZN(n6879) );
  OAI21_X1 U8741 ( .B1(n6922), .B2(n9476), .A(n6879), .ZN(P1_U3338) );
  XNOR2_X1 U8742 ( .A(n6880), .B(n7849), .ZN(n6882) );
  OAI22_X1 U8743 ( .A1(n7305), .A2(n8396), .B1(n7476), .B2(n8394), .ZN(n6881)
         );
  AOI21_X1 U8744 ( .B1(n6882), .B2(n8433), .A(n6881), .ZN(n9931) );
  OAI22_X1 U8745 ( .A1(n8413), .A2(n7415), .B1(n7308), .B2(n9863), .ZN(n6883)
         );
  AOI21_X1 U8746 ( .B1(n9925), .B2(n8438), .A(n6883), .ZN(n6888) );
  NAND2_X1 U8747 ( .A1(n6884), .A2(n7849), .ZN(n6885) );
  NAND2_X1 U8748 ( .A1(n6886), .A2(n6885), .ZN(n9928) );
  INV_X1 U8749 ( .A(n8441), .ZN(n8405) );
  NAND2_X1 U8750 ( .A1(n9928), .A2(n8405), .ZN(n6887) );
  OAI211_X1 U8751 ( .C1(n9931), .C2(n6677), .A(n6888), .B(n6887), .ZN(P2_U3223) );
  OAI21_X1 U8752 ( .B1(n6890), .B2(n6896), .A(n6889), .ZN(n7144) );
  AOI21_X1 U8753 ( .B1(n6891), .B2(n6964), .A(n9317), .ZN(n6892) );
  AND2_X1 U8754 ( .A1(n6892), .A2(n7345), .ZN(n7151) );
  INV_X1 U8755 ( .A(n8916), .ZN(n6895) );
  INV_X1 U8756 ( .A(n6893), .ZN(n6894) );
  AOI21_X1 U8757 ( .B1(n6895), .B2(n4812), .A(n6894), .ZN(n6897) );
  NOR2_X1 U8758 ( .A1(n6897), .A2(n6896), .ZN(n7338) );
  AOI21_X1 U8759 ( .B1(n6897), .B2(n6896), .A(n7338), .ZN(n6900) );
  OAI22_X1 U8760 ( .A1(n6980), .A2(n8798), .B1(n6898), .B2(n8800), .ZN(n6972)
         );
  INV_X1 U8761 ( .A(n6972), .ZN(n6899) );
  OAI21_X1 U8762 ( .B1(n6900), .B2(n9314), .A(n6899), .ZN(n7145) );
  AOI211_X1 U8763 ( .C1(n9673), .C2(n7144), .A(n7151), .B(n7145), .ZN(n6906)
         );
  INV_X1 U8764 ( .A(n6964), .ZN(n7149) );
  OAI22_X1 U8765 ( .A1(n7149), .A2(n9387), .B1(n9678), .B2(n5871), .ZN(n6901)
         );
  INV_X1 U8766 ( .A(n6901), .ZN(n6902) );
  OAI21_X1 U8767 ( .B1(n6906), .B2(n9676), .A(n6902), .ZN(P1_U3530) );
  INV_X1 U8768 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6903) );
  OAI22_X1 U8769 ( .A1(n7149), .A2(n9442), .B1(n9464), .B2(n6903), .ZN(n6904)
         );
  INV_X1 U8770 ( .A(n6904), .ZN(n6905) );
  OAI21_X1 U8771 ( .B1(n6906), .B2(n9674), .A(n6905), .ZN(P1_U3477) );
  XNOR2_X1 U8772 ( .A(n6908), .B(n6907), .ZN(n7695) );
  NAND2_X1 U8773 ( .A1(n7695), .A2(n7696), .ZN(n7694) );
  OAI21_X1 U8774 ( .B1(n6909), .B2(n6908), .A(n7694), .ZN(n6914) );
  OAI21_X1 U8775 ( .B1(n6912), .B2(n6911), .A(n6910), .ZN(n6913) );
  XNOR2_X1 U8776 ( .A(n6914), .B(n6913), .ZN(n6920) );
  AOI22_X1 U8777 ( .A1(n6915), .A2(n8805), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6916) );
  OAI21_X1 U8778 ( .B1(n7110), .B2(n8803), .A(n6916), .ZN(n6917) );
  AOI21_X1 U8779 ( .B1(n6918), .B2(n8790), .A(n6917), .ZN(n6919) );
  OAI21_X1 U8780 ( .B1(n6920), .B2(n8792), .A(n6919), .ZN(P1_U3239) );
  INV_X1 U8781 ( .A(n9843), .ZN(n8244) );
  OAI222_X1 U8782 ( .A1(n8562), .A2(n6922), .B1(n8244), .B2(P2_U3151), .C1(
        n6921), .C2(n8555), .ZN(P2_U3278) );
  INV_X1 U8783 ( .A(n6923), .ZN(n6975) );
  AOI22_X1 U8784 ( .A1(n9613), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10045), .ZN(n6924) );
  OAI21_X1 U8785 ( .B1(n6975), .B2(n9476), .A(n6924), .ZN(P1_U3337) );
  INV_X1 U8786 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6935) );
  INV_X1 U8787 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U8788 ( .A1(n6925), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6928) );
  INV_X1 U8789 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8443) );
  OR2_X1 U8790 ( .A1(n6926), .A2(n8443), .ZN(n6927) );
  OAI211_X1 U8791 ( .C1(n6929), .C2(n8276), .A(n6928), .B(n6927), .ZN(n6930)
         );
  INV_X1 U8792 ( .A(n6930), .ZN(n6931) );
  INV_X1 U8793 ( .A(n8273), .ZN(n6933) );
  NAND2_X1 U8794 ( .A1(n6933), .A2(P2_U3893), .ZN(n6934) );
  OAI21_X1 U8795 ( .B1(P2_U3893), .B2(n6935), .A(n6934), .ZN(P2_U3522) );
  AOI21_X1 U8796 ( .B1(n8172), .B2(n8196), .A(n6936), .ZN(n6939) );
  OR2_X1 U8797 ( .A1(n8170), .A2(n6937), .ZN(n6938) );
  OAI211_X1 U8798 ( .C1(n8174), .C2(n6940), .A(n6939), .B(n6938), .ZN(n6947)
         );
  XNOR2_X1 U8799 ( .A(n7735), .B(n9906), .ZN(n6951) );
  XNOR2_X1 U8800 ( .A(n8195), .B(n6951), .ZN(n6945) );
  OAI22_X1 U8801 ( .A1(n6943), .A2(n6942), .B1(n6941), .B2(n8196), .ZN(n6944)
         );
  AOI211_X1 U8802 ( .C1(n6945), .C2(n6944), .A(n8177), .B(n6950), .ZN(n6946)
         );
  AOI211_X1 U8803 ( .C1(n6948), .C2(n8182), .A(n6947), .B(n6946), .ZN(n6949)
         );
  INV_X1 U8804 ( .A(n6949), .ZN(P2_U3179) );
  INV_X1 U8805 ( .A(n6952), .ZN(n9910) );
  AOI21_X1 U8806 ( .B1(n6951), .B2(n8195), .A(n6950), .ZN(n6954) );
  XNOR2_X1 U8807 ( .A(n6952), .B(n7735), .ZN(n7004) );
  XNOR2_X1 U8808 ( .A(n7004), .B(n8194), .ZN(n6953) );
  NAND2_X1 U8809 ( .A1(n6954), .A2(n6953), .ZN(n7005) );
  OAI21_X1 U8810 ( .B1(n6954), .B2(n6953), .A(n7005), .ZN(n6955) );
  NAND2_X1 U8811 ( .A1(n6955), .A2(n8160), .ZN(n6960) );
  AND2_X1 U8812 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9714) );
  AOI21_X1 U8813 ( .B1(n8172), .B2(n8195), .A(n9714), .ZN(n6956) );
  OAI21_X1 U8814 ( .B1(n7055), .B2(n8170), .A(n6956), .ZN(n6957) );
  AOI21_X1 U8815 ( .B1(n6958), .B2(n8164), .A(n6957), .ZN(n6959) );
  OAI211_X1 U8816 ( .C1(n9910), .C2(n8167), .A(n6960), .B(n6959), .ZN(P2_U3153) );
  AOI22_X1 U8817 ( .A1(n9068), .A2(n8635), .B1(n6964), .B2(n6773), .ZN(n6969)
         );
  INV_X1 U8818 ( .A(n6961), .ZN(n6962) );
  NAND2_X1 U8819 ( .A1(n6963), .A2(n6962), .ZN(n6992) );
  NAND2_X1 U8820 ( .A1(n6964), .A2(n4574), .ZN(n6965) );
  OAI21_X1 U8821 ( .B1(n6966), .B2(n8629), .A(n6965), .ZN(n6967) );
  XNOR2_X1 U8822 ( .A(n6967), .B(n6422), .ZN(n6990) );
  XNOR2_X1 U8823 ( .A(n6992), .B(n6990), .ZN(n6968) );
  NAND2_X1 U8824 ( .A1(n6968), .A2(n6969), .ZN(n6997) );
  OAI21_X1 U8825 ( .B1(n6969), .B2(n6968), .A(n6997), .ZN(n6970) );
  NAND2_X1 U8826 ( .A1(n6970), .A2(n8797), .ZN(n6974) );
  NOR2_X1 U8827 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5872), .ZN(n9516) );
  NOR2_X1 U8828 ( .A1(n8803), .A2(n7146), .ZN(n6971) );
  AOI211_X1 U8829 ( .C1(n8805), .C2(n6972), .A(n9516), .B(n6971), .ZN(n6973)
         );
  OAI211_X1 U8830 ( .C1(n7149), .C2(n8807), .A(n6974), .B(n6973), .ZN(P1_U3221) );
  INV_X1 U8831 ( .A(n8262), .ZN(n8252) );
  OAI222_X1 U8832 ( .A1(n8555), .A2(n6976), .B1(n8252), .B2(P2_U3151), .C1(
        n8562), .C2(n6975), .ZN(P2_U3277) );
  OAI21_X1 U8833 ( .B1(n6978), .B2(n8851), .A(n6977), .ZN(n7367) );
  INV_X1 U8834 ( .A(n7367), .ZN(n6989) );
  XNOR2_X1 U8835 ( .A(n6979), .B(n8851), .ZN(n6981) );
  OAI22_X1 U8836 ( .A1(n6980), .A2(n8800), .B1(n7227), .B2(n8798), .ZN(n7130)
         );
  AOI21_X1 U8837 ( .B1(n6981), .B2(n9329), .A(n7130), .ZN(n7376) );
  INV_X1 U8838 ( .A(n6982), .ZN(n7032) );
  OAI211_X1 U8839 ( .C1(n7128), .C2(n6983), .A(n7032), .B(n9342), .ZN(n7370)
         );
  NAND2_X1 U8840 ( .A1(n7376), .A2(n7370), .ZN(n6987) );
  OAI22_X1 U8841 ( .A1(n7128), .A2(n9387), .B1(n9678), .B2(n6485), .ZN(n6984)
         );
  AOI21_X1 U8842 ( .B1(n6987), .B2(n9678), .A(n6984), .ZN(n6985) );
  OAI21_X1 U8843 ( .B1(n6989), .B2(n9407), .A(n6985), .ZN(P1_U3532) );
  OAI22_X1 U8844 ( .A1(n7128), .A2(n9442), .B1(n9464), .B2(n5902), .ZN(n6986)
         );
  AOI21_X1 U8845 ( .B1(n6987), .B2(n9464), .A(n6986), .ZN(n6988) );
  OAI21_X1 U8846 ( .B1(n6989), .B2(n9462), .A(n6988), .ZN(P1_U3483) );
  INV_X1 U8847 ( .A(n6990), .ZN(n6991) );
  NAND2_X1 U8848 ( .A1(n6992), .A2(n6991), .ZN(n6996) );
  AND2_X1 U8849 ( .A1(n6997), .A2(n6996), .ZN(n6999) );
  NAND2_X1 U8850 ( .A1(n7352), .A2(n4574), .ZN(n6994) );
  NAND2_X1 U8851 ( .A1(n9067), .A2(n6773), .ZN(n6993) );
  NAND2_X1 U8852 ( .A1(n6994), .A2(n6993), .ZN(n6995) );
  XNOR2_X1 U8853 ( .A(n6995), .B(n6466), .ZN(n7117) );
  AOI22_X1 U8854 ( .A1(n7352), .A2(n6773), .B1(n9067), .B2(n8635), .ZN(n7118)
         );
  XNOR2_X1 U8855 ( .A(n7117), .B(n7118), .ZN(n6998) );
  OAI211_X1 U8856 ( .C1(n6999), .C2(n6998), .A(n8797), .B(n7125), .ZN(n7003)
         );
  INV_X1 U8857 ( .A(n8803), .ZN(n8767) );
  INV_X1 U8858 ( .A(n7349), .ZN(n7001) );
  NOR2_X1 U8859 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10200), .ZN(n9131) );
  NAND2_X1 U8860 ( .A1(n9066), .A2(n8784), .ZN(n7346) );
  NAND2_X1 U8861 ( .A1(n9068), .A2(n9042), .ZN(n7340) );
  AOI21_X1 U8862 ( .B1(n7346), .B2(n7340), .A(n8775), .ZN(n7000) );
  AOI211_X1 U8863 ( .C1(n8767), .C2(n7001), .A(n9131), .B(n7000), .ZN(n7002)
         );
  OAI211_X1 U8864 ( .C1(n5894), .C2(n8807), .A(n7003), .B(n7002), .ZN(P1_U3231) );
  XNOR2_X1 U8865 ( .A(n9917), .B(n7735), .ZN(n7047) );
  XNOR2_X1 U8866 ( .A(n7047), .B(n8193), .ZN(n7048) );
  XOR2_X1 U8867 ( .A(n7049), .B(n7048), .Z(n7012) );
  INV_X1 U8868 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7006) );
  NOR2_X1 U8869 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7006), .ZN(n9728) );
  AOI21_X1 U8870 ( .B1(n8172), .B2(n8194), .A(n9728), .ZN(n7008) );
  OR2_X1 U8871 ( .A1(n8170), .A2(n7305), .ZN(n7007) );
  OAI211_X1 U8872 ( .C1(n8174), .C2(n7009), .A(n7008), .B(n7007), .ZN(n7010)
         );
  AOI21_X1 U8873 ( .B1(n9917), .B2(n8182), .A(n7010), .ZN(n7011) );
  OAI21_X1 U8874 ( .B1(n7012), .B2(n8177), .A(n7011), .ZN(P2_U3161) );
  NAND2_X1 U8875 ( .A1(n7014), .A2(n7013), .ZN(n7016) );
  AND2_X1 U8876 ( .A1(n7016), .A2(n7015), .ZN(n7019) );
  INV_X1 U8877 ( .A(n7017), .ZN(n7018) );
  AOI21_X1 U8878 ( .B1(n7019), .B2(n7021), .A(n7018), .ZN(n9923) );
  INV_X1 U8879 ( .A(n9923), .ZN(n7028) );
  XNOR2_X1 U8880 ( .A(n7020), .B(n4673), .ZN(n7024) );
  NAND2_X1 U8881 ( .A1(n9923), .A2(n9927), .ZN(n7023) );
  AOI22_X1 U8882 ( .A1(n9866), .A2(n8193), .B1(n8192), .B2(n9869), .ZN(n7022)
         );
  OAI211_X1 U8883 ( .C1(n9873), .C2(n7024), .A(n7023), .B(n7022), .ZN(n9921)
         );
  NAND2_X1 U8884 ( .A1(n9921), .A2(n9876), .ZN(n7027) );
  OAI22_X1 U8885 ( .A1(n8413), .A2(n5227), .B1(n7054), .B2(n9863), .ZN(n7025)
         );
  AOI21_X1 U8886 ( .B1(n7050), .B2(n8438), .A(n7025), .ZN(n7026) );
  OAI211_X1 U8887 ( .C1(n7028), .C2(n8286), .A(n7027), .B(n7026), .ZN(P2_U3224) );
  OAI21_X1 U8888 ( .B1(n7030), .B2(n8849), .A(n7029), .ZN(n7156) );
  INV_X1 U8889 ( .A(n7031), .ZN(n7168) );
  AOI211_X1 U8890 ( .C1(n7229), .C2(n7032), .A(n9317), .B(n7168), .ZN(n7160)
         );
  INV_X1 U8891 ( .A(n7033), .ZN(n7034) );
  AOI211_X1 U8892 ( .C1(n8849), .C2(n7035), .A(n9314), .B(n7034), .ZN(n7036)
         );
  OAI22_X1 U8893 ( .A1(n7276), .A2(n8798), .B1(n7127), .B2(n8800), .ZN(n7243)
         );
  OR2_X1 U8894 ( .A1(n7036), .A2(n7243), .ZN(n7155) );
  AOI211_X1 U8895 ( .C1(n7156), .C2(n9673), .A(n7160), .B(n7155), .ZN(n7039)
         );
  AOI22_X1 U8896 ( .A1(n7229), .A2(n9405), .B1(n9676), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7037) );
  OAI21_X1 U8897 ( .B1(n7039), .B2(n9676), .A(n7037), .ZN(P1_U3533) );
  INV_X1 U8898 ( .A(n9442), .ZN(n9460) );
  AOI22_X1 U8899 ( .A1(n7229), .A2(n9460), .B1(n9674), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7038) );
  OAI21_X1 U8900 ( .B1(n7039), .B2(n9674), .A(n7038), .ZN(P1_U3486) );
  XNOR2_X1 U8901 ( .A(n7040), .B(n7929), .ZN(n9933) );
  XNOR2_X1 U8902 ( .A(n7041), .B(n7929), .ZN(n7042) );
  OAI222_X1 U8903 ( .A1(n8394), .A2(n7458), .B1(n8396), .B2(n7449), .C1(n9873), 
        .C2(n7042), .ZN(n9934) );
  NAND2_X1 U8904 ( .A1(n9934), .A2(n9876), .ZN(n7046) );
  OAI22_X1 U8905 ( .A1(n8413), .A2(n7043), .B1(n7402), .B2(n9863), .ZN(n7044)
         );
  AOI21_X1 U8906 ( .B1(n9936), .B2(n8438), .A(n7044), .ZN(n7045) );
  OAI211_X1 U8907 ( .C1(n9933), .C2(n8441), .A(n7046), .B(n7045), .ZN(P2_U3222) );
  INV_X1 U8908 ( .A(n7050), .ZN(n9920) );
  XNOR2_X1 U8909 ( .A(n7050), .B(n7735), .ZN(n7301) );
  XNOR2_X1 U8910 ( .A(n7301), .B(n7051), .ZN(n7052) );
  OAI211_X1 U8911 ( .C1(n7053), .C2(n7052), .A(n7303), .B(n8160), .ZN(n7060)
         );
  INV_X1 U8912 ( .A(n7054), .ZN(n7058) );
  OR2_X1 U8913 ( .A1(n8143), .A2(n7055), .ZN(n7056) );
  NAND2_X1 U8914 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3151), .ZN(n9758) );
  OAI211_X1 U8915 ( .C1(n8170), .C2(n7449), .A(n7056), .B(n9758), .ZN(n7057)
         );
  AOI21_X1 U8916 ( .B1(n8164), .B2(n7058), .A(n7057), .ZN(n7059) );
  OAI211_X1 U8917 ( .C1(n9920), .C2(n8167), .A(n7060), .B(n7059), .ZN(P2_U3171) );
  INV_X1 U8918 ( .A(n7061), .ZN(n7062) );
  OAI222_X1 U8919 ( .A1(n8265), .A2(P2_U3151), .B1(n8562), .B2(n7062), .C1(
        n8555), .C2(n5418), .ZN(P2_U3276) );
  OAI222_X1 U8920 ( .A1(n9478), .A2(n10110), .B1(n9476), .B2(n7062), .C1(
        P1_U3086), .C2(n4431), .ZN(P1_U3336) );
  INV_X1 U8921 ( .A(n7063), .ZN(n7079) );
  NAND2_X1 U8922 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  NAND2_X1 U8923 ( .A1(n7069), .A2(n7135), .ZN(n7070) );
  MUX2_X1 U8924 ( .A(n7071), .B(n10152), .S(n9321), .Z(n7078) );
  INV_X2 U8925 ( .A(n9624), .ZN(n9321) );
  INV_X1 U8926 ( .A(n7072), .ZN(n7076) );
  OAI22_X1 U8927 ( .A1(n9324), .A2(n7074), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9621), .ZN(n7075) );
  AOI21_X1 U8928 ( .B1(n9318), .B2(n7076), .A(n7075), .ZN(n7077) );
  OAI211_X1 U8929 ( .C1(n7079), .C2(n9328), .A(n7078), .B(n7077), .ZN(P1_U3290) );
  XNOR2_X1 U8930 ( .A(n7080), .B(n7930), .ZN(n7081) );
  OAI222_X1 U8931 ( .A1(n8394), .A2(n7568), .B1(n8396), .B2(n7476), .C1(n7081), 
        .C2(n9873), .ZN(n9940) );
  INV_X1 U8932 ( .A(n9940), .ZN(n7087) );
  OAI22_X1 U8933 ( .A1(n8413), .A2(n7082), .B1(n7479), .B2(n9863), .ZN(n7083)
         );
  AOI21_X1 U8934 ( .B1(n9942), .B2(n8438), .A(n7083), .ZN(n7086) );
  NAND2_X1 U8935 ( .A1(n7084), .A2(n7930), .ZN(n9937) );
  NAND3_X1 U8936 ( .A1(n9939), .A2(n9937), .A3(n8405), .ZN(n7085) );
  OAI211_X1 U8937 ( .C1(n7087), .C2(n6677), .A(n7086), .B(n7085), .ZN(P2_U3221) );
  INV_X1 U8938 ( .A(n9621), .ZN(n9319) );
  AOI21_X1 U8939 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9319), .A(n7088), .ZN(
        n7096) );
  INV_X1 U8940 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7089) );
  OAI22_X1 U8941 ( .A1(n9324), .A2(n7090), .B1(n9624), .B2(n7089), .ZN(n7091)
         );
  AOI21_X1 U8942 ( .B1(n7092), .B2(n9318), .A(n7091), .ZN(n7095) );
  NAND2_X1 U8943 ( .A1(n7093), .A2(n9338), .ZN(n7094) );
  OAI211_X1 U8944 ( .C1(n7096), .C2(n9321), .A(n7095), .B(n7094), .ZN(P1_U3291) );
  INV_X1 U8945 ( .A(n7097), .ZN(n7105) );
  MUX2_X1 U8946 ( .A(n6383), .B(n7098), .S(n9624), .Z(n7104) );
  INV_X1 U8947 ( .A(n7099), .ZN(n7102) );
  OAI22_X1 U8948 ( .A1(n9324), .A2(n7100), .B1(n9621), .B2(n8755), .ZN(n7101)
         );
  AOI21_X1 U8949 ( .B1(n7102), .B2(n9318), .A(n7101), .ZN(n7103) );
  OAI211_X1 U8950 ( .C1(n7105), .C2(n9328), .A(n7104), .B(n7103), .ZN(P1_U3289) );
  INV_X1 U8951 ( .A(n7106), .ZN(n7116) );
  INV_X1 U8952 ( .A(n7107), .ZN(n7108) );
  MUX2_X1 U8953 ( .A(n7109), .B(n7108), .S(n9624), .Z(n7115) );
  OAI22_X1 U8954 ( .A1(n9324), .A2(n7111), .B1(n9621), .B2(n7110), .ZN(n7112)
         );
  AOI21_X1 U8955 ( .B1(n7113), .B2(n9318), .A(n7112), .ZN(n7114) );
  OAI211_X1 U8956 ( .C1(n7116), .C2(n9328), .A(n7115), .B(n7114), .ZN(P1_U3287) );
  INV_X1 U8957 ( .A(n7117), .ZN(n7119) );
  OR2_X1 U8958 ( .A1(n7119), .A2(n7118), .ZN(n7123) );
  NAND2_X1 U8959 ( .A1(n7373), .A2(n4574), .ZN(n7121) );
  NAND2_X1 U8960 ( .A1(n9066), .A2(n6773), .ZN(n7120) );
  NAND2_X1 U8961 ( .A1(n7121), .A2(n7120), .ZN(n7122) );
  XNOR2_X1 U8962 ( .A(n7122), .B(n8681), .ZN(n7124) );
  INV_X1 U8963 ( .A(n7235), .ZN(n7126) );
  NOR2_X1 U8964 ( .A1(n7234), .A2(n7126), .ZN(n7129) );
  OAI22_X1 U8965 ( .A1(n7128), .A2(n8629), .B1(n7127), .B2(n6361), .ZN(n7236)
         );
  XNOR2_X1 U8966 ( .A(n7129), .B(n7236), .ZN(n7134) );
  AOI22_X1 U8967 ( .A1(n7130), .A2(n8805), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7131) );
  OAI21_X1 U8968 ( .B1(n7368), .B2(n8803), .A(n7131), .ZN(n7132) );
  AOI21_X1 U8969 ( .B1(n7373), .B2(n8790), .A(n7132), .ZN(n7133) );
  OAI21_X1 U8970 ( .B1(n7134), .B2(n8792), .A(n7133), .ZN(P1_U3217) );
  NOR2_X1 U8971 ( .A1(n9321), .A2(n7135), .ZN(n9632) );
  INV_X1 U8972 ( .A(n9632), .ZN(n7142) );
  NAND2_X1 U8973 ( .A1(n7136), .A2(n9624), .ZN(n7141) );
  AOI22_X1 U8974 ( .A1(n9321), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9319), .ZN(n7137) );
  OAI21_X1 U8975 ( .B1(n9324), .B2(n8820), .A(n7137), .ZN(n7138) );
  AOI21_X1 U8976 ( .B1(n7139), .B2(n9318), .A(n7138), .ZN(n7140) );
  OAI211_X1 U8977 ( .C1(n7143), .C2(n7142), .A(n7141), .B(n7140), .ZN(P1_U3292) );
  INV_X1 U8978 ( .A(n7144), .ZN(n7154) );
  NAND2_X1 U8979 ( .A1(n7145), .A2(n9624), .ZN(n7153) );
  NOR2_X1 U8980 ( .A1(n9621), .A2(n7146), .ZN(n7147) );
  AOI21_X1 U8981 ( .B1(n9321), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7147), .ZN(
        n7148) );
  OAI21_X1 U8982 ( .B1(n9324), .B2(n7149), .A(n7148), .ZN(n7150) );
  AOI21_X1 U8983 ( .B1(n7151), .B2(n9318), .A(n7150), .ZN(n7152) );
  OAI211_X1 U8984 ( .C1(n7154), .C2(n9328), .A(n7153), .B(n7152), .ZN(P1_U3285) );
  INV_X1 U8985 ( .A(n7155), .ZN(n7163) );
  NAND2_X1 U8986 ( .A1(n7156), .A2(n9338), .ZN(n7162) );
  NOR2_X1 U8987 ( .A1(n7246), .A2(n9324), .ZN(n7159) );
  OAI22_X1 U8988 ( .A1(n9624), .A2(n7157), .B1(n7240), .B2(n9621), .ZN(n7158)
         );
  AOI211_X1 U8989 ( .C1(n7160), .C2(n9318), .A(n7159), .B(n7158), .ZN(n7161)
         );
  OAI211_X1 U8990 ( .C1(n9321), .C2(n7163), .A(n7162), .B(n7161), .ZN(P1_U3282) );
  OAI21_X1 U8991 ( .B1(n7165), .B2(n8867), .A(n7164), .ZN(n7357) );
  INV_X1 U8992 ( .A(n7357), .ZN(n7175) );
  XNOR2_X1 U8993 ( .A(n7166), .B(n8867), .ZN(n7167) );
  OAI22_X1 U8994 ( .A1(n7490), .A2(n8798), .B1(n7227), .B2(n8800), .ZN(n7287)
         );
  AOI21_X1 U8995 ( .B1(n7167), .B2(n9329), .A(n7287), .ZN(n7366) );
  INV_X1 U8996 ( .A(n7363), .ZN(n7290) );
  OAI211_X1 U8997 ( .C1(n7168), .C2(n7290), .A(n9342), .B(n7263), .ZN(n7360)
         );
  NAND2_X1 U8998 ( .A1(n7366), .A2(n7360), .ZN(n7173) );
  OAI22_X1 U8999 ( .A1(n7290), .A2(n9387), .B1(n9678), .B2(n7181), .ZN(n7169)
         );
  AOI21_X1 U9000 ( .B1(n7173), .B2(n9678), .A(n7169), .ZN(n7170) );
  OAI21_X1 U9001 ( .B1(n7175), .B2(n9407), .A(n7170), .ZN(P1_U3534) );
  INV_X1 U9002 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7171) );
  OAI22_X1 U9003 ( .A1(n7290), .A2(n9442), .B1(n9464), .B2(n7171), .ZN(n7172)
         );
  AOI21_X1 U9004 ( .B1(n7173), .B2(n9464), .A(n7172), .ZN(n7174) );
  OAI21_X1 U9005 ( .B1(n7175), .B2(n9462), .A(n7174), .ZN(P1_U3489) );
  NAND2_X1 U9006 ( .A1(n7178), .A2(n10046), .ZN(n7176) );
  OAI211_X1 U9007 ( .C1(n7177), .C2(n9478), .A(n7176), .B(n9034), .ZN(P1_U3335) );
  INV_X1 U9008 ( .A(n7178), .ZN(n7179) );
  OAI222_X1 U9009 ( .A1(n8555), .A2(n7180), .B1(n8562), .B2(n7179), .C1(
        P2_U3151), .C2(n8024), .ZN(P2_U3275) );
  INV_X1 U9010 ( .A(n9597), .ZN(n9609) );
  XNOR2_X1 U9011 ( .A(n9147), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U9012 ( .A1(n7195), .A2(n7181), .ZN(n7182) );
  NAND2_X1 U9013 ( .A1(n7183), .A2(n7182), .ZN(n9550) );
  INV_X1 U9014 ( .A(n9550), .ZN(n7185) );
  INV_X1 U9015 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7184) );
  XNOR2_X1 U9016 ( .A(n9553), .B(n7184), .ZN(n9548) );
  NAND2_X1 U9017 ( .A1(n7185), .A2(n9548), .ZN(n9552) );
  NAND2_X1 U9018 ( .A1(n9553), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7186) );
  AND2_X1 U9019 ( .A1(n9552), .A2(n7186), .ZN(n9569) );
  XNOR2_X1 U9020 ( .A(n9566), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9568) );
  NOR2_X1 U9021 ( .A1(n9569), .A2(n9568), .ZN(n9567) );
  AOI21_X1 U9022 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9566), .A(n9567), .ZN(
        n7187) );
  NOR2_X1 U9023 ( .A1(n7187), .A2(n7199), .ZN(n7188) );
  XNOR2_X1 U9024 ( .A(n7199), .B(n7187), .ZN(n9580) );
  NOR2_X1 U9025 ( .A1(n9579), .A2(n9580), .ZN(n9578) );
  NOR2_X1 U9026 ( .A1(n7188), .A2(n9578), .ZN(n9596) );
  XNOR2_X1 U9027 ( .A(n9599), .B(n7189), .ZN(n9595) );
  AOI22_X1 U9028 ( .A1(n9596), .A2(n9595), .B1(n7190), .B2(n7189), .ZN(n9149)
         );
  XOR2_X1 U9029 ( .A(n9148), .B(n9149), .Z(n7212) );
  OR2_X1 U9030 ( .A1(n9147), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U9031 ( .A1(n9147), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7191) );
  AND2_X1 U9032 ( .A1(n9141), .A2(n7191), .ZN(n7206) );
  NAND2_X1 U9033 ( .A1(n9553), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U9034 ( .B1(n9553), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7192), .ZN(
        n9544) );
  NAND2_X1 U9035 ( .A1(n7194), .A2(n7193), .ZN(n7197) );
  NAND2_X1 U9036 ( .A1(n7195), .A2(n7359), .ZN(n7196) );
  NAND2_X1 U9037 ( .A1(n7197), .A2(n7196), .ZN(n9543) );
  NOR2_X1 U9038 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  AOI21_X1 U9039 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9553), .A(n9545), .ZN(
        n9561) );
  NAND2_X1 U9040 ( .A1(n9566), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7198) );
  OAI21_X1 U9041 ( .B1(n9566), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7198), .ZN(
        n9562) );
  NOR2_X1 U9042 ( .A1(n9561), .A2(n9562), .ZN(n9563) );
  AOI21_X1 U9043 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9566), .A(n9563), .ZN(
        n7200) );
  NOR2_X1 U9044 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  INV_X1 U9045 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9583) );
  XOR2_X1 U9046 ( .A(n9587), .B(n7200), .Z(n9584) );
  NOR2_X1 U9047 ( .A1(n9583), .A2(n9584), .ZN(n9582) );
  NOR2_X1 U9048 ( .A1(n7201), .A2(n9582), .ZN(n9592) );
  INV_X1 U9049 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7604) );
  OR2_X1 U9050 ( .A1(n9599), .A2(n7604), .ZN(n7203) );
  NAND2_X1 U9051 ( .A1(n9599), .A2(n7604), .ZN(n7202) );
  AND2_X1 U9052 ( .A1(n7203), .A2(n7202), .ZN(n9591) );
  OR2_X1 U9053 ( .A1(n9592), .A2(n9591), .ZN(n9594) );
  NAND2_X1 U9054 ( .A1(n9599), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7204) );
  AND2_X1 U9055 ( .A1(n9594), .A2(n7204), .ZN(n7205) );
  NAND2_X1 U9056 ( .A1(n7205), .A2(n7206), .ZN(n9142) );
  OAI21_X1 U9057 ( .B1(n7206), .B2(n7205), .A(n9142), .ZN(n7207) );
  NAND2_X1 U9058 ( .A1(n7207), .A2(n9605), .ZN(n7211) );
  INV_X1 U9059 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7208) );
  NAND2_X1 U9060 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8733) );
  OAI21_X1 U9061 ( .B1(n9620), .B2(n7208), .A(n8733), .ZN(n7209) );
  AOI21_X1 U9062 ( .B1(n9147), .B2(n9612), .A(n7209), .ZN(n7210) );
  OAI211_X1 U9063 ( .C1(n9609), .C2(n7212), .A(n7211), .B(n7210), .ZN(P1_U3260) );
  XNOR2_X1 U9064 ( .A(n7213), .B(n7851), .ZN(n9520) );
  NAND2_X1 U9065 ( .A1(n7214), .A2(n7851), .ZN(n7215) );
  NAND3_X1 U9066 ( .A1(n7216), .A2(n8433), .A3(n7215), .ZN(n7218) );
  AOI22_X1 U9067 ( .A1(n8431), .A2(n9869), .B1(n9866), .B2(n8190), .ZN(n7217)
         );
  NAND2_X1 U9068 ( .A1(n7218), .A2(n7217), .ZN(n9522) );
  INV_X1 U9069 ( .A(n9523), .ZN(n7219) );
  NOR2_X1 U9070 ( .A1(n7219), .A2(n9864), .ZN(n7220) );
  OAI21_X1 U9071 ( .B1(n9522), .B2(n7220), .A(n8413), .ZN(n7223) );
  INV_X1 U9072 ( .A(n7465), .ZN(n7221) );
  AOI22_X1 U9073 ( .A1(n6677), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8437), .B2(
        n7221), .ZN(n7222) );
  OAI211_X1 U9074 ( .C1(n9520), .C2(n8441), .A(n7223), .B(n7222), .ZN(P2_U3220) );
  NAND2_X1 U9075 ( .A1(n7229), .A2(n4574), .ZN(n7225) );
  NAND2_X1 U9076 ( .A1(n9065), .A2(n6773), .ZN(n7224) );
  NAND2_X1 U9077 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  XNOR2_X1 U9078 ( .A(n7226), .B(n8681), .ZN(n7231) );
  INV_X1 U9079 ( .A(n7231), .ZN(n7233) );
  NOR2_X1 U9080 ( .A1(n7227), .A2(n6361), .ZN(n7228) );
  AOI21_X1 U9081 ( .B1(n7229), .B2(n6773), .A(n7228), .ZN(n7230) );
  INV_X1 U9082 ( .A(n7230), .ZN(n7232) );
  AND2_X1 U9083 ( .A1(n7231), .A2(n7230), .ZN(n7272) );
  AOI21_X1 U9084 ( .B1(n7233), .B2(n7232), .A(n7272), .ZN(n7238) );
  OAI21_X1 U9085 ( .B1(n7238), .B2(n7237), .A(n7283), .ZN(n7239) );
  NAND2_X1 U9086 ( .A1(n7239), .A2(n8797), .ZN(n7245) );
  NAND2_X1 U9087 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9540) );
  INV_X1 U9088 ( .A(n9540), .ZN(n7242) );
  NOR2_X1 U9089 ( .A1(n8803), .A2(n7240), .ZN(n7241) );
  AOI211_X1 U9090 ( .C1(n8805), .C2(n7243), .A(n7242), .B(n7241), .ZN(n7244)
         );
  OAI211_X1 U9091 ( .C1(n7246), .C2(n8807), .A(n7245), .B(n7244), .ZN(P1_U3236) );
  INV_X1 U9092 ( .A(n7247), .ZN(n7255) );
  NAND2_X1 U9093 ( .A1(n7248), .A2(n9318), .ZN(n7251) );
  INV_X1 U9094 ( .A(n7249), .ZN(n7701) );
  AOI22_X1 U9095 ( .A1(n9321), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7701), .B2(
        n9319), .ZN(n7250) );
  OAI211_X1 U9096 ( .C1(n7704), .C2(n9324), .A(n7251), .B(n7250), .ZN(n7252)
         );
  AOI21_X1 U9097 ( .B1(n7253), .B2(n9338), .A(n7252), .ZN(n7254) );
  OAI21_X1 U9098 ( .B1(n7255), .B2(n9321), .A(n7254), .ZN(P1_U3288) );
  OAI21_X1 U9099 ( .B1(n7257), .B2(n7258), .A(n7256), .ZN(n7297) );
  INV_X1 U9100 ( .A(n7297), .ZN(n7269) );
  INV_X1 U9101 ( .A(n7258), .ZN(n8869) );
  XNOR2_X1 U9102 ( .A(n7259), .B(n8869), .ZN(n7260) );
  NAND2_X1 U9103 ( .A1(n7260), .A2(n9329), .ZN(n7261) );
  AOI22_X1 U9104 ( .A1(n9064), .A2(n9042), .B1(n8784), .B2(n9062), .ZN(n7390)
         );
  NAND2_X1 U9105 ( .A1(n7261), .A2(n7390), .ZN(n7292) );
  INV_X1 U9106 ( .A(n7382), .ZN(n7395) );
  INV_X1 U9107 ( .A(n7494), .ZN(n7262) );
  AOI211_X1 U9108 ( .C1(n7382), .C2(n7263), .A(n9317), .B(n7262), .ZN(n7291)
         );
  NAND2_X1 U9109 ( .A1(n7291), .A2(n9318), .ZN(n7266) );
  INV_X1 U9110 ( .A(n7264), .ZN(n7392) );
  AOI22_X1 U9111 ( .A1(n9321), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7392), .B2(
        n9319), .ZN(n7265) );
  OAI211_X1 U9112 ( .C1(n7395), .C2(n9324), .A(n7266), .B(n7265), .ZN(n7267)
         );
  AOI21_X1 U9113 ( .B1(n7292), .B2(n9624), .A(n7267), .ZN(n7268) );
  OAI21_X1 U9114 ( .B1(n7269), .B2(n9328), .A(n7268), .ZN(P1_U3280) );
  INV_X1 U9115 ( .A(n7270), .ZN(n7312) );
  OAI222_X1 U9116 ( .A1(n8562), .A2(n7312), .B1(n7837), .B2(P2_U3151), .C1(
        n7271), .C2(n8555), .ZN(P2_U3274) );
  INV_X1 U9117 ( .A(n7272), .ZN(n7282) );
  NAND2_X1 U9118 ( .A1(n7363), .A2(n4574), .ZN(n7274) );
  NAND2_X1 U9119 ( .A1(n9064), .A2(n6773), .ZN(n7273) );
  NAND2_X1 U9120 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  XNOR2_X1 U9121 ( .A(n7275), .B(n8681), .ZN(n7279) );
  NOR2_X1 U9122 ( .A1(n7276), .A2(n6361), .ZN(n7277) );
  AOI21_X1 U9123 ( .B1(n7363), .B2(n6773), .A(n7277), .ZN(n7278) );
  NAND2_X1 U9124 ( .A1(n7279), .A2(n7278), .ZN(n7377) );
  OR2_X1 U9125 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  NAND2_X1 U9126 ( .A1(n7377), .A2(n7280), .ZN(n7281) );
  AND3_X1 U9127 ( .A1(n7283), .A2(n7282), .A3(n7281), .ZN(n7284) );
  OAI21_X1 U9128 ( .B1(n7388), .B2(n7284), .A(n8797), .ZN(n7289) );
  NOR2_X1 U9129 ( .A1(n8803), .A2(n7358), .ZN(n7285) );
  AOI211_X1 U9130 ( .C1(n8805), .C2(n7287), .A(n7286), .B(n7285), .ZN(n7288)
         );
  OAI211_X1 U9131 ( .C1(n7290), .C2(n8807), .A(n7289), .B(n7288), .ZN(P1_U3224) );
  NOR2_X1 U9132 ( .A1(n7292), .A2(n7291), .ZN(n7300) );
  NAND2_X1 U9133 ( .A1(n7297), .A2(n7293), .ZN(n7295) );
  AOI22_X1 U9134 ( .A1(n7382), .A2(n9405), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9676), .ZN(n7294) );
  OAI211_X1 U9135 ( .C1(n7300), .C2(n9676), .A(n7295), .B(n7294), .ZN(P1_U3535) );
  NAND2_X1 U9136 ( .A1(n7297), .A2(n7296), .ZN(n7299) );
  AOI22_X1 U9137 ( .A1(n7382), .A2(n9460), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9674), .ZN(n7298) );
  OAI211_X1 U9138 ( .C1(n7300), .C2(n9674), .A(n7299), .B(n7298), .ZN(P1_U3492) );
  XNOR2_X1 U9139 ( .A(n7457), .B(n8192), .ZN(n7396) );
  XNOR2_X1 U9140 ( .A(n9925), .B(n7726), .ZN(n7450) );
  INV_X1 U9141 ( .A(n7450), .ZN(n7452) );
  XNOR2_X1 U9142 ( .A(n7396), .B(n7452), .ZN(n7311) );
  INV_X1 U9143 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7304) );
  NOR2_X1 U9144 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7304), .ZN(n7442) );
  NOR2_X1 U9145 ( .A1(n8143), .A2(n7305), .ZN(n7306) );
  AOI211_X1 U9146 ( .C1(n8141), .C2(n8191), .A(n7442), .B(n7306), .ZN(n7307)
         );
  OAI21_X1 U9147 ( .B1(n7308), .B2(n8174), .A(n7307), .ZN(n7309) );
  AOI21_X1 U9148 ( .B1(n9925), .B2(n8182), .A(n7309), .ZN(n7310) );
  OAI21_X1 U9149 ( .B1(n7311), .B2(n8177), .A(n7310), .ZN(P2_U3157) );
  OAI222_X1 U9150 ( .A1(n9478), .A2(n7313), .B1(n9476), .B2(n7312), .C1(n9035), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  OAI21_X1 U9151 ( .B1(n9629), .B2(n9317), .A(n9324), .ZN(n7323) );
  OAI22_X1 U9152 ( .A1(n9624), .A2(n7315), .B1(n7314), .B2(n9621), .ZN(n7322)
         );
  NAND3_X1 U9153 ( .A1(n7318), .A2(n7317), .A3(n7316), .ZN(n7320) );
  AOI21_X1 U9154 ( .B1(n7320), .B2(n7319), .A(n9321), .ZN(n7321) );
  AOI211_X1 U9155 ( .C1(n7324), .C2(n7323), .A(n7322), .B(n7321), .ZN(n7325)
         );
  INV_X1 U9156 ( .A(n7325), .ZN(P1_U3293) );
  INV_X1 U9157 ( .A(n7853), .ZN(n7946) );
  XNOR2_X1 U9158 ( .A(n7326), .B(n7946), .ZN(n7472) );
  OAI21_X1 U9159 ( .B1(n7328), .B2(n7853), .A(n8433), .ZN(n7329) );
  OR2_X1 U9160 ( .A1(n7330), .A2(n7329), .ZN(n7332) );
  AOI22_X1 U9161 ( .A1(n8189), .A2(n9866), .B1(n9869), .B2(n8422), .ZN(n7331)
         );
  NAND2_X1 U9162 ( .A1(n7332), .A2(n7331), .ZN(n7471) );
  INV_X1 U9163 ( .A(n7570), .ZN(n7579) );
  NOR2_X1 U9164 ( .A1(n7579), .A2(n9864), .ZN(n7333) );
  OAI21_X1 U9165 ( .B1(n7471), .B2(n7333), .A(n8413), .ZN(n7336) );
  INV_X1 U9166 ( .A(n7334), .ZN(n7576) );
  AOI22_X1 U9167 ( .A1(n6677), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8437), .B2(
        n7576), .ZN(n7335) );
  OAI211_X1 U9168 ( .C1(n7472), .C2(n8441), .A(n7336), .B(n7335), .ZN(P2_U3219) );
  NOR2_X1 U9169 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
  XOR2_X1 U9170 ( .A(n7343), .B(n7339), .Z(n7341) );
  OAI21_X1 U9171 ( .B1(n7341), .B2(n9314), .A(n7340), .ZN(n9670) );
  INV_X1 U9172 ( .A(n9670), .ZN(n7356) );
  OAI21_X1 U9173 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n9672) );
  XNOR2_X1 U9174 ( .A(n7345), .B(n5894), .ZN(n7348) );
  INV_X1 U9175 ( .A(n7346), .ZN(n7347) );
  AOI21_X1 U9176 ( .B1(n7348), .B2(n9342), .A(n7347), .ZN(n9668) );
  OAI22_X1 U9177 ( .A1(n9624), .A2(n7350), .B1(n7349), .B2(n9621), .ZN(n7351)
         );
  AOI21_X1 U9178 ( .B1(n9627), .B2(n7352), .A(n7351), .ZN(n7353) );
  OAI21_X1 U9179 ( .B1(n9668), .B2(n9629), .A(n7353), .ZN(n7354) );
  AOI21_X1 U9180 ( .B1(n9672), .B2(n9338), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9181 ( .B1(n7356), .B2(n9321), .A(n7355), .ZN(P1_U3284) );
  NAND2_X1 U9182 ( .A1(n7357), .A2(n9338), .ZN(n7365) );
  OAI22_X1 U9183 ( .A1(n9624), .A2(n7359), .B1(n7358), .B2(n9621), .ZN(n7362)
         );
  NOR2_X1 U9184 ( .A1(n7360), .A2(n9629), .ZN(n7361) );
  AOI211_X1 U9185 ( .C1(n9627), .C2(n7363), .A(n7362), .B(n7361), .ZN(n7364)
         );
  OAI211_X1 U9186 ( .C1(n9321), .C2(n7366), .A(n7365), .B(n7364), .ZN(P1_U3281) );
  NAND2_X1 U9187 ( .A1(n7367), .A2(n9338), .ZN(n7375) );
  OAI22_X1 U9188 ( .A1(n9624), .A2(n7369), .B1(n7368), .B2(n9621), .ZN(n7372)
         );
  NOR2_X1 U9189 ( .A1(n7370), .A2(n9629), .ZN(n7371) );
  AOI211_X1 U9190 ( .C1(n9627), .C2(n7373), .A(n7372), .B(n7371), .ZN(n7374)
         );
  OAI211_X1 U9191 ( .C1(n9321), .C2(n7376), .A(n7375), .B(n7374), .ZN(P1_U3283) );
  INV_X1 U9192 ( .A(n7377), .ZN(n7387) );
  NAND2_X1 U9193 ( .A1(n7382), .A2(n4574), .ZN(n7379) );
  NAND2_X1 U9194 ( .A1(n9063), .A2(n6773), .ZN(n7378) );
  NAND2_X1 U9195 ( .A1(n7379), .A2(n7378), .ZN(n7380) );
  XNOR2_X1 U9196 ( .A(n7380), .B(n8681), .ZN(n7384) );
  NOR2_X1 U9197 ( .A1(n7490), .A2(n6361), .ZN(n7381) );
  AOI21_X1 U9198 ( .B1(n7382), .B2(n6773), .A(n7381), .ZN(n7383) );
  NAND2_X1 U9199 ( .A1(n7384), .A2(n7383), .ZN(n7527) );
  OR2_X1 U9200 ( .A1(n7384), .A2(n7383), .ZN(n7385) );
  AND2_X1 U9201 ( .A1(n7527), .A2(n7385), .ZN(n7386) );
  NOR3_X1 U9202 ( .A1(n7388), .A2(n7387), .A3(n7386), .ZN(n7389) );
  OAI21_X1 U9203 ( .B1(n4502), .B2(n7389), .A(n8797), .ZN(n7394) );
  NAND2_X1 U9204 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9558) );
  OAI21_X1 U9205 ( .B1(n7390), .B2(n8775), .A(n9558), .ZN(n7391) );
  AOI21_X1 U9206 ( .B1(n7392), .B2(n8767), .A(n7391), .ZN(n7393) );
  OAI211_X1 U9207 ( .C1(n7395), .C2(n8807), .A(n7394), .B(n7393), .ZN(P1_U3234) );
  OAI22_X1 U9208 ( .A1(n7396), .A2(n7450), .B1(n8192), .B2(n7457), .ZN(n7398)
         );
  XNOR2_X1 U9209 ( .A(n9936), .B(n7735), .ZN(n7453) );
  XNOR2_X1 U9210 ( .A(n7453), .B(n7476), .ZN(n7397) );
  XNOR2_X1 U9211 ( .A(n7398), .B(n7397), .ZN(n7405) );
  NAND2_X1 U9212 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9773) );
  INV_X1 U9213 ( .A(n9773), .ZN(n7400) );
  NOR2_X1 U9214 ( .A1(n8143), .A2(n7449), .ZN(n7399) );
  AOI211_X1 U9215 ( .C1(n8141), .C2(n8190), .A(n7400), .B(n7399), .ZN(n7401)
         );
  OAI21_X1 U9216 ( .B1(n7402), .B2(n8174), .A(n7401), .ZN(n7403) );
  AOI21_X1 U9217 ( .B1(n9936), .B2(n8182), .A(n7403), .ZN(n7404) );
  OAI21_X1 U9218 ( .B1(n7405), .B2(n8177), .A(n7404), .ZN(P2_U3176) );
  NOR2_X1 U9219 ( .A1(n7432), .A2(n7406), .ZN(n7407) );
  AND2_X1 U9220 ( .A1(n7409), .A2(n7433), .ZN(n7410) );
  MUX2_X1 U9221 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7412), .S(n9729), .Z(n9739)
         );
  NOR2_X1 U9222 ( .A1(n9746), .A2(n7413), .ZN(n7414) );
  NOR2_X1 U9223 ( .A1(n7414), .A2(n9754), .ZN(n7419) );
  OR2_X1 U9224 ( .A1(n7438), .A2(n7415), .ZN(n7617) );
  NAND2_X1 U9225 ( .A1(n7438), .A2(n7415), .ZN(n7416) );
  NAND2_X1 U9226 ( .A1(n7617), .A2(n7416), .ZN(n7418) );
  INV_X1 U9227 ( .A(n7618), .ZN(n7417) );
  AOI21_X1 U9228 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n7448) );
  INV_X1 U9229 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U9230 ( .A1(n7632), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7625) );
  INV_X1 U9231 ( .A(n7625), .ZN(n7420) );
  AOI21_X1 U9232 ( .B1(n7438), .B2(n9959), .A(n7420), .ZN(n7427) );
  AOI22_X1 U9233 ( .A1(n9729), .A2(n5202), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7428), .ZN(n9735) );
  OR2_X1 U9234 ( .A1(n7432), .A2(n6684), .ZN(n7421) );
  NAND2_X1 U9235 ( .A1(n7422), .A2(n7421), .ZN(n7423) );
  XNOR2_X1 U9236 ( .A(n7423), .B(n9715), .ZN(n9716) );
  OAI21_X1 U9237 ( .B1(n9729), .B2(n5202), .A(n9734), .ZN(n7424) );
  NAND2_X1 U9238 ( .A1(n7436), .A2(n7424), .ZN(n7425) );
  NAND2_X1 U9239 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n9748), .ZN(n9747) );
  NAND2_X1 U9240 ( .A1(n7425), .A2(n9747), .ZN(n7426) );
  NAND2_X1 U9241 ( .A1(n7426), .A2(n7427), .ZN(n7624) );
  OAI21_X1 U9242 ( .B1(n7427), .B2(n7426), .A(n7624), .ZN(n7446) );
  MUX2_X1 U9243 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8257), .Z(n7437) );
  XNOR2_X1 U9244 ( .A(n7437), .B(n9746), .ZN(n9751) );
  MUX2_X1 U9245 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8257), .Z(n7429) );
  OR2_X1 U9246 ( .A1(n7429), .A2(n7428), .ZN(n7435) );
  XNOR2_X1 U9247 ( .A(n7429), .B(n9729), .ZN(n9731) );
  MUX2_X1 U9248 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8257), .Z(n7434) );
  XOR2_X1 U9249 ( .A(n9715), .B(n7434), .Z(n9723) );
  NAND2_X1 U9250 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  OAI21_X1 U9251 ( .B1(n7437), .B2(n7436), .A(n9749), .ZN(n7440) );
  MUX2_X1 U9252 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8213), .Z(n7633) );
  XNOR2_X1 U9253 ( .A(n7633), .B(n7438), .ZN(n7439) );
  NAND2_X1 U9254 ( .A1(n7439), .A2(n7440), .ZN(n7634) );
  OAI21_X1 U9255 ( .B1(n7440), .B2(n7439), .A(n7634), .ZN(n7443) );
  INV_X1 U9256 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U9257 ( .A1(n9713), .A2(n10196), .ZN(n7441) );
  AOI211_X1 U9258 ( .C1(n9851), .C2(n7443), .A(n7442), .B(n7441), .ZN(n7444)
         );
  OAI21_X1 U9259 ( .B1(n7632), .B2(n9708), .A(n7444), .ZN(n7445) );
  AOI21_X1 U9260 ( .B1(n7446), .B2(n9852), .A(n7445), .ZN(n7447) );
  OAI21_X1 U9261 ( .B1(n7448), .B2(n9856), .A(n7447), .ZN(P2_U3192) );
  XNOR2_X1 U9262 ( .A(n9942), .B(n7735), .ZN(n7459) );
  INV_X1 U9263 ( .A(n7459), .ZN(n7460) );
  AOI22_X1 U9264 ( .A1(n7453), .A2(n7476), .B1(n7449), .B2(n7452), .ZN(n7456)
         );
  AOI21_X1 U9265 ( .B1(n7450), .B2(n8192), .A(n8191), .ZN(n7454) );
  NAND2_X1 U9266 ( .A1(n8191), .A2(n8192), .ZN(n7451) );
  OAI22_X1 U9267 ( .A1(n7454), .A2(n7453), .B1(n7452), .B2(n7451), .ZN(n7455)
         );
  XNOR2_X1 U9268 ( .A(n7459), .B(n7458), .ZN(n7482) );
  XOR2_X1 U9269 ( .A(n7735), .B(n9523), .Z(n7569) );
  XNOR2_X1 U9270 ( .A(n7569), .B(n8189), .ZN(n7461) );
  XNOR2_X1 U9271 ( .A(n4507), .B(n7461), .ZN(n7468) );
  AND2_X1 U9272 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7642) );
  NOR2_X1 U9273 ( .A1(n8170), .A2(n7462), .ZN(n7463) );
  AOI211_X1 U9274 ( .C1(n8172), .C2(n8190), .A(n7642), .B(n7463), .ZN(n7464)
         );
  OAI21_X1 U9275 ( .B1(n7465), .B2(n8174), .A(n7464), .ZN(n7466) );
  AOI21_X1 U9276 ( .B1(n9523), .B2(n8182), .A(n7466), .ZN(n7467) );
  OAI21_X1 U9277 ( .B1(n7468), .B2(n8177), .A(n7467), .ZN(P2_U3174) );
  MUX2_X1 U9278 ( .A(n7471), .B(P2_REG1_REG_14__SCAN_IN), .S(n5726), .Z(n7470)
         );
  OAI22_X1 U9279 ( .A1(n7472), .A2(n8479), .B1(n7579), .B2(n8471), .ZN(n7469)
         );
  OR2_X1 U9280 ( .A1(n7470), .A2(n7469), .ZN(P2_U3473) );
  MUX2_X1 U9281 ( .A(n7471), .B(P2_REG0_REG_14__SCAN_IN), .S(n9944), .Z(n7474)
         );
  INV_X1 U9282 ( .A(n9938), .ZN(n9932) );
  OAI22_X1 U9283 ( .A1(n7472), .A2(n8550), .B1(n7579), .B2(n8530), .ZN(n7473)
         );
  OR2_X1 U9284 ( .A1(n7474), .A2(n7473), .ZN(P2_U3432) );
  NOR2_X1 U9285 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7475), .ZN(n9785) );
  NOR2_X1 U9286 ( .A1(n8143), .A2(n7476), .ZN(n7477) );
  AOI211_X1 U9287 ( .C1(n8141), .C2(n8189), .A(n9785), .B(n7477), .ZN(n7478)
         );
  OAI21_X1 U9288 ( .B1(n7479), .B2(n8174), .A(n7478), .ZN(n7484) );
  AOI211_X1 U9289 ( .C1(n7482), .C2(n7480), .A(n8177), .B(n7481), .ZN(n7483)
         );
  AOI211_X1 U9290 ( .C1(n9942), .C2(n8182), .A(n7484), .B(n7483), .ZN(n7485)
         );
  INV_X1 U9291 ( .A(n7485), .ZN(P2_U3164) );
  XNOR2_X1 U9292 ( .A(n7486), .B(n8937), .ZN(n9408) );
  NAND2_X1 U9293 ( .A1(n7487), .A2(n8937), .ZN(n7488) );
  AOI21_X1 U9294 ( .B1(n7489), .B2(n7488), .A(n9314), .ZN(n7492) );
  OAI22_X1 U9295 ( .A1(n7491), .A2(n8798), .B1(n7490), .B2(n8800), .ZN(n7548)
         );
  AOI211_X1 U9296 ( .C1(n9408), .C2(n7493), .A(n7492), .B(n7548), .ZN(n9413)
         );
  AOI211_X1 U9297 ( .C1(n9410), .C2(n7494), .A(n9317), .B(n7506), .ZN(n9409)
         );
  NOR2_X1 U9298 ( .A1(n7530), .A2(n9324), .ZN(n7497) );
  OAI22_X1 U9299 ( .A1(n9624), .A2(n7495), .B1(n7550), .B2(n9621), .ZN(n7496)
         );
  AOI211_X1 U9300 ( .C1(n9409), .C2(n9318), .A(n7497), .B(n7496), .ZN(n7499)
         );
  NAND2_X1 U9301 ( .A1(n9408), .A2(n9632), .ZN(n7498) );
  OAI211_X1 U9302 ( .C1(n9413), .C2(n9321), .A(n7499), .B(n7498), .ZN(P1_U3279) );
  INV_X1 U9303 ( .A(n10047), .ZN(n7501) );
  OAI222_X1 U9304 ( .A1(n8555), .A2(n7502), .B1(n8562), .B2(n7501), .C1(
        P2_U3151), .C2(n7500), .ZN(P2_U3273) );
  XOR2_X1 U9305 ( .A(n8870), .B(n7503), .Z(n7520) );
  OAI211_X1 U9306 ( .C1(n8870), .C2(n7504), .A(n7555), .B(n9329), .ZN(n7505)
         );
  AOI22_X1 U9307 ( .A1(n9060), .A2(n8784), .B1(n9042), .B2(n9062), .ZN(n7538)
         );
  NAND2_X1 U9308 ( .A1(n7505), .A2(n7538), .ZN(n7514) );
  INV_X1 U9309 ( .A(n7506), .ZN(n7507) );
  AOI211_X1 U9310 ( .C1(n7541), .C2(n7507), .A(n9317), .B(n7561), .ZN(n7515)
         );
  NAND2_X1 U9311 ( .A1(n7515), .A2(n9318), .ZN(n7510) );
  INV_X1 U9312 ( .A(n7537), .ZN(n7508) );
  AOI22_X1 U9313 ( .A1(n9321), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7508), .B2(
        n9319), .ZN(n7509) );
  OAI211_X1 U9314 ( .C1(n7511), .C2(n9324), .A(n7510), .B(n7509), .ZN(n7512)
         );
  AOI21_X1 U9315 ( .B1(n7514), .B2(n9624), .A(n7512), .ZN(n7513) );
  OAI21_X1 U9316 ( .B1(n7520), .B2(n9328), .A(n7513), .ZN(P1_U3278) );
  INV_X1 U9317 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7516) );
  AOI211_X1 U9318 ( .C1(n9411), .C2(n7541), .A(n7515), .B(n7514), .ZN(n7518)
         );
  MUX2_X1 U9319 ( .A(n7516), .B(n7518), .S(n9464), .Z(n7517) );
  OAI21_X1 U9320 ( .B1(n7520), .B2(n9462), .A(n7517), .ZN(P1_U3498) );
  MUX2_X1 U9321 ( .A(n9579), .B(n7518), .S(n9678), .Z(n7519) );
  OAI21_X1 U9322 ( .B1(n7520), .B2(n9407), .A(n7519), .ZN(P1_U3537) );
  NAND2_X1 U9323 ( .A1(n7524), .A2(n7521), .ZN(n7523) );
  NAND2_X1 U9324 ( .A1(n7522), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8032) );
  OAI211_X1 U9325 ( .C1(n10258), .C2(n8555), .A(n7523), .B(n8032), .ZN(
        P2_U3272) );
  NAND2_X1 U9326 ( .A1(n7524), .A2(n10046), .ZN(n7525) );
  OR2_X1 U9327 ( .A1(n9036), .A2(P1_U3086), .ZN(n9044) );
  OAI211_X1 U9328 ( .C1(n7526), .C2(n9478), .A(n7525), .B(n9044), .ZN(P1_U3332) );
  AOI22_X1 U9329 ( .A1(n9410), .A2(n4574), .B1(n6773), .B2(n9062), .ZN(n7528)
         );
  XNOR2_X1 U9330 ( .A(n7528), .B(n6422), .ZN(n7532) );
  NAND2_X1 U9331 ( .A1(n7531), .A2(n7532), .ZN(n7544) );
  OAI22_X1 U9332 ( .A1(n7530), .A2(n8629), .B1(n7529), .B2(n6361), .ZN(n7547)
         );
  NAND2_X1 U9333 ( .A1(n7544), .A2(n7547), .ZN(n7535) );
  INV_X1 U9334 ( .A(n7531), .ZN(n7534) );
  INV_X1 U9335 ( .A(n7532), .ZN(n7533) );
  NAND2_X1 U9336 ( .A1(n7534), .A2(n7533), .ZN(n7545) );
  AOI22_X1 U9337 ( .A1(n7541), .A2(n4574), .B1(n6773), .B2(n9061), .ZN(n7536)
         );
  XNOR2_X1 U9338 ( .A(n7536), .B(n6466), .ZN(n8565) );
  AOI22_X1 U9339 ( .A1(n7541), .A2(n6773), .B1(n8635), .B2(n9061), .ZN(n8566)
         );
  NOR2_X1 U9340 ( .A1(n8803), .A2(n7537), .ZN(n7540) );
  OAI22_X1 U9341 ( .A1(n7538), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10272), .ZN(n7539) );
  AOI211_X1 U9342 ( .C1(n7541), .C2(n8790), .A(n7540), .B(n7539), .ZN(n7542)
         );
  OAI21_X1 U9343 ( .B1(n7543), .B2(n8792), .A(n7542), .ZN(P1_U3241) );
  NAND2_X1 U9344 ( .A1(n7545), .A2(n7544), .ZN(n7546) );
  XOR2_X1 U9345 ( .A(n7547), .B(n7546), .Z(n7553) );
  AOI22_X1 U9346 ( .A1(n7548), .A2(n8805), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7549) );
  OAI21_X1 U9347 ( .B1(n7550), .B2(n8803), .A(n7549), .ZN(n7551) );
  AOI21_X1 U9348 ( .B1(n9410), .B2(n8790), .A(n7551), .ZN(n7552) );
  OAI21_X1 U9349 ( .B1(n7553), .B2(n8792), .A(n7552), .ZN(P1_U3215) );
  XNOR2_X1 U9350 ( .A(n7554), .B(n8872), .ZN(n7602) );
  NAND2_X1 U9351 ( .A1(n7555), .A2(n8957), .ZN(n7556) );
  NAND2_X1 U9352 ( .A1(n7556), .A2(n8872), .ZN(n7557) );
  NAND2_X1 U9353 ( .A1(n7557), .A2(n7581), .ZN(n7560) );
  NAND2_X1 U9354 ( .A1(n9061), .A2(n9042), .ZN(n7559) );
  NAND2_X1 U9355 ( .A1(n9059), .A2(n8784), .ZN(n7558) );
  NAND2_X1 U9356 ( .A1(n7559), .A2(n7558), .ZN(n8722) );
  AOI21_X1 U9357 ( .B1(n7560), .B2(n9329), .A(n8722), .ZN(n7610) );
  OAI211_X1 U9358 ( .C1(n7562), .C2(n7561), .A(n4447), .B(n9342), .ZN(n7605)
         );
  NAND2_X1 U9359 ( .A1(n7610), .A2(n7605), .ZN(n7565) );
  MUX2_X1 U9360 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7565), .S(n9678), .Z(n7563)
         );
  AOI21_X1 U9361 ( .B1(n9405), .B2(n8726), .A(n7563), .ZN(n7564) );
  OAI21_X1 U9362 ( .B1(n7602), .B2(n9407), .A(n7564), .ZN(P1_U3538) );
  MUX2_X1 U9363 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n7565), .S(n9464), .Z(n7566)
         );
  AOI21_X1 U9364 ( .B1(n9460), .B2(n8726), .A(n7566), .ZN(n7567) );
  OAI21_X1 U9365 ( .B1(n7602), .B2(n9462), .A(n7567), .ZN(P1_U3501) );
  XNOR2_X1 U9366 ( .A(n7570), .B(n7735), .ZN(n7722) );
  XNOR2_X1 U9367 ( .A(n7722), .B(n8431), .ZN(n7571) );
  NAND2_X1 U9368 ( .A1(n7572), .A2(n7571), .ZN(n7724) );
  OAI21_X1 U9369 ( .B1(n7572), .B2(n7571), .A(n7724), .ZN(n7573) );
  NAND2_X1 U9370 ( .A1(n7573), .A2(n8160), .ZN(n7578) );
  AOI22_X1 U9371 ( .A1(n8172), .A2(n8189), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7574) );
  OAI21_X1 U9372 ( .B1(n8120), .B2(n8170), .A(n7574), .ZN(n7575) );
  AOI21_X1 U9373 ( .B1(n7576), .B2(n8164), .A(n7575), .ZN(n7577) );
  OAI211_X1 U9374 ( .C1(n7579), .C2(n8167), .A(n7578), .B(n7577), .ZN(P2_U3155) );
  INV_X1 U9375 ( .A(n7582), .ZN(n8964) );
  XNOR2_X1 U9376 ( .A(n7580), .B(n8964), .ZN(n7598) );
  AOI211_X1 U9377 ( .C1(n8575), .C2(n4447), .A(n9317), .B(n4499), .ZN(n7588)
         );
  INV_X1 U9378 ( .A(n7581), .ZN(n7583) );
  OAI21_X1 U9379 ( .B1(n7583), .B2(n8835), .A(n7582), .ZN(n7585) );
  NAND3_X1 U9380 ( .A1(n7585), .A2(n7584), .A3(n9329), .ZN(n7586) );
  AOI22_X1 U9381 ( .A1(n9060), .A2(n9042), .B1(n8784), .B2(n9058), .ZN(n8734)
         );
  NAND2_X1 U9382 ( .A1(n7586), .A2(n8734), .ZN(n7593) );
  AOI211_X1 U9383 ( .C1(n9411), .C2(n8575), .A(n7588), .B(n7593), .ZN(n7595)
         );
  MUX2_X1 U9384 ( .A(n10077), .B(n7595), .S(n9678), .Z(n7587) );
  OAI21_X1 U9385 ( .B1(n7598), .B2(n9407), .A(n7587), .ZN(P1_U3539) );
  NAND2_X1 U9386 ( .A1(n7588), .A2(n9318), .ZN(n7591) );
  INV_X1 U9387 ( .A(n7589), .ZN(n8736) );
  AOI22_X1 U9388 ( .A1(n9321), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8736), .B2(
        n9319), .ZN(n7590) );
  OAI211_X1 U9389 ( .C1(n8739), .C2(n9324), .A(n7591), .B(n7590), .ZN(n7592)
         );
  AOI21_X1 U9390 ( .B1(n7593), .B2(n9624), .A(n7592), .ZN(n7594) );
  OAI21_X1 U9391 ( .B1(n7598), .B2(n9328), .A(n7594), .ZN(P1_U3276) );
  INV_X1 U9392 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7596) );
  MUX2_X1 U9393 ( .A(n7596), .B(n7595), .S(n9464), .Z(n7597) );
  OAI21_X1 U9394 ( .B1(n7598), .B2(n9462), .A(n7597), .ZN(P1_U3504) );
  INV_X1 U9395 ( .A(n7599), .ZN(n7650) );
  OAI222_X1 U9396 ( .A1(P1_U3086), .A2(n7601), .B1(n9476), .B2(n7650), .C1(
        n7600), .C2(n9478), .ZN(P1_U3331) );
  INV_X1 U9397 ( .A(n7602), .ZN(n7603) );
  NAND2_X1 U9398 ( .A1(n7603), .A2(n9338), .ZN(n7609) );
  OAI22_X1 U9399 ( .A1(n9624), .A2(n7604), .B1(n8724), .B2(n9621), .ZN(n7607)
         );
  NOR2_X1 U9400 ( .A1(n7605), .A2(n9629), .ZN(n7606) );
  AOI211_X1 U9401 ( .C1(n9627), .C2(n8726), .A(n7607), .B(n7606), .ZN(n7608)
         );
  OAI211_X1 U9402 ( .C1(n9321), .C2(n7610), .A(n7609), .B(n7608), .ZN(P1_U3277) );
  INV_X1 U9403 ( .A(n6156), .ZN(n7613) );
  INV_X1 U9404 ( .A(n7611), .ZN(n7668) );
  OAI222_X1 U9405 ( .A1(P1_U3086), .A2(n7613), .B1(n9476), .B2(n7668), .C1(
        n7612), .C2(n9478), .ZN(P1_U3329) );
  INV_X1 U9406 ( .A(n7614), .ZN(n8034) );
  OAI222_X1 U9407 ( .A1(P1_U3086), .A2(n7616), .B1(n9476), .B2(n8034), .C1(
        n7615), .C2(n9478), .ZN(P1_U3330) );
  INV_X1 U9408 ( .A(n7620), .ZN(n7619) );
  NOR2_X1 U9409 ( .A1(n9761), .A2(n7619), .ZN(n7621) );
  NAND2_X1 U9410 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7637), .ZN(n7622) );
  OAI21_X1 U9411 ( .B1(n7637), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7622), .ZN(
        n9787) );
  AOI21_X1 U9412 ( .B1(n5306), .B2(n7623), .A(n8203), .ZN(n7648) );
  NAND2_X1 U9413 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7637), .ZN(n7628) );
  AOI22_X1 U9414 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7637), .B1(n9776), .B2(
        n5287), .ZN(n9779) );
  NAND2_X1 U9415 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U9416 ( .A1(n7630), .A2(n7626), .ZN(n7627) );
  XNOR2_X1 U9417 ( .A(n7626), .B(n9761), .ZN(n9763) );
  NAND2_X1 U9418 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9763), .ZN(n9762) );
  NAND2_X1 U9419 ( .A1(n7627), .A2(n9762), .ZN(n9778) );
  NAND2_X1 U9420 ( .A1(n9779), .A2(n9778), .ZN(n9777) );
  NAND2_X1 U9421 ( .A1(n7628), .A2(n9777), .ZN(n8235) );
  XNOR2_X1 U9422 ( .A(n8235), .B(n8202), .ZN(n7629) );
  NAND2_X1 U9423 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7629), .ZN(n8237) );
  OAI21_X1 U9424 ( .B1(n7629), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8237), .ZN(
        n7646) );
  MUX2_X1 U9425 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8257), .Z(n7638) );
  XNOR2_X1 U9426 ( .A(n7638), .B(n9776), .ZN(n9782) );
  MUX2_X1 U9427 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8257), .Z(n7631) );
  OR2_X1 U9428 ( .A1(n7631), .A2(n7630), .ZN(n7636) );
  XNOR2_X1 U9429 ( .A(n7631), .B(n9761), .ZN(n9766) );
  OR2_X1 U9430 ( .A1(n7633), .A2(n7632), .ZN(n7635) );
  NAND2_X1 U9431 ( .A1(n7635), .A2(n7634), .ZN(n9765) );
  NAND2_X1 U9432 ( .A1(n9766), .A2(n9765), .ZN(n9764) );
  NAND2_X1 U9433 ( .A1(n7636), .A2(n9764), .ZN(n9781) );
  NAND2_X1 U9434 ( .A1(n9782), .A2(n9781), .ZN(n9780) );
  OAI21_X1 U9435 ( .B1(n7638), .B2(n7637), .A(n9780), .ZN(n7640) );
  MUX2_X1 U9436 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8257), .Z(n8215) );
  XNOR2_X1 U9437 ( .A(n8215), .B(n8202), .ZN(n7639) );
  NAND2_X1 U9438 ( .A1(n7639), .A2(n7640), .ZN(n8216) );
  OAI21_X1 U9439 ( .B1(n7640), .B2(n7639), .A(n8216), .ZN(n7643) );
  INV_X1 U9440 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U9441 ( .A1(n9713), .A2(n10228), .ZN(n7641) );
  AOI211_X1 U9442 ( .C1(n9851), .C2(n7643), .A(n7642), .B(n7641), .ZN(n7644)
         );
  OAI21_X1 U9443 ( .B1(n8236), .B2(n9708), .A(n7644), .ZN(n7645) );
  AOI21_X1 U9444 ( .B1(n7646), .B2(n9852), .A(n7645), .ZN(n7647) );
  OAI21_X1 U9445 ( .B1(n7648), .B2(n9856), .A(n7647), .ZN(P2_U3195) );
  INV_X1 U9446 ( .A(n7681), .ZN(n9475) );
  OAI222_X1 U9447 ( .A1(n8562), .A2(n9475), .B1(n7652), .B2(P2_U3151), .C1(
        n7651), .C2(n8555), .ZN(P2_U3266) );
  INV_X1 U9448 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7824) );
  INV_X1 U9449 ( .A(SI_29_), .ZN(n7653) );
  OR2_X1 U9450 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  MUX2_X1 U9451 ( .A(n10213), .B(n7824), .S(n7671), .Z(n7659) );
  INV_X1 U9452 ( .A(SI_30_), .ZN(n7658) );
  NAND2_X1 U9453 ( .A1(n7659), .A2(n7658), .ZN(n7669) );
  INV_X1 U9454 ( .A(n7659), .ZN(n7660) );
  NAND2_X1 U9455 ( .A1(n7660), .A2(SI_30_), .ZN(n7661) );
  NAND2_X1 U9456 ( .A1(n7669), .A2(n7661), .ZN(n7662) );
  NAND2_X1 U9457 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  NAND2_X1 U9458 ( .A1(n7670), .A2(n7664), .ZN(n7823) );
  INV_X1 U9459 ( .A(n7823), .ZN(n9473) );
  OAI222_X1 U9460 ( .A1(n8555), .A2(n7824), .B1(n8562), .B2(n9473), .C1(
        P2_U3151), .C2(n7665), .ZN(P2_U3265) );
  OAI222_X1 U9461 ( .A1(n8562), .A2(n7668), .B1(P2_U3151), .B2(n7667), .C1(
        n7666), .C2(n8555), .ZN(P2_U3269) );
  NAND2_X1 U9462 ( .A1(n7670), .A2(n7669), .ZN(n7675) );
  MUX2_X1 U9463 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7671), .Z(n7673) );
  INV_X1 U9464 ( .A(SI_31_), .ZN(n7672) );
  XNOR2_X1 U9465 ( .A(n7673), .B(n7672), .ZN(n7674) );
  MUX2_X1 U9466 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8552), .S(n7676), .Z(n7678) );
  NAND2_X1 U9467 ( .A1(n7823), .A2(n5855), .ZN(n7680) );
  OR2_X1 U9468 ( .A1(n7682), .A2(n10213), .ZN(n7679) );
  NAND2_X1 U9469 ( .A1(n7681), .A2(n5855), .ZN(n7684) );
  OR2_X1 U9470 ( .A1(n7682), .A2(n9477), .ZN(n7683) );
  INV_X1 U9471 ( .A(n7719), .ZN(n9174) );
  NAND2_X1 U9472 ( .A1(n5007), .A2(n9342), .ZN(n7691) );
  INV_X1 U9473 ( .A(P1_B_REG_SCAN_IN), .ZN(n10053) );
  NOR2_X1 U9474 ( .A1(n7819), .A2(n10053), .ZN(n7685) );
  NOR2_X1 U9475 ( .A1(n8798), .A2(n7685), .ZN(n7717) );
  INV_X1 U9476 ( .A(n7717), .ZN(n7686) );
  INV_X1 U9477 ( .A(n9352), .ZN(n7687) );
  NAND2_X1 U9478 ( .A1(n7687), .A2(n9624), .ZN(n9165) );
  NAND2_X1 U9479 ( .A1(n9321), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9480 ( .A1(n9165), .A2(n7688), .ZN(n7689) );
  AOI21_X1 U9481 ( .B1(n8844), .B2(n9627), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9482 ( .B1(n7691), .B2(n9629), .A(n7690), .ZN(P1_U3263) );
  INV_X1 U9483 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7692) );
  MUX2_X1 U9484 ( .A(n7692), .B(n9349), .S(n9464), .Z(n7693) );
  OAI21_X1 U9485 ( .B1(n4685), .B2(n9442), .A(n7693), .ZN(P1_U3521) );
  OAI21_X1 U9486 ( .B1(n7696), .B2(n7695), .A(n7694), .ZN(n7697) );
  NAND2_X1 U9487 ( .A1(n7697), .A2(n8797), .ZN(n7703) );
  OAI22_X1 U9488 ( .A1(n7699), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7698), .ZN(n7700) );
  AOI21_X1 U9489 ( .B1(n7701), .B2(n8767), .A(n7700), .ZN(n7702) );
  OAI211_X1 U9490 ( .C1(n7704), .C2(n8807), .A(n7703), .B(n7702), .ZN(P1_U3227) );
  OAI21_X1 U9491 ( .B1(n7705), .B2(n8684), .A(n4450), .ZN(n7707) );
  NAND2_X1 U9492 ( .A1(n7719), .A2(n7706), .ZN(n9017) );
  NAND2_X1 U9493 ( .A1(n9016), .A2(n9017), .ZN(n9014) );
  XNOR2_X1 U9494 ( .A(n7707), .B(n9014), .ZN(n9178) );
  AOI211_X1 U9495 ( .C1(n7708), .C2(n7719), .A(n9317), .B(n9162), .ZN(n9169)
         );
  NAND2_X1 U9496 ( .A1(n7710), .A2(n8809), .ZN(n7712) );
  INV_X1 U9497 ( .A(n9014), .ZN(n7711) );
  NAND2_X1 U9498 ( .A1(n5804), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U9499 ( .A1(n7713), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U9500 ( .A1(n6293), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7714) );
  NAND3_X1 U9501 ( .A1(n7716), .A2(n7715), .A3(n7714), .ZN(n9049) );
  AOI22_X1 U9502 ( .A1(n9050), .A2(n9042), .B1(n7717), .B2(n9049), .ZN(n7718)
         );
  MUX2_X1 U9503 ( .A(n7720), .B(n7790), .S(n9464), .Z(n7721) );
  OAI21_X1 U9504 ( .B1(n9178), .B2(n9462), .A(n7721), .ZN(P1_U3519) );
  NAND2_X1 U9505 ( .A1(n7722), .A2(n7462), .ZN(n7723) );
  NAND2_X1 U9506 ( .A1(n7724), .A2(n7723), .ZN(n8178) );
  XNOR2_X1 U9507 ( .A(n8547), .B(n7735), .ZN(n7728) );
  XNOR2_X1 U9508 ( .A(n7728), .B(n8120), .ZN(n8179) );
  INV_X1 U9509 ( .A(n8179), .ZN(n7725) );
  XNOR2_X1 U9510 ( .A(n8540), .B(n7726), .ZN(n7727) );
  NOR2_X1 U9511 ( .A1(n7727), .A2(n8430), .ZN(n8126) );
  AOI21_X1 U9512 ( .B1(n7727), .B2(n8430), .A(n8126), .ZN(n8115) );
  INV_X1 U9513 ( .A(n7728), .ZN(n7729) );
  NAND2_X1 U9514 ( .A1(n7729), .A2(n8422), .ZN(n8116) );
  XNOR2_X1 U9515 ( .A(n8534), .B(n7735), .ZN(n7731) );
  NAND2_X1 U9516 ( .A1(n7731), .A2(n8395), .ZN(n8147) );
  INV_X1 U9517 ( .A(n7731), .ZN(n7732) );
  INV_X1 U9518 ( .A(n8395), .ZN(n8421) );
  NAND2_X1 U9519 ( .A1(n7732), .A2(n8421), .ZN(n7733) );
  AND2_X1 U9520 ( .A1(n8147), .A2(n7733), .ZN(n8125) );
  NAND2_X1 U9521 ( .A1(n7734), .A2(n8125), .ZN(n8127) );
  NAND2_X1 U9522 ( .A1(n8127), .A2(n8147), .ZN(n7739) );
  XNOR2_X1 U9523 ( .A(n8531), .B(n7726), .ZN(n7736) );
  NAND2_X1 U9524 ( .A1(n7736), .A2(n8382), .ZN(n8082) );
  INV_X1 U9525 ( .A(n7736), .ZN(n7737) );
  NAND2_X1 U9526 ( .A1(n7737), .A2(n8411), .ZN(n7738) );
  AND2_X1 U9527 ( .A1(n8082), .A2(n7738), .ZN(n8148) );
  NAND2_X1 U9528 ( .A1(n7739), .A2(n8148), .ZN(n8081) );
  NAND2_X1 U9529 ( .A1(n8081), .A2(n8082), .ZN(n7743) );
  XNOR2_X1 U9530 ( .A(n8523), .B(n4432), .ZN(n7740) );
  NAND2_X1 U9531 ( .A1(n7740), .A2(n8393), .ZN(n8135) );
  INV_X1 U9532 ( .A(n7740), .ZN(n7741) );
  NAND2_X1 U9533 ( .A1(n7741), .A2(n8372), .ZN(n7742) );
  AND2_X1 U9534 ( .A1(n8135), .A2(n7742), .ZN(n8083) );
  NAND2_X1 U9535 ( .A1(n7743), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U9536 ( .A1(n8085), .A2(n8135), .ZN(n7802) );
  XNOR2_X1 U9537 ( .A(n8518), .B(n7735), .ZN(n7744) );
  NAND2_X1 U9538 ( .A1(n7744), .A2(n8383), .ZN(n7803) );
  INV_X1 U9539 ( .A(n7744), .ZN(n7745) );
  NAND2_X1 U9540 ( .A1(n7745), .A2(n8360), .ZN(n7746) );
  XNOR2_X1 U9541 ( .A(n8513), .B(n4432), .ZN(n7747) );
  NAND2_X1 U9542 ( .A1(n7747), .A2(n7796), .ZN(n7805) );
  INV_X1 U9543 ( .A(n7747), .ZN(n7748) );
  NAND2_X1 U9544 ( .A1(n7748), .A2(n5471), .ZN(n7749) );
  XNOR2_X1 U9545 ( .A(n8350), .B(n7735), .ZN(n7755) );
  XNOR2_X1 U9546 ( .A(n7755), .B(n7750), .ZN(n7753) );
  AND2_X1 U9547 ( .A1(n8093), .A2(n7753), .ZN(n7752) );
  AND2_X1 U9548 ( .A1(n8136), .A2(n7752), .ZN(n7751) );
  NAND2_X1 U9549 ( .A1(n7802), .A2(n7751), .ZN(n7808) );
  INV_X1 U9550 ( .A(n7803), .ZN(n8094) );
  NAND2_X1 U9551 ( .A1(n7752), .A2(n8094), .ZN(n7809) );
  INV_X1 U9552 ( .A(n7753), .ZN(n7806) );
  NOR2_X1 U9553 ( .A1(n7806), .A2(n7805), .ZN(n7810) );
  INV_X1 U9554 ( .A(n7810), .ZN(n7754) );
  NAND2_X1 U9555 ( .A1(n7808), .A2(n7757), .ZN(n7761) );
  INV_X1 U9556 ( .A(n7761), .ZN(n7759) );
  XNOR2_X1 U9557 ( .A(n8507), .B(n4432), .ZN(n7760) );
  INV_X1 U9558 ( .A(n7760), .ZN(n7758) );
  INV_X1 U9559 ( .A(n7767), .ZN(n8073) );
  INV_X1 U9560 ( .A(n7766), .ZN(n7765) );
  XNOR2_X1 U9561 ( .A(n8501), .B(n7726), .ZN(n7762) );
  NAND2_X1 U9562 ( .A1(n7762), .A2(n8077), .ZN(n8102) );
  INV_X1 U9563 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U9564 ( .A1(n7763), .A2(n8341), .ZN(n7764) );
  AND2_X1 U9565 ( .A1(n8102), .A2(n7764), .ZN(n7768) );
  NOR3_X1 U9566 ( .A1(n8073), .A2(n7765), .A3(n7768), .ZN(n7770) );
  NAND2_X1 U9567 ( .A1(n7767), .A2(n7766), .ZN(n7769) );
  NAND2_X1 U9568 ( .A1(n7769), .A2(n7768), .ZN(n8037) );
  INV_X1 U9569 ( .A(n8037), .ZN(n8105) );
  OAI21_X1 U9570 ( .B1(n7770), .B2(n8105), .A(n8160), .ZN(n7774) );
  AOI22_X1 U9571 ( .A1(n8321), .A2(n8141), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7771) );
  OAI21_X1 U9572 ( .B1(n8332), .B2(n8143), .A(n7771), .ZN(n7772) );
  AOI21_X1 U9573 ( .B1(n8333), .B2(n8164), .A(n7772), .ZN(n7773) );
  OAI211_X1 U9574 ( .C1(n8501), .C2(n8167), .A(n7774), .B(n7773), .ZN(P2_U3169) );
  XOR2_X1 U9575 ( .A(n7995), .B(n7775), .Z(n7789) );
  INV_X1 U9576 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n7778) );
  XNOR2_X1 U9577 ( .A(n7776), .B(n7995), .ZN(n7777) );
  AOI222_X1 U9578 ( .A1(n8433), .A2(n7777), .B1(n8341), .B2(n9866), .C1(n8187), 
        .C2(n9869), .ZN(n7783) );
  MUX2_X1 U9579 ( .A(n7778), .B(n7783), .S(n9946), .Z(n7780) );
  NAND2_X1 U9580 ( .A1(n8038), .A2(n8546), .ZN(n7779) );
  OAI211_X1 U9581 ( .C1(n7789), .C2(n8550), .A(n7780), .B(n7779), .ZN(P2_U3452) );
  MUX2_X1 U9582 ( .A(n10089), .B(n7783), .S(n9963), .Z(n7782) );
  NAND2_X1 U9583 ( .A1(n8038), .A2(n5724), .ZN(n7781) );
  OAI211_X1 U9584 ( .C1(n7789), .C2(n8479), .A(n7782), .B(n7781), .ZN(P2_U3484) );
  INV_X1 U9585 ( .A(n7783), .ZN(n7786) );
  INV_X1 U9586 ( .A(n8111), .ZN(n7784) );
  OAI22_X1 U9587 ( .A1(n8114), .A2(n9864), .B1(n7784), .B2(n9863), .ZN(n7785)
         );
  OAI21_X1 U9588 ( .B1(n7786), .B2(n7785), .A(n8413), .ZN(n7788) );
  NAND2_X1 U9589 ( .A1(n6677), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7787) );
  OAI211_X1 U9590 ( .C1(n7789), .C2(n8441), .A(n7788), .B(n7787), .ZN(P2_U3208) );
  MUX2_X1 U9591 ( .A(n7791), .B(n7790), .S(n9678), .Z(n7792) );
  OAI21_X1 U9592 ( .B1(n9178), .B2(n9407), .A(n7792), .ZN(P1_U3551) );
  XNOR2_X1 U9593 ( .A(n7793), .B(n7984), .ZN(n8352) );
  XNOR2_X1 U9594 ( .A(n7794), .B(n7984), .ZN(n7795) );
  OAI222_X1 U9595 ( .A1(n8396), .A2(n7796), .B1(n8394), .B2(n8332), .C1(n9873), 
        .C2(n7795), .ZN(n8347) );
  AOI21_X1 U9596 ( .B1(n9938), .B2(n8352), .A(n8347), .ZN(n7799) );
  MUX2_X1 U9597 ( .A(n7797), .B(n7799), .S(n9946), .Z(n7798) );
  OAI21_X1 U9598 ( .B1(n8350), .B2(n8530), .A(n7798), .ZN(P2_U3449) );
  INV_X1 U9599 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7800) );
  MUX2_X1 U9600 ( .A(n7800), .B(n7799), .S(n9963), .Z(n7801) );
  OAI21_X1 U9601 ( .B1(n8350), .B2(n8471), .A(n7801), .ZN(P2_U3481) );
  NAND2_X1 U9602 ( .A1(n7802), .A2(n8136), .ZN(n8092) );
  NAND2_X1 U9603 ( .A1(n8092), .A2(n7803), .ZN(n7804) );
  INV_X1 U9604 ( .A(n7805), .ZN(n7807) );
  NOR3_X1 U9605 ( .A1(n8095), .A2(n7807), .A3(n7753), .ZN(n7813) );
  NAND2_X1 U9606 ( .A1(n7808), .A2(n7809), .ZN(n7811) );
  OR2_X1 U9607 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  OAI21_X1 U9608 ( .B1(n7813), .B2(n7812), .A(n8160), .ZN(n7817) );
  AOI22_X1 U9609 ( .A1(n5471), .A2(n8172), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7814) );
  OAI21_X1 U9610 ( .B1(n8332), .B2(n8170), .A(n7814), .ZN(n7815) );
  AOI21_X1 U9611 ( .B1(n8348), .B2(n8164), .A(n7815), .ZN(n7816) );
  OAI211_X1 U9612 ( .C1(n8350), .C2(n8167), .A(n7817), .B(n7816), .ZN(P2_U3175) );
  INV_X1 U9613 ( .A(n7818), .ZN(n8035) );
  OAI222_X1 U9614 ( .A1(P1_U3086), .A2(n7819), .B1(n9476), .B2(n8035), .C1(
        n9478), .C2(n6073), .ZN(P1_U3328) );
  OR2_X1 U9615 ( .A1(n7825), .A2(n6298), .ZN(n7820) );
  NAND2_X1 U9616 ( .A1(n7823), .A2(n7822), .ZN(n7827) );
  OR2_X1 U9617 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  INV_X1 U9618 ( .A(n8185), .ZN(n8293) );
  NAND2_X1 U9619 ( .A1(n7828), .A2(n8293), .ZN(n8011) );
  INV_X1 U9620 ( .A(n8184), .ZN(n7829) );
  AND2_X1 U9621 ( .A1(n8485), .A2(n7829), .ZN(n8009) );
  INV_X1 U9622 ( .A(n8009), .ZN(n7866) );
  OAI211_X1 U9623 ( .C1(n8481), .C2(n8446), .A(n8011), .B(n7866), .ZN(n7830)
         );
  INV_X1 U9624 ( .A(n8022), .ZN(n7834) );
  NAND2_X1 U9625 ( .A1(n8481), .A2(n8006), .ZN(n7832) );
  INV_X1 U9626 ( .A(n8006), .ZN(n7868) );
  INV_X1 U9627 ( .A(n7978), .ZN(n7987) );
  NOR2_X1 U9628 ( .A1(n7976), .A2(n7987), .ZN(n8340) );
  INV_X1 U9629 ( .A(n8370), .ZN(n8367) );
  INV_X1 U9630 ( .A(n8390), .ZN(n8399) );
  NAND2_X1 U9631 ( .A1(n7836), .A2(n7880), .ZN(n7873) );
  INV_X1 U9632 ( .A(n7873), .ZN(n7841) );
  NAND2_X1 U9633 ( .A1(n6185), .A2(n7837), .ZN(n7882) );
  NOR2_X1 U9634 ( .A1(n7838), .A2(n7882), .ZN(n7840) );
  NAND4_X1 U9635 ( .A1(n7841), .A2(n5103), .A3(n7840), .A4(n7839), .ZN(n7845)
         );
  INV_X1 U9636 ( .A(n7842), .ZN(n7844) );
  NOR3_X1 U9637 ( .A1(n7845), .A2(n7844), .A3(n7843), .ZN(n7847) );
  NAND4_X1 U9638 ( .A1(n4673), .A2(n7847), .A3(n7916), .A4(n7846), .ZN(n7848)
         );
  NOR2_X1 U9639 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  NAND4_X1 U9640 ( .A1(n7851), .A2(n5640), .A3(n7850), .A4(n4700), .ZN(n7852)
         );
  NOR2_X1 U9641 ( .A1(n7853), .A2(n7852), .ZN(n7857) );
  INV_X1 U9642 ( .A(n7854), .ZN(n7855) );
  AND4_X1 U9643 ( .A1(n8409), .A2(n8419), .A3(n7857), .A4(n8429), .ZN(n7858)
         );
  NAND4_X1 U9644 ( .A1(n8367), .A2(n8381), .A3(n8399), .A4(n7858), .ZN(n7859)
         );
  NOR2_X1 U9645 ( .A1(n8358), .A2(n7859), .ZN(n7860) );
  NAND4_X1 U9646 ( .A1(n8329), .A2(n7861), .A3(n8340), .A4(n7860), .ZN(n7862)
         );
  NOR2_X1 U9647 ( .A1(n7862), .A2(n7995), .ZN(n7863) );
  NAND3_X1 U9648 ( .A1(n8318), .A2(n7863), .A3(n8308), .ZN(n7864) );
  NOR2_X1 U9649 ( .A1(n8291), .A2(n7864), .ZN(n7865) );
  NAND2_X1 U9650 ( .A1(n8011), .A2(n8007), .ZN(n8008) );
  INV_X1 U9651 ( .A(n8008), .ZN(n7870) );
  NAND2_X1 U9652 ( .A1(n8281), .A2(n8185), .ZN(n8010) );
  INV_X1 U9653 ( .A(n8010), .ZN(n7869) );
  NOR3_X1 U9654 ( .A1(n8006), .A2(n7870), .A3(n7869), .ZN(n8020) );
  NAND2_X1 U9655 ( .A1(n8198), .A2(n9884), .ZN(n7871) );
  AND2_X1 U9656 ( .A1(n7904), .A2(n7871), .ZN(n7877) );
  NAND2_X1 U9657 ( .A1(n7879), .A2(n8007), .ZN(n7872) );
  AND2_X1 U9658 ( .A1(n7873), .A2(n7872), .ZN(n7878) );
  NAND2_X1 U9659 ( .A1(n7889), .A2(n7874), .ZN(n7875) );
  AOI21_X1 U9660 ( .B1(n7878), .B2(n7839), .A(n7875), .ZN(n7876) );
  MUX2_X1 U9661 ( .A(n7877), .B(n7876), .S(n8007), .Z(n7888) );
  INV_X1 U9662 ( .A(n7878), .ZN(n7885) );
  INV_X1 U9663 ( .A(n7879), .ZN(n7884) );
  NAND4_X1 U9664 ( .A1(n7882), .A2(n8007), .A3(n7881), .A4(n7880), .ZN(n7883)
         );
  OAI21_X1 U9665 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7886) );
  NAND2_X1 U9666 ( .A1(n7886), .A2(n7839), .ZN(n7887) );
  NAND2_X1 U9667 ( .A1(n7888), .A2(n7887), .ZN(n7906) );
  NAND3_X1 U9668 ( .A1(n7906), .A2(n7905), .A3(n7889), .ZN(n7891) );
  NAND3_X1 U9669 ( .A1(n7891), .A2(n7890), .A3(n7910), .ZN(n7892) );
  NAND2_X1 U9670 ( .A1(n7892), .A2(n7908), .ZN(n7893) );
  NAND3_X1 U9671 ( .A1(n7893), .A2(n7916), .A3(n7914), .ZN(n7895) );
  NAND3_X1 U9672 ( .A1(n7895), .A2(n7896), .A3(n7894), .ZN(n7900) );
  AND2_X1 U9673 ( .A1(n7901), .A2(n7896), .ZN(n7899) );
  AND2_X1 U9674 ( .A1(n7922), .A2(n7897), .ZN(n7898) );
  MUX2_X1 U9675 ( .A(n7899), .B(n7898), .S(n8005), .Z(n7918) );
  NAND2_X1 U9676 ( .A1(n7900), .A2(n7918), .ZN(n7902) );
  NAND3_X1 U9677 ( .A1(n7902), .A2(n7924), .A3(n7901), .ZN(n7903) );
  NAND2_X1 U9678 ( .A1(n7903), .A2(n7923), .ZN(n7928) );
  NAND3_X1 U9679 ( .A1(n7906), .A2(n7905), .A3(n7904), .ZN(n7909) );
  NAND3_X1 U9680 ( .A1(n7909), .A2(n7908), .A3(n7907), .ZN(n7915) );
  INV_X1 U9681 ( .A(n7910), .ZN(n7912) );
  NAND2_X1 U9682 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  NAND3_X1 U9683 ( .A1(n7915), .A2(n7914), .A3(n7913), .ZN(n7917) );
  NAND2_X1 U9684 ( .A1(n7917), .A2(n7916), .ZN(n7921) );
  INV_X1 U9685 ( .A(n7918), .ZN(n7919) );
  AOI21_X1 U9686 ( .B1(n7921), .B2(n7920), .A(n7919), .ZN(n7926) );
  NAND2_X1 U9687 ( .A1(n7923), .A2(n7922), .ZN(n7925) );
  OAI21_X1 U9688 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7927) );
  MUX2_X1 U9689 ( .A(n7928), .B(n7927), .S(n8007), .Z(n7942) );
  INV_X1 U9690 ( .A(n7935), .ZN(n7941) );
  NAND2_X1 U9691 ( .A1(n7932), .A2(n7931), .ZN(n7934) );
  NAND2_X1 U9692 ( .A1(n7934), .A2(n7933), .ZN(n7937) );
  NAND2_X1 U9693 ( .A1(n7936), .A2(n7944), .ZN(n7939) );
  NAND2_X1 U9694 ( .A1(n7943), .A2(n7937), .ZN(n7938) );
  AOI21_X1 U9695 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7951) );
  MUX2_X1 U9696 ( .A(n7944), .B(n7943), .S(n8005), .Z(n7945) );
  NAND2_X1 U9697 ( .A1(n7946), .A2(n7945), .ZN(n7950) );
  MUX2_X1 U9698 ( .A(n7948), .B(n7947), .S(n8005), .Z(n7949) );
  OAI211_X1 U9699 ( .C1(n7951), .C2(n7950), .A(n8429), .B(n7949), .ZN(n7955)
         );
  MUX2_X1 U9700 ( .A(n7953), .B(n7952), .S(n8005), .Z(n7954) );
  OAI211_X1 U9701 ( .C1(n8005), .C2(n7957), .A(n8409), .B(n7956), .ZN(n7963)
         );
  INV_X1 U9702 ( .A(n7960), .ZN(n7962) );
  NAND2_X1 U9703 ( .A1(n7969), .A2(n7972), .ZN(n7965) );
  NAND2_X1 U9704 ( .A1(n7965), .A2(n7970), .ZN(n7975) );
  INV_X1 U9705 ( .A(n7966), .ZN(n7968) );
  OAI21_X1 U9706 ( .B1(n7969), .B2(n7968), .A(n7967), .ZN(n7973) );
  INV_X1 U9707 ( .A(n7970), .ZN(n7971) );
  AOI21_X1 U9708 ( .B1(n7973), .B2(n7972), .A(n7971), .ZN(n7974) );
  INV_X1 U9709 ( .A(n7976), .ZN(n7985) );
  NAND2_X1 U9710 ( .A1(n7978), .A2(n7977), .ZN(n7981) );
  INV_X1 U9711 ( .A(n7979), .ZN(n7980) );
  MUX2_X1 U9712 ( .A(n7981), .B(n7980), .S(n8005), .Z(n7982) );
  INV_X1 U9713 ( .A(n7982), .ZN(n7983) );
  AND2_X1 U9714 ( .A1(n7989), .A2(n7985), .ZN(n7986) );
  NOR2_X1 U9715 ( .A1(n7988), .A2(n7987), .ZN(n7991) );
  INV_X1 U9716 ( .A(n7989), .ZN(n7990) );
  MUX2_X1 U9717 ( .A(n4473), .B(n7992), .S(n8005), .Z(n7993) );
  INV_X1 U9718 ( .A(n7993), .ZN(n7994) );
  OAI21_X1 U9719 ( .B1(n7996), .B2(n7995), .A(n7994), .ZN(n7997) );
  MUX2_X1 U9720 ( .A(n7998), .B(n4495), .S(n8007), .Z(n7999) );
  MUX2_X1 U9721 ( .A(n8320), .B(n8452), .S(n8005), .Z(n8001) );
  NAND2_X1 U9722 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  MUX2_X1 U9723 ( .A(n8186), .B(n8448), .S(n8007), .Z(n8004) );
  MUX2_X1 U9724 ( .A(n8011), .B(n8010), .S(n8007), .Z(n8003) );
  OAI21_X1 U9725 ( .B1(n8017), .B2(n8004), .A(n8003), .ZN(n8019) );
  NOR4_X1 U9726 ( .A1(n8019), .A2(n8006), .A3(n8005), .A4(n8186), .ZN(n8018)
         );
  NOR3_X1 U9727 ( .A1(n8009), .A2(n8306), .A3(n8007), .ZN(n8016) );
  NAND2_X1 U9728 ( .A1(n8010), .A2(n8448), .ZN(n8012) );
  NAND3_X1 U9729 ( .A1(n8012), .A2(n8011), .A3(n8184), .ZN(n8014) );
  AOI21_X1 U9730 ( .B1(n8012), .B2(n8011), .A(n8184), .ZN(n8013) );
  AOI21_X1 U9731 ( .B1(n8485), .B2(n8014), .A(n8013), .ZN(n8015) );
  NAND3_X1 U9732 ( .A1(n8028), .A2(n8027), .A3(n8257), .ZN(n8029) );
  OAI211_X1 U9733 ( .C1(n8030), .C2(n8032), .A(n8029), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8031) );
  OAI222_X1 U9734 ( .A1(n8562), .A2(n8034), .B1(P2_U3151), .B2(n8033), .C1(
        n10247), .C2(n8555), .ZN(P2_U3270) );
  OAI222_X1 U9735 ( .A1(n8555), .A2(n8036), .B1(n8562), .B2(n8035), .C1(
        P2_U3151), .C2(n8257), .ZN(P2_U3268) );
  NAND2_X1 U9736 ( .A1(n8037), .A2(n8102), .ZN(n8039) );
  XNOR2_X1 U9737 ( .A(n8038), .B(n7735), .ZN(n8040) );
  XNOR2_X1 U9738 ( .A(n8040), .B(n8321), .ZN(n8103) );
  NAND2_X1 U9739 ( .A1(n8040), .A2(n8331), .ZN(n8041) );
  XNOR2_X1 U9740 ( .A(n8496), .B(n4432), .ZN(n8158) );
  XNOR2_X1 U9741 ( .A(n8452), .B(n7726), .ZN(n8042) );
  NAND2_X1 U9742 ( .A1(n8042), .A2(n8320), .ZN(n8043) );
  OAI21_X1 U9743 ( .B1(n8042), .B2(n8320), .A(n8043), .ZN(n8065) );
  NAND2_X1 U9744 ( .A1(n8063), .A2(n8043), .ZN(n8045) );
  XNOR2_X1 U9745 ( .A(n8291), .B(n7735), .ZN(n8044) );
  XNOR2_X1 U9746 ( .A(n8045), .B(n8044), .ZN(n8046) );
  NAND2_X1 U9747 ( .A1(n8046), .A2(n8160), .ZN(n8052) );
  INV_X1 U9748 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8047) );
  OAI22_X1 U9749 ( .A1(n8294), .A2(n8143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8047), .ZN(n8050) );
  INV_X1 U9750 ( .A(n8048), .ZN(n8300) );
  OAI22_X1 U9751 ( .A1(n8293), .A2(n8170), .B1(n8300), .B2(n8174), .ZN(n8049)
         );
  AOI211_X1 U9752 ( .C1(n8448), .C2(n8182), .A(n8050), .B(n8049), .ZN(n8051)
         );
  NAND2_X1 U9753 ( .A1(n8052), .A2(n8051), .ZN(P2_U3160) );
  INV_X1 U9754 ( .A(n8053), .ZN(n8563) );
  OAI222_X1 U9755 ( .A1(n9478), .A2(n8055), .B1(n9476), .B2(n8563), .C1(n8054), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  OAI21_X1 U9756 ( .B1(n8690), .B2(n9621), .A(n8056), .ZN(n8060) );
  AOI22_X1 U9757 ( .A1(n8692), .A2(n9627), .B1(n9321), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n8057) );
  OAI21_X1 U9758 ( .B1(n8058), .B2(n9629), .A(n8057), .ZN(n8059) );
  AOI21_X1 U9759 ( .B1(n8060), .B2(n9624), .A(n8059), .ZN(n8061) );
  OAI21_X1 U9760 ( .B1(n8062), .B2(n9328), .A(n8061), .ZN(P1_U3265) );
  INV_X1 U9761 ( .A(n8452), .ZN(n8072) );
  NAND2_X1 U9762 ( .A1(n8064), .A2(n8065), .ZN(n8066) );
  NAND3_X1 U9763 ( .A1(n8063), .A2(n8160), .A3(n8066), .ZN(n8071) );
  INV_X1 U9764 ( .A(n8312), .ZN(n8068) );
  AOI22_X1 U9765 ( .A1(n8187), .A2(n8172), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8067) );
  OAI21_X1 U9766 ( .B1(n8068), .B2(n8174), .A(n8067), .ZN(n8069) );
  AOI21_X1 U9767 ( .B1(n8141), .B2(n8186), .A(n8069), .ZN(n8070) );
  OAI211_X1 U9768 ( .C1(n8072), .C2(n8167), .A(n8071), .B(n8070), .ZN(P2_U3154) );
  AOI21_X1 U9769 ( .B1(n8188), .B2(n8074), .A(n8073), .ZN(n8080) );
  AOI22_X1 U9770 ( .A1(n8361), .A2(n8172), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8076) );
  NAND2_X1 U9771 ( .A1(n8344), .A2(n8164), .ZN(n8075) );
  OAI211_X1 U9772 ( .C1(n8077), .C2(n8170), .A(n8076), .B(n8075), .ZN(n8078)
         );
  AOI21_X1 U9773 ( .B1(n8507), .B2(n8182), .A(n8078), .ZN(n8079) );
  OAI21_X1 U9774 ( .B1(n8080), .B2(n8177), .A(n8079), .ZN(P2_U3156) );
  INV_X1 U9775 ( .A(n8523), .ZN(n8091) );
  INV_X1 U9776 ( .A(n8081), .ZN(n8151) );
  INV_X1 U9777 ( .A(n8082), .ZN(n8084) );
  NOR3_X1 U9778 ( .A1(n8151), .A2(n8084), .A3(n8083), .ZN(n8086) );
  INV_X1 U9779 ( .A(n8085), .ZN(n8138) );
  OAI21_X1 U9780 ( .B1(n8086), .B2(n8138), .A(n8160), .ZN(n8090) );
  NOR2_X1 U9781 ( .A1(n10241), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8267) );
  AOI21_X1 U9782 ( .B1(n8360), .B2(n8141), .A(n8267), .ZN(n8087) );
  OAI21_X1 U9783 ( .B1(n8382), .B2(n8143), .A(n8087), .ZN(n8088) );
  AOI21_X1 U9784 ( .B1(n8387), .B2(n8164), .A(n8088), .ZN(n8089) );
  OAI211_X1 U9785 ( .C1(n8091), .C2(n8167), .A(n8090), .B(n8089), .ZN(P2_U3159) );
  INV_X1 U9786 ( .A(n8092), .ZN(n8139) );
  NOR3_X1 U9787 ( .A1(n8139), .A2(n8094), .A3(n8093), .ZN(n8096) );
  OAI21_X1 U9788 ( .B1(n8096), .B2(n8095), .A(n8160), .ZN(n8100) );
  AOI22_X1 U9789 ( .A1(n8361), .A2(n8141), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8097) );
  OAI21_X1 U9790 ( .B1(n8383), .B2(n8143), .A(n8097), .ZN(n8098) );
  AOI21_X1 U9791 ( .B1(n8364), .B2(n8164), .A(n8098), .ZN(n8099) );
  OAI211_X1 U9792 ( .C1(n8101), .C2(n8167), .A(n8100), .B(n8099), .ZN(P2_U3163) );
  INV_X1 U9793 ( .A(n8102), .ZN(n8104) );
  NOR3_X1 U9794 ( .A1(n8105), .A2(n8104), .A3(n8103), .ZN(n8108) );
  INV_X1 U9795 ( .A(n8106), .ZN(n8107) );
  OAI21_X1 U9796 ( .B1(n8108), .B2(n8107), .A(n8160), .ZN(n8113) );
  AOI22_X1 U9797 ( .A1(n8341), .A2(n8172), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8109) );
  OAI21_X1 U9798 ( .B1(n8307), .B2(n8170), .A(n8109), .ZN(n8110) );
  AOI21_X1 U9799 ( .B1(n8111), .B2(n8164), .A(n8110), .ZN(n8112) );
  OAI211_X1 U9800 ( .C1(n8114), .C2(n8167), .A(n8113), .B(n8112), .ZN(P2_U3165) );
  INV_X1 U9801 ( .A(n8540), .ZN(n8124) );
  AOI21_X1 U9802 ( .B1(n8175), .B2(n8116), .A(n8115), .ZN(n8117) );
  OAI21_X1 U9803 ( .B1(n4498), .B2(n8117), .A(n8160), .ZN(n8123) );
  INV_X1 U9804 ( .A(n8118), .ZN(n8424) );
  AOI22_X1 U9805 ( .A1(n8141), .A2(n8421), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8119) );
  OAI21_X1 U9806 ( .B1(n8120), .B2(n8143), .A(n8119), .ZN(n8121) );
  AOI21_X1 U9807 ( .B1(n8424), .B2(n8164), .A(n8121), .ZN(n8122) );
  OAI211_X1 U9808 ( .C1(n8124), .C2(n8167), .A(n8123), .B(n8122), .ZN(P2_U3166) );
  NOR3_X1 U9809 ( .A1(n4498), .A2(n8126), .A3(n8125), .ZN(n8128) );
  INV_X1 U9810 ( .A(n8127), .ZN(n8150) );
  OAI21_X1 U9811 ( .B1(n8128), .B2(n8150), .A(n8160), .ZN(n8133) );
  INV_X1 U9812 ( .A(n8129), .ZN(n8415) );
  NAND2_X1 U9813 ( .A1(n8141), .A2(n8411), .ZN(n8130) );
  NAND2_X1 U9814 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9859) );
  OAI211_X1 U9815 ( .C1(n8169), .C2(n8143), .A(n8130), .B(n9859), .ZN(n8131)
         );
  AOI21_X1 U9816 ( .B1(n8164), .B2(n8415), .A(n8131), .ZN(n8132) );
  OAI211_X1 U9817 ( .C1(n8134), .C2(n8167), .A(n8133), .B(n8132), .ZN(P2_U3168) );
  INV_X1 U9818 ( .A(n8135), .ZN(n8137) );
  NOR3_X1 U9819 ( .A1(n8138), .A2(n8137), .A3(n8136), .ZN(n8140) );
  OAI21_X1 U9820 ( .B1(n8140), .B2(n8139), .A(n8160), .ZN(n8146) );
  AOI22_X1 U9821 ( .A1(n5471), .A2(n8141), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8142) );
  OAI21_X1 U9822 ( .B1(n8393), .B2(n8143), .A(n8142), .ZN(n8144) );
  AOI21_X1 U9823 ( .B1(n8375), .B2(n8164), .A(n8144), .ZN(n8145) );
  OAI211_X1 U9824 ( .C1(n5459), .C2(n8167), .A(n8146), .B(n8145), .ZN(P2_U3173) );
  INV_X1 U9825 ( .A(n8147), .ZN(n8149) );
  NOR3_X1 U9826 ( .A1(n8150), .A2(n8149), .A3(n8148), .ZN(n8152) );
  OAI21_X1 U9827 ( .B1(n8152), .B2(n8151), .A(n8160), .ZN(n8156) );
  NAND2_X1 U9828 ( .A1(n8172), .A2(n8421), .ZN(n8153) );
  NAND2_X1 U9829 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8227) );
  OAI211_X1 U9830 ( .C1(n8393), .C2(n8170), .A(n8153), .B(n8227), .ZN(n8154)
         );
  AOI21_X1 U9831 ( .B1(n8164), .B2(n8401), .A(n8154), .ZN(n8155) );
  OAI211_X1 U9832 ( .C1(n8531), .C2(n8167), .A(n8156), .B(n8155), .ZN(P2_U3178) );
  XNOR2_X1 U9833 ( .A(n8158), .B(n8187), .ZN(n8159) );
  XNOR2_X1 U9834 ( .A(n8157), .B(n8159), .ZN(n8161) );
  NAND2_X1 U9835 ( .A1(n8161), .A2(n8160), .ZN(n8166) );
  AOI22_X1 U9836 ( .A1(n8321), .A2(n8172), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8162) );
  OAI21_X1 U9837 ( .B1(n8294), .B2(n8170), .A(n8162), .ZN(n8163) );
  AOI21_X1 U9838 ( .B1(n8324), .B2(n8164), .A(n8163), .ZN(n8165) );
  OAI211_X1 U9839 ( .C1(n8168), .C2(n8167), .A(n8166), .B(n8165), .ZN(P2_U3180) );
  NOR2_X1 U9840 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10147), .ZN(n9817) );
  NOR2_X1 U9841 ( .A1(n8170), .A2(n8169), .ZN(n8171) );
  AOI211_X1 U9842 ( .C1(n8172), .C2(n8431), .A(n9817), .B(n8171), .ZN(n8173)
         );
  OAI21_X1 U9843 ( .B1(n8435), .B2(n8174), .A(n8173), .ZN(n8181) );
  INV_X1 U9844 ( .A(n8175), .ZN(n8176) );
  AOI211_X1 U9845 ( .C1(n8179), .C2(n8178), .A(n8177), .B(n8176), .ZN(n8180)
         );
  AOI211_X1 U9846 ( .C1(n8547), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8183)
         );
  INV_X1 U9847 ( .A(n8183), .ZN(P2_U3181) );
  MUX2_X1 U9848 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8184), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9849 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8185), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8186), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8187), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9852 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8321), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9853 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8341), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9854 ( .A(n8188), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8225), .Z(
        P2_U3514) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8361), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9856 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n5471), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8360), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8372), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8411), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8421), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8430), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9862 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8422), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9863 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8431), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9864 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8189), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9865 ( .A(n8190), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8225), .Z(
        P2_U3503) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8191), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9867 ( .A(n8192), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8225), .Z(
        P2_U3501) );
  MUX2_X1 U9868 ( .A(n8193), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8225), .Z(
        P2_U3499) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8194), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9870 ( .A(n8195), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8225), .Z(
        P2_U3497) );
  MUX2_X1 U9871 ( .A(n8196), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8225), .Z(
        P2_U3496) );
  MUX2_X1 U9872 ( .A(n8197), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8225), .Z(
        P2_U3495) );
  MUX2_X1 U9873 ( .A(n9868), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8225), .Z(
        P2_U3494) );
  MUX2_X1 U9874 ( .A(n8198), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8225), .Z(
        P2_U3493) );
  MUX2_X1 U9875 ( .A(n9867), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8225), .Z(
        P2_U3492) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n5632), .S(P2_U3893), .Z(
        P2_U3491) );
  NOR2_X1 U9877 ( .A1(n8252), .A2(n8199), .ZN(n8200) );
  AOI21_X1 U9878 ( .B1(n8199), .B2(n8252), .A(n8200), .ZN(n8210) );
  NOR2_X1 U9879 ( .A1(n8202), .A2(n8201), .ZN(n8204) );
  NAND2_X1 U9880 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8234), .ZN(n8205) );
  OAI21_X1 U9881 ( .B1(n8234), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8205), .ZN(
        n9803) );
  NOR2_X1 U9882 ( .A1(n9809), .A2(n8206), .ZN(n8207) );
  XNOR2_X1 U9883 ( .A(n9809), .B(n8206), .ZN(n9819) );
  NOR2_X1 U9884 ( .A1(n8434), .A2(n9819), .ZN(n9818) );
  XNOR2_X1 U9885 ( .A(n8232), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U9886 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  NOR2_X1 U9887 ( .A1(n9843), .A2(n8208), .ZN(n8209) );
  XNOR2_X1 U9888 ( .A(n9843), .B(n8208), .ZN(n9855) );
  AOI21_X1 U9889 ( .B1(n8210), .B2(n4496), .A(n8250), .ZN(n8249) );
  MUX2_X1 U9890 ( .A(n8414), .B(n10123), .S(n8257), .Z(n8221) );
  XNOR2_X1 U9891 ( .A(n8244), .B(n8221), .ZN(n9849) );
  MUX2_X1 U9892 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8213), .Z(n8211) );
  OR2_X1 U9893 ( .A1(n8232), .A2(n8211), .ZN(n8220) );
  XNOR2_X1 U9894 ( .A(n8211), .B(n9825), .ZN(n9831) );
  MUX2_X1 U9895 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8257), .Z(n8212) );
  OR2_X1 U9896 ( .A1(n8212), .A2(n8241), .ZN(n8219) );
  XNOR2_X1 U9897 ( .A(n9809), .B(n8212), .ZN(n9814) );
  MUX2_X1 U9898 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8213), .Z(n8214) );
  OR2_X1 U9899 ( .A1(n8214), .A2(n8234), .ZN(n8218) );
  XNOR2_X1 U9900 ( .A(n8214), .B(n9793), .ZN(n9799) );
  OR2_X1 U9901 ( .A1(n8215), .A2(n8236), .ZN(n8217) );
  NAND2_X1 U9902 ( .A1(n8217), .A2(n8216), .ZN(n9798) );
  NAND2_X1 U9903 ( .A1(n9799), .A2(n9798), .ZN(n9797) );
  NAND2_X1 U9904 ( .A1(n8218), .A2(n9797), .ZN(n9813) );
  NAND2_X1 U9905 ( .A1(n9814), .A2(n9813), .ZN(n9812) );
  NAND2_X1 U9906 ( .A1(n8219), .A2(n9812), .ZN(n9830) );
  NAND2_X1 U9907 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  MUX2_X1 U9908 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8257), .Z(n8222) );
  NOR2_X1 U9909 ( .A1(n8223), .A2(n8222), .ZN(n8260) );
  NAND2_X1 U9910 ( .A1(n8223), .A2(n8222), .ZN(n8261) );
  INV_X1 U9911 ( .A(n8261), .ZN(n8224) );
  NOR2_X1 U9912 ( .A1(n8260), .A2(n8224), .ZN(n8228) );
  INV_X1 U9913 ( .A(n8228), .ZN(n8226) );
  OAI21_X1 U9914 ( .B1(n8226), .B2(n8225), .A(n9708), .ZN(n8231) );
  INV_X1 U9915 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9971) );
  OAI21_X1 U9916 ( .B1(n9713), .B2(n9971), .A(n8227), .ZN(n8230) );
  NOR3_X1 U9917 ( .A1(n8228), .A2(n8262), .A3(n9692), .ZN(n8229) );
  AOI211_X1 U9918 ( .C1(n8262), .C2(n8231), .A(n8230), .B(n8229), .ZN(n8248)
         );
  AOI22_X1 U9919 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8232), .B1(n9825), .B2(
        n10255), .ZN(n9828) );
  NAND2_X1 U9920 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8234), .ZN(n8239) );
  AOI22_X1 U9921 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8234), .B1(n9793), .B2(
        n8233), .ZN(n9796) );
  NAND2_X1 U9922 ( .A1(n8236), .A2(n8235), .ZN(n8238) );
  NAND2_X1 U9923 ( .A1(n8238), .A2(n8237), .ZN(n9795) );
  NAND2_X1 U9924 ( .A1(n9796), .A2(n9795), .ZN(n9794) );
  NAND2_X1 U9925 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U9926 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9811), .ZN(n9810) );
  NAND2_X1 U9927 ( .A1(n8242), .A2(n9810), .ZN(n9827) );
  NAND2_X1 U9928 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  OAI21_X1 U9929 ( .B1(n9825), .B2(n10255), .A(n9826), .ZN(n8243) );
  NAND2_X1 U9930 ( .A1(n8244), .A2(n8243), .ZN(n8245) );
  NAND2_X1 U9931 ( .A1(n8245), .A2(n9845), .ZN(n8254) );
  XNOR2_X1 U9932 ( .A(n8262), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8253) );
  XNOR2_X1 U9933 ( .A(n8254), .B(n8253), .ZN(n8246) );
  NAND2_X1 U9934 ( .A1(n8246), .A2(n9852), .ZN(n8247) );
  OAI211_X1 U9935 ( .C1(n8249), .C2(n9856), .A(n8248), .B(n8247), .ZN(P2_U3200) );
  MUX2_X1 U9936 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8386), .S(n8255), .Z(n8259)
         );
  AOI22_X1 U9937 ( .A1(n8254), .A2(n8253), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8252), .ZN(n8256) );
  XNOR2_X1 U9938 ( .A(n8255), .B(n8465), .ZN(n8258) );
  XNOR2_X1 U9939 ( .A(n8256), .B(n8258), .ZN(n8269) );
  MUX2_X1 U9940 ( .A(n8259), .B(n8258), .S(n8257), .Z(n8264) );
  AOI21_X1 U9941 ( .B1(n8262), .B2(n8261), .A(n8260), .ZN(n8263) );
  NOR2_X1 U9942 ( .A1(n9708), .A2(n8265), .ZN(n8266) );
  AOI211_X1 U9943 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n9842), .A(n8267), .B(
        n8266), .ZN(n8268) );
  NAND2_X1 U9944 ( .A1(n8481), .A2(n8438), .ZN(n8275) );
  INV_X1 U9945 ( .A(n8271), .ZN(n8272) );
  NOR2_X1 U9946 ( .A1(n8273), .A2(n8272), .ZN(n8482) );
  NOR2_X1 U9947 ( .A1(n8274), .A2(n9863), .ZN(n8283) );
  AOI21_X1 U9948 ( .B1(n8482), .B2(n9876), .A(n8283), .ZN(n8278) );
  OAI211_X1 U9949 ( .C1(n8413), .C2(n8276), .A(n8275), .B(n8278), .ZN(P2_U3202) );
  NAND2_X1 U9950 ( .A1(n6677), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8277) );
  OAI211_X1 U9951 ( .C1(n8446), .C2(n8403), .A(n8278), .B(n8277), .ZN(P2_U3203) );
  INV_X1 U9952 ( .A(n8279), .ZN(n8287) );
  NAND2_X1 U9953 ( .A1(n8280), .A2(n8413), .ZN(n8285) );
  NOR2_X1 U9954 ( .A1(n8281), .A2(n8403), .ZN(n8282) );
  AOI211_X1 U9955 ( .C1(n6677), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8283), .B(
        n8282), .ZN(n8284) );
  OAI211_X1 U9956 ( .C1(n8287), .C2(n8286), .A(n8285), .B(n8284), .ZN(P2_U3204) );
  INV_X1 U9957 ( .A(n8288), .ZN(n8289) );
  AOI21_X1 U9958 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n8490) );
  NAND2_X1 U9959 ( .A1(n8447), .A2(n9876), .ZN(n8303) );
  INV_X1 U9960 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8299) );
  OAI22_X1 U9961 ( .A1(n8300), .A2(n9863), .B1(n8413), .B2(n8299), .ZN(n8301)
         );
  AOI21_X1 U9962 ( .B1(n8448), .B2(n8438), .A(n8301), .ZN(n8302) );
  OAI211_X1 U9963 ( .C1(n8490), .C2(n8441), .A(n8303), .B(n8302), .ZN(P2_U3205) );
  XNOR2_X1 U9964 ( .A(n8304), .B(n8308), .ZN(n8305) );
  OAI222_X1 U9965 ( .A1(n8396), .A2(n8307), .B1(n8394), .B2(n8306), .C1(n8305), 
        .C2(n9873), .ZN(n8451) );
  OR2_X1 U9966 ( .A1(n8309), .A2(n8308), .ZN(n8311) );
  NAND2_X1 U9967 ( .A1(n8311), .A2(n8310), .ZN(n8494) );
  AOI22_X1 U9968 ( .A1(n8312), .A2(n8437), .B1(n6677), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U9969 ( .A1(n8452), .A2(n8438), .ZN(n8313) );
  OAI211_X1 U9970 ( .C1(n8494), .C2(n8441), .A(n8314), .B(n8313), .ZN(n8315)
         );
  AOI21_X1 U9971 ( .B1(n8451), .B2(n9876), .A(n8315), .ZN(n8316) );
  INV_X1 U9972 ( .A(n8316), .ZN(P2_U3206) );
  XOR2_X1 U9973 ( .A(n8318), .B(n8317), .Z(n8499) );
  INV_X1 U9974 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8323) );
  XNOR2_X1 U9975 ( .A(n8319), .B(n8318), .ZN(n8322) );
  AOI222_X1 U9976 ( .A1(n8433), .A2(n8322), .B1(n8321), .B2(n9866), .C1(n8320), 
        .C2(n9869), .ZN(n8495) );
  MUX2_X1 U9977 ( .A(n8323), .B(n8495), .S(n9876), .Z(n8326) );
  AOI22_X1 U9978 ( .A1(n8496), .A2(n8438), .B1(n8437), .B2(n8324), .ZN(n8325)
         );
  OAI211_X1 U9979 ( .C1(n8499), .C2(n8441), .A(n8326), .B(n8325), .ZN(P2_U3207) );
  XOR2_X1 U9980 ( .A(n8327), .B(n8329), .Z(n8502) );
  XOR2_X1 U9981 ( .A(n8329), .B(n8328), .Z(n8330) );
  OAI222_X1 U9982 ( .A1(n8396), .A2(n8332), .B1(n8394), .B2(n8331), .C1(n8330), 
        .C2(n9873), .ZN(n8500) );
  INV_X1 U9983 ( .A(n8333), .ZN(n8334) );
  OAI22_X1 U9984 ( .A1(n8501), .A2(n9864), .B1(n8334), .B2(n9863), .ZN(n8335)
         );
  OAI21_X1 U9985 ( .B1(n8500), .B2(n8335), .A(n8413), .ZN(n8337) );
  NAND2_X1 U9986 ( .A1(n6677), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8336) );
  OAI211_X1 U9987 ( .C1(n8502), .C2(n8441), .A(n8337), .B(n8336), .ZN(P2_U3209) );
  XNOR2_X1 U9988 ( .A(n8338), .B(n8340), .ZN(n8510) );
  INV_X1 U9989 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8343) );
  XOR2_X1 U9990 ( .A(n8340), .B(n8339), .Z(n8342) );
  AOI222_X1 U9991 ( .A1(n8433), .A2(n8342), .B1(n8341), .B2(n9869), .C1(n8361), 
        .C2(n9866), .ZN(n8505) );
  MUX2_X1 U9992 ( .A(n8343), .B(n8505), .S(n9876), .Z(n8346) );
  AOI22_X1 U9993 ( .A1(n8507), .A2(n8438), .B1(n8437), .B2(n8344), .ZN(n8345)
         );
  OAI211_X1 U9994 ( .C1(n8510), .C2(n8441), .A(n8346), .B(n8345), .ZN(P2_U3210) );
  INV_X1 U9995 ( .A(n8347), .ZN(n8354) );
  AOI22_X1 U9996 ( .A1(n8348), .A2(n8437), .B1(n6677), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8349) );
  OAI21_X1 U9997 ( .B1(n8350), .B2(n8403), .A(n8349), .ZN(n8351) );
  AOI21_X1 U9998 ( .B1(n8352), .B2(n8405), .A(n8351), .ZN(n8353) );
  OAI21_X1 U9999 ( .B1(n8354), .B2(n6677), .A(n8353), .ZN(P2_U3211) );
  NAND2_X1 U10000 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  XNOR2_X1 U10001 ( .A(n8357), .B(n8358), .ZN(n8516) );
  INV_X1 U10002 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U10003 ( .A(n8359), .B(n8358), .ZN(n8362) );
  AOI222_X1 U10004 ( .A1(n8433), .A2(n8362), .B1(n8361), .B2(n9869), .C1(n8360), .C2(n9866), .ZN(n8511) );
  MUX2_X1 U10005 ( .A(n8363), .B(n8511), .S(n9876), .Z(n8366) );
  AOI22_X1 U10006 ( .A1(n8513), .A2(n8438), .B1(n8437), .B2(n8364), .ZN(n8365)
         );
  OAI211_X1 U10007 ( .C1(n8516), .C2(n8441), .A(n8366), .B(n8365), .ZN(
        P2_U3212) );
  XNOR2_X1 U10008 ( .A(n8368), .B(n8367), .ZN(n8521) );
  INV_X1 U10009 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8374) );
  OAI21_X1 U10010 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8373) );
  AOI222_X1 U10011 ( .A1(n8433), .A2(n8373), .B1(n5471), .B2(n9869), .C1(n8372), .C2(n9866), .ZN(n8517) );
  MUX2_X1 U10012 ( .A(n8374), .B(n8517), .S(n9876), .Z(n8377) );
  AOI22_X1 U10013 ( .A1(n8518), .A2(n8438), .B1(n8437), .B2(n8375), .ZN(n8376)
         );
  OAI211_X1 U10014 ( .C1(n8521), .C2(n8441), .A(n8377), .B(n8376), .ZN(
        P2_U3213) );
  XNOR2_X1 U10015 ( .A(n8378), .B(n8381), .ZN(n8526) );
  AOI211_X1 U10016 ( .C1(n8381), .C2(n8380), .A(n9873), .B(n8379), .ZN(n8385)
         );
  OAI22_X1 U10017 ( .A1(n8383), .A2(n8394), .B1(n8382), .B2(n8396), .ZN(n8384)
         );
  NOR2_X1 U10018 ( .A1(n8385), .A2(n8384), .ZN(n8522) );
  MUX2_X1 U10019 ( .A(n8386), .B(n8522), .S(n9876), .Z(n8389) );
  AOI22_X1 U10020 ( .A1(n8523), .A2(n8438), .B1(n8437), .B2(n8387), .ZN(n8388)
         );
  OAI211_X1 U10021 ( .C1(n8526), .C2(n8441), .A(n8389), .B(n8388), .ZN(
        P2_U3214) );
  XNOR2_X1 U10022 ( .A(n8391), .B(n8390), .ZN(n8392) );
  OAI222_X1 U10023 ( .A1(n8396), .A2(n8395), .B1(n8394), .B2(n8393), .C1(n8392), .C2(n9873), .ZN(n8468) );
  INV_X1 U10024 ( .A(n8468), .ZN(n8407) );
  NAND2_X1 U10025 ( .A1(n8398), .A2(n8397), .ZN(n8400) );
  XNOR2_X1 U10026 ( .A(n8400), .B(n8399), .ZN(n8469) );
  AOI22_X1 U10027 ( .A1(n6677), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8437), .B2(
        n8401), .ZN(n8402) );
  OAI21_X1 U10028 ( .B1(n8531), .B2(n8403), .A(n8402), .ZN(n8404) );
  AOI21_X1 U10029 ( .B1(n8469), .B2(n8405), .A(n8404), .ZN(n8406) );
  OAI21_X1 U10030 ( .B1(n8407), .B2(n6677), .A(n8406), .ZN(P2_U3215) );
  XNOR2_X1 U10031 ( .A(n8408), .B(n8409), .ZN(n8537) );
  XOR2_X1 U10032 ( .A(n8410), .B(n8409), .Z(n8412) );
  AOI222_X1 U10033 ( .A1(n8433), .A2(n8412), .B1(n8430), .B2(n9866), .C1(n8411), .C2(n9869), .ZN(n8532) );
  MUX2_X1 U10034 ( .A(n8414), .B(n8532), .S(n8413), .Z(n8417) );
  AOI22_X1 U10035 ( .A1(n8534), .A2(n8438), .B1(n8437), .B2(n8415), .ZN(n8416)
         );
  OAI211_X1 U10036 ( .C1(n8537), .C2(n8441), .A(n8417), .B(n8416), .ZN(
        P2_U3216) );
  XNOR2_X1 U10037 ( .A(n8418), .B(n8419), .ZN(n8543) );
  XNOR2_X1 U10038 ( .A(n8420), .B(n8419), .ZN(n8423) );
  AOI222_X1 U10039 ( .A1(n8433), .A2(n8423), .B1(n8422), .B2(n9866), .C1(n8421), .C2(n9869), .ZN(n8538) );
  MUX2_X1 U10040 ( .A(n10197), .B(n8538), .S(n9876), .Z(n8426) );
  AOI22_X1 U10041 ( .A1(n8540), .A2(n8438), .B1(n8437), .B2(n8424), .ZN(n8425)
         );
  OAI211_X1 U10042 ( .C1(n8543), .C2(n8441), .A(n8426), .B(n8425), .ZN(
        P2_U3217) );
  XNOR2_X1 U10043 ( .A(n8427), .B(n8429), .ZN(n8551) );
  XOR2_X1 U10044 ( .A(n8429), .B(n8428), .Z(n8432) );
  AOI222_X1 U10045 ( .A1(n8433), .A2(n8432), .B1(n8431), .B2(n9866), .C1(n8430), .C2(n9869), .ZN(n8544) );
  MUX2_X1 U10046 ( .A(n8434), .B(n8544), .S(n9876), .Z(n8440) );
  INV_X1 U10047 ( .A(n8435), .ZN(n8436) );
  AOI22_X1 U10048 ( .A1(n8547), .A2(n8438), .B1(n8437), .B2(n8436), .ZN(n8439)
         );
  OAI211_X1 U10049 ( .C1(n8551), .C2(n8441), .A(n8440), .B(n8439), .ZN(
        P2_U3218) );
  NAND2_X1 U10050 ( .A1(n8481), .A2(n5724), .ZN(n8442) );
  NAND2_X1 U10051 ( .A1(n8482), .A2(n9963), .ZN(n8444) );
  OAI211_X1 U10052 ( .C1(n9963), .C2(n8443), .A(n8442), .B(n8444), .ZN(
        P2_U3490) );
  NAND2_X1 U10053 ( .A1(n5726), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8445) );
  OAI211_X1 U10054 ( .C1(n8446), .C2(n8471), .A(n8445), .B(n8444), .ZN(
        P2_U3489) );
  INV_X1 U10055 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8449) );
  AOI21_X1 U10056 ( .B1(n9943), .B2(n8448), .A(n8447), .ZN(n8488) );
  MUX2_X1 U10057 ( .A(n8449), .B(n8488), .S(n9963), .Z(n8450) );
  OAI21_X1 U10058 ( .B1(n8490), .B2(n8479), .A(n8450), .ZN(P2_U3487) );
  MUX2_X1 U10059 ( .A(n10067), .B(n8491), .S(n9963), .Z(n8453) );
  OAI21_X1 U10060 ( .B1(n8479), .B2(n8494), .A(n8453), .ZN(P2_U3486) );
  MUX2_X1 U10061 ( .A(n10266), .B(n8495), .S(n9963), .Z(n8455) );
  NAND2_X1 U10062 ( .A1(n8496), .A2(n5724), .ZN(n8454) );
  OAI211_X1 U10063 ( .C1(n8479), .C2(n8499), .A(n8455), .B(n8454), .ZN(
        P2_U3485) );
  MUX2_X1 U10064 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8500), .S(n9963), .Z(n8457) );
  OAI22_X1 U10065 ( .A1(n8502), .A2(n8479), .B1(n8501), .B2(n8471), .ZN(n8456)
         );
  OR2_X1 U10066 ( .A1(n8457), .A2(n8456), .ZN(P2_U3483) );
  MUX2_X1 U10067 ( .A(n10065), .B(n8505), .S(n9963), .Z(n8459) );
  NAND2_X1 U10068 ( .A1(n8507), .A2(n5724), .ZN(n8458) );
  OAI211_X1 U10069 ( .C1(n8510), .C2(n8479), .A(n8459), .B(n8458), .ZN(
        P2_U3482) );
  MUX2_X1 U10070 ( .A(n10178), .B(n8511), .S(n9963), .Z(n8461) );
  NAND2_X1 U10071 ( .A1(n8513), .A2(n5724), .ZN(n8460) );
  OAI211_X1 U10072 ( .C1(n8479), .C2(n8516), .A(n8461), .B(n8460), .ZN(
        P2_U3480) );
  INV_X1 U10073 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8462) );
  MUX2_X1 U10074 ( .A(n8462), .B(n8517), .S(n9963), .Z(n8464) );
  NAND2_X1 U10075 ( .A1(n8518), .A2(n5724), .ZN(n8463) );
  OAI211_X1 U10076 ( .C1(n8521), .C2(n8479), .A(n8464), .B(n8463), .ZN(
        P2_U3479) );
  MUX2_X1 U10077 ( .A(n8465), .B(n8522), .S(n9963), .Z(n8467) );
  NAND2_X1 U10078 ( .A1(n8523), .A2(n5724), .ZN(n8466) );
  OAI211_X1 U10079 ( .C1(n8526), .C2(n8479), .A(n8467), .B(n8466), .ZN(
        P2_U3478) );
  AOI21_X1 U10080 ( .B1(n8469), .B2(n9938), .A(n8468), .ZN(n8527) );
  MUX2_X1 U10081 ( .A(n10165), .B(n8527), .S(n9963), .Z(n8470) );
  OAI21_X1 U10082 ( .B1(n8531), .B2(n8471), .A(n8470), .ZN(P2_U3477) );
  MUX2_X1 U10083 ( .A(n10123), .B(n8532), .S(n9963), .Z(n8473) );
  NAND2_X1 U10084 ( .A1(n8534), .A2(n5724), .ZN(n8472) );
  OAI211_X1 U10085 ( .C1(n8537), .C2(n8479), .A(n8473), .B(n8472), .ZN(
        P2_U3476) );
  MUX2_X1 U10086 ( .A(n10255), .B(n8538), .S(n9963), .Z(n8475) );
  NAND2_X1 U10087 ( .A1(n8540), .A2(n5724), .ZN(n8474) );
  OAI211_X1 U10088 ( .C1(n8543), .C2(n8479), .A(n8475), .B(n8474), .ZN(
        P2_U3475) );
  MUX2_X1 U10089 ( .A(n8476), .B(n8544), .S(n9963), .Z(n8478) );
  NAND2_X1 U10090 ( .A1(n8547), .A2(n5724), .ZN(n8477) );
  OAI211_X1 U10091 ( .C1(n8479), .C2(n8551), .A(n8478), .B(n8477), .ZN(
        P2_U3474) );
  MUX2_X1 U10092 ( .A(n8480), .B(P2_REG1_REG_0__SCAN_IN), .S(n5726), .Z(
        P2_U3459) );
  INV_X1 U10093 ( .A(n8481), .ZN(n8484) );
  NAND2_X1 U10094 ( .A1(n8482), .A2(n9946), .ZN(n8486) );
  NAND2_X1 U10095 ( .A1(n9944), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8483) );
  OAI211_X1 U10096 ( .C1(n8484), .C2(n8530), .A(n8486), .B(n8483), .ZN(
        P2_U3458) );
  NAND2_X1 U10097 ( .A1(n8485), .A2(n8546), .ZN(n8487) );
  OAI211_X1 U10098 ( .C1(n5666), .C2(n9946), .A(n8487), .B(n8486), .ZN(
        P2_U3457) );
  MUX2_X1 U10099 ( .A(n10237), .B(n8488), .S(n9946), .Z(n8489) );
  OAI21_X1 U10100 ( .B1(n8490), .B2(n8550), .A(n8489), .ZN(P2_U3455) );
  INV_X1 U10101 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8492) );
  MUX2_X1 U10102 ( .A(n8492), .B(n8491), .S(n9946), .Z(n8493) );
  MUX2_X1 U10103 ( .A(n10243), .B(n8495), .S(n9946), .Z(n8498) );
  NAND2_X1 U10104 ( .A1(n8496), .A2(n8546), .ZN(n8497) );
  OAI211_X1 U10105 ( .C1(n8499), .C2(n8550), .A(n8498), .B(n8497), .ZN(
        P2_U3453) );
  MUX2_X1 U10106 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8500), .S(n9946), .Z(n8504) );
  OAI22_X1 U10107 ( .A1(n8502), .A2(n8550), .B1(n8501), .B2(n8530), .ZN(n8503)
         );
  OR2_X1 U10108 ( .A1(n8504), .A2(n8503), .ZN(P2_U3451) );
  INV_X1 U10109 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8506) );
  MUX2_X1 U10110 ( .A(n8506), .B(n8505), .S(n9946), .Z(n8509) );
  NAND2_X1 U10111 ( .A1(n8507), .A2(n8546), .ZN(n8508) );
  OAI211_X1 U10112 ( .C1(n8510), .C2(n8550), .A(n8509), .B(n8508), .ZN(
        P2_U3450) );
  INV_X1 U10113 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8512) );
  MUX2_X1 U10114 ( .A(n8512), .B(n8511), .S(n9946), .Z(n8515) );
  NAND2_X1 U10115 ( .A1(n8513), .A2(n8546), .ZN(n8514) );
  OAI211_X1 U10116 ( .C1(n8516), .C2(n8550), .A(n8515), .B(n8514), .ZN(
        P2_U3448) );
  MUX2_X1 U10117 ( .A(n10127), .B(n8517), .S(n9946), .Z(n8520) );
  NAND2_X1 U10118 ( .A1(n8518), .A2(n8546), .ZN(n8519) );
  OAI211_X1 U10119 ( .C1(n8521), .C2(n8550), .A(n8520), .B(n8519), .ZN(
        P2_U3447) );
  MUX2_X1 U10120 ( .A(n10170), .B(n8522), .S(n9946), .Z(n8525) );
  NAND2_X1 U10121 ( .A1(n8523), .A2(n8546), .ZN(n8524) );
  OAI211_X1 U10122 ( .C1(n8526), .C2(n8550), .A(n8525), .B(n8524), .ZN(
        P2_U3446) );
  MUX2_X1 U10123 ( .A(n8528), .B(n8527), .S(n9946), .Z(n8529) );
  OAI21_X1 U10124 ( .B1(n8531), .B2(n8530), .A(n8529), .ZN(P2_U3444) );
  INV_X1 U10125 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8533) );
  MUX2_X1 U10126 ( .A(n8533), .B(n8532), .S(n9946), .Z(n8536) );
  NAND2_X1 U10127 ( .A1(n8534), .A2(n8546), .ZN(n8535) );
  OAI211_X1 U10128 ( .C1(n8537), .C2(n8550), .A(n8536), .B(n8535), .ZN(
        P2_U3441) );
  INV_X1 U10129 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U10130 ( .A(n8539), .B(n8538), .S(n9946), .Z(n8542) );
  NAND2_X1 U10131 ( .A1(n8540), .A2(n8546), .ZN(n8541) );
  OAI211_X1 U10132 ( .C1(n8543), .C2(n8550), .A(n8542), .B(n8541), .ZN(
        P2_U3438) );
  INV_X1 U10133 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8545) );
  MUX2_X1 U10134 ( .A(n8545), .B(n8544), .S(n9946), .Z(n8549) );
  NAND2_X1 U10135 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  OAI211_X1 U10136 ( .C1(n8551), .C2(n8550), .A(n8549), .B(n8548), .ZN(
        P2_U3435) );
  INV_X1 U10137 ( .A(n8552), .ZN(n9471) );
  NAND3_X1 U10138 ( .A1(n8554), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8556) );
  OAI22_X1 U10139 ( .A1(n8553), .A2(n8556), .B1(n6298), .B2(n8555), .ZN(n8557)
         );
  INV_X1 U10140 ( .A(n8557), .ZN(n8558) );
  OAI21_X1 U10141 ( .B1(n9471), .B2(n8562), .A(n8558), .ZN(P2_U3264) );
  AOI21_X1 U10142 ( .B1(n8560), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8559), .ZN(
        n8561) );
  OAI21_X1 U10143 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(P2_U3267) );
  MUX2_X1 U10144 ( .A(n8564), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10145 ( .A1(n8726), .A2(n4574), .ZN(n8568) );
  NAND2_X1 U10146 ( .A1(n9060), .A2(n6773), .ZN(n8567) );
  NAND2_X1 U10147 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  XNOR2_X1 U10148 ( .A(n8569), .B(n8681), .ZN(n8573) );
  NOR2_X1 U10149 ( .A1(n8570), .A2(n6361), .ZN(n8571) );
  AOI21_X1 U10150 ( .B1(n8726), .B2(n6773), .A(n8571), .ZN(n8572) );
  NAND2_X1 U10151 ( .A1(n8573), .A2(n8572), .ZN(n8720) );
  AND2_X1 U10152 ( .A1(n9059), .A2(n8635), .ZN(n8574) );
  AOI21_X1 U10153 ( .B1(n8575), .B2(n6773), .A(n8574), .ZN(n8577) );
  AOI22_X1 U10154 ( .A1(n8575), .A2(n4574), .B1(n6773), .B2(n9059), .ZN(n8576)
         );
  XNOR2_X1 U10155 ( .A(n8576), .B(n6422), .ZN(n8578) );
  XOR2_X1 U10156 ( .A(n8577), .B(n8578), .Z(n8731) );
  AOI22_X1 U10157 ( .A1(n9459), .A2(n4574), .B1(n6773), .B2(n9058), .ZN(n8579)
         );
  XNOR2_X1 U10158 ( .A(n8579), .B(n6466), .ZN(n8781) );
  INV_X1 U10159 ( .A(n8781), .ZN(n8581) );
  AOI22_X1 U10160 ( .A1(n9459), .A2(n6773), .B1(n8635), .B2(n9058), .ZN(n8780)
         );
  OAI21_X1 U10161 ( .B1(n8582), .B2(n8581), .A(n8580), .ZN(n8673) );
  AND2_X1 U10162 ( .A1(n8785), .A2(n8635), .ZN(n8583) );
  AOI21_X1 U10163 ( .B1(n9399), .B2(n6773), .A(n8583), .ZN(n8587) );
  NAND2_X1 U10164 ( .A1(n9399), .A2(n4574), .ZN(n8585) );
  NAND2_X1 U10165 ( .A1(n8785), .A2(n6773), .ZN(n8584) );
  NAND2_X1 U10166 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  XNOR2_X1 U10167 ( .A(n8586), .B(n6422), .ZN(n8589) );
  XOR2_X1 U10168 ( .A(n8587), .B(n8589), .Z(n8672) );
  INV_X1 U10169 ( .A(n8587), .ZN(n8588) );
  NAND2_X1 U10170 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  OAI22_X1 U10171 ( .A1(n9301), .A2(n8629), .B1(n8591), .B2(n6361), .ZN(n8593)
         );
  AOI22_X1 U10172 ( .A1(n9450), .A2(n4574), .B1(n6773), .B2(n9057), .ZN(n8592)
         );
  XNOR2_X1 U10173 ( .A(n8592), .B(n6466), .ZN(n8595) );
  XOR2_X1 U10174 ( .A(n8593), .B(n8595), .Z(n8762) );
  INV_X1 U10175 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U10176 ( .A1(n9390), .A2(n4574), .ZN(n8597) );
  NAND2_X1 U10177 ( .A1(n9056), .A2(n6773), .ZN(n8596) );
  NAND2_X1 U10178 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  XNOR2_X1 U10179 ( .A(n8598), .B(n8681), .ZN(n8701) );
  INV_X1 U10180 ( .A(n8701), .ZN(n8601) );
  AND2_X1 U10181 ( .A1(n9056), .A2(n8635), .ZN(n8599) );
  AOI21_X1 U10182 ( .B1(n9390), .B2(n6773), .A(n8599), .ZN(n8700) );
  INV_X1 U10183 ( .A(n8700), .ZN(n8600) );
  NAND2_X1 U10184 ( .A1(n8601), .A2(n8600), .ZN(n8614) );
  OAI22_X1 U10185 ( .A1(n9443), .A2(n8630), .B1(n8668), .B2(n8629), .ZN(n8602)
         );
  XNOR2_X1 U10186 ( .A(n8602), .B(n6422), .ZN(n8613) );
  NAND2_X1 U10187 ( .A1(n8701), .A2(n8700), .ZN(n8612) );
  NAND2_X1 U10188 ( .A1(n9379), .A2(n4574), .ZN(n8604) );
  NAND2_X1 U10189 ( .A1(n9054), .A2(n6773), .ZN(n8603) );
  NAND2_X1 U10190 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  XNOR2_X1 U10191 ( .A(n8605), .B(n8681), .ZN(n8607) );
  AND2_X1 U10192 ( .A1(n9054), .A2(n8635), .ZN(n8606) );
  AOI21_X1 U10193 ( .B1(n9379), .B2(n6773), .A(n8606), .ZN(n8608) );
  NAND2_X1 U10194 ( .A1(n8607), .A2(n8608), .ZN(n8743) );
  INV_X1 U10195 ( .A(n8607), .ZN(n8610) );
  INV_X1 U10196 ( .A(n8608), .ZN(n8609) );
  NAND2_X1 U10197 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U10198 ( .A1(n8743), .A2(n8611), .ZN(n8663) );
  INV_X1 U10199 ( .A(n8612), .ZN(n8616) );
  INV_X1 U10200 ( .A(n8613), .ZN(n8615) );
  OAI22_X1 U10201 ( .A1(n9443), .A2(n8629), .B1(n8668), .B2(n6361), .ZN(n8772)
         );
  NAND2_X1 U10202 ( .A1(n8744), .A2(n8743), .ZN(n8625) );
  OAI22_X1 U10203 ( .A1(n9242), .A2(n8630), .B1(n8713), .B2(n8629), .ZN(n8617)
         );
  XNOR2_X1 U10204 ( .A(n8617), .B(n8681), .ZN(n8620) );
  OR2_X1 U10205 ( .A1(n9242), .A2(n8629), .ZN(n8619) );
  NAND2_X1 U10206 ( .A1(n9053), .A2(n8635), .ZN(n8618) );
  AND2_X1 U10207 ( .A1(n8619), .A2(n8618), .ZN(n8621) );
  NAND2_X1 U10208 ( .A1(n8620), .A2(n8621), .ZN(n8626) );
  INV_X1 U10209 ( .A(n8620), .ZN(n8623) );
  INV_X1 U10210 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U10211 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  AND2_X1 U10212 ( .A1(n8626), .A2(n8624), .ZN(n8741) );
  NAND2_X1 U10213 ( .A1(n8625), .A2(n8741), .ZN(n8746) );
  OR2_X1 U10214 ( .A1(n9428), .A2(n8629), .ZN(n8628) );
  OR2_X1 U10215 ( .A1(n8801), .A2(n6361), .ZN(n8627) );
  NAND2_X1 U10216 ( .A1(n8628), .A2(n8627), .ZN(n8637) );
  OAI22_X1 U10217 ( .A1(n9428), .A2(n8630), .B1(n8801), .B2(n8629), .ZN(n8631)
         );
  XNOR2_X1 U10218 ( .A(n8631), .B(n6466), .ZN(n8638) );
  XOR2_X1 U10219 ( .A(n8637), .B(n8638), .Z(n8710) );
  NAND2_X1 U10220 ( .A1(n9362), .A2(n4574), .ZN(n8633) );
  NAND2_X1 U10221 ( .A1(n9051), .A2(n6773), .ZN(n8632) );
  NAND2_X1 U10222 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  XNOR2_X1 U10223 ( .A(n8634), .B(n8681), .ZN(n8640) );
  AND2_X1 U10224 ( .A1(n9051), .A2(n8635), .ZN(n8636) );
  AOI21_X1 U10225 ( .B1(n9362), .B2(n6773), .A(n8636), .ZN(n8641) );
  XNOR2_X1 U10226 ( .A(n8640), .B(n8641), .ZN(n8794) );
  NOR2_X1 U10227 ( .A1(n8638), .A2(n8637), .ZN(n8795) );
  NOR2_X1 U10228 ( .A1(n8794), .A2(n8795), .ZN(n8639) );
  INV_X1 U10229 ( .A(n8640), .ZN(n8643) );
  INV_X1 U10230 ( .A(n8641), .ZN(n8642) );
  NAND2_X1 U10231 ( .A1(n8643), .A2(n8642), .ZN(n8654) );
  NAND2_X1 U10232 ( .A1(n9188), .A2(n4574), .ZN(n8646) );
  NAND2_X1 U10233 ( .A1(n8644), .A2(n6773), .ZN(n8645) );
  NAND2_X1 U10234 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  XNOR2_X1 U10235 ( .A(n8647), .B(n8681), .ZN(n8650) );
  INV_X1 U10236 ( .A(n8650), .ZN(n8652) );
  NOR2_X1 U10237 ( .A1(n8799), .A2(n6361), .ZN(n8648) );
  AOI21_X1 U10238 ( .B1(n9188), .B2(n6773), .A(n8648), .ZN(n8649) );
  INV_X1 U10239 ( .A(n8649), .ZN(n8651) );
  AOI21_X1 U10240 ( .B1(n8652), .B2(n8651), .A(n8693), .ZN(n8653) );
  AOI21_X1 U10241 ( .B1(n8796), .B2(n8654), .A(n8653), .ZN(n8657) );
  INV_X1 U10242 ( .A(n8653), .ZN(n8656) );
  INV_X1 U10243 ( .A(n8654), .ZN(n8655) );
  OAI21_X1 U10244 ( .B1(n8657), .B2(n8687), .A(n8797), .ZN(n8662) );
  NOR2_X1 U10245 ( .A1(n8803), .A2(n9189), .ZN(n8660) );
  AOI22_X1 U10246 ( .A1(n9050), .A2(n8784), .B1(n9042), .B2(n9051), .ZN(n9184)
         );
  OAI22_X1 U10247 ( .A1(n9184), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8658), .ZN(n8659) );
  AOI211_X1 U10248 ( .C1(n9188), .C2(n8790), .A(n8660), .B(n8659), .ZN(n8661)
         );
  NAND2_X1 U10249 ( .A1(n8662), .A2(n8661), .ZN(P1_U3214) );
  INV_X1 U10250 ( .A(n8744), .ZN(n8667) );
  INV_X1 U10251 ( .A(n8663), .ZN(n8664) );
  AOI21_X1 U10252 ( .B1(n8665), .B2(n4434), .A(n8664), .ZN(n8666) );
  OAI21_X1 U10253 ( .B1(n8667), .B2(n8666), .A(n8797), .ZN(n8671) );
  OAI22_X1 U10254 ( .A1(n8713), .A2(n8798), .B1(n8668), .B2(n8800), .ZN(n9250)
         );
  OAI22_X1 U10255 ( .A1(n8803), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10052), .ZN(n8669) );
  AOI21_X1 U10256 ( .B1(n9250), .B2(n8805), .A(n8669), .ZN(n8670) );
  OAI211_X1 U10257 ( .C1(n9259), .C2(n8807), .A(n8671), .B(n8670), .ZN(
        P1_U3216) );
  AOI21_X1 U10258 ( .B1(n8673), .B2(n8672), .A(n8792), .ZN(n8675) );
  NAND2_X1 U10259 ( .A1(n8675), .A2(n8674), .ZN(n8678) );
  AOI22_X1 U10260 ( .A1(n9057), .A2(n8784), .B1(n9042), .B2(n9058), .ZN(n9313)
         );
  OAI22_X1 U10261 ( .A1(n9313), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10167), .ZN(n8676) );
  AOI21_X1 U10262 ( .B1(n9320), .B2(n8767), .A(n8676), .ZN(n8677) );
  OAI211_X1 U10263 ( .C1(n9325), .C2(n8807), .A(n8678), .B(n8677), .ZN(
        P1_U3219) );
  NAND2_X1 U10264 ( .A1(n8692), .A2(n4574), .ZN(n8680) );
  NAND2_X1 U10265 ( .A1(n9050), .A2(n6773), .ZN(n8679) );
  NAND2_X1 U10266 ( .A1(n8680), .A2(n8679), .ZN(n8682) );
  XNOR2_X1 U10267 ( .A(n8682), .B(n8681), .ZN(n8686) );
  NAND2_X1 U10268 ( .A1(n8692), .A2(n6773), .ZN(n8683) );
  OAI21_X1 U10269 ( .B1(n8684), .B2(n6361), .A(n8683), .ZN(n8685) );
  XNOR2_X1 U10270 ( .A(n8686), .B(n8685), .ZN(n8694) );
  NAND3_X1 U10271 ( .A1(n8687), .A2(n8797), .A3(n8694), .ZN(n8697) );
  AOI22_X1 U10272 ( .A1(n8688), .A2(n8805), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8689) );
  OAI21_X1 U10273 ( .B1(n8690), .B2(n8803), .A(n8689), .ZN(n8691) );
  AOI21_X1 U10274 ( .B1(n8692), .B2(n8790), .A(n8691), .ZN(n8696) );
  NAND3_X1 U10275 ( .A1(n8694), .A2(n8797), .A3(n8693), .ZN(n8695) );
  NAND4_X1 U10276 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(
        P1_U3220) );
  XNOR2_X1 U10277 ( .A(n8701), .B(n8700), .ZN(n8702) );
  XNOR2_X1 U10278 ( .A(n8699), .B(n8702), .ZN(n8707) );
  NOR2_X1 U10279 ( .A1(n8803), .A2(n9286), .ZN(n8705) );
  AOI22_X1 U10280 ( .A1(n9055), .A2(n8784), .B1(n9042), .B2(n9057), .ZN(n9281)
         );
  INV_X1 U10281 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8703) );
  OAI22_X1 U10282 ( .A1(n9281), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8703), .ZN(n8704) );
  AOI211_X1 U10283 ( .C1(n9390), .C2(n8790), .A(n8705), .B(n8704), .ZN(n8706)
         );
  OAI21_X1 U10284 ( .B1(n8707), .B2(n8792), .A(n8706), .ZN(P1_U3223) );
  OAI21_X1 U10285 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8711) );
  NAND2_X1 U10286 ( .A1(n8711), .A2(n8797), .ZN(n8716) );
  OAI22_X1 U10287 ( .A1(n8713), .A2(n8800), .B1(n8712), .B2(n8798), .ZN(n9216)
         );
  OAI22_X1 U10288 ( .A1(n9223), .A2(n8803), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10093), .ZN(n8714) );
  AOI21_X1 U10289 ( .B1(n9216), .B2(n8805), .A(n8714), .ZN(n8715) );
  OAI211_X1 U10290 ( .C1(n9428), .C2(n8807), .A(n8716), .B(n8715), .ZN(
        P1_U3225) );
  INV_X1 U10291 ( .A(n8717), .ZN(n8721) );
  NAND2_X1 U10292 ( .A1(n4508), .A2(n8720), .ZN(n8718) );
  AOI22_X1 U10293 ( .A1(n8721), .A2(n8720), .B1(n8719), .B2(n8718), .ZN(n8728)
         );
  AOI22_X1 U10294 ( .A1(n8805), .A2(n8722), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n8723) );
  OAI21_X1 U10295 ( .B1(n8724), .B2(n8803), .A(n8723), .ZN(n8725) );
  AOI21_X1 U10296 ( .B1(n8726), .B2(n8790), .A(n8725), .ZN(n8727) );
  OAI21_X1 U10297 ( .B1(n8728), .B2(n8792), .A(n8727), .ZN(P1_U3226) );
  OAI21_X1 U10298 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n8732) );
  NAND2_X1 U10299 ( .A1(n8732), .A2(n8797), .ZN(n8738) );
  OAI21_X1 U10300 ( .B1(n8734), .B2(n8775), .A(n8733), .ZN(n8735) );
  AOI21_X1 U10301 ( .B1(n8736), .B2(n8767), .A(n8735), .ZN(n8737) );
  OAI211_X1 U10302 ( .C1(n8739), .C2(n8807), .A(n8738), .B(n8737), .ZN(
        P1_U3228) );
  INV_X1 U10303 ( .A(n8801), .ZN(n9052) );
  AOI22_X1 U10304 ( .A1(n9052), .A2(n8784), .B1(n9042), .B2(n9054), .ZN(n9235)
         );
  AOI22_X1 U10305 ( .A1(n9239), .A2(n8767), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8740) );
  OAI21_X1 U10306 ( .B1(n9235), .B2(n8775), .A(n8740), .ZN(n8748) );
  INV_X1 U10307 ( .A(n8741), .ZN(n8742) );
  NAND3_X1 U10308 ( .A1(n8744), .A2(n8743), .A3(n8742), .ZN(n8745) );
  AOI21_X1 U10309 ( .B1(n8746), .B2(n8745), .A(n8792), .ZN(n8747) );
  AOI211_X1 U10310 ( .C1(n9432), .C2(n8790), .A(n8748), .B(n8747), .ZN(n8749)
         );
  INV_X1 U10311 ( .A(n8749), .ZN(P1_U3229) );
  OAI211_X1 U10312 ( .C1(n8752), .C2(n8751), .A(n8750), .B(n8797), .ZN(n8760)
         );
  AOI21_X1 U10313 ( .B1(n8790), .B2(n8754), .A(n8753), .ZN(n8759) );
  OR2_X1 U10314 ( .A1(n8803), .A2(n8755), .ZN(n8758) );
  NAND2_X1 U10315 ( .A1(n8756), .A2(n8805), .ZN(n8757) );
  NAND4_X1 U10316 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), .ZN(
        P1_U3230) );
  AOI21_X1 U10317 ( .B1(n8762), .B2(n8761), .A(n4505), .ZN(n8769) );
  AND2_X1 U10318 ( .A1(n8785), .A2(n9042), .ZN(n8763) );
  AOI21_X1 U10319 ( .B1(n9056), .B2(n8784), .A(n8763), .ZN(n9296) );
  OAI22_X1 U10320 ( .A1(n9296), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8764), .ZN(n8766) );
  NOR2_X1 U10321 ( .A1(n9301), .A2(n8807), .ZN(n8765) );
  AOI211_X1 U10322 ( .C1(n8767), .C2(n9302), .A(n8766), .B(n8765), .ZN(n8768)
         );
  OAI21_X1 U10323 ( .B1(n8769), .B2(n8792), .A(n8768), .ZN(P1_U3233) );
  NAND2_X1 U10324 ( .A1(n4434), .A2(n8770), .ZN(n8771) );
  XOR2_X1 U10325 ( .A(n8772), .B(n8771), .Z(n8779) );
  NOR2_X1 U10326 ( .A1(n8803), .A2(n9270), .ZN(n8777) );
  AND2_X1 U10327 ( .A1(n9056), .A2(n9042), .ZN(n8773) );
  AOI21_X1 U10328 ( .B1(n9054), .B2(n8784), .A(n8773), .ZN(n9266) );
  OAI22_X1 U10329 ( .A1(n9266), .A2(n8775), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8774), .ZN(n8776) );
  AOI211_X1 U10330 ( .C1(n9269), .C2(n8790), .A(n8777), .B(n8776), .ZN(n8778)
         );
  OAI21_X1 U10331 ( .B1(n8779), .B2(n8792), .A(n8778), .ZN(P1_U3235) );
  XNOR2_X1 U10332 ( .A(n8781), .B(n8780), .ZN(n8782) );
  XNOR2_X1 U10333 ( .A(n8783), .B(n8782), .ZN(n8793) );
  NAND2_X1 U10334 ( .A1(n9059), .A2(n9042), .ZN(n8787) );
  NAND2_X1 U10335 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NAND2_X1 U10336 ( .A1(n8787), .A2(n8786), .ZN(n9332) );
  AOI22_X1 U10337 ( .A1(n8805), .A2(n9332), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8788) );
  OAI21_X1 U10338 ( .B1(n9340), .B2(n8803), .A(n8788), .ZN(n8789) );
  AOI21_X1 U10339 ( .B1(n9459), .B2(n8790), .A(n8789), .ZN(n8791) );
  OAI21_X1 U10340 ( .B1(n8793), .B2(n8792), .A(n8791), .ZN(P1_U3238) );
  INV_X1 U10341 ( .A(n9362), .ZN(n9204) );
  OAI22_X1 U10342 ( .A1(n8801), .A2(n8800), .B1(n8799), .B2(n8798), .ZN(n9209)
         );
  INV_X1 U10343 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8802) );
  OAI22_X1 U10344 ( .A1(n8803), .A2(n9201), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8802), .ZN(n8804) );
  AOI21_X1 U10345 ( .B1(n9209), .B2(n8805), .A(n8804), .ZN(n8806) );
  NAND2_X1 U10346 ( .A1(n4685), .A2(n9021), .ZN(n9039) );
  NAND2_X1 U10347 ( .A1(n8809), .A2(n8808), .ZN(n9010) );
  NAND2_X1 U10348 ( .A1(n9009), .A2(n9002), .ZN(n8891) );
  NAND2_X1 U10349 ( .A1(n8993), .A2(n8810), .ZN(n8991) );
  NAND2_X1 U10350 ( .A1(n8991), .A2(n9234), .ZN(n8811) );
  NAND2_X1 U10351 ( .A1(n8997), .A2(n8811), .ZN(n8812) );
  NAND2_X1 U10352 ( .A1(n8812), .A2(n8998), .ZN(n8813) );
  AND2_X1 U10353 ( .A1(n9205), .A2(n8813), .ZN(n8836) );
  NOR2_X1 U10354 ( .A1(n9390), .A2(n8814), .ZN(n8837) );
  AND2_X1 U10355 ( .A1(n8987), .A2(n8966), .ZN(n8979) );
  AND2_X1 U10356 ( .A1(n9234), .A2(n8815), .ZN(n8990) );
  OAI211_X1 U10357 ( .C1(n8837), .C2(n8979), .A(n8998), .B(n8990), .ZN(n8816)
         );
  AOI21_X1 U10358 ( .B1(n8836), .B2(n8816), .A(n4632), .ZN(n8817) );
  NOR2_X1 U10359 ( .A1(n8891), .A2(n8817), .ZN(n8818) );
  NOR2_X1 U10360 ( .A1(n9010), .A2(n8818), .ZN(n8890) );
  NAND2_X1 U10361 ( .A1(n8970), .A2(n8819), .ZN(n8848) );
  AOI21_X1 U10362 ( .B1(n8965), .B2(n8848), .A(n4869), .ZN(n8967) );
  NAND2_X1 U10363 ( .A1(n9074), .A2(n8820), .ZN(n8821) );
  AND4_X1 U10364 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n8827)
         );
  NAND4_X1 U10365 ( .A1(n8827), .A2(n8826), .A3(n8911), .A4(n8825), .ZN(n8828)
         );
  AOI211_X1 U10366 ( .C1(n4448), .C2(n8828), .A(n4607), .B(n4501), .ZN(n8829)
         );
  NAND2_X1 U10367 ( .A1(n8931), .A2(n8928), .ZN(n8947) );
  NOR2_X1 U10368 ( .A1(n8829), .A2(n8947), .ZN(n8830) );
  NAND2_X1 U10369 ( .A1(n8933), .A2(n8929), .ZN(n8948) );
  OAI211_X1 U10370 ( .C1(n8830), .C2(n8948), .A(n8951), .B(n8955), .ZN(n8831)
         );
  NAND3_X1 U10371 ( .A1(n8831), .A2(n8952), .A3(n8958), .ZN(n8833) );
  AND2_X1 U10372 ( .A1(n8960), .A2(n8832), .ZN(n8938) );
  AOI211_X1 U10373 ( .C1(n8833), .C2(n8938), .A(n8941), .B(n4586), .ZN(n8834)
         );
  OAI211_X1 U10374 ( .C1(n8835), .C2(n8834), .A(n8965), .B(n8969), .ZN(n8839)
         );
  INV_X1 U10375 ( .A(n8836), .ZN(n8838) );
  INV_X1 U10376 ( .A(n8837), .ZN(n8986) );
  NAND2_X1 U10377 ( .A1(n8986), .A2(n8978), .ZN(n8981) );
  OR2_X1 U10378 ( .A1(n8838), .A2(n8981), .ZN(n8888) );
  AOI21_X1 U10379 ( .B1(n8967), .B2(n8839), .A(n8888), .ZN(n8841) );
  INV_X1 U10380 ( .A(n8891), .ZN(n8840) );
  OAI21_X1 U10381 ( .B1(n8841), .B2(n4859), .A(n8840), .ZN(n8842) );
  NAND2_X1 U10382 ( .A1(n9016), .A2(n9012), .ZN(n8887) );
  AOI21_X1 U10383 ( .B1(n8890), .B2(n8842), .A(n8887), .ZN(n8843) );
  INV_X1 U10384 ( .A(n9049), .ZN(n9025) );
  NAND2_X1 U10385 ( .A1(n9167), .A2(n9025), .ZN(n8882) );
  NAND2_X1 U10386 ( .A1(n8882), .A2(n9017), .ZN(n8893) );
  OR2_X1 U10387 ( .A1(n9167), .A2(n9025), .ZN(n8897) );
  OAI21_X1 U10388 ( .B1(n8843), .B2(n8893), .A(n8897), .ZN(n8845) );
  AND2_X1 U10389 ( .A1(n8844), .A2(n8896), .ZN(n8847) );
  AOI21_X1 U10390 ( .B1(n9039), .B2(n8845), .A(n8847), .ZN(n8846) );
  XNOR2_X1 U10391 ( .A(n8846), .B(n4431), .ZN(n8908) );
  NAND2_X1 U10392 ( .A1(n8977), .A2(n8971), .ZN(n9308) );
  INV_X1 U10393 ( .A(n9308), .ZN(n9311) );
  INV_X1 U10394 ( .A(n8848), .ZN(n8875) );
  INV_X1 U10395 ( .A(n8850), .ZN(n8865) );
  AND4_X1 U10396 ( .A1(n8854), .A2(n9035), .A3(n8853), .A4(n8852), .ZN(n8861)
         );
  INV_X1 U10397 ( .A(n8856), .ZN(n8860) );
  NOR2_X1 U10398 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND4_X1 U10399 ( .A1(n8861), .A2(n4808), .A3(n8860), .A4(n8859), .ZN(n8863)
         );
  NOR2_X1 U10400 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  NAND4_X1 U10401 ( .A1(n4817), .A2(n8865), .A3(n4640), .A4(n8864), .ZN(n8866)
         );
  NOR2_X1 U10402 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  NAND4_X1 U10403 ( .A1(n8870), .A2(n4651), .A3(n8869), .A4(n8868), .ZN(n8871)
         );
  NOR2_X1 U10404 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  AND2_X1 U10405 ( .A1(n8873), .A2(n8969), .ZN(n8874) );
  NAND4_X1 U10406 ( .A1(n9311), .A2(n8875), .A3(n8874), .A4(n9310), .ZN(n8876)
         );
  NOR2_X1 U10407 ( .A1(n9294), .A2(n8876), .ZN(n8877) );
  INV_X1 U10408 ( .A(n9277), .ZN(n9279) );
  NAND4_X1 U10409 ( .A1(n9248), .A2(n9262), .A3(n8877), .A4(n9279), .ZN(n8878)
         );
  NOR2_X1 U10410 ( .A1(n9230), .A2(n8878), .ZN(n8879) );
  AND4_X1 U10411 ( .A1(n9182), .A2(n6129), .A3(n9221), .A4(n8879), .ZN(n8880)
         );
  NAND4_X1 U10412 ( .A1(n8897), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n8883)
         );
  NOR2_X1 U10413 ( .A1(n8883), .A2(n9014), .ZN(n8884) );
  NAND3_X1 U10414 ( .A1(n9033), .A2(n9039), .A3(n8884), .ZN(n8903) );
  INV_X1 U10415 ( .A(n8903), .ZN(n8886) );
  NOR2_X1 U10416 ( .A1(n4431), .A2(n8885), .ZN(n9030) );
  AOI21_X1 U10417 ( .B1(n8886), .B2(n9030), .A(n9044), .ZN(n8906) );
  INV_X1 U10418 ( .A(n8887), .ZN(n8895) );
  INV_X1 U10419 ( .A(n8888), .ZN(n8889) );
  AOI21_X1 U10420 ( .B1(n8889), .B2(n9295), .A(n4859), .ZN(n8892) );
  OAI21_X1 U10421 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8894) );
  AOI21_X1 U10422 ( .B1(n8895), .B2(n8894), .A(n8893), .ZN(n8899) );
  NOR2_X1 U10423 ( .A1(n8897), .A2(n8896), .ZN(n8898) );
  OAI22_X1 U10424 ( .A1(n8899), .A2(n8898), .B1(n9420), .B2(n9021), .ZN(n8902)
         );
  INV_X1 U10425 ( .A(n9039), .ZN(n8901) );
  OAI211_X1 U10426 ( .C1(n8902), .C2(n8901), .A(n8900), .B(n9033), .ZN(n8904)
         );
  NAND4_X1 U10427 ( .A1(n8904), .A2(n8907), .A3(n8903), .A4(n4431), .ZN(n8905)
         );
  OAI211_X1 U10428 ( .C1(n8908), .C2(n8907), .A(n8906), .B(n8905), .ZN(n9048)
         );
  INV_X1 U10429 ( .A(n8909), .ZN(n8912) );
  OAI211_X1 U10430 ( .C1(n8913), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8915)
         );
  NAND2_X1 U10431 ( .A1(n8915), .A2(n8914), .ZN(n8917) );
  MUX2_X1 U10432 ( .A(n8917), .B(n8916), .S(n9020), .Z(n8918) );
  INV_X1 U10433 ( .A(n8919), .ZN(n8922) );
  NAND2_X1 U10434 ( .A1(n8926), .A2(n8920), .ZN(n8921) );
  INV_X1 U10435 ( .A(n8923), .ZN(n8924) );
  INV_X1 U10436 ( .A(n8926), .ZN(n8927) );
  AOI21_X1 U10437 ( .B1(n8946), .B2(n8944), .A(n8927), .ZN(n8930) );
  OAI211_X1 U10438 ( .C1(n8930), .C2(n4637), .A(n8945), .B(n8929), .ZN(n8932)
         );
  NAND3_X1 U10439 ( .A1(n8932), .A2(n8951), .A3(n8931), .ZN(n8934) );
  NAND2_X1 U10440 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  NAND2_X1 U10441 ( .A1(n8935), .A2(n8955), .ZN(n8940) );
  INV_X1 U10442 ( .A(n8952), .ZN(n8936) );
  NOR2_X1 U10443 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  NAND2_X1 U10444 ( .A1(n8963), .A2(n8941), .ZN(n8942) );
  NAND2_X1 U10445 ( .A1(n8942), .A2(n8962), .ZN(n8943) );
  INV_X1 U10446 ( .A(n8947), .ZN(n8949) );
  AOI21_X1 U10447 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8954) );
  INV_X1 U10448 ( .A(n8951), .ZN(n8953) );
  OAI21_X1 U10449 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(n8956) );
  NAND3_X1 U10450 ( .A1(n8956), .A2(n4651), .A3(n8955), .ZN(n8959) );
  NAND3_X1 U10451 ( .A1(n8959), .A2(n8958), .A3(n8957), .ZN(n8961) );
  INV_X1 U10452 ( .A(n8965), .ZN(n8968) );
  OAI211_X1 U10453 ( .C1(n8974), .C2(n8968), .A(n8967), .B(n8966), .ZN(n8976)
         );
  AND2_X1 U10454 ( .A1(n9310), .A2(n8969), .ZN(n8973) );
  NAND2_X1 U10455 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  AOI21_X1 U10456 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8975) );
  MUX2_X1 U10457 ( .A(n8976), .B(n8975), .S(n9020), .Z(n8985) );
  AOI21_X1 U10458 ( .B1(n8978), .B2(n8977), .A(n4616), .ZN(n8984) );
  INV_X1 U10459 ( .A(n8979), .ZN(n8980) );
  MUX2_X1 U10460 ( .A(n8981), .B(n8980), .S(n9020), .Z(n8982) );
  INV_X1 U10461 ( .A(n8982), .ZN(n8983) );
  OAI21_X1 U10462 ( .B1(n8985), .B2(n8984), .A(n8983), .ZN(n8989) );
  MUX2_X1 U10463 ( .A(n8987), .B(n8986), .S(n9020), .Z(n8988) );
  AOI21_X1 U10464 ( .B1(n8989), .B2(n8988), .A(n9264), .ZN(n8996) );
  INV_X1 U10465 ( .A(n8990), .ZN(n8992) );
  MUX2_X1 U10466 ( .A(n8992), .B(n8991), .S(n9020), .Z(n8995) );
  INV_X1 U10467 ( .A(n9230), .ZN(n9233) );
  MUX2_X1 U10468 ( .A(n8993), .B(n9234), .S(n9020), .Z(n8994) );
  MUX2_X1 U10469 ( .A(n8998), .B(n8997), .S(n9020), .Z(n8999) );
  NAND2_X1 U10470 ( .A1(n9003), .A2(n9000), .ZN(n9001) );
  NAND2_X1 U10471 ( .A1(n9001), .A2(n9002), .ZN(n9006) );
  NAND2_X1 U10472 ( .A1(n9002), .A2(n9205), .ZN(n9004) );
  NAND2_X1 U10473 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  MUX2_X1 U10474 ( .A(n9006), .B(n9005), .S(n4616), .Z(n9008) );
  INV_X1 U10475 ( .A(n9009), .ZN(n9007) );
  OAI21_X1 U10476 ( .B1(n9010), .B2(n9009), .A(n9012), .ZN(n9011) );
  AOI22_X1 U10477 ( .A1(n9013), .A2(n9012), .B1(n4616), .B2(n9011), .ZN(n9015)
         );
  OR2_X1 U10478 ( .A1(n9015), .A2(n9014), .ZN(n9019) );
  MUX2_X1 U10479 ( .A(n9017), .B(n9016), .S(n4616), .Z(n9018) );
  NAND2_X1 U10480 ( .A1(n9019), .A2(n9018), .ZN(n9024) );
  MUX2_X1 U10481 ( .A(n9024), .B(n9020), .S(n9167), .Z(n9023) );
  OAI21_X1 U10482 ( .B1(n4685), .B2(n9049), .A(n9021), .ZN(n9022) );
  NAND2_X1 U10483 ( .A1(n9023), .A2(n9022), .ZN(n9029) );
  MUX2_X1 U10484 ( .A(n4616), .B(n9024), .S(n9167), .Z(n9027) );
  NOR2_X1 U10485 ( .A1(n4685), .A2(n9025), .ZN(n9026) );
  NAND2_X1 U10486 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  NAND3_X1 U10487 ( .A1(n9029), .A2(n9028), .A3(n9033), .ZN(n9032) );
  INV_X1 U10488 ( .A(n9030), .ZN(n9031) );
  AOI211_X1 U10489 ( .C1(n9032), .C2(n10044), .A(n9035), .B(n9031), .ZN(n9047)
         );
  OAI21_X1 U10490 ( .B1(n9033), .B2(n4616), .A(n9032), .ZN(n9038) );
  NOR4_X1 U10491 ( .A1(n9036), .A2(n10044), .A3(n9035), .A4(n9034), .ZN(n9037)
         );
  OAI211_X1 U10492 ( .C1(n9039), .C2(n4431), .A(n9038), .B(n9037), .ZN(n9046)
         );
  NAND4_X1 U10493 ( .A1(n9042), .A2(n9667), .A3(n9041), .A4(n9040), .ZN(n9043)
         );
  OAI211_X1 U10494 ( .C1(n10044), .C2(n9044), .A(n9043), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9045) );
  OAI211_X1 U10495 ( .C1(n9048), .C2(n9047), .A(n9046), .B(n9045), .ZN(
        P1_U3242) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9049), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9050), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10498 ( .A(n9051), .B(P1_DATAO_REG_26__SCAN_IN), .S(n6670), .Z(
        P1_U3580) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9052), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10500 ( .A(n9053), .B(P1_DATAO_REG_24__SCAN_IN), .S(n6670), .Z(
        P1_U3578) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9054), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9055), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9056), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9057), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10505 ( .A(n9058), .B(P1_DATAO_REG_18__SCAN_IN), .S(n6670), .Z(
        P1_U3572) );
  MUX2_X1 U10506 ( .A(n9059), .B(P1_DATAO_REG_17__SCAN_IN), .S(n6670), .Z(
        P1_U3571) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9060), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10508 ( .A(n9061), .B(P1_DATAO_REG_15__SCAN_IN), .S(n6670), .Z(
        P1_U3569) );
  MUX2_X1 U10509 ( .A(n9062), .B(P1_DATAO_REG_14__SCAN_IN), .S(n6670), .Z(
        P1_U3568) );
  MUX2_X1 U10510 ( .A(n9063), .B(P1_DATAO_REG_13__SCAN_IN), .S(n6670), .Z(
        P1_U3567) );
  MUX2_X1 U10511 ( .A(n9064), .B(P1_DATAO_REG_12__SCAN_IN), .S(n6670), .Z(
        P1_U3566) );
  MUX2_X1 U10512 ( .A(n9065), .B(P1_DATAO_REG_11__SCAN_IN), .S(n6670), .Z(
        P1_U3565) );
  MUX2_X1 U10513 ( .A(n9066), .B(P1_DATAO_REG_10__SCAN_IN), .S(n6670), .Z(
        P1_U3564) );
  MUX2_X1 U10514 ( .A(n9067), .B(P1_DATAO_REG_9__SCAN_IN), .S(n6670), .Z(
        P1_U3563) );
  MUX2_X1 U10515 ( .A(n9068), .B(P1_DATAO_REG_8__SCAN_IN), .S(n6670), .Z(
        P1_U3562) );
  MUX2_X1 U10516 ( .A(n9069), .B(P1_DATAO_REG_7__SCAN_IN), .S(n6670), .Z(
        P1_U3561) );
  MUX2_X1 U10517 ( .A(n9070), .B(P1_DATAO_REG_6__SCAN_IN), .S(n6670), .Z(
        P1_U3560) );
  MUX2_X1 U10518 ( .A(n9071), .B(P1_DATAO_REG_5__SCAN_IN), .S(n6670), .Z(
        P1_U3559) );
  MUX2_X1 U10519 ( .A(n9072), .B(P1_DATAO_REG_3__SCAN_IN), .S(n6670), .Z(
        P1_U3557) );
  MUX2_X1 U10520 ( .A(n9073), .B(P1_DATAO_REG_2__SCAN_IN), .S(n6670), .Z(
        P1_U3556) );
  MUX2_X1 U10521 ( .A(n9074), .B(P1_DATAO_REG_1__SCAN_IN), .S(n6670), .Z(
        P1_U3555) );
  OAI211_X1 U10522 ( .C1(n9077), .C2(n9076), .A(n9605), .B(n9075), .ZN(n9085)
         );
  AOI22_X1 U10523 ( .A1(n9518), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9084) );
  NAND2_X1 U10524 ( .A1(n9612), .A2(n9078), .ZN(n9083) );
  OAI211_X1 U10525 ( .C1(n9081), .C2(n9080), .A(n9597), .B(n9079), .ZN(n9082)
         );
  NAND4_X1 U10526 ( .A1(n9085), .A2(n9084), .A3(n9083), .A4(n9082), .ZN(
        P1_U3244) );
  INV_X1 U10527 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U10528 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9086) );
  OAI21_X1 U10529 ( .B1(n9620), .B2(n9087), .A(n9086), .ZN(n9088) );
  AOI21_X1 U10530 ( .B1(n9089), .B2(n9612), .A(n9088), .ZN(n9098) );
  OAI211_X1 U10531 ( .C1(n9092), .C2(n9091), .A(n9597), .B(n9090), .ZN(n9097)
         );
  OAI211_X1 U10532 ( .C1(n9095), .C2(n9094), .A(n9605), .B(n9093), .ZN(n9096)
         );
  NAND3_X1 U10533 ( .A1(n9098), .A2(n9097), .A3(n9096), .ZN(P1_U3246) );
  INV_X1 U10534 ( .A(n9099), .ZN(n9103) );
  INV_X1 U10535 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U10536 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9100) );
  OAI21_X1 U10537 ( .B1(n9620), .B2(n9101), .A(n9100), .ZN(n9102) );
  AOI21_X1 U10538 ( .B1(n9103), .B2(n9612), .A(n9102), .ZN(n9112) );
  OAI211_X1 U10539 ( .C1(n9106), .C2(n9105), .A(n9597), .B(n9104), .ZN(n9111)
         );
  OAI211_X1 U10540 ( .C1(n9109), .C2(n9108), .A(n9605), .B(n9107), .ZN(n9110)
         );
  NAND3_X1 U10541 ( .A1(n9112), .A2(n9111), .A3(n9110), .ZN(P1_U3248) );
  INV_X1 U10542 ( .A(n9113), .ZN(n9117) );
  INV_X1 U10543 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U10544 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9114) );
  OAI21_X1 U10545 ( .B1(n9620), .B2(n9115), .A(n9114), .ZN(n9116) );
  AOI21_X1 U10546 ( .B1(n9117), .B2(n9612), .A(n9116), .ZN(n9126) );
  OAI211_X1 U10547 ( .C1(n9120), .C2(n9119), .A(n9597), .B(n9118), .ZN(n9125)
         );
  OAI211_X1 U10548 ( .C1(n9123), .C2(n9122), .A(n9605), .B(n9121), .ZN(n9124)
         );
  NAND3_X1 U10549 ( .A1(n9126), .A2(n9125), .A3(n9124), .ZN(P1_U3249) );
  OAI21_X1 U10550 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10551 ( .A1(n9130), .A2(n9597), .ZN(n9140) );
  AOI21_X1 U10552 ( .B1(n9518), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9131), .ZN(
        n9139) );
  OAI21_X1 U10553 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9135) );
  NAND2_X1 U10554 ( .A1(n9135), .A2(n9605), .ZN(n9138) );
  NAND2_X1 U10555 ( .A1(n9612), .A2(n9136), .ZN(n9137) );
  NAND4_X1 U10556 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(
        P1_U3252) );
  INV_X1 U10557 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9161) );
  AND2_X1 U10558 ( .A1(n9142), .A2(n9141), .ZN(n9608) );
  INV_X1 U10559 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9341) );
  OR2_X1 U10560 ( .A1(n9613), .A2(n9341), .ZN(n9144) );
  NAND2_X1 U10561 ( .A1(n9613), .A2(n9341), .ZN(n9143) );
  NAND2_X1 U10562 ( .A1(n9144), .A2(n9143), .ZN(n9607) );
  NAND2_X1 U10563 ( .A1(n9608), .A2(n9607), .ZN(n9606) );
  NAND2_X1 U10564 ( .A1(n9613), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U10565 ( .A1(n9606), .A2(n9145), .ZN(n9146) );
  XNOR2_X1 U10566 ( .A(n9146), .B(n6006), .ZN(n9153) );
  OAI22_X1 U10567 ( .A1(n9149), .A2(n9148), .B1(n9147), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U10568 ( .A1(n9613), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9150) );
  OAI21_X1 U10569 ( .B1(n9613), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9150), .ZN(
        n9610) );
  OR2_X1 U10570 ( .A1(n9611), .A2(n9610), .ZN(n9614) );
  NAND2_X1 U10571 ( .A1(n9614), .A2(n9150), .ZN(n9151) );
  XNOR2_X1 U10572 ( .A(n9151), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9155) );
  INV_X1 U10573 ( .A(n9155), .ZN(n9152) );
  AOI22_X1 U10574 ( .A1(n9153), .A2(n9605), .B1(n9597), .B2(n9152), .ZN(n9158)
         );
  NOR2_X1 U10575 ( .A1(n9153), .A2(n9581), .ZN(n9154) );
  AOI211_X1 U10576 ( .C1(n9597), .C2(n9155), .A(n9612), .B(n9154), .ZN(n9157)
         );
  MUX2_X1 U10577 ( .A(n9158), .B(n9157), .S(n9156), .Z(n9160) );
  NAND2_X1 U10578 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9159) );
  OAI211_X1 U10579 ( .C1(n9161), .C2(n9620), .A(n9160), .B(n9159), .ZN(
        P1_U3262) );
  NOR2_X1 U10580 ( .A1(n9420), .A2(n9162), .ZN(n9163) );
  OAI21_X1 U10581 ( .B1(n9624), .B2(n10193), .A(n9165), .ZN(n9166) );
  AOI21_X1 U10582 ( .B1(n9167), .B2(n9627), .A(n9166), .ZN(n9168) );
  OAI21_X1 U10583 ( .B1(n9353), .B2(n9629), .A(n9168), .ZN(P1_U3264) );
  NAND2_X1 U10584 ( .A1(n9169), .A2(n9318), .ZN(n9173) );
  INV_X1 U10585 ( .A(n9170), .ZN(n9171) );
  AOI22_X1 U10586 ( .A1(n9321), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9171), .B2(
        n9319), .ZN(n9172) );
  OAI211_X1 U10587 ( .C1(n9174), .C2(n9324), .A(n9173), .B(n9172), .ZN(n9175)
         );
  AOI21_X1 U10588 ( .B1(n9176), .B2(n9624), .A(n9175), .ZN(n9177) );
  OAI21_X1 U10589 ( .B1(n9178), .B2(n9328), .A(n9177), .ZN(P1_U3356) );
  XNOR2_X1 U10590 ( .A(n9179), .B(n9182), .ZN(n9358) );
  INV_X1 U10591 ( .A(n9358), .ZN(n9195) );
  OAI21_X1 U10592 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9183) );
  NAND2_X1 U10593 ( .A1(n9183), .A2(n9329), .ZN(n9185) );
  NAND2_X1 U10594 ( .A1(n9185), .A2(n9184), .ZN(n9356) );
  AOI211_X1 U10595 ( .C1(n9188), .C2(n9200), .A(n9317), .B(n9187), .ZN(n9357)
         );
  NAND2_X1 U10596 ( .A1(n9357), .A2(n9318), .ZN(n9192) );
  INV_X1 U10597 ( .A(n9189), .ZN(n9190) );
  AOI22_X1 U10598 ( .A1(n9321), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9190), .B2(
        n9319), .ZN(n9191) );
  OAI211_X1 U10599 ( .C1(n6139), .C2(n9324), .A(n9192), .B(n9191), .ZN(n9193)
         );
  AOI21_X1 U10600 ( .B1(n9356), .B2(n9624), .A(n9193), .ZN(n9194) );
  OAI21_X1 U10601 ( .B1(n9195), .B2(n9328), .A(n9194), .ZN(P1_U3266) );
  NAND2_X1 U10602 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  XOR2_X1 U10603 ( .A(n9199), .B(n9198), .Z(n9365) );
  AOI211_X1 U10604 ( .C1(n9362), .C2(n9224), .A(n9317), .B(n9186), .ZN(n9361)
         );
  INV_X1 U10605 ( .A(n9201), .ZN(n9202) );
  AOI22_X1 U10606 ( .A1(n9321), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9202), .B2(
        n9319), .ZN(n9203) );
  OAI21_X1 U10607 ( .B1(n9204), .B2(n9324), .A(n9203), .ZN(n9212) );
  AND2_X1 U10608 ( .A1(n9206), .A2(n9205), .ZN(n9208) );
  OAI21_X1 U10609 ( .B1(n9208), .B2(n6129), .A(n9207), .ZN(n9210) );
  AOI21_X1 U10610 ( .B1(n9210), .B2(n9329), .A(n9209), .ZN(n9364) );
  NOR2_X1 U10611 ( .A1(n9364), .A2(n9321), .ZN(n9211) );
  AOI211_X1 U10612 ( .C1(n9361), .C2(n9318), .A(n9212), .B(n9211), .ZN(n9213)
         );
  OAI21_X1 U10613 ( .B1(n9365), .B2(n9328), .A(n9213), .ZN(P1_U3267) );
  INV_X1 U10614 ( .A(n9221), .ZN(n9214) );
  XNOR2_X1 U10615 ( .A(n9215), .B(n9214), .ZN(n9217) );
  AOI21_X1 U10616 ( .B1(n9217), .B2(n9329), .A(n9216), .ZN(n9367) );
  NAND2_X1 U10617 ( .A1(n9219), .A2(n9218), .ZN(n9220) );
  XOR2_X1 U10618 ( .A(n9221), .B(n9220), .Z(n9369) );
  OR2_X1 U10619 ( .A1(n9369), .A2(n9328), .ZN(n9229) );
  OAI22_X1 U10620 ( .A1(n9223), .A2(n9621), .B1(n9222), .B2(n9624), .ZN(n9226)
         );
  OAI211_X1 U10621 ( .C1(n9428), .C2(n9238), .A(n9342), .B(n9224), .ZN(n9366)
         );
  NOR2_X1 U10622 ( .A1(n9366), .A2(n9629), .ZN(n9225) );
  AOI211_X1 U10623 ( .C1(n9627), .C2(n9227), .A(n9226), .B(n9225), .ZN(n9228)
         );
  OAI211_X1 U10624 ( .C1(n9321), .C2(n9367), .A(n9229), .B(n9228), .ZN(
        P1_U3268) );
  XNOR2_X1 U10625 ( .A(n9230), .B(n9231), .ZN(n9434) );
  NAND2_X1 U10626 ( .A1(n9232), .A2(n9329), .ZN(n9237) );
  AOI21_X1 U10627 ( .B1(n9246), .B2(n9234), .A(n9233), .ZN(n9236) );
  OAI21_X1 U10628 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9373) );
  AOI211_X1 U10629 ( .C1(n9432), .C2(n9253), .A(n9317), .B(n9238), .ZN(n9372)
         );
  NAND2_X1 U10630 ( .A1(n9372), .A2(n9318), .ZN(n9241) );
  AOI22_X1 U10631 ( .A1(n9239), .A2(n9319), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9321), .ZN(n9240) );
  OAI211_X1 U10632 ( .C1(n9242), .C2(n9324), .A(n9241), .B(n9240), .ZN(n9243)
         );
  AOI21_X1 U10633 ( .B1(n9373), .B2(n9624), .A(n9243), .ZN(n9244) );
  OAI21_X1 U10634 ( .B1(n9434), .B2(n9328), .A(n9244), .ZN(P1_U3269) );
  XNOR2_X1 U10635 ( .A(n9245), .B(n9248), .ZN(n9438) );
  OAI21_X1 U10636 ( .B1(n9248), .B2(n9247), .A(n9246), .ZN(n9249) );
  NAND2_X1 U10637 ( .A1(n9249), .A2(n9329), .ZN(n9252) );
  INV_X1 U10638 ( .A(n9250), .ZN(n9251) );
  NAND2_X1 U10639 ( .A1(n9252), .A2(n9251), .ZN(n9377) );
  INV_X1 U10640 ( .A(n9253), .ZN(n9254) );
  AOI211_X1 U10641 ( .C1(n9379), .C2(n4683), .A(n9317), .B(n9254), .ZN(n9378)
         );
  NAND2_X1 U10642 ( .A1(n9378), .A2(n9318), .ZN(n9258) );
  INV_X1 U10643 ( .A(n9255), .ZN(n9256) );
  AOI22_X1 U10644 ( .A1(n9256), .A2(n9319), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9321), .ZN(n9257) );
  OAI211_X1 U10645 ( .C1(n9259), .C2(n9324), .A(n9258), .B(n9257), .ZN(n9260)
         );
  AOI21_X1 U10646 ( .B1(n9377), .B2(n9624), .A(n9260), .ZN(n9261) );
  OAI21_X1 U10647 ( .B1(n9438), .B2(n9328), .A(n9261), .ZN(P1_U3270) );
  XNOR2_X1 U10648 ( .A(n9263), .B(n9262), .ZN(n9384) );
  INV_X1 U10649 ( .A(n9384), .ZN(n9276) );
  XNOR2_X1 U10650 ( .A(n9265), .B(n9264), .ZN(n9267) );
  OAI21_X1 U10651 ( .B1(n9267), .B2(n9314), .A(n9266), .ZN(n9382) );
  AOI211_X1 U10652 ( .C1(n9269), .C2(n9284), .A(n9317), .B(n9268), .ZN(n9383)
         );
  NAND2_X1 U10653 ( .A1(n9383), .A2(n9318), .ZN(n9273) );
  INV_X1 U10654 ( .A(n9270), .ZN(n9271) );
  AOI22_X1 U10655 ( .A1(n9271), .A2(n9319), .B1(n9321), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9272) );
  OAI211_X1 U10656 ( .C1(n9443), .C2(n9324), .A(n9273), .B(n9272), .ZN(n9274)
         );
  AOI21_X1 U10657 ( .B1(n9382), .B2(n9624), .A(n9274), .ZN(n9275) );
  OAI21_X1 U10658 ( .B1(n9276), .B2(n9328), .A(n9275), .ZN(P1_U3271) );
  XNOR2_X1 U10659 ( .A(n9278), .B(n9277), .ZN(n9447) );
  XNOR2_X1 U10660 ( .A(n9280), .B(n9279), .ZN(n9282) );
  OAI21_X1 U10661 ( .B1(n9282), .B2(n9314), .A(n9281), .ZN(n9388) );
  INV_X1 U10662 ( .A(n9283), .ZN(n9300) );
  INV_X1 U10663 ( .A(n9284), .ZN(n9285) );
  AOI211_X1 U10664 ( .C1(n9390), .C2(n9300), .A(n9317), .B(n9285), .ZN(n9389)
         );
  NAND2_X1 U10665 ( .A1(n9389), .A2(n9318), .ZN(n9289) );
  INV_X1 U10666 ( .A(n9286), .ZN(n9287) );
  AOI22_X1 U10667 ( .A1(n9321), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9287), .B2(
        n9319), .ZN(n9288) );
  OAI211_X1 U10668 ( .C1(n9290), .C2(n9324), .A(n9289), .B(n9288), .ZN(n9291)
         );
  AOI21_X1 U10669 ( .B1(n9388), .B2(n9624), .A(n9291), .ZN(n9292) );
  OAI21_X1 U10670 ( .B1(n9447), .B2(n9328), .A(n9292), .ZN(P1_U3272) );
  XNOR2_X1 U10671 ( .A(n9293), .B(n9294), .ZN(n9452) );
  AOI21_X1 U10672 ( .B1(n9295), .B2(n9294), .A(n9314), .ZN(n9299) );
  INV_X1 U10673 ( .A(n9296), .ZN(n9297) );
  AOI21_X1 U10674 ( .B1(n9299), .B2(n9298), .A(n9297), .ZN(n9394) );
  INV_X1 U10675 ( .A(n9394), .ZN(n9306) );
  OAI211_X1 U10676 ( .C1(n9301), .C2(n9316), .A(n9300), .B(n9342), .ZN(n9393)
         );
  AOI22_X1 U10677 ( .A1(n9321), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9302), .B2(
        n9319), .ZN(n9304) );
  NAND2_X1 U10678 ( .A1(n9450), .A2(n9627), .ZN(n9303) );
  OAI211_X1 U10679 ( .C1(n9393), .C2(n9629), .A(n9304), .B(n9303), .ZN(n9305)
         );
  AOI21_X1 U10680 ( .B1(n9306), .B2(n9624), .A(n9305), .ZN(n9307) );
  OAI21_X1 U10681 ( .B1(n9452), .B2(n9328), .A(n9307), .ZN(P1_U3273) );
  XNOR2_X1 U10682 ( .A(n9309), .B(n9308), .ZN(n9456) );
  NAND2_X1 U10683 ( .A1(n9330), .A2(n9310), .ZN(n9312) );
  XNOR2_X1 U10684 ( .A(n9312), .B(n9311), .ZN(n9315) );
  OAI21_X1 U10685 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9397) );
  AOI211_X1 U10686 ( .C1(n9399), .C2(n9343), .A(n9317), .B(n9316), .ZN(n9398)
         );
  NAND2_X1 U10687 ( .A1(n9398), .A2(n9318), .ZN(n9323) );
  AOI22_X1 U10688 ( .A1(n9321), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9320), .B2(
        n9319), .ZN(n9322) );
  OAI211_X1 U10689 ( .C1(n9325), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9326)
         );
  AOI21_X1 U10690 ( .B1(n9397), .B2(n9624), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10691 ( .B1(n9456), .B2(n9328), .A(n9327), .ZN(P1_U3274) );
  OAI211_X1 U10692 ( .C1(n9336), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9334)
         );
  INV_X1 U10693 ( .A(n9332), .ZN(n9333) );
  INV_X1 U10694 ( .A(n9335), .ZN(n9337) );
  XOR2_X1 U10695 ( .A(n9337), .B(n9336), .Z(n9463) );
  INV_X1 U10696 ( .A(n9463), .ZN(n9339) );
  NAND2_X1 U10697 ( .A1(n9339), .A2(n9338), .ZN(n9348) );
  OAI22_X1 U10698 ( .A1(n9624), .A2(n9341), .B1(n9340), .B2(n9621), .ZN(n9346)
         );
  OAI211_X1 U10699 ( .C1(n4499), .C2(n9344), .A(n9343), .B(n9342), .ZN(n9402)
         );
  NOR2_X1 U10700 ( .A1(n9402), .A2(n9629), .ZN(n9345) );
  AOI211_X1 U10701 ( .C1(n9627), .C2(n9459), .A(n9346), .B(n9345), .ZN(n9347)
         );
  OAI211_X1 U10702 ( .C1(n9321), .C2(n9403), .A(n9348), .B(n9347), .ZN(
        P1_U3275) );
  INV_X1 U10703 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9350) );
  MUX2_X1 U10704 ( .A(n9350), .B(n9349), .S(n9678), .Z(n9351) );
  OAI21_X1 U10705 ( .B1(n4685), .B2(n9387), .A(n9351), .ZN(P1_U3553) );
  NAND2_X1 U10706 ( .A1(n9353), .A2(n9352), .ZN(n9417) );
  MUX2_X1 U10707 ( .A(n9417), .B(P1_REG1_REG_30__SCAN_IN), .S(n9676), .Z(n9354) );
  INV_X1 U10708 ( .A(n9354), .ZN(n9355) );
  OAI21_X1 U10709 ( .B1(n9420), .B2(n9387), .A(n9355), .ZN(P1_U3552) );
  MUX2_X1 U10710 ( .A(n9359), .B(n9421), .S(n9678), .Z(n9360) );
  AOI21_X1 U10711 ( .B1(n9411), .B2(n9362), .A(n9361), .ZN(n9363) );
  OAI211_X1 U10712 ( .C1(n9365), .C2(n9368), .A(n9364), .B(n9363), .ZN(n9424)
         );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9424), .S(n9678), .Z(
        P1_U3548) );
  OAI211_X1 U10714 ( .C1(n9369), .C2(n9368), .A(n9367), .B(n9366), .ZN(n9425)
         );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9425), .S(n9678), .Z(n9370) );
  INV_X1 U10716 ( .A(n9370), .ZN(n9371) );
  OAI21_X1 U10717 ( .B1(n9428), .B2(n9387), .A(n9371), .ZN(P1_U3547) );
  NOR2_X1 U10718 ( .A1(n9373), .A2(n9372), .ZN(n9429) );
  MUX2_X1 U10719 ( .A(n9374), .B(n9429), .S(n9678), .Z(n9376) );
  NAND2_X1 U10720 ( .A1(n9432), .A2(n9405), .ZN(n9375) );
  OAI211_X1 U10721 ( .C1(n9434), .C2(n9407), .A(n9376), .B(n9375), .ZN(
        P1_U3546) );
  AOI211_X1 U10722 ( .C1(n9411), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9435)
         );
  MUX2_X1 U10723 ( .A(n9380), .B(n9435), .S(n9678), .Z(n9381) );
  OAI21_X1 U10724 ( .B1(n9438), .B2(n9407), .A(n9381), .ZN(P1_U3545) );
  INV_X1 U10725 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9385) );
  AOI211_X1 U10726 ( .C1(n9384), .C2(n9673), .A(n9383), .B(n9382), .ZN(n9439)
         );
  MUX2_X1 U10727 ( .A(n9385), .B(n9439), .S(n9678), .Z(n9386) );
  OAI21_X1 U10728 ( .B1(n9443), .B2(n9387), .A(n9386), .ZN(P1_U3544) );
  INV_X1 U10729 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9391) );
  AOI211_X1 U10730 ( .C1(n9411), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9444)
         );
  MUX2_X1 U10731 ( .A(n9391), .B(n9444), .S(n9678), .Z(n9392) );
  OAI21_X1 U10732 ( .B1(n9447), .B2(n9407), .A(n9392), .ZN(P1_U3543) );
  NAND2_X1 U10733 ( .A1(n9394), .A2(n9393), .ZN(n9448) );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9448), .S(n9678), .Z(n9395) );
  AOI21_X1 U10735 ( .B1(n9405), .B2(n9450), .A(n9395), .ZN(n9396) );
  OAI21_X1 U10736 ( .B1(n9452), .B2(n9407), .A(n9396), .ZN(P1_U3542) );
  INV_X1 U10737 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9400) );
  AOI211_X1 U10738 ( .C1(n9411), .C2(n9399), .A(n9398), .B(n9397), .ZN(n9453)
         );
  MUX2_X1 U10739 ( .A(n9400), .B(n9453), .S(n9678), .Z(n9401) );
  OAI21_X1 U10740 ( .B1(n9456), .B2(n9407), .A(n9401), .ZN(P1_U3541) );
  NAND2_X1 U10741 ( .A1(n9403), .A2(n9402), .ZN(n9457) );
  MUX2_X1 U10742 ( .A(n9457), .B(P1_REG1_REG_18__SCAN_IN), .S(n9676), .Z(n9404) );
  AOI21_X1 U10743 ( .B1(n9405), .B2(n9459), .A(n9404), .ZN(n9406) );
  OAI21_X1 U10744 ( .B1(n9463), .B2(n9407), .A(n9406), .ZN(P1_U3540) );
  INV_X1 U10745 ( .A(n9408), .ZN(n9415) );
  AOI21_X1 U10746 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9412) );
  OAI211_X1 U10747 ( .C1(n9415), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9465)
         );
  MUX2_X1 U10748 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9465), .S(n9678), .Z(
        P1_U3536) );
  MUX2_X1 U10749 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9416), .S(n9678), .Z(
        P1_U3522) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9417), .S(n9464), .Z(n9418) );
  INV_X1 U10751 ( .A(n9418), .ZN(n9419) );
  OAI21_X1 U10752 ( .B1(n9420), .B2(n9442), .A(n9419), .ZN(P1_U3520) );
  MUX2_X1 U10753 ( .A(n9422), .B(n9421), .S(n9464), .Z(n9423) );
  OAI21_X1 U10754 ( .B1(n6139), .B2(n9442), .A(n9423), .ZN(P1_U3517) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9424), .S(n9464), .Z(
        P1_U3516) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9425), .S(n9464), .Z(n9426) );
  INV_X1 U10757 ( .A(n9426), .ZN(n9427) );
  OAI21_X1 U10758 ( .B1(n9428), .B2(n9442), .A(n9427), .ZN(P1_U3515) );
  INV_X1 U10759 ( .A(n9429), .ZN(n9430) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9430), .S(n9464), .Z(n9431) );
  AOI21_X1 U10761 ( .B1(n9460), .B2(n9432), .A(n9431), .ZN(n9433) );
  OAI21_X1 U10762 ( .B1(n9434), .B2(n9462), .A(n9433), .ZN(P1_U3514) );
  INV_X1 U10763 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9436) );
  MUX2_X1 U10764 ( .A(n9436), .B(n9435), .S(n9464), .Z(n9437) );
  OAI21_X1 U10765 ( .B1(n9438), .B2(n9462), .A(n9437), .ZN(P1_U3513) );
  INV_X1 U10766 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9440) );
  MUX2_X1 U10767 ( .A(n9440), .B(n9439), .S(n9464), .Z(n9441) );
  OAI21_X1 U10768 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(P1_U3512) );
  INV_X1 U10769 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U10770 ( .A(n9445), .B(n9444), .S(n9464), .Z(n9446) );
  OAI21_X1 U10771 ( .B1(n9447), .B2(n9462), .A(n9446), .ZN(P1_U3511) );
  MUX2_X1 U10772 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9448), .S(n9464), .Z(n9449) );
  AOI21_X1 U10773 ( .B1(n9460), .B2(n9450), .A(n9449), .ZN(n9451) );
  OAI21_X1 U10774 ( .B1(n9452), .B2(n9462), .A(n9451), .ZN(P1_U3510) );
  INV_X1 U10775 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9454) );
  MUX2_X1 U10776 ( .A(n9454), .B(n9453), .S(n9464), .Z(n9455) );
  OAI21_X1 U10777 ( .B1(n9456), .B2(n9462), .A(n9455), .ZN(P1_U3509) );
  MUX2_X1 U10778 ( .A(n9457), .B(P1_REG0_REG_18__SCAN_IN), .S(n9674), .Z(n9458) );
  AOI21_X1 U10779 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9461) );
  OAI21_X1 U10780 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(P1_U3507) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9465), .S(n9464), .Z(
        P1_U3495) );
  MUX2_X1 U10782 ( .A(P1_D_REG_1__SCAN_IN), .B(n9466), .S(n9667), .Z(P1_U3440)
         );
  INV_X1 U10783 ( .A(n9467), .ZN(n9468) );
  NOR4_X1 U10784 ( .A1(n9468), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5745), .A4(
        P1_U3086), .ZN(n9469) );
  AOI21_X1 U10785 ( .B1(n10045), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9469), 
        .ZN(n9470) );
  OAI21_X1 U10786 ( .B1(n9471), .B2(n9476), .A(n9470), .ZN(P1_U3324) );
  OAI222_X1 U10787 ( .A1(n9478), .A2(n10213), .B1(n9476), .B2(n9473), .C1(
        P1_U3086), .C2(n9472), .ZN(P1_U3325) );
  OAI222_X1 U10788 ( .A1(n9478), .A2(n9477), .B1(n9476), .B2(n9475), .C1(n9474), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U10789 ( .A(n9479), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10790 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9491) );
  AOI211_X1 U10791 ( .C1(n9482), .C2(n9481), .A(n9480), .B(n9609), .ZN(n9487)
         );
  AOI211_X1 U10792 ( .C1(n9485), .C2(n9484), .A(n9483), .B(n9581), .ZN(n9486)
         );
  AOI211_X1 U10793 ( .C1(n9612), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9490)
         );
  NAND2_X1 U10794 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9489) );
  OAI211_X1 U10795 ( .C1(n9620), .C2(n9491), .A(n9490), .B(n9489), .ZN(
        P1_U3253) );
  INV_X1 U10796 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9505) );
  OAI21_X1 U10797 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9501) );
  OAI211_X1 U10798 ( .C1(n9497), .C2(n9496), .A(n9597), .B(n9495), .ZN(n9500)
         );
  NAND2_X1 U10799 ( .A1(n9612), .A2(n9498), .ZN(n9499) );
  OAI211_X1 U10800 ( .C1(n9501), .C2(n9581), .A(n9500), .B(n9499), .ZN(n9502)
         );
  INV_X1 U10801 ( .A(n9502), .ZN(n9504) );
  OAI211_X1 U10802 ( .C1(n9620), .C2(n9505), .A(n9504), .B(n9503), .ZN(
        P1_U3250) );
  OAI21_X1 U10803 ( .B1(n9507), .B2(n9506), .A(n9597), .ZN(n9514) );
  AOI211_X1 U10804 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9581), .ZN(n9511)
         );
  AOI21_X1 U10805 ( .B1(n9612), .B2(n9512), .A(n9511), .ZN(n9513) );
  OAI21_X1 U10806 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(n9517) );
  AOI211_X1 U10807 ( .C1(n9518), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9517), .B(
        n9516), .ZN(n9519) );
  INV_X1 U10808 ( .A(n9519), .ZN(P1_U3251) );
  NOR2_X1 U10809 ( .A1(n9520), .A2(n9932), .ZN(n9521) );
  AOI211_X1 U10810 ( .C1(n9943), .C2(n9523), .A(n9522), .B(n9521), .ZN(n9525)
         );
  AOI22_X1 U10811 ( .A1(n9963), .A2(n9525), .B1(n5305), .B2(n5726), .ZN(
        P2_U3472) );
  INV_X1 U10812 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U10813 ( .A1(n9946), .A2(n9525), .B1(n9524), .B2(n9944), .ZN(
        P2_U3429) );
  XNOR2_X1 U10814 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10815 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U10816 ( .A1(n9527), .A2(n9526), .ZN(n9530) );
  INV_X1 U10817 ( .A(n9528), .ZN(n9529) );
  NAND2_X1 U10818 ( .A1(n9530), .A2(n9529), .ZN(n9538) );
  NAND2_X1 U10819 ( .A1(n9612), .A2(n9531), .ZN(n9537) );
  AOI21_X1 U10820 ( .B1(n9534), .B2(n9533), .A(n9532), .ZN(n9535) );
  NAND2_X1 U10821 ( .A1(n9597), .A2(n9535), .ZN(n9536) );
  OAI211_X1 U10822 ( .C1(n9581), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9539)
         );
  INV_X1 U10823 ( .A(n9539), .ZN(n9541) );
  OAI211_X1 U10824 ( .C1(n9620), .C2(n9542), .A(n9541), .B(n9540), .ZN(
        P1_U3254) );
  INV_X1 U10825 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U10826 ( .A1(n9544), .A2(n9543), .ZN(n9547) );
  INV_X1 U10827 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U10828 ( .A1(n9547), .A2(n9546), .ZN(n9556) );
  INV_X1 U10829 ( .A(n9548), .ZN(n9549) );
  NAND2_X1 U10830 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  NAND3_X1 U10831 ( .A1(n9597), .A2(n9552), .A3(n9551), .ZN(n9555) );
  NAND2_X1 U10832 ( .A1(n9612), .A2(n9553), .ZN(n9554) );
  OAI211_X1 U10833 ( .C1(n9581), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9557)
         );
  INV_X1 U10834 ( .A(n9557), .ZN(n9559) );
  OAI211_X1 U10835 ( .C1(n9620), .C2(n9560), .A(n9559), .B(n9558), .ZN(
        P1_U3256) );
  INV_X1 U10836 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U10837 ( .A1(n9562), .A2(n9561), .ZN(n9565) );
  INV_X1 U10838 ( .A(n9563), .ZN(n9564) );
  NAND2_X1 U10839 ( .A1(n9565), .A2(n9564), .ZN(n9573) );
  NAND2_X1 U10840 ( .A1(n9612), .A2(n9566), .ZN(n9572) );
  AOI21_X1 U10841 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9570) );
  NAND2_X1 U10842 ( .A1(n9597), .A2(n9570), .ZN(n9571) );
  OAI211_X1 U10843 ( .C1(n9581), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9574)
         );
  INV_X1 U10844 ( .A(n9574), .ZN(n9576) );
  NAND2_X1 U10845 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9575) );
  OAI211_X1 U10846 ( .C1(n9620), .C2(n9577), .A(n9576), .B(n9575), .ZN(
        P1_U3257) );
  INV_X1 U10847 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9590) );
  AOI211_X1 U10848 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9609), .ZN(n9586)
         );
  AOI211_X1 U10849 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9585)
         );
  AOI211_X1 U10850 ( .C1(n9612), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9589)
         );
  NAND2_X1 U10851 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9588) );
  OAI211_X1 U10852 ( .C1(n9620), .C2(n9590), .A(n9589), .B(n9588), .ZN(
        P1_U3258) );
  NAND2_X1 U10853 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  NAND3_X1 U10854 ( .A1(n9594), .A2(n9605), .A3(n9593), .ZN(n9602) );
  XNOR2_X1 U10855 ( .A(n9596), .B(n9595), .ZN(n9598) );
  NAND2_X1 U10856 ( .A1(n9598), .A2(n9597), .ZN(n9601) );
  NAND2_X1 U10857 ( .A1(n9612), .A2(n9599), .ZN(n9600) );
  AND3_X1 U10858 ( .A1(n9602), .A2(n9601), .A3(n9600), .ZN(n9604) );
  NAND2_X1 U10859 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9603) );
  OAI211_X1 U10860 ( .C1(n10068), .C2(n9620), .A(n9604), .B(n9603), .ZN(
        P1_U3259) );
  OAI211_X1 U10861 ( .C1(n9608), .C2(n9607), .A(n9606), .B(n9605), .ZN(n9617)
         );
  AOI21_X1 U10862 ( .B1(n9611), .B2(n9610), .A(n9609), .ZN(n9615) );
  AOI22_X1 U10863 ( .A1(n9615), .A2(n9614), .B1(n9613), .B2(n9612), .ZN(n9616)
         );
  AND2_X1 U10864 ( .A1(n9617), .A2(n9616), .ZN(n9619) );
  NAND2_X1 U10865 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9618) );
  OAI211_X1 U10866 ( .C1(n9620), .C2(n9969), .A(n9619), .B(n9618), .ZN(
        P1_U3261) );
  OAI22_X1 U10867 ( .A1(n9624), .A2(n9623), .B1(n9622), .B2(n9621), .ZN(n9625)
         );
  AOI21_X1 U10868 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9628) );
  OAI21_X1 U10869 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9631) );
  AOI21_X1 U10870 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9634) );
  OAI21_X1 U10871 ( .B1(n9321), .B2(n9635), .A(n9634), .ZN(P1_U3286) );
  INV_X1 U10872 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9638) );
  NOR2_X1 U10873 ( .A1(n9655), .A2(n9638), .ZN(P1_U3294) );
  INV_X1 U10874 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9639) );
  NOR2_X1 U10875 ( .A1(n9655), .A2(n9639), .ZN(P1_U3295) );
  INV_X1 U10876 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9640) );
  NOR2_X1 U10877 ( .A1(n9655), .A2(n9640), .ZN(P1_U3296) );
  INV_X1 U10878 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U10879 ( .A1(n9655), .A2(n9641), .ZN(P1_U3297) );
  INV_X1 U10880 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9642) );
  NOR2_X1 U10881 ( .A1(n9655), .A2(n9642), .ZN(P1_U3298) );
  INV_X1 U10882 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9643) );
  NOR2_X1 U10883 ( .A1(n9655), .A2(n9643), .ZN(P1_U3299) );
  INV_X1 U10884 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9644) );
  NOR2_X1 U10885 ( .A1(n9655), .A2(n9644), .ZN(P1_U3300) );
  INV_X1 U10886 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9645) );
  NOR2_X1 U10887 ( .A1(n9655), .A2(n9645), .ZN(P1_U3301) );
  INV_X1 U10888 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9646) );
  NOR2_X1 U10889 ( .A1(n9655), .A2(n9646), .ZN(P1_U3302) );
  INV_X1 U10890 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9647) );
  NOR2_X1 U10891 ( .A1(n9655), .A2(n9647), .ZN(P1_U3303) );
  INV_X1 U10892 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9648) );
  NOR2_X1 U10893 ( .A1(n9655), .A2(n9648), .ZN(P1_U3304) );
  INV_X1 U10894 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U10895 ( .A1(n9655), .A2(n9649), .ZN(P1_U3305) );
  INV_X1 U10896 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9650) );
  NOR2_X1 U10897 ( .A1(n9655), .A2(n9650), .ZN(P1_U3306) );
  INV_X1 U10898 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9651) );
  NOR2_X1 U10899 ( .A1(n9655), .A2(n9651), .ZN(P1_U3307) );
  INV_X1 U10900 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9652) );
  NOR2_X1 U10901 ( .A1(n9655), .A2(n9652), .ZN(P1_U3308) );
  INV_X1 U10902 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U10903 ( .A1(n9655), .A2(n9653), .ZN(P1_U3309) );
  INV_X1 U10904 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U10905 ( .A1(n9655), .A2(n10191), .ZN(P1_U3310) );
  INV_X1 U10906 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U10907 ( .A1(n9655), .A2(n10079), .ZN(P1_U3311) );
  INV_X1 U10908 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9654) );
  NOR2_X1 U10909 ( .A1(n9655), .A2(n9654), .ZN(P1_U3312) );
  INV_X1 U10910 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9656) );
  NOR2_X1 U10911 ( .A1(n9664), .A2(n9656), .ZN(P1_U3313) );
  INV_X1 U10912 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9657) );
  NOR2_X1 U10913 ( .A1(n9664), .A2(n9657), .ZN(P1_U3314) );
  INV_X1 U10914 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10154) );
  NOR2_X1 U10915 ( .A1(n9664), .A2(n10154), .ZN(P1_U3315) );
  INV_X1 U10916 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9658) );
  NOR2_X1 U10917 ( .A1(n9664), .A2(n9658), .ZN(P1_U3316) );
  INV_X1 U10918 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U10919 ( .A1(n9664), .A2(n10138), .ZN(P1_U3317) );
  INV_X1 U10920 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9659) );
  NOR2_X1 U10921 ( .A1(n9664), .A2(n9659), .ZN(P1_U3318) );
  INV_X1 U10922 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9660) );
  NOR2_X1 U10923 ( .A1(n9664), .A2(n9660), .ZN(P1_U3319) );
  INV_X1 U10924 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9661) );
  NOR2_X1 U10925 ( .A1(n9664), .A2(n9661), .ZN(P1_U3320) );
  INV_X1 U10926 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9662) );
  NOR2_X1 U10927 ( .A1(n9664), .A2(n9662), .ZN(P1_U3321) );
  INV_X1 U10928 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9663) );
  NOR2_X1 U10929 ( .A1(n9664), .A2(n9663), .ZN(P1_U3322) );
  INV_X1 U10930 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10155) );
  NOR2_X1 U10931 ( .A1(n9664), .A2(n10155), .ZN(P1_U3323) );
  INV_X1 U10932 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9666) );
  OAI21_X1 U10933 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(P1_U3439) );
  OAI21_X1 U10934 ( .B1(n5894), .B2(n9669), .A(n9668), .ZN(n9671) );
  AOI211_X1 U10935 ( .C1(n9673), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9677)
         );
  INV_X1 U10936 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U10937 ( .A1(n9464), .A2(n9677), .B1(n9675), .B2(n9674), .ZN(
        P1_U3480) );
  AOI22_X1 U10938 ( .A1(n9678), .A2(n9677), .B1(n5886), .B2(n9676), .ZN(
        P1_U3531) );
  INV_X1 U10939 ( .A(n9679), .ZN(n9680) );
  AOI21_X1 U10940 ( .B1(n6767), .B2(n9681), .A(n9680), .ZN(n9686) );
  XNOR2_X1 U10941 ( .A(n9682), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9684) );
  AOI21_X1 U10942 ( .B1(n9852), .B2(n9684), .A(n9683), .ZN(n9685) );
  OAI21_X1 U10943 ( .B1(n9686), .B2(n9856), .A(n9685), .ZN(n9687) );
  AOI21_X1 U10944 ( .B1(n9688), .B2(n9844), .A(n9687), .ZN(n9696) );
  AOI21_X1 U10945 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9693) );
  NOR2_X1 U10946 ( .A1(n9693), .A2(n9692), .ZN(n9694) );
  AOI21_X1 U10947 ( .B1(n9842), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9694), .ZN(
        n9695) );
  NAND2_X1 U10948 ( .A1(n9696), .A2(n9695), .ZN(P2_U3185) );
  INV_X1 U10949 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9712) );
  XNOR2_X1 U10950 ( .A(n9697), .B(n6686), .ZN(n9701) );
  OAI21_X1 U10951 ( .B1(n9699), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9698), .ZN(
        n9700) );
  AOI22_X1 U10952 ( .A1(n9718), .A2(n9701), .B1(n9852), .B2(n9700), .ZN(n9711)
         );
  OAI211_X1 U10953 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9851), .ZN(n9706)
         );
  OAI211_X1 U10954 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9709)
         );
  INV_X1 U10955 ( .A(n9709), .ZN(n9710) );
  OAI211_X1 U10956 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(
        P2_U3187) );
  AOI21_X1 U10957 ( .B1(n9844), .B2(n9715), .A(n9714), .ZN(n9722) );
  XNOR2_X1 U10958 ( .A(n9716), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U10959 ( .A1(n9717), .A2(n9852), .ZN(n9721) );
  NAND2_X1 U10960 ( .A1(n9719), .A2(n9718), .ZN(n9720) );
  AND3_X1 U10961 ( .A1(n9722), .A2(n9721), .A3(n9720), .ZN(n9727) );
  XNOR2_X1 U10962 ( .A(n9724), .B(n9723), .ZN(n9725) );
  AOI22_X1 U10963 ( .A1(n9725), .A2(n9851), .B1(n9842), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U10964 ( .A1(n9727), .A2(n9726), .ZN(P2_U3189) );
  AOI21_X1 U10965 ( .B1(n9844), .B2(n9729), .A(n9728), .ZN(n9745) );
  OAI21_X1 U10966 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  AOI22_X1 U10967 ( .A1(n9733), .A2(n9851), .B1(n9842), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n9744) );
  OAI21_X1 U10968 ( .B1(n9736), .B2(n9735), .A(n9734), .ZN(n9737) );
  NAND2_X1 U10969 ( .A1(n9737), .A2(n9852), .ZN(n9743) );
  AOI21_X1 U10970 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9741) );
  OR2_X1 U10971 ( .A1(n9741), .A2(n9856), .ZN(n9742) );
  NAND4_X1 U10972 ( .A1(n9745), .A2(n9744), .A3(n9743), .A4(n9742), .ZN(
        P2_U3190) );
  AOI22_X1 U10973 ( .A1(n9844), .A2(n9746), .B1(n9842), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n9760) );
  OAI21_X1 U10974 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n9748), .A(n9747), .ZN(
        n9753) );
  OAI21_X1 U10975 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9752) );
  AOI22_X1 U10976 ( .A1(n9753), .A2(n9852), .B1(n9851), .B2(n9752), .ZN(n9759)
         );
  AOI21_X1 U10977 ( .B1(n9755), .B2(n5227), .A(n9754), .ZN(n9756) );
  OR2_X1 U10978 ( .A1(n9856), .A2(n9756), .ZN(n9757) );
  NAND4_X1 U10979 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), .ZN(
        P2_U3191) );
  AOI22_X1 U10980 ( .A1(n9844), .A2(n9761), .B1(n9842), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n9775) );
  OAI21_X1 U10981 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9763), .A(n9762), .ZN(
        n9768) );
  OAI21_X1 U10982 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9767) );
  AOI22_X1 U10983 ( .A1(n9768), .A2(n9852), .B1(n9851), .B2(n9767), .ZN(n9774)
         );
  AOI21_X1 U10984 ( .B1(n9770), .B2(n7043), .A(n9769), .ZN(n9771) );
  OR2_X1 U10985 ( .A1(n9771), .A2(n9856), .ZN(n9772) );
  NAND4_X1 U10986 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(
        P2_U3193) );
  AOI22_X1 U10987 ( .A1(n9844), .A2(n9776), .B1(n9842), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9792) );
  OAI21_X1 U10988 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9784) );
  OAI21_X1 U10989 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9783) );
  AOI22_X1 U10990 ( .A1(n9784), .A2(n9852), .B1(n9851), .B2(n9783), .ZN(n9791)
         );
  INV_X1 U10991 ( .A(n9785), .ZN(n9790) );
  AOI21_X1 U10992 ( .B1(n4503), .B2(n9787), .A(n9786), .ZN(n9788) );
  OR2_X1 U10993 ( .A1(n9788), .A2(n9856), .ZN(n9789) );
  NAND4_X1 U10994 ( .A1(n9792), .A2(n9791), .A3(n9790), .A4(n9789), .ZN(
        P2_U3194) );
  AOI22_X1 U10995 ( .A1(n9844), .A2(n9793), .B1(n9842), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9808) );
  OAI21_X1 U10996 ( .B1(n9796), .B2(n9795), .A(n9794), .ZN(n9801) );
  OAI21_X1 U10997 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n9800) );
  AOI22_X1 U10998 ( .A1(n9801), .A2(n9852), .B1(n9851), .B2(n9800), .ZN(n9807)
         );
  NAND2_X1 U10999 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9806) );
  AOI21_X1 U11000 ( .B1(n4504), .B2(n9803), .A(n9802), .ZN(n9804) );
  OR2_X1 U11001 ( .A1(n9804), .A2(n9856), .ZN(n9805) );
  NAND4_X1 U11002 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(
        P2_U3196) );
  AOI22_X1 U11003 ( .A1(n9844), .A2(n9809), .B1(n9842), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9824) );
  OAI21_X1 U11004 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9811), .A(n9810), .ZN(
        n9816) );
  OAI21_X1 U11005 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  AOI22_X1 U11006 ( .A1(n9816), .A2(n9852), .B1(n9851), .B2(n9815), .ZN(n9823)
         );
  INV_X1 U11007 ( .A(n9817), .ZN(n9822) );
  AOI21_X1 U11008 ( .B1(n9819), .B2(n8434), .A(n9818), .ZN(n9820) );
  OR2_X1 U11009 ( .A1(n9856), .A2(n9820), .ZN(n9821) );
  NAND4_X1 U11010 ( .A1(n9824), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(
        P2_U3197) );
  AOI22_X1 U11011 ( .A1(n9844), .A2(n9825), .B1(n9842), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n9841) );
  OAI21_X1 U11012 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9833) );
  OAI21_X1 U11013 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9832) );
  AOI22_X1 U11014 ( .A1(n9833), .A2(n9852), .B1(n9851), .B2(n9832), .ZN(n9840)
         );
  NAND2_X1 U11015 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9839) );
  AOI21_X1 U11016 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9837) );
  OR2_X1 U11017 ( .A1(n9837), .A2(n9856), .ZN(n9838) );
  NAND4_X1 U11018 ( .A1(n9841), .A2(n9840), .A3(n9839), .A4(n9838), .ZN(
        P2_U3198) );
  AOI22_X1 U11019 ( .A1(n9844), .A2(n9843), .B1(n9842), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9861) );
  OAI21_X1 U11020 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9846), .A(n9845), .ZN(
        n9853) );
  OAI21_X1 U11021 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9850) );
  AOI22_X1 U11022 ( .A1(n9853), .A2(n9852), .B1(n9851), .B2(n9850), .ZN(n9860)
         );
  AOI21_X1 U11023 ( .B1(n9855), .B2(n8414), .A(n9854), .ZN(n9857) );
  OR2_X1 U11024 ( .A1(n9857), .A2(n9856), .ZN(n9858) );
  NAND4_X1 U11025 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(
        P2_U3199) );
  XNOR2_X1 U11026 ( .A(n9862), .B(n7839), .ZN(n9887) );
  OAI22_X1 U11027 ( .A1(n9884), .A2(n9864), .B1(n6321), .B2(n9863), .ZN(n9874)
         );
  XNOR2_X1 U11028 ( .A(n9865), .B(n7839), .ZN(n9872) );
  NAND2_X1 U11029 ( .A1(n9887), .A2(n9927), .ZN(n9871) );
  AOI22_X1 U11030 ( .A1(n9869), .A2(n9868), .B1(n9867), .B2(n9866), .ZN(n9870)
         );
  OAI211_X1 U11031 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9885)
         );
  AOI211_X1 U11032 ( .C1(n9875), .C2(n9887), .A(n9874), .B(n9885), .ZN(n9877)
         );
  AOI22_X1 U11033 ( .A1(n6677), .A2(n9878), .B1(n9877), .B2(n9876), .ZN(
        P2_U3231) );
  NOR2_X1 U11034 ( .A1(n9879), .A2(n9919), .ZN(n9881) );
  AOI211_X1 U11035 ( .C1(n9926), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9948)
         );
  INV_X1 U11036 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U11037 ( .A1(n9946), .A2(n9948), .B1(n9883), .B2(n9944), .ZN(
        P2_U3393) );
  NOR2_X1 U11038 ( .A1(n9884), .A2(n9919), .ZN(n9886) );
  AOI211_X1 U11039 ( .C1(n9926), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9949)
         );
  INV_X1 U11040 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U11041 ( .A1(n9946), .A2(n9949), .B1(n9888), .B2(n9944), .ZN(
        P2_U3396) );
  AOI22_X1 U11042 ( .A1(n9890), .A2(n9938), .B1(n9943), .B2(n9889), .ZN(n9891)
         );
  AND2_X1 U11043 ( .A1(n9892), .A2(n9891), .ZN(n9951) );
  INV_X1 U11044 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U11045 ( .A1(n9946), .A2(n9951), .B1(n9893), .B2(n9944), .ZN(
        P2_U3399) );
  INV_X1 U11046 ( .A(n9894), .ZN(n9898) );
  OAI21_X1 U11047 ( .B1(n9896), .B2(n9919), .A(n9895), .ZN(n9897) );
  AOI21_X1 U11048 ( .B1(n9898), .B2(n9938), .A(n9897), .ZN(n9952) );
  AOI22_X1 U11049 ( .A1(n9946), .A2(n9952), .B1(n5107), .B2(n9944), .ZN(
        P2_U3402) );
  NOR2_X1 U11050 ( .A1(n9899), .A2(n9919), .ZN(n9901) );
  AOI211_X1 U11051 ( .C1(n9926), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9953)
         );
  INV_X1 U11052 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U11053 ( .A1(n9946), .A2(n9953), .B1(n9903), .B2(n9944), .ZN(
        P2_U3405) );
  INV_X1 U11054 ( .A(n9904), .ZN(n9908) );
  OAI21_X1 U11055 ( .B1(n9906), .B2(n9919), .A(n9905), .ZN(n9907) );
  AOI21_X1 U11056 ( .B1(n9908), .B2(n9938), .A(n9907), .ZN(n9954) );
  INV_X1 U11057 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U11058 ( .A1(n9946), .A2(n9954), .B1(n10064), .B2(n9944), .ZN(
        P2_U3408) );
  INV_X1 U11059 ( .A(n9909), .ZN(n9913) );
  OAI22_X1 U11060 ( .A1(n9911), .A2(n9932), .B1(n9910), .B2(n9919), .ZN(n9912)
         );
  NOR2_X1 U11061 ( .A1(n9913), .A2(n9912), .ZN(n9956) );
  AOI22_X1 U11062 ( .A1(n9946), .A2(n9956), .B1(n5165), .B2(n9944), .ZN(
        P2_U3411) );
  NOR2_X1 U11063 ( .A1(n9914), .A2(n9932), .ZN(n9916) );
  AOI211_X1 U11064 ( .C1(n9943), .C2(n9917), .A(n9916), .B(n9915), .ZN(n9957)
         );
  INV_X1 U11065 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U11066 ( .A1(n9946), .A2(n9957), .B1(n9918), .B2(n9944), .ZN(
        P2_U3414) );
  NOR2_X1 U11067 ( .A1(n9920), .A2(n9919), .ZN(n9922) );
  AOI211_X1 U11068 ( .C1(n9923), .C2(n9926), .A(n9922), .B(n9921), .ZN(n9958)
         );
  INV_X1 U11069 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U11070 ( .A1(n9946), .A2(n9958), .B1(n9924), .B2(n9944), .ZN(
        P2_U3417) );
  AOI22_X1 U11071 ( .A1(n9928), .A2(n9926), .B1(n9943), .B2(n9925), .ZN(n9930)
         );
  NAND2_X1 U11072 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  AOI22_X1 U11073 ( .A1(n9946), .A2(n9960), .B1(n5247), .B2(n9944), .ZN(
        P2_U3420) );
  NOR2_X1 U11074 ( .A1(n9933), .A2(n9932), .ZN(n9935) );
  AOI211_X1 U11075 ( .C1(n9943), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9961)
         );
  INV_X1 U11076 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U11077 ( .A1(n9946), .A2(n9961), .B1(n10225), .B2(n9944), .ZN(
        P2_U3423) );
  AND3_X1 U11078 ( .A1(n9939), .A2(n9938), .A3(n9937), .ZN(n9941) );
  AOI211_X1 U11079 ( .C1(n9943), .C2(n9942), .A(n9941), .B(n9940), .ZN(n9962)
         );
  INV_X1 U11080 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9945) );
  AOI22_X1 U11081 ( .A1(n9946), .A2(n9962), .B1(n9945), .B2(n9944), .ZN(
        P2_U3426) );
  INV_X1 U11082 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11083 ( .A1(n9963), .A2(n9948), .B1(n9947), .B2(n5726), .ZN(
        P2_U3460) );
  AOI22_X1 U11084 ( .A1(n9963), .A2(n9949), .B1(n6310), .B2(n5726), .ZN(
        P2_U3461) );
  INV_X1 U11085 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11086 ( .A1(n9963), .A2(n9951), .B1(n9950), .B2(n5726), .ZN(
        P2_U3462) );
  AOI22_X1 U11087 ( .A1(n9963), .A2(n9952), .B1(n6542), .B2(n5726), .ZN(
        P2_U3463) );
  AOI22_X1 U11088 ( .A1(n9963), .A2(n9953), .B1(n6685), .B2(n5726), .ZN(
        P2_U3464) );
  AOI22_X1 U11089 ( .A1(n9963), .A2(n9954), .B1(n6684), .B2(n5726), .ZN(
        P2_U3465) );
  INV_X1 U11090 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11091 ( .A1(n9963), .A2(n9956), .B1(n9955), .B2(n5726), .ZN(
        P2_U3466) );
  AOI22_X1 U11092 ( .A1(n9963), .A2(n9957), .B1(n5202), .B2(n5726), .ZN(
        P2_U3467) );
  AOI22_X1 U11093 ( .A1(n9963), .A2(n9958), .B1(n5228), .B2(n5726), .ZN(
        P2_U3468) );
  AOI22_X1 U11094 ( .A1(n9963), .A2(n9960), .B1(n9959), .B2(n5726), .ZN(
        P2_U3469) );
  AOI22_X1 U11095 ( .A1(n9963), .A2(n9961), .B1(n5273), .B2(n5726), .ZN(
        P2_U3470) );
  AOI22_X1 U11096 ( .A1(n9963), .A2(n9962), .B1(n5287), .B2(n5726), .ZN(
        P2_U3471) );
  OAI222_X1 U11097 ( .A1(n10246), .A2(n9967), .B1(n10246), .B2(n9966), .C1(
        n9965), .C2(n9964), .ZN(ADD_1068_U5) );
  XOR2_X1 U11098 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11099 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9972) );
  XNOR2_X1 U11100 ( .A(n9972), .B(n9971), .ZN(ADD_1068_U55) );
  OAI21_X1 U11101 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(ADD_1068_U56) );
  OAI21_X1 U11102 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(ADD_1068_U57) );
  OAI21_X1 U11103 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(ADD_1068_U58) );
  OAI21_X1 U11104 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(ADD_1068_U59) );
  OAI21_X1 U11105 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(ADD_1068_U60) );
  OAI21_X1 U11106 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(ADD_1068_U61) );
  OAI21_X1 U11107 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(ADD_1068_U62) );
  OAI21_X1 U11108 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(ADD_1068_U63) );
  NOR4_X1 U11109 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG2_REG_19__SCAN_IN), 
        .A3(P2_REG0_REG_19__SCAN_IN), .A4(P2_REG2_REG_12__SCAN_IN), .ZN(n9997)
         );
  NAND3_X1 U11110 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .A3(n9997), .ZN(n10006) );
  NOR4_X1 U11111 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .A3(P2_REG1_REG_16__SCAN_IN), .A4(P2_REG0_REG_14__SCAN_IN), .ZN(n10004) );
  NOR4_X1 U11112 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(SI_31_), .A4(P1_REG2_REG_30__SCAN_IN), .ZN(n10003) );
  NAND4_X1 U11113 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_REG0_REG_28__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P2_REG0_REG_20__SCAN_IN), .ZN(n10001) );
  NAND4_X1 U11114 ( .A1(P2_D_REG_0__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(P2_REG3_REG_15__SCAN_IN), .A4(P2_ADDR_REG_13__SCAN_IN), .ZN(n10000) );
  NAND4_X1 U11115 ( .A1(SI_25_), .A2(P1_DATAO_REG_25__SCAN_IN), .A3(
        P2_REG1_REG_13__SCAN_IN), .A4(P2_REG2_REG_0__SCAN_IN), .ZN(n9999) );
  NAND4_X1 U11116 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), 
        .A3(P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9998) );
  NOR4_X1 U11117 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10002) );
  NAND3_X1 U11118 ( .A1(n10004), .A2(n10003), .A3(n10002), .ZN(n10005) );
  NOR4_X1 U11119 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P2_REG1_REG_17__SCAN_IN), 
        .A3(n10006), .A4(n10005), .ZN(n10043) );
  NAND4_X1 U11120 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P1_REG0_REG_16__SCAN_IN), .A4(P1_REG2_REG_16__SCAN_IN), .ZN(n10010) );
  NAND4_X1 U11121 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_1__SCAN_IN), .A4(P1_ADDR_REG_16__SCAN_IN), .ZN(n10009)
         );
  NAND4_X1 U11122 ( .A1(P1_B_REG_SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), .A3(
        P2_REG1_REG_18__SCAN_IN), .A4(P2_REG2_REG_14__SCAN_IN), .ZN(n10008) );
  NAND4_X1 U11123 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P1_REG2_REG_17__SCAN_IN), 
        .A3(P2_REG3_REG_21__SCAN_IN), .A4(P2_REG2_REG_16__SCAN_IN), .ZN(n10007) );
  NOR4_X1 U11124 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n10042) );
  NAND4_X1 U11125 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_REG3_REG_19__SCAN_IN), .A4(P2_REG3_REG_3__SCAN_IN), .ZN(n10014) );
  NAND4_X1 U11126 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(P2_REG1_REG_8__SCAN_IN), 
        .A3(P2_REG2_REG_8__SCAN_IN), .A4(P2_REG2_REG_7__SCAN_IN), .ZN(n10013)
         );
  NAND4_X1 U11127 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(P1_REG1_REG_7__SCAN_IN), 
        .A3(P1_REG2_REG_2__SCAN_IN), .A4(P1_REG0_REG_1__SCAN_IN), .ZN(n10012)
         );
  NAND4_X1 U11128 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG0_REG_4__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n10011)
         );
  NOR4_X1 U11129 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10041) );
  NAND3_X1 U11130 ( .A1(n10016), .A2(n10015), .A3(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10017) );
  NOR3_X1 U11131 ( .A1(n10017), .A2(P1_RD_REG_SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n10019) );
  NAND3_X1 U11132 ( .A1(n10019), .A2(n10018), .A3(n10246), .ZN(n10039) );
  INV_X1 U11133 ( .A(SI_15_), .ZN(n10106) );
  NAND4_X1 U11134 ( .A1(SI_16_), .A2(SI_12_), .A3(n10257), .A4(n10106), .ZN(
        n10020) );
  NOR3_X1 U11135 ( .A1(SI_19_), .A2(n10110), .A3(n10020), .ZN(n10027) );
  NOR4_X1 U11136 ( .A1(P1_D_REG_10__SCAN_IN), .A2(SI_27_), .A3(
        P1_REG3_REG_8__SCAN_IN), .A4(P2_REG0_REG_29__SCAN_IN), .ZN(n10021) );
  NAND3_X1 U11137 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(n10021), .A3(n10241), .ZN(
        n10025) );
  NOR2_X1 U11138 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n10023) );
  NOR4_X1 U11139 ( .A1(SI_22_), .A2(P1_DATAO_REG_8__SCAN_IN), .A3(SI_6_), .A4(
        P1_DATAO_REG_1__SCAN_IN), .ZN(n10022) );
  NAND4_X1 U11140 ( .A1(n10155), .A2(P1_IR_REG_5__SCAN_IN), .A3(n10023), .A4(
        n10022), .ZN(n10024) );
  NOR4_X1 U11141 ( .A1(n10025), .A2(P2_DATAO_REG_30__SCAN_IN), .A3(
        P1_IR_REG_2__SCAN_IN), .A4(n10024), .ZN(n10026) );
  NAND4_X1 U11142 ( .A1(SI_17_), .A2(n10027), .A3(n10026), .A4(n5418), .ZN(
        n10038) );
  NOR4_X1 U11143 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), 
        .A3(P2_REG3_REG_1__SCAN_IN), .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n10031)
         );
  NOR4_X1 U11144 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG0_REG_11__SCAN_IN), 
        .A3(P2_REG0_REG_10__SCAN_IN), .A4(P2_REG0_REG_6__SCAN_IN), .ZN(n10030)
         );
  NOR4_X1 U11145 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(SI_28_), .A3(
        P1_REG2_REG_5__SCAN_IN), .A4(P1_REG2_REG_3__SCAN_IN), .ZN(n10029) );
  NOR4_X1 U11146 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .A3(P1_REG3_REG_9__SCAN_IN), .A4(P1_REG0_REG_5__SCAN_IN), .ZN(n10028)
         );
  NAND4_X1 U11147 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10037) );
  NOR4_X1 U11148 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(P2_REG1_REG_27__SCAN_IN), 
        .A3(P2_REG0_REG_26__SCAN_IN), .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n10035) );
  NOR4_X1 U11149 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_ADDR_REG_10__SCAN_IN), .ZN(n10034) );
  NOR4_X1 U11150 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .A3(P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n10033) );
  NOR4_X1 U11151 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(P2_REG1_REG_25__SCAN_IN), 
        .A3(P2_REG0_REG_24__SCAN_IN), .A4(P2_REG1_REG_21__SCAN_IN), .ZN(n10032) );
  NAND4_X1 U11152 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10036) );
  NOR4_X1 U11153 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n10040) );
  NAND4_X1 U11154 ( .A1(n10043), .A2(n10042), .A3(n10041), .A4(n10040), .ZN(
        n10290) );
  AOI222_X1 U11155 ( .A1(n10047), .A2(n10046), .B1(P2_DATAO_REG_22__SCAN_IN), 
        .B2(n10045), .C1(P1_STATE_REG_SCAN_IN), .C2(n10044), .ZN(n10288) );
  INV_X1 U11156 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U11157 ( .A1(n10050), .A2(keyinput110), .B1(n10049), .B2(keyinput79), .ZN(n10048) );
  OAI221_X1 U11158 ( .B1(n10050), .B2(keyinput110), .C1(n10049), .C2(
        keyinput79), .A(n10048), .ZN(n10060) );
  AOI22_X1 U11159 ( .A1(n10053), .A2(keyinput103), .B1(keyinput114), .B2(
        n10052), .ZN(n10051) );
  OAI221_X1 U11160 ( .B1(n10053), .B2(keyinput103), .C1(n10052), .C2(
        keyinput114), .A(n10051), .ZN(n10059) );
  XOR2_X1 U11161 ( .A(n8386), .B(keyinput101), .Z(n10057) );
  XNOR2_X1 U11162 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput59), .ZN(n10056) );
  XNOR2_X1 U11163 ( .A(SI_12_), .B(keyinput39), .ZN(n10055) );
  XNOR2_X1 U11164 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput25), .ZN(n10054) );
  NAND4_X1 U11165 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10058) );
  NOR3_X1 U11166 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(n10104) );
  AOI22_X1 U11167 ( .A1(n10062), .A2(keyinput68), .B1(n9341), .B2(keyinput4), 
        .ZN(n10061) );
  OAI221_X1 U11168 ( .B1(n10062), .B2(keyinput68), .C1(n9341), .C2(keyinput4), 
        .A(n10061), .ZN(n10074) );
  AOI22_X1 U11169 ( .A1(n10065), .A2(keyinput86), .B1(keyinput44), .B2(n10064), 
        .ZN(n10063) );
  OAI221_X1 U11170 ( .B1(n10065), .B2(keyinput86), .C1(n10064), .C2(keyinput44), .A(n10063), .ZN(n10073) );
  AOI22_X1 U11171 ( .A1(n10068), .A2(keyinput54), .B1(n10067), .B2(keyinput49), 
        .ZN(n10066) );
  OAI221_X1 U11172 ( .B1(n10068), .B2(keyinput54), .C1(n10067), .C2(keyinput49), .A(n10066), .ZN(n10072) );
  XNOR2_X1 U11173 ( .A(P2_REG0_REG_14__SCAN_IN), .B(keyinput105), .ZN(n10070)
         );
  XNOR2_X1 U11174 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput98), .ZN(n10069) );
  NAND2_X1 U11175 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  NOR4_X1 U11176 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10103) );
  AOI22_X1 U11177 ( .A1(n10077), .A2(keyinput2), .B1(keyinput38), .B2(n10076), 
        .ZN(n10075) );
  OAI221_X1 U11178 ( .B1(n10077), .B2(keyinput2), .C1(n10076), .C2(keyinput38), 
        .A(n10075), .ZN(n10086) );
  AOI22_X1 U11179 ( .A1(n10079), .A2(keyinput121), .B1(keyinput47), .B2(n5305), 
        .ZN(n10078) );
  OAI221_X1 U11180 ( .B1(n10079), .B2(keyinput121), .C1(n5305), .C2(keyinput47), .A(n10078), .ZN(n10085) );
  AOI22_X1 U11181 ( .A1(n7672), .A2(keyinput111), .B1(n5886), .B2(keyinput53), 
        .ZN(n10080) );
  OAI221_X1 U11182 ( .B1(n7672), .B2(keyinput111), .C1(n5886), .C2(keyinput53), 
        .A(n10080), .ZN(n10084) );
  INV_X1 U11183 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U11184 ( .A1(n5418), .A2(keyinput0), .B1(keyinput9), .B2(n10082), 
        .ZN(n10081) );
  OAI221_X1 U11185 ( .B1(n5418), .B2(keyinput0), .C1(n10082), .C2(keyinput9), 
        .A(n10081), .ZN(n10083) );
  NOR4_X1 U11186 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10102) );
  AOI22_X1 U11187 ( .A1(n10089), .A2(keyinput75), .B1(n10088), .B2(keyinput62), 
        .ZN(n10087) );
  OAI221_X1 U11188 ( .B1(n10089), .B2(keyinput75), .C1(n10088), .C2(keyinput62), .A(n10087), .ZN(n10100) );
  AOI22_X1 U11189 ( .A1(n5836), .A2(keyinput34), .B1(keyinput66), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11190 ( .B1(n5836), .B2(keyinput34), .C1(n10091), .C2(keyinput66), 
        .A(n10090), .ZN(n10099) );
  INV_X1 U11191 ( .A(SI_6_), .ZN(n10094) );
  AOI22_X1 U11192 ( .A1(n5759), .A2(keyinput6), .B1(keyinput96), .B2(n10096), 
        .ZN(n10095) );
  OAI221_X1 U11193 ( .B1(n5759), .B2(keyinput6), .C1(n10096), .C2(keyinput96), 
        .A(n10095), .ZN(n10097) );
  NOR4_X1 U11194 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10101) );
  NAND4_X1 U11195 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10286) );
  AOI22_X1 U11196 ( .A1(n10106), .A2(keyinput123), .B1(keyinput32), .B2(n5975), 
        .ZN(n10105) );
  OAI221_X1 U11197 ( .B1(n10106), .B2(keyinput123), .C1(n5975), .C2(keyinput32), .A(n10105), .ZN(n10118) );
  AOI22_X1 U11198 ( .A1(n10108), .A2(keyinput89), .B1(keyinput124), .B2(n7604), 
        .ZN(n10107) );
  OAI221_X1 U11199 ( .B1(n10108), .B2(keyinput89), .C1(n7604), .C2(keyinput124), .A(n10107), .ZN(n10117) );
  INV_X1 U11200 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U11201 ( .A1(n10111), .A2(keyinput92), .B1(n10110), .B2(keyinput18), 
        .ZN(n10109) );
  OAI221_X1 U11202 ( .B1(n10111), .B2(keyinput92), .C1(n10110), .C2(keyinput18), .A(n10109), .ZN(n10116) );
  AOI22_X1 U11203 ( .A1(n10114), .A2(keyinput113), .B1(n10113), .B2(
        keyinput106), .ZN(n10112) );
  OAI221_X1 U11204 ( .B1(n10114), .B2(keyinput113), .C1(n10113), .C2(
        keyinput106), .A(n10112), .ZN(n10115) );
  NOR4_X1 U11205 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10163) );
  AOI22_X1 U11206 ( .A1(n10121), .A2(keyinput107), .B1(n10120), .B2(keyinput41), .ZN(n10119) );
  OAI221_X1 U11207 ( .B1(n10121), .B2(keyinput107), .C1(n10120), .C2(
        keyinput41), .A(n10119), .ZN(n10133) );
  AOI22_X1 U11208 ( .A1(n10124), .A2(keyinput112), .B1(keyinput56), .B2(n10123), .ZN(n10122) );
  OAI221_X1 U11209 ( .B1(n10124), .B2(keyinput112), .C1(n10123), .C2(
        keyinput56), .A(n10122), .ZN(n10132) );
  AOI22_X1 U11210 ( .A1(n10127), .A2(keyinput82), .B1(n10126), .B2(keyinput109), .ZN(n10125) );
  OAI221_X1 U11211 ( .B1(n10127), .B2(keyinput82), .C1(n10126), .C2(
        keyinput109), .A(n10125), .ZN(n10131) );
  XOR2_X1 U11212 ( .A(n7109), .B(keyinput99), .Z(n10129) );
  XNOR2_X1 U11213 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput57), .ZN(n10128) );
  NAND2_X1 U11214 ( .A1(n10129), .A2(n10128), .ZN(n10130) );
  NOR4_X1 U11215 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10162) );
  AOI22_X1 U11216 ( .A1(n10135), .A2(keyinput55), .B1(n6479), .B2(keyinput36), 
        .ZN(n10134) );
  OAI221_X1 U11217 ( .B1(n10135), .B2(keyinput55), .C1(n6479), .C2(keyinput36), 
        .A(n10134), .ZN(n10145) );
  INV_X1 U11218 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U11219 ( .A1(n5862), .A2(keyinput87), .B1(keyinput50), .B2(n10137), 
        .ZN(n10136) );
  OAI221_X1 U11220 ( .B1(n5862), .B2(keyinput87), .C1(n10137), .C2(keyinput50), 
        .A(n10136), .ZN(n10144) );
  XNOR2_X1 U11221 ( .A(n10138), .B(keyinput116), .ZN(n10143) );
  XOR2_X1 U11222 ( .A(n5872), .B(keyinput10), .Z(n10141) );
  XNOR2_X1 U11223 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput8), .ZN(n10140) );
  XNOR2_X1 U11224 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput45), .ZN(n10139) );
  NAND3_X1 U11225 ( .A1(n10141), .A2(n10140), .A3(n10139), .ZN(n10142) );
  NOR4_X1 U11226 ( .A1(n10145), .A2(n10144), .A3(n10143), .A4(n10142), .ZN(
        n10161) );
  AOI22_X1 U11227 ( .A1(n10147), .A2(keyinput126), .B1(n5043), .B2(keyinput64), 
        .ZN(n10146) );
  OAI221_X1 U11228 ( .B1(n10147), .B2(keyinput126), .C1(n5043), .C2(keyinput64), .A(n10146), .ZN(n10159) );
  INV_X1 U11229 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U11230 ( .A1(n10150), .A2(keyinput84), .B1(keyinput90), .B2(n10149), 
        .ZN(n10148) );
  OAI221_X1 U11231 ( .B1(n10150), .B2(keyinput84), .C1(n10149), .C2(keyinput90), .A(n10148), .ZN(n10158) );
  AOI22_X1 U11232 ( .A1(n10152), .A2(keyinput70), .B1(n6006), .B2(keyinput14), 
        .ZN(n10151) );
  OAI221_X1 U11233 ( .B1(n10152), .B2(keyinput70), .C1(n6006), .C2(keyinput14), 
        .A(n10151), .ZN(n10157) );
  AOI22_X1 U11234 ( .A1(n10155), .A2(keyinput88), .B1(keyinput67), .B2(n10154), 
        .ZN(n10153) );
  OAI221_X1 U11235 ( .B1(n10155), .B2(keyinput88), .C1(n10154), .C2(keyinput67), .A(n10153), .ZN(n10156) );
  NOR4_X1 U11236 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  NAND4_X1 U11237 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10285) );
  AOI22_X1 U11238 ( .A1(n6818), .A2(keyinput74), .B1(n10165), .B2(keyinput16), 
        .ZN(n10164) );
  OAI221_X1 U11239 ( .B1(n6818), .B2(keyinput74), .C1(n10165), .C2(keyinput16), 
        .A(n10164), .ZN(n10176) );
  AOI22_X1 U11240 ( .A1(n10167), .A2(keyinput102), .B1(keyinput22), .B2(n5681), 
        .ZN(n10166) );
  OAI221_X1 U11241 ( .B1(n10167), .B2(keyinput102), .C1(n5681), .C2(keyinput22), .A(n10166), .ZN(n10175) );
  AOI22_X1 U11242 ( .A1(n10170), .A2(keyinput119), .B1(n10169), .B2(keyinput78), .ZN(n10168) );
  OAI221_X1 U11243 ( .B1(n10170), .B2(keyinput119), .C1(n10169), .C2(
        keyinput78), .A(n10168), .ZN(n10174) );
  XOR2_X1 U11244 ( .A(n5202), .B(keyinput125), .Z(n10172) );
  XNOR2_X1 U11245 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput11), .ZN(n10171) );
  NAND2_X1 U11246 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  NOR4_X1 U11247 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10223) );
  AOI22_X1 U11248 ( .A1(n10178), .A2(keyinput31), .B1(keyinput52), .B2(n7082), 
        .ZN(n10177) );
  OAI221_X1 U11249 ( .B1(n10178), .B2(keyinput31), .C1(n7082), .C2(keyinput52), 
        .A(n10177), .ZN(n10188) );
  AOI22_X1 U11250 ( .A1(n10180), .A2(keyinput72), .B1(keyinput71), .B2(n5676), 
        .ZN(n10179) );
  OAI221_X1 U11251 ( .B1(n10180), .B2(keyinput72), .C1(n5676), .C2(keyinput71), 
        .A(n10179), .ZN(n10187) );
  AOI22_X1 U11252 ( .A1(n6073), .A2(keyinput5), .B1(keyinput63), .B2(n10182), 
        .ZN(n10181) );
  OAI221_X1 U11253 ( .B1(n6073), .B2(keyinput5), .C1(n10182), .C2(keyinput63), 
        .A(n10181), .ZN(n10186) );
  XOR2_X1 U11254 ( .A(n5105), .B(keyinput97), .Z(n10184) );
  XNOR2_X1 U11255 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput42), .ZN(n10183) );
  NAND2_X1 U11256 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NOR4_X1 U11257 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10222) );
  AOI22_X1 U11258 ( .A1(n10191), .A2(keyinput46), .B1(keyinput83), .B2(n10190), 
        .ZN(n10189) );
  OAI221_X1 U11259 ( .B1(n10191), .B2(keyinput46), .C1(n10190), .C2(keyinput83), .A(n10189), .ZN(n10204) );
  INV_X1 U11260 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11261 ( .A1(n10194), .A2(keyinput91), .B1(keyinput115), .B2(n10193), .ZN(n10192) );
  OAI221_X1 U11262 ( .B1(n10194), .B2(keyinput91), .C1(n10193), .C2(
        keyinput115), .A(n10192), .ZN(n10203) );
  AOI22_X1 U11263 ( .A1(n10197), .A2(keyinput81), .B1(keyinput65), .B2(n10196), 
        .ZN(n10195) );
  OAI221_X1 U11264 ( .B1(n10197), .B2(keyinput81), .C1(n10196), .C2(keyinput65), .A(n10195), .ZN(n10202) );
  AOI22_X1 U11265 ( .A1(n10200), .A2(keyinput12), .B1(n10199), .B2(keyinput127), .ZN(n10198) );
  OAI221_X1 U11266 ( .B1(n10200), .B2(keyinput12), .C1(n10199), .C2(
        keyinput127), .A(n10198), .ZN(n10201) );
  NOR4_X1 U11267 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        n10221) );
  AOI22_X1 U11268 ( .A1(n10207), .A2(keyinput104), .B1(keyinput120), .B2(
        n10206), .ZN(n10205) );
  OAI221_X1 U11269 ( .B1(n10207), .B2(keyinput104), .C1(n10206), .C2(
        keyinput120), .A(n10205), .ZN(n10219) );
  AOI22_X1 U11270 ( .A1(n10210), .A2(keyinput29), .B1(keyinput40), .B2(n10209), 
        .ZN(n10208) );
  OAI221_X1 U11271 ( .B1(n10210), .B2(keyinput29), .C1(n10209), .C2(keyinput40), .A(n10208), .ZN(n10218) );
  AOI22_X1 U11272 ( .A1(n10213), .A2(keyinput48), .B1(n10212), .B2(keyinput94), 
        .ZN(n10211) );
  OAI221_X1 U11273 ( .B1(n10213), .B2(keyinput48), .C1(n10212), .C2(keyinput94), .A(n10211), .ZN(n10217) );
  XNOR2_X1 U11274 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput93), .ZN(n10215)
         );
  XNOR2_X1 U11275 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput60), .ZN(n10214) );
  NAND2_X1 U11276 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  NOR4_X1 U11277 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  NAND4_X1 U11278 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10284) );
  AOI22_X1 U11279 ( .A1(n4591), .A2(keyinput20), .B1(keyinput85), .B2(n10225), 
        .ZN(n10224) );
  OAI221_X1 U11280 ( .B1(n4591), .B2(keyinput20), .C1(n10225), .C2(keyinput85), 
        .A(n10224), .ZN(n10235) );
  AOI22_X1 U11281 ( .A1(n10228), .A2(keyinput76), .B1(n10227), .B2(keyinput24), 
        .ZN(n10226) );
  OAI221_X1 U11282 ( .B1(n10228), .B2(keyinput76), .C1(n10227), .C2(keyinput24), .A(n10226), .ZN(n10234) );
  XOR2_X1 U11283 ( .A(n5247), .B(keyinput73), .Z(n10232) );
  XNOR2_X1 U11284 ( .A(SI_17_), .B(keyinput3), .ZN(n10231) );
  XNOR2_X1 U11285 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput17), .ZN(n10230) );
  XNOR2_X1 U11286 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput26), .ZN(n10229) );
  NAND4_X1 U11287 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10233) );
  NOR3_X1 U11288 ( .A1(n10235), .A2(n10234), .A3(n10233), .ZN(n10282) );
  AOI22_X1 U11289 ( .A1(n10238), .A2(keyinput118), .B1(keyinput80), .B2(n10237), .ZN(n10236) );
  OAI221_X1 U11290 ( .B1(n10238), .B2(keyinput118), .C1(n10237), .C2(
        keyinput80), .A(n10236), .ZN(n10251) );
  INV_X1 U11291 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11292 ( .A1(n10241), .A2(keyinput95), .B1(n10240), .B2(keyinput61), 
        .ZN(n10239) );
  OAI221_X1 U11293 ( .B1(n10241), .B2(keyinput95), .C1(n10240), .C2(keyinput61), .A(n10239), .ZN(n10250) );
  AOI22_X1 U11294 ( .A1(n10244), .A2(keyinput69), .B1(keyinput7), .B2(n10243), 
        .ZN(n10242) );
  OAI221_X1 U11295 ( .B1(n10244), .B2(keyinput69), .C1(n10243), .C2(keyinput7), 
        .A(n10242), .ZN(n10249) );
  AOI22_X1 U11296 ( .A1(n10247), .A2(keyinput108), .B1(keyinput100), .B2(
        n10246), .ZN(n10245) );
  OAI221_X1 U11297 ( .B1(n10247), .B2(keyinput108), .C1(n10246), .C2(
        keyinput100), .A(n10245), .ZN(n10248) );
  NOR4_X1 U11298 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10281) );
  AOI22_X1 U11299 ( .A1(n7412), .A2(keyinput37), .B1(keyinput43), .B2(n10253), 
        .ZN(n10252) );
  OAI221_X1 U11300 ( .B1(n7412), .B2(keyinput37), .C1(n10253), .C2(keyinput43), 
        .A(n10252), .ZN(n10264) );
  AOI22_X1 U11301 ( .A1(n10255), .A2(keyinput117), .B1(keyinput1), .B2(n5333), 
        .ZN(n10254) );
  OAI221_X1 U11302 ( .B1(n10255), .B2(keyinput117), .C1(n5333), .C2(keyinput1), 
        .A(n10254), .ZN(n10263) );
  AOI22_X1 U11303 ( .A1(n10258), .A2(keyinput27), .B1(keyinput122), .B2(n10257), .ZN(n10256) );
  OAI221_X1 U11304 ( .B1(n10258), .B2(keyinput27), .C1(n10257), .C2(
        keyinput122), .A(n10256), .ZN(n10262) );
  XOR2_X1 U11305 ( .A(n5174), .B(keyinput77), .Z(n10260) );
  XNOR2_X1 U11306 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput30), .ZN(n10259) );
  NAND2_X1 U11307 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  NOR4_X1 U11308 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10280) );
  AOI22_X1 U11309 ( .A1(n10267), .A2(keyinput23), .B1(keyinput19), .B2(n10266), 
        .ZN(n10265) );
  OAI221_X1 U11310 ( .B1(n10267), .B2(keyinput23), .C1(n10266), .C2(keyinput19), .A(n10265), .ZN(n10278) );
  AOI22_X1 U11311 ( .A1(n9222), .A2(keyinput15), .B1(keyinput13), .B2(n10269), 
        .ZN(n10268) );
  OAI221_X1 U11312 ( .B1(n9222), .B2(keyinput15), .C1(n10269), .C2(keyinput13), 
        .A(n10268), .ZN(n10277) );
  INV_X1 U11313 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U11314 ( .A1(n10272), .A2(keyinput35), .B1(keyinput28), .B2(n10271), 
        .ZN(n10270) );
  OAI221_X1 U11315 ( .B1(n10272), .B2(keyinput35), .C1(n10271), .C2(keyinput28), .A(n10270), .ZN(n10276) );
  XNOR2_X1 U11316 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput33), .ZN(n10274)
         );
  XNOR2_X1 U11317 ( .A(P1_REG2_REG_26__SCAN_IN), .B(keyinput51), .ZN(n10273)
         );
  NAND2_X1 U11318 ( .A1(n10274), .A2(n10273), .ZN(n10275) );
  NOR4_X1 U11319 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10279) );
  NAND4_X1 U11320 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10283) );
  NOR4_X1 U11321 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10287) );
  XNOR2_X1 U11322 ( .A(n10288), .B(n10287), .ZN(n10289) );
  XNOR2_X1 U11323 ( .A(n10290), .B(n10289), .ZN(P1_U3333) );
  OAI21_X1 U11324 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(ADD_1068_U50) );
  OAI21_X1 U11325 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(ADD_1068_U51) );
  OAI21_X1 U11326 ( .B1(n10299), .B2(n10298), .A(n10297), .ZN(ADD_1068_U47) );
  OAI21_X1 U11327 ( .B1(n10302), .B2(n10301), .A(n10300), .ZN(ADD_1068_U49) );
  OAI21_X1 U11328 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(ADD_1068_U48) );
  AOI21_X1 U11329 ( .B1(n10308), .B2(n10307), .A(n10306), .ZN(ADD_1068_U54) );
  AOI21_X1 U11330 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(ADD_1068_U53) );
  OAI21_X1 U11331 ( .B1(n10314), .B2(n10313), .A(n10312), .ZN(ADD_1068_U52) );
  AND3_X1 U5974 ( .A1(n5083), .A2(n5082), .A3(n5081), .ZN(n9884) );
  CLKBUF_X1 U5978 ( .A(n6422), .Z(n6466) );
  CLKBUF_X1 U6596 ( .A(n5805), .Z(n7682) );
endmodule

