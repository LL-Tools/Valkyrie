

module b20_C_SARLock_k_64_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133;

  NAND2_X1 U4795 ( .A1(n8180), .A2(n8232), .ZN(n8235) );
  NAND2_X1 U4796 ( .A1(n8497), .A2(n8498), .ZN(n8804) );
  CLKBUF_X2 U4797 ( .A(n6214), .Z(n6264) );
  AND3_X1 U4798 ( .A1(n4937), .A2(n4936), .A3(n4935), .ZN(n7321) );
  INV_X1 U4799 ( .A(n7048), .ZN(n9855) );
  INV_X2 U4800 ( .A(n8715), .ZN(n6091) );
  NAND2_X1 U4801 ( .A1(n4322), .A2(n4894), .ZN(n5517) );
  INV_X1 U4802 ( .A(n5738), .ZN(n6046) );
  CLKBUF_X2 U4803 ( .A(n5726), .Z(n6069) );
  AND2_X1 U4804 ( .A1(n6378), .A2(n6379), .ZN(n5671) );
  INV_X2 U4805 ( .A(n4315), .ZN(n5726) );
  NAND2_X1 U4806 ( .A1(n6102), .A2(n6101), .ZN(n7803) );
  CLKBUF_X1 U4807 ( .A(n6725), .Z(n4289) );
  OR2_X1 U4808 ( .A1(n6100), .A2(n4300), .ZN(n6101) );
  NAND2_X1 U4809 ( .A1(n6642), .A2(n4907), .ZN(n5827) );
  NAND2_X1 U4810 ( .A1(n5686), .A2(n9033), .ZN(n8309) );
  INV_X2 U4812 ( .A(n9092), .ZN(n6234) );
  NAND2_X1 U4813 ( .A1(n5704), .A2(n5703), .ZN(n8366) );
  OAI211_X1 U4814 ( .C1(n4310), .C2(n6727), .A(n5737), .B(n5736), .ZN(n6835)
         );
  OAI211_X1 U4815 ( .C1(n6590), .C2(n5074), .A(n4918), .B(n4917), .ZN(n7259)
         );
  XNOR2_X1 U4816 ( .A(n8316), .B(n4572), .ZN(n6558) );
  INV_X1 U4817 ( .A(n8825), .ZN(n8796) );
  INV_X1 U4818 ( .A(n8333), .ZN(n8386) );
  AND2_X1 U4819 ( .A1(n4528), .A2(n4321), .ZN(n5851) );
  INV_X2 U4820 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U4821 ( .A1(n6624), .A2(n6189), .ZN(n9085) );
  INV_X1 U4822 ( .A(n7458), .ZN(n7568) );
  AND3_X1 U4823 ( .A1(n4977), .A2(n4976), .A3(n4975), .ZN(n7433) );
  INV_X1 U4824 ( .A(n7259), .ZN(n10097) );
  AND3_X2 U4825 ( .A1(n4891), .A2(n4890), .A3(n4889), .ZN(n7103) );
  AND4_X1 U4826 ( .A1(n5692), .A2(n5691), .A3(n5690), .A4(n5689), .ZN(n6800)
         );
  NAND2_X1 U4827 ( .A1(n6141), .A2(n8465), .ZN(n8886) );
  OAI21_X1 U4828 ( .B1(n6605), .B2(n5827), .A(n5826), .ZN(n9878) );
  NAND2_X1 U4829 ( .A1(n6106), .A2(n6107), .ZN(n6110) );
  NAND2_X1 U4830 ( .A1(n9023), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5682) );
  CLKBUF_X2 U4831 ( .A(n4926), .Z(n5495) );
  INV_X1 U4832 ( .A(n4939), .ZN(n5462) );
  NAND2_X1 U4833 ( .A1(n5671), .A2(n6383), .ZN(n6624) );
  INV_X1 U4834 ( .A(n7103), .ZN(n9770) );
  NAND4_X2 U4835 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8563)
         );
  INV_X1 U4836 ( .A(n9837), .ZN(n9839) );
  INV_X1 U4837 ( .A(n5687), .ZN(n9033) );
  XNOR2_X1 U4838 ( .A(n5746), .B(n5745), .ZN(n6859) );
  INV_X1 U4839 ( .A(n5545), .ZN(n7419) );
  NAND2_X1 U4840 ( .A1(n4309), .A2(n6572), .ZN(n4288) );
  OAI21_X2 U4841 ( .B1(n9156), .B2(n4589), .A(n4319), .ZN(n6434) );
  AND3_X1 U4842 ( .A1(n4895), .A2(n4438), .A3(n4439), .ZN(n4322) );
  NOR2_X2 U4843 ( .A1(n5693), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5683) );
  OAI21_X2 U4844 ( .B1(n8188), .B2(n8187), .A(n8189), .ZN(n8211) );
  NAND2_X2 U4845 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  NAND2_X4 U4846 ( .A1(n5686), .A2(n5687), .ZN(n5940) );
  XNOR2_X1 U4848 ( .A(n5721), .B(n9983), .ZN(n6725) );
  XNOR2_X2 U4849 ( .A(n4539), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8715) );
  NAND2_X4 U4850 ( .A1(n4311), .A2(n6196), .ZN(n9092) );
  XNOR2_X2 U4851 ( .A(n5682), .B(n9024), .ZN(n5688) );
  OAI21_X2 U4852 ( .B1(n6110), .B2(P2_D_REG_0__SCAN_IN), .A(n6601), .ZN(n6797)
         );
  OAI21_X1 U4853 ( .B1(n6558), .B2(n9833), .A(n4292), .ZN(n4291) );
  NAND2_X1 U4854 ( .A1(n8833), .A2(n8837), .ZN(n8835) );
  NAND2_X1 U4855 ( .A1(n4633), .A2(n4327), .ZN(n8851) );
  NAND2_X1 U4856 ( .A1(n8886), .A2(n8471), .ZN(n4633) );
  NAND2_X1 U4857 ( .A1(n4457), .A2(n5966), .ZN(n5985) );
  NAND2_X1 U4858 ( .A1(n7043), .A2(n7042), .ZN(n7271) );
  AND2_X1 U4859 ( .A1(n6225), .A2(n6224), .ZN(n7200) );
  NAND2_X1 U4860 ( .A1(n4304), .A2(n8328), .ZN(n7182) );
  OR3_X1 U4861 ( .A1(n5797), .A2(n5796), .A3(n5795), .ZN(n8418) );
  NAND2_X1 U4862 ( .A1(n8396), .A2(n8389), .ZN(n8333) );
  NAND2_X1 U4863 ( .A1(n6134), .A2(n7176), .ZN(n8331) );
  INV_X1 U4864 ( .A(n8560), .ZN(n8431) );
  NAND2_X1 U4865 ( .A1(n5750), .A2(n7005), .ZN(n8389) );
  INV_X1 U4866 ( .A(n8946), .ZN(n5703) );
  INV_X2 U4868 ( .A(n5971), .ZN(n5738) );
  NAND2_X2 U4869 ( .A1(n4866), .A2(n4867), .ZN(n4939) );
  CLKBUF_X1 U4870 ( .A(n4920), .Z(n5472) );
  INV_X1 U4871 ( .A(n9726), .ZN(n4867) );
  NAND2_X2 U4872 ( .A1(n4866), .A2(n9726), .ZN(n4979) );
  NAND2_X1 U4873 ( .A1(n4310), .A2(n6572), .ZN(n4313) );
  AND2_X1 U4874 ( .A1(n5669), .A2(n4352), .ZN(n6379) );
  INV_X1 U4875 ( .A(n4997), .ZN(n4998) );
  OAI21_X1 U4876 ( .B1(n4973), .B2(n4887), .A(n4886), .ZN(n4909) );
  INV_X2 U4877 ( .A(n4907), .ZN(n4973) );
  NOR2_X1 U4879 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4574) );
  INV_X1 U4880 ( .A(n4291), .ZN(n8163) );
  AND2_X1 U4881 ( .A1(n4567), .A2(n4568), .ZN(n4848) );
  AOI21_X1 U4882 ( .B1(n4341), .B2(n8209), .A(n8208), .ZN(n8210) );
  AND2_X1 U4883 ( .A1(n6557), .A2(n6551), .ZN(n4292) );
  NAND2_X1 U4884 ( .A1(n4301), .A2(n8511), .ZN(n8749) );
  AOI211_X1 U4885 ( .C1(n8728), .C2(n8727), .A(n8726), .B(n8725), .ZN(n8729)
         );
  AND2_X1 U4886 ( .A1(n8255), .A2(n4748), .ZN(n4744) );
  NAND2_X1 U4887 ( .A1(n6150), .A2(n4647), .ZN(n4301) );
  AOI211_X1 U4888 ( .C1(n8676), .C2(n8692), .A(n8675), .B(n8674), .ZN(n8677)
         );
  NAND2_X1 U4889 ( .A1(n8766), .A2(n8503), .ZN(n6150) );
  NOR2_X1 U4890 ( .A1(n8672), .A2(n8938), .ZN(n8685) );
  NAND2_X1 U4891 ( .A1(n8835), .A2(n8479), .ZN(n8813) );
  AOI21_X1 U4892 ( .B1(n9503), .B2(n6490), .A(n6489), .ZN(n9491) );
  AOI21_X1 U4893 ( .B1(n9524), .B2(n6488), .A(n6487), .ZN(n9503) );
  AOI21_X1 U4894 ( .B1(n9535), .B2(n6486), .A(n4840), .ZN(n9524) );
  AOI21_X1 U4895 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8622), .A(n8621), .ZN(
        n8645) );
  NAND2_X1 U4896 ( .A1(n8851), .A2(n6144), .ZN(n8855) );
  AND2_X1 U4897 ( .A1(n4611), .A2(n4609), .ZN(n4608) );
  AOI21_X1 U4898 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8622), .A(n8610), .ZN(
        n8630) );
  NOR2_X1 U4899 ( .A1(n7956), .A2(n5886), .ZN(n8599) );
  NAND2_X1 U4900 ( .A1(n7667), .A2(n7666), .ZN(n7679) );
  NAND2_X1 U4901 ( .A1(n7829), .A2(n7830), .ZN(n7954) );
  NAND2_X1 U4902 ( .A1(n7482), .A2(n8446), .ZN(n7749) );
  NAND2_X1 U4903 ( .A1(n4684), .A2(n4344), .ZN(n7829) );
  OR2_X1 U4904 ( .A1(n7535), .A2(n5855), .ZN(n4684) );
  AND2_X1 U4905 ( .A1(n8496), .A2(n8488), .ZN(n8819) );
  NAND2_X1 U4906 ( .A1(n7442), .A2(n6138), .ZN(n7482) );
  NOR2_X1 U4907 ( .A1(n7596), .A2(n4397), .ZN(n7824) );
  NAND2_X1 U4908 ( .A1(n5978), .A2(n5977), .ZN(n8830) );
  NAND2_X1 U4909 ( .A1(n6243), .A2(n4828), .ZN(n6246) );
  NAND2_X1 U4910 ( .A1(n7271), .A2(n4369), .ZN(n7283) );
  NAND2_X1 U4911 ( .A1(n4293), .A2(n8400), .ZN(n7158) );
  NOR2_X1 U4912 ( .A1(n7496), .A2(n4660), .ZN(n7532) );
  NAND2_X1 U4913 ( .A1(n4296), .A2(n4294), .ZN(n4293) );
  NAND2_X1 U4914 ( .A1(n5126), .A2(n5125), .ZN(n9124) );
  NOR2_X1 U4915 ( .A1(n7220), .A2(n7219), .ZN(n7496) );
  AND2_X1 U4916 ( .A1(n4624), .A2(n4622), .ZN(n4297) );
  NAND2_X1 U4917 ( .A1(n7182), .A2(n6133), .ZN(n7149) );
  XNOR2_X1 U4918 ( .A(n6213), .B(n6355), .ZN(n7365) );
  XNOR2_X1 U4919 ( .A(n6217), .B(n6355), .ZN(n7363) );
  OR2_X1 U4920 ( .A1(n5120), .A2(n5119), .ZN(n4734) );
  INV_X1 U4921 ( .A(n8335), .ZN(n4295) );
  NAND2_X1 U4922 ( .A1(n6805), .A2(n6806), .ZN(n6821) );
  AND2_X1 U4923 ( .A1(n5090), .A2(n4573), .ZN(n6605) );
  INV_X1 U4924 ( .A(n8401), .ZN(n4294) );
  NAND2_X1 U4925 ( .A1(n8373), .A2(n8366), .ZN(n9820) );
  OR2_X1 U4926 ( .A1(n7078), .A2(n7205), .ZN(n7077) );
  NAND2_X1 U4927 ( .A1(n7055), .A2(n8368), .ZN(n8373) );
  NAND2_X1 U4928 ( .A1(n6132), .A2(n6813), .ZN(n7055) );
  CLKBUF_X1 U4929 ( .A(n6131), .Z(n8566) );
  NAND2_X1 U4930 ( .A1(n6123), .A2(n8320), .ZN(n9829) );
  OR2_X1 U4931 ( .A1(n8376), .A2(n6839), .ZN(n6134) );
  AND4_X1 U4932 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n8419)
         );
  AND4_X2 U4933 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n5750)
         );
  AND3_X1 U4934 ( .A1(n5717), .A2(n4303), .A3(n5718), .ZN(n4302) );
  INV_X1 U4935 ( .A(n6835), .ZN(n6839) );
  AND4_X2 U4936 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n8376)
         );
  NAND2_X1 U4937 ( .A1(n4681), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4680) );
  AND4_X1 U4938 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n7305)
         );
  OR2_X1 U4939 ( .A1(n4307), .A2(n6715), .ZN(n4303) );
  NAND4_X1 U4940 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n9270)
         );
  CLKBUF_X3 U4941 ( .A(n8309), .Z(n4306) );
  CLKBUF_X3 U4942 ( .A(n8309), .Z(n4307) );
  INV_X1 U4943 ( .A(n8377), .ZN(n9841) );
  AND2_X2 U4944 ( .A1(n5004), .A2(n5663), .ZN(n6508) );
  CLKBUF_X1 U4945 ( .A(n5038), .Z(n5298) );
  AOI21_X1 U4946 ( .B1(n4450), .B2(n4452), .A(n4448), .ZN(n4447) );
  XNOR2_X1 U4947 ( .A(n5963), .B(n5962), .ZN(n6127) );
  OAI211_X1 U4948 ( .C1(n4310), .C2(n4289), .A(n5723), .B(n5722), .ZN(n8377)
         );
  OAI211_X1 U4949 ( .C1(n6642), .C2(n6704), .A(n5702), .B(n5701), .ZN(n8946)
         );
  OR2_X1 U4950 ( .A1(n4313), .A2(n6574), .ZN(n5737) );
  NAND2_X1 U4951 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  INV_X1 U4952 ( .A(n5971), .ZN(n4290) );
  XNOR2_X1 U4953 ( .A(n6099), .B(n4298), .ZN(n7879) );
  NAND2_X1 U4954 ( .A1(n5091), .A2(n4907), .ZN(n5038) );
  AOI21_X1 U4955 ( .B1(n4719), .B2(n5039), .A(n4451), .ZN(n4450) );
  NAND2_X1 U4956 ( .A1(n4864), .A2(n4433), .ZN(n9726) );
  NOR2_X1 U4957 ( .A1(n5049), .A2(n4720), .ZN(n4719) );
  MUX2_X1 U4958 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4863), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4864) );
  XNOR2_X1 U4959 ( .A(n5507), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U4960 ( .A1(n5620), .A2(n7402), .ZN(n6504) );
  NAND2_X1 U4961 ( .A1(n4339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  NAND2_X2 U4962 ( .A1(n6090), .A2(n6659), .ZN(n6642) );
  NAND2_X1 U4963 ( .A1(n4998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5507) );
  XNOR2_X1 U4964 ( .A(n5695), .B(n5694), .ZN(n6090) );
  INV_X1 U4965 ( .A(n5619), .ZN(n5620) );
  INV_X1 U4966 ( .A(n8715), .ZN(n6659) );
  MUX2_X1 U4967 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4877), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4878) );
  XNOR2_X1 U4968 ( .A(n5548), .B(n5547), .ZN(n7402) );
  OR2_X1 U4969 ( .A1(n5780), .A2(n5779), .ZN(n7074) );
  NAND2_X1 U4970 ( .A1(n4876), .A2(n4861), .ZN(n4879) );
  NAND2_X1 U4971 ( .A1(n4873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U4972 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U4973 ( .A1(n6104), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5696) );
  AND2_X1 U4974 ( .A1(n4325), .A2(n4391), .ZN(n4818) );
  NAND2_X1 U4975 ( .A1(n5734), .A2(n5761), .ZN(n6727) );
  NOR2_X1 U4976 ( .A1(n5761), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5764) );
  NOR2_X1 U4977 ( .A1(n4655), .A2(n4354), .ZN(n4654) );
  NAND2_X1 U4978 ( .A1(n4882), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4469) );
  AND2_X1 U4979 ( .A1(n4349), .A2(n4321), .ZN(n4531) );
  AND2_X1 U4980 ( .A1(n4772), .A2(n4530), .ZN(n4529) );
  OR2_X1 U4981 ( .A1(n5733), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5761) );
  AND2_X1 U4982 ( .A1(n4767), .A2(n4772), .ZN(n4528) );
  AND2_X1 U4983 ( .A1(n4816), .A2(n4814), .ZN(n4813) );
  INV_X1 U4984 ( .A(n4656), .ZN(n4655) );
  AND4_X1 U4985 ( .A1(n4856), .A2(n4855), .A3(n4857), .A4(n4854), .ZN(n4837)
         );
  AND4_X1 U4986 ( .A1(n4770), .A2(n9983), .A3(n4768), .A4(n4769), .ZN(n4767)
         );
  AND2_X1 U4987 ( .A1(n5777), .A2(n5763), .ZN(n4772) );
  AND4_X1 U4988 ( .A1(n4771), .A2(n6649), .A3(n5793), .A4(n5745), .ZN(n4321)
         );
  AND2_X1 U4989 ( .A1(n5679), .A2(n5680), .ZN(n4656) );
  AND2_X1 U4990 ( .A1(n4853), .A2(n4817), .ZN(n4816) );
  NOR2_X1 U4991 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4853) );
  NOR2_X1 U4992 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5920) );
  INV_X1 U4993 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4854) );
  NOR2_X1 U4994 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4857) );
  NOR2_X1 U4995 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4855) );
  INV_X1 U4996 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4298) );
  NOR2_X1 U4997 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4856) );
  INV_X1 U4998 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5850) );
  INV_X1 U4999 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5962) );
  INV_X1 U5000 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5950) );
  INV_X1 U5001 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4769) );
  INV_X1 U5002 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4771) );
  INV_X1 U5003 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4299) );
  INV_X1 U5004 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4300) );
  NOR3_X1 U5005 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n4858) );
  NOR2_X2 U5006 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4912) );
  INV_X4 U5007 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5008 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  XNOR2_X1 U5009 ( .A(n4296), .B(n4295), .ZN(n9859) );
  NAND2_X1 U5010 ( .A1(n4621), .A2(n4297), .ZN(n4296) );
  NAND3_X1 U5011 ( .A1(n4300), .A2(n4299), .A3(n4298), .ZN(n4354) );
  NAND2_X2 U5012 ( .A1(n6147), .A2(n8493), .ZN(n8766) );
  OAI21_X2 U5013 ( .B1(n7808), .B2(n8460), .A(n8458), .ZN(n7962) );
  OAI21_X2 U5014 ( .B1(n7749), .B2(n6140), .A(n6139), .ZN(n7808) );
  XNOR2_X1 U5015 ( .A(n8565), .B(n8377), .ZN(n8328) );
  NAND2_X2 U5016 ( .A1(n4302), .A2(n5716), .ZN(n8565) );
  INV_X1 U5017 ( .A(n9820), .ZN(n4304) );
  OAI21_X2 U5018 ( .B1(n8803), .B2(n6146), .A(n8497), .ZN(n8791) );
  OAI21_X2 U5019 ( .B1(n8813), .B2(n4657), .A(n8488), .ZN(n8803) );
  NAND2_X2 U5020 ( .A1(n9033), .A2(n5688), .ZN(n4315) );
  NAND2_X1 U5021 ( .A1(n4866), .A2(n4867), .ZN(n4305) );
  AND3_X1 U5022 ( .A1(n4340), .A2(n4767), .A3(n4529), .ZN(n4527) );
  NOR2_X2 U5023 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5719) );
  INV_X4 U5024 ( .A(n9088), .ZN(n6355) );
  NAND2_X1 U5025 ( .A1(n6090), .A2(n6659), .ZN(n4309) );
  NAND2_X2 U5026 ( .A1(n6090), .A2(n6659), .ZN(n4310) );
  NAND2_X1 U5027 ( .A1(n6624), .A2(n6189), .ZN(n4311) );
  NAND2_X1 U5028 ( .A1(n6624), .A2(n6189), .ZN(n4312) );
  OAI211_X2 U5029 ( .C1(n6246), .C2(n4601), .A(n4600), .B(n4599), .ZN(n7856)
         );
  OAI22_X2 U5030 ( .A1(n7032), .A2(n7031), .B1(n6210), .B2(n6209), .ZN(n7364)
         );
  INV_X1 U5031 ( .A(n6800), .ZN(n5704) );
  NAND2_X4 U5032 ( .A1(n6799), .A2(n6798), .ZN(n6803) );
  OAI21_X2 U5033 ( .B1(n7193), .B2(n7188), .A(n8420), .ZN(n7344) );
  OAI21_X2 U5034 ( .B1(n8749), .B2(n8361), .A(n8327), .ZN(n8739) );
  OR2_X1 U5035 ( .A1(n5750), .A2(n7005), .ZN(n8396) );
  NAND2_X1 U5037 ( .A1(n4309), .A2(n6572), .ZN(n4314) );
  OAI21_X1 U5038 ( .B1(n4491), .B2(n4489), .A(n4379), .ZN(n4488) );
  INV_X1 U5039 ( .A(n6492), .ZN(n4489) );
  INV_X1 U5040 ( .A(n9261), .ZN(n7721) );
  INV_X1 U5041 ( .A(SI_15_), .ZN(n5178) );
  INV_X1 U5042 ( .A(n5043), .ZN(n4720) );
  NAND2_X1 U5043 ( .A1(n5006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U5044 ( .A1(n4424), .A2(n4422), .ZN(n5213) );
  NAND2_X1 U5045 ( .A1(n4426), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U5046 ( .A1(n5030), .A2(n4374), .ZN(n4424) );
  INV_X1 U5047 ( .A(n5078), .ZN(n4423) );
  OR2_X1 U5048 ( .A1(n8474), .A2(n8522), .ZN(n4560) );
  NOR3_X1 U5049 ( .A1(n5311), .A2(n5262), .A3(n5261), .ZN(n5320) );
  OAI21_X1 U5050 ( .B1(n4563), .B2(n8536), .A(n4562), .ZN(n4561) );
  NAND2_X1 U5051 ( .A1(n8494), .A2(n8536), .ZN(n4562) );
  AOI21_X1 U5052 ( .B1(n8495), .B2(n4360), .A(n4564), .ZN(n4563) );
  AND2_X1 U5053 ( .A1(n8958), .A2(n8751), .ZN(n6062) );
  OAI21_X1 U5054 ( .B1(n5447), .B2(n4808), .A(n5556), .ZN(n4446) );
  NAND2_X1 U5055 ( .A1(n5455), .A2(n5454), .ZN(n5474) );
  INV_X1 U5056 ( .A(n4733), .ZN(n4732) );
  OAI21_X1 U5057 ( .B1(n4735), .B2(n5153), .A(n5157), .ZN(n4733) );
  INV_X1 U5058 ( .A(n5137), .ZN(n5141) );
  OR2_X1 U5059 ( .A1(n7687), .A2(n7794), .ZN(n8434) );
  INV_X1 U5060 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4530) );
  INV_X1 U5061 ( .A(n8389), .ZN(n4623) );
  OR2_X1 U5062 ( .A1(n8774), .A2(n8244), .ZN(n4644) );
  AND2_X1 U5063 ( .A1(n8364), .A2(n8768), .ZN(n8503) );
  OR2_X1 U5064 ( .A1(n8975), .A2(n8760), .ZN(n8502) );
  OR2_X1 U5065 ( .A1(n8923), .A2(n8238), .ZN(n8493) );
  OR2_X1 U5066 ( .A1(n9380), .A2(n6525), .ZN(n4522) );
  OR2_X1 U5067 ( .A1(n6525), .A2(n8105), .ZN(n5556) );
  OR2_X1 U5068 ( .A1(n9618), .A2(n9195), .ZN(n6511) );
  OR2_X1 U5069 ( .A1(n5463), .A2(n8103), .ZN(n5578) );
  INV_X1 U5070 ( .A(n9249), .ZN(n5509) );
  AND2_X1 U5071 ( .A1(n9190), .A2(n9260), .ZN(n6483) );
  INV_X1 U5072 ( .A(n9262), .ZN(n6477) );
  INV_X1 U5073 ( .A(n7107), .ZN(n6453) );
  AND2_X1 U5074 ( .A1(n5385), .A2(n5369), .ZN(n5383) );
  NAND2_X1 U5075 ( .A1(n5325), .A2(n5324), .ZN(n5342) );
  NAND2_X1 U5076 ( .A1(n4742), .A2(n4407), .ZN(n5325) );
  OAI21_X1 U5077 ( .B1(n5297), .B2(n5296), .A(n5272), .ZN(n5287) );
  OAI21_X1 U5078 ( .B1(n5245), .B2(n5244), .A(n5246), .ZN(n5267) );
  NAND2_X1 U5079 ( .A1(n5174), .A2(n5173), .ZN(n5177) );
  NAND2_X1 U5080 ( .A1(n5107), .A2(n5106), .ZN(n5120) );
  NAND2_X1 U5081 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5082 ( .A1(n4766), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U5083 ( .A1(n8220), .A2(n4764), .ZN(n4761) );
  NAND2_X1 U5084 ( .A1(n8201), .A2(n4764), .ZN(n4763) );
  INV_X1 U5085 ( .A(n7002), .ZN(n7000) );
  INV_X1 U5086 ( .A(n5940), .ZN(n6085) );
  OAI21_X1 U5087 ( .B1(n7208), .B2(n7207), .A(n4398), .ZN(n7210) );
  OR3_X1 U5088 ( .A1(n7879), .A2(n7981), .A3(n7803), .ZN(n6680) );
  INV_X1 U5089 ( .A(n8712), .ZN(n8696) );
  AND2_X1 U5090 ( .A1(n8533), .A2(n8742), .ZN(n6552) );
  OR2_X1 U5091 ( .A1(n5955), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U5092 ( .A1(n9884), .A2(n7681), .ZN(n4653) );
  INV_X1 U5093 ( .A(n9884), .ZN(n4652) );
  NAND2_X1 U5094 ( .A1(n6814), .A2(n6154), .ZN(n9833) );
  OR2_X1 U5095 ( .A1(n8757), .A2(n8758), .ZN(n4645) );
  INV_X1 U5096 ( .A(n9829), .ZN(n8862) );
  OR2_X1 U5097 ( .A1(n6792), .A2(n8522), .ZN(n8864) );
  OAI21_X1 U5098 ( .B1(n7476), .B2(n4628), .A(n4625), .ZN(n7964) );
  AOI21_X1 U5099 ( .B1(n4627), .B2(n4626), .A(n4402), .ZN(n4625) );
  INV_X1 U5100 ( .A(n4631), .ZN(n4626) );
  INV_X1 U5101 ( .A(n4314), .ZN(n5965) );
  INV_X1 U5102 ( .A(n6642), .ZN(n5964) );
  OR2_X1 U5103 ( .A1(n6176), .A2(n8550), .ZN(n9874) );
  NAND2_X1 U5104 ( .A1(n9129), .A2(n6364), .ZN(n4588) );
  INV_X1 U5105 ( .A(n9129), .ZN(n4589) );
  AND2_X1 U5106 ( .A1(n6531), .A2(n6398), .ZN(n6415) );
  AND2_X1 U5107 ( .A1(n6626), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6567) );
  AND2_X1 U5108 ( .A1(n4475), .A2(n4474), .ZN(n6932) );
  NAND2_X1 U5109 ( .A1(n6914), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4474) );
  OR2_X1 U5110 ( .A1(n9408), .A2(n9669), .ZN(n9409) );
  AOI21_X1 U5111 ( .B1(n4493), .B2(n4492), .A(n4377), .ZN(n4491) );
  INV_X1 U5112 ( .A(n6491), .ZN(n4492) );
  NAND2_X1 U5113 ( .A1(n7772), .A2(n4363), .ZN(n4805) );
  INV_X1 U5114 ( .A(n5589), .ZN(n4806) );
  NAND2_X1 U5115 ( .A1(n7422), .A2(n6468), .ZN(n4484) );
  NOR2_X1 U5116 ( .A1(n4500), .A2(n4401), .ZN(n4498) );
  CLKBUF_X1 U5117 ( .A(n5091), .Z(n6629) );
  INV_X1 U5118 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5119 ( .A1(n4433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U5120 ( .A1(n4715), .A2(n5416), .ZN(n5422) );
  NAND2_X1 U5121 ( .A1(n5090), .A2(n5089), .ZN(n5102) );
  INV_X1 U5122 ( .A(n5063), .ZN(n4451) );
  INV_X1 U5123 ( .A(n4719), .ZN(n4452) );
  NAND2_X1 U5124 ( .A1(n4555), .A2(n5022), .ZN(n5041) );
  INV_X1 U5125 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5126 ( .A1(n5616), .A2(n4846), .ZN(n5618) );
  NAND2_X1 U5127 ( .A1(n5613), .A2(n5612), .ZN(n5616) );
  INV_X1 U5128 ( .A(n5611), .ZN(n5612) );
  AOI21_X1 U5129 ( .B1(n4425), .B2(n5633), .A(n5632), .ZN(n5214) );
  OAI21_X1 U5130 ( .B1(n5213), .B2(n5212), .A(n5630), .ZN(n4425) );
  NAND2_X1 U5131 ( .A1(n4559), .A2(n4557), .ZN(n4556) );
  AND2_X1 U5132 ( .A1(n4558), .A2(n8484), .ZN(n4557) );
  AND2_X1 U5133 ( .A1(n8473), .A2(n8522), .ZN(n4558) );
  AOI21_X1 U5134 ( .B1(n4437), .B2(n4434), .A(n9534), .ZN(n5311) );
  AOI21_X1 U5135 ( .B1(n4435), .B2(n5614), .A(n4365), .ZN(n4434) );
  OR2_X1 U5136 ( .A1(n5220), .A2(n5614), .ZN(n4437) );
  OAI21_X1 U5137 ( .B1(n8506), .B2(n4561), .A(n8505), .ZN(n8507) );
  INV_X1 U5138 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5865) );
  AND2_X1 U5139 ( .A1(n8119), .A2(n5556), .ZN(n4442) );
  AOI21_X1 U5140 ( .B1(n8905), .B2(n8318), .A(n8358), .ZN(n8314) );
  OR2_X1 U5141 ( .A1(n8318), .A2(n8317), .ZN(n8356) );
  NAND2_X1 U5142 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5143 ( .A1(n8534), .A2(n8531), .ZN(n4571) );
  INV_X1 U5144 ( .A(n7953), .ZN(n4664) );
  INV_X1 U5145 ( .A(n6084), .ZN(n8164) );
  NAND2_X1 U5146 ( .A1(n4641), .A2(n4336), .ZN(n4640) );
  INV_X1 U5147 ( .A(n6062), .ZN(n4641) );
  NAND2_X1 U5148 ( .A1(n4639), .A2(n4336), .ZN(n4638) );
  OR2_X1 U5149 ( .A1(n8964), .A2(n8199), .ZN(n8327) );
  OR2_X1 U5150 ( .A1(n8958), .A2(n8291), .ZN(n8515) );
  AND2_X1 U5151 ( .A1(n8964), .A2(n8199), .ZN(n8361) );
  OR2_X1 U5152 ( .A1(n8991), .A2(n8796), .ZN(n8497) );
  NOR2_X1 U5153 ( .A1(n8817), .A2(n8819), .ZN(n4620) );
  OR2_X1 U5154 ( .A1(n8830), .A2(n8843), .ZN(n8496) );
  INV_X1 U5155 ( .A(n8522), .ZN(n8536) );
  OR2_X1 U5156 ( .A1(n8935), .A2(n8842), .ZN(n8484) );
  NAND2_X1 U5157 ( .A1(n5869), .A2(n5676), .ZN(n4786) );
  INV_X1 U5158 ( .A(n6302), .ZN(n4596) );
  INV_X1 U5159 ( .A(n9136), .ZN(n4593) );
  NOR2_X1 U5160 ( .A1(n5463), .A2(n4522), .ZN(n4521) );
  OR2_X1 U5161 ( .A1(n9614), .A2(n9109), .ZN(n6513) );
  NAND2_X1 U5162 ( .A1(n5595), .A2(n9553), .ZN(n4803) );
  NAND2_X1 U5163 ( .A1(n7778), .A2(n7723), .ZN(n4510) );
  NAND2_X1 U5164 ( .A1(n4323), .A2(n4376), .ZN(n4419) );
  INV_X1 U5165 ( .A(n7333), .ZN(n4421) );
  NAND2_X1 U5166 ( .A1(n7340), .A2(n7433), .ZN(n4506) );
  OR2_X1 U5167 ( .A1(n9644), .A2(n9236), .ZN(n5643) );
  AND2_X1 U5168 ( .A1(n7653), .A2(n9805), .ZN(n7527) );
  INV_X1 U5169 ( .A(n4926), .ZN(n5074) );
  OAI21_X1 U5170 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5490) );
  OR2_X1 U5171 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  INV_X1 U5172 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5173 ( .B1(n5414), .B2(n4718), .A(n5421), .ZN(n4717) );
  AOI21_X1 U5174 ( .B1(n5348), .B2(n4725), .A(n4723), .ZN(n4722) );
  NAND2_X1 U5175 ( .A1(n4724), .A2(n5385), .ZN(n4723) );
  NAND2_X1 U5176 ( .A1(n4725), .A2(n4727), .ZN(n4724) );
  NAND2_X1 U5177 ( .A1(n5273), .A2(n5284), .ZN(n4741) );
  OR2_X1 U5178 ( .A1(n5273), .A2(n5284), .ZN(n4743) );
  OAI21_X1 U5179 ( .B1(n5267), .B2(n4458), .A(n5266), .ZN(n5297) );
  INV_X1 U5180 ( .A(n5263), .ZN(n4458) );
  OAI21_X1 U5181 ( .B1(n5225), .B2(n5224), .A(n5227), .ZN(n5245) );
  INV_X1 U5182 ( .A(n5223), .ZN(n5226) );
  INV_X1 U5183 ( .A(n4731), .ZN(n4461) );
  NAND2_X1 U5184 ( .A1(n4731), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U5185 ( .A1(n4455), .A2(n4989), .ZN(n4453) );
  NAND2_X1 U5186 ( .A1(n5041), .A2(n5040), .ZN(n4721) );
  INV_X1 U5187 ( .A(n8246), .ZN(n4751) );
  OR2_X1 U5188 ( .A1(n8309), .A2(n7060), .ZN(n5692) );
  OR2_X1 U5189 ( .A1(n4315), .A2(n5685), .ZN(n5691) );
  OR2_X1 U5190 ( .A1(n4306), .A2(n5705), .ZN(n5710) );
  NAND2_X1 U5191 ( .A1(n4692), .A2(n4691), .ZN(n4690) );
  INV_X1 U5192 ( .A(n6717), .ZN(n4692) );
  NAND2_X1 U5193 ( .A1(n6717), .A2(n6727), .ZN(n6742) );
  NAND2_X1 U5194 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5195 ( .A1(n4693), .A2(n6977), .ZN(n6979) );
  INV_X1 U5196 ( .A(n4694), .ZN(n4693) );
  NAND2_X1 U5197 ( .A1(n4696), .A2(n4682), .ZN(n4695) );
  NAND2_X1 U5198 ( .A1(n6855), .A2(n6963), .ZN(n6977) );
  NAND2_X1 U5199 ( .A1(n6862), .A2(n6963), .ZN(n6971) );
  NAND2_X1 U5200 ( .A1(n4704), .A2(n4703), .ZN(n4702) );
  INV_X1 U5201 ( .A(n7072), .ZN(n4704) );
  NAND2_X1 U5202 ( .A1(n4702), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4701) );
  AOI21_X1 U5203 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7497), .A(n7485), .ZN(
        n7544) );
  NAND2_X1 U5204 ( .A1(n7488), .A2(n7489), .ZN(n7490) );
  AND2_X1 U5205 ( .A1(n7497), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4660) );
  NOR2_X1 U5206 ( .A1(n8681), .A2(n8680), .ZN(n8683) );
  AOI21_X1 U5207 ( .B1(n8686), .B2(n4672), .A(n4665), .ZN(n4671) );
  INV_X1 U5208 ( .A(n8711), .ZN(n4665) );
  NAND2_X1 U5209 ( .A1(n4618), .A2(n4318), .ZN(n4613) );
  NAND2_X1 U5210 ( .A1(n4612), .A2(n4318), .ZN(n4611) );
  INV_X1 U5211 ( .A(n4614), .ZN(n4612) );
  AOI21_X1 U5212 ( .B1(n4618), .B2(n4616), .A(n4615), .ZN(n4614) );
  INV_X1 U5213 ( .A(n5987), .ZN(n4616) );
  NAND2_X1 U5214 ( .A1(n5968), .A2(n5967), .ZN(n5979) );
  INV_X1 U5215 ( .A(n5969), .ZN(n5968) );
  INV_X1 U5216 ( .A(n5888), .ZN(n5887) );
  AND2_X1 U5217 ( .A1(n5881), .A2(n4632), .ZN(n4631) );
  AOI21_X1 U5218 ( .B1(n5882), .B2(n4631), .A(n4357), .ZN(n4630) );
  OR2_X1 U5219 ( .A1(n5856), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5875) );
  INV_X1 U5220 ( .A(n8435), .ZN(n4650) );
  OR2_X1 U5221 ( .A1(n5841), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5856) );
  OR2_X1 U5222 ( .A1(n5800), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U5223 ( .A1(n8547), .A2(n8539), .ZN(n6176) );
  NOR2_X1 U5224 ( .A1(n6050), .A2(n4643), .ZN(n4642) );
  INV_X1 U5225 ( .A(n4644), .ZN(n4643) );
  AND2_X1 U5226 ( .A1(n8515), .A2(n8516), .ZN(n8740) );
  NAND2_X1 U5227 ( .A1(n8751), .A2(n9824), .ZN(n4464) );
  AND2_X1 U5228 ( .A1(n8365), .A2(n8510), .ZN(n4647) );
  AOI21_X1 U5229 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(n8757) );
  NAND2_X1 U5230 ( .A1(n8975), .A2(n8785), .ZN(n6025) );
  NOR2_X1 U5231 ( .A1(n8975), .A2(n8785), .ZN(n6024) );
  OR2_X1 U5232 ( .A1(n8981), .A2(n8795), .ZN(n8767) );
  NAND2_X1 U5233 ( .A1(n8814), .A2(n5987), .ZN(n4619) );
  NAND2_X1 U5234 ( .A1(n6792), .A2(n8536), .ZN(n8866) );
  INV_X1 U5235 ( .A(n7964), .ZN(n5918) );
  AND2_X1 U5236 ( .A1(n8465), .A2(n8467), .ZN(n8463) );
  AND2_X1 U5237 ( .A1(n7804), .A2(n8458), .ZN(n8348) );
  INV_X1 U5238 ( .A(n8866), .ZN(n9824) );
  NAND2_X1 U5239 ( .A1(n7437), .A2(n8343), .ZN(n5864) );
  NAND2_X1 U5240 ( .A1(n6109), .A2(n6108), .ZN(n6175) );
  NAND2_X1 U5241 ( .A1(n6098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6100) );
  INV_X1 U5242 ( .A(n6080), .ZN(n6082) );
  NAND2_X1 U5243 ( .A1(n5951), .A2(n5950), .ZN(n5961) );
  AND2_X1 U5244 ( .A1(n5764), .A2(n5763), .ZN(n5778) );
  INV_X1 U5245 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6078) );
  INV_X1 U5246 ( .A(n4579), .ZN(n4578) );
  OAI21_X1 U5247 ( .B1(n9117), .B2(n4580), .A(n9184), .ZN(n4579) );
  INV_X1 U5248 ( .A(n6278), .ZN(n4580) );
  OR2_X1 U5249 ( .A1(n7321), .A2(n6234), .ZN(n6211) );
  XNOR2_X1 U5250 ( .A(n6197), .B(n6196), .ZN(n6209) );
  OAI21_X1 U5251 ( .B1(n9037), .B2(n9039), .A(n9038), .ZN(n6287) );
  OR2_X1 U5252 ( .A1(n5031), .A2(n7635), .ZN(n5057) );
  OR2_X1 U5253 ( .A1(n6277), .A2(n6276), .ZN(n6278) );
  NOR2_X1 U5254 ( .A1(n5540), .A2(n5539), .ZN(n5604) );
  OR2_X1 U5255 ( .A1(n5544), .A2(n5658), .ZN(n5607) );
  OR4_X1 U5256 ( .A1(n8094), .A2(n8101), .A3(n9403), .A4(n5537), .ZN(n5538) );
  INV_X1 U5257 ( .A(n5472), .ZN(n5466) );
  INV_X1 U5258 ( .A(n4938), .ZN(n5469) );
  AND4_X1 U5259 ( .A1(n4988), .A2(n4987), .A3(n4986), .A4(n4985), .ZN(n7575)
         );
  NAND2_X1 U5260 ( .A1(n4938), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4438) );
  OR2_X1 U5261 ( .A1(n4920), .A2(n4893), .ZN(n4439) );
  NAND2_X1 U5262 ( .A1(n9319), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U5263 ( .A1(n9318), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U5264 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  INV_X1 U5265 ( .A(n6885), .ZN(n4552) );
  NOR2_X1 U5266 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  NOR2_X1 U5267 ( .A1(n7702), .A2(n4547), .ZN(n7729) );
  AND2_X1 U5268 ( .A1(n7703), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U5269 ( .A1(n6503), .A2(n6502), .ZN(n8095) );
  OR2_X1 U5270 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  AND2_X1 U5271 ( .A1(n5407), .A2(n5427), .ZN(n9411) );
  NAND2_X1 U5272 ( .A1(n9433), .A2(n6515), .ZN(n9419) );
  NAND2_X1 U5273 ( .A1(n5372), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5406) );
  INV_X1 U5274 ( .A(n5374), .ZN(n5372) );
  AOI21_X1 U5275 ( .B1(n4792), .B2(n4794), .A(n4790), .ZN(n4789) );
  AND2_X1 U5276 ( .A1(n6513), .A2(n5359), .ZN(n9466) );
  NAND2_X1 U5277 ( .A1(n9491), .A2(n6491), .ZN(n4495) );
  NAND2_X1 U5278 ( .A1(n9511), .A2(n9510), .ZN(n4791) );
  OR2_X1 U5279 ( .A1(n5238), .A2(n5237), .ZN(n5254) );
  NOR2_X1 U5280 ( .A1(n9580), .A2(n9644), .ZN(n9555) );
  OR2_X1 U5281 ( .A1(n8070), .A2(n9585), .ZN(n9580) );
  AND2_X1 U5282 ( .A1(n5215), .A2(n5635), .ZN(n4804) );
  OR2_X1 U5283 ( .A1(n9124), .A2(n7721), .ZN(n5589) );
  NAND2_X1 U5284 ( .A1(n4484), .A2(n4481), .ZN(n7753) );
  NAND2_X1 U5285 ( .A1(n4421), .A2(n4337), .ZN(n4800) );
  XNOR2_X1 U5286 ( .A(n9270), .B(n7321), .ZN(n7303) );
  AND2_X1 U5287 ( .A1(n7125), .A2(n7103), .ZN(n7257) );
  NAND2_X1 U5288 ( .A1(n5578), .A2(n5600), .ZN(n8121) );
  AOI22_X1 U5289 ( .A1(n8095), .A2(n8094), .B1(n8105), .B2(n9393), .ZN(n8096)
         );
  INV_X1 U5290 ( .A(n9427), .ZN(n9600) );
  AND2_X1 U5291 ( .A1(n6516), .A2(n5510), .ZN(n9418) );
  OAI21_X1 U5292 ( .B1(n9435), .B2(n4370), .A(n6497), .ZN(n9398) );
  INV_X1 U5293 ( .A(n4486), .ZN(n9446) );
  NAND2_X1 U5294 ( .A1(n4493), .A2(n6492), .ZN(n4490) );
  INV_X1 U5295 ( .A(n4488), .ZN(n4487) );
  INV_X1 U5296 ( .A(n9463), .ZN(n9614) );
  NAND2_X1 U5297 ( .A1(n6481), .A2(n6480), .ZN(n7871) );
  NAND2_X1 U5298 ( .A1(n4836), .A2(n4501), .ZN(n4500) );
  AND2_X1 U5299 ( .A1(n5589), .A2(n5526), .ZN(n7773) );
  INV_X1 U5300 ( .A(n6531), .ZN(n7113) );
  AND3_X1 U5301 ( .A1(n6456), .A2(n6455), .A3(n6454), .ZN(n6532) );
  NAND2_X1 U5302 ( .A1(n6521), .A2(n6520), .ZN(n9575) );
  INV_X1 U5303 ( .A(n7110), .ZN(n7108) );
  XNOR2_X1 U5304 ( .A(n5490), .B(n5489), .ZN(n8298) );
  XNOR2_X1 U5305 ( .A(n5670), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U5306 ( .A1(n5365), .A2(n5364), .ZN(n5384) );
  NAND2_X1 U5307 ( .A1(n5663), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5665) );
  XNOR2_X1 U5308 ( .A(n5297), .B(n5296), .ZN(n7247) );
  INV_X1 U5309 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4814) );
  OR2_X1 U5310 ( .A1(n5158), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U5311 ( .A1(n4738), .A2(n4735), .ZN(n5155) );
  NAND2_X1 U5312 ( .A1(n5120), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5313 ( .A1(n4449), .A2(n4447), .ZN(n5090) );
  NAND2_X1 U5314 ( .A1(n5041), .A2(n4450), .ZN(n4449) );
  INV_X1 U5315 ( .A(n5069), .ZN(n4448) );
  NAND2_X1 U5316 ( .A1(n4549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4915) );
  INV_X1 U5317 ( .A(n4912), .ZN(n4549) );
  NAND2_X1 U5318 ( .A1(n8958), .A2(n8228), .ZN(n8207) );
  AOI21_X1 U5319 ( .B1(n8797), .B2(n6085), .A(n6001), .ZN(n8238) );
  NAND2_X1 U5320 ( .A1(n4290), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5743) );
  NAND3_X1 U5321 ( .A1(n4773), .A2(n6833), .A3(n6832), .ZN(n6996) );
  AOI21_X1 U5322 ( .B1(n4776), .B2(n4778), .A(n4359), .ZN(n4775) );
  NOR2_X1 U5323 ( .A1(n4757), .A2(n8272), .ZN(n4755) );
  NOR2_X1 U5324 ( .A1(n4758), .A2(n4372), .ZN(n4757) );
  INV_X1 U5325 ( .A(n4760), .ZN(n4758) );
  NAND2_X1 U5326 ( .A1(n4760), .A2(n4765), .ZN(n4759) );
  OR2_X1 U5327 ( .A1(n4766), .A2(n8201), .ZN(n4765) );
  NAND2_X1 U5328 ( .A1(n6066), .A2(n6065), .ZN(n8533) );
  INV_X1 U5329 ( .A(n4316), .ZN(n8547) );
  XNOR2_X1 U5330 ( .A(n6075), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8550) );
  INV_X1 U5331 ( .A(n8524), .ZN(n8742) );
  NOR2_X1 U5332 ( .A1(n6737), .A2(n4526), .ZN(n6740) );
  AND2_X1 U5333 ( .A1(n6738), .A2(n4691), .ZN(n4526) );
  NAND2_X1 U5334 ( .A1(n6740), .A2(n6739), .ZN(n6846) );
  INV_X1 U5335 ( .A(n8719), .ZN(n8664) );
  OAI21_X1 U5336 ( .B1(n8698), .B2(n8697), .A(n8724), .ZN(n4535) );
  NOR2_X1 U5337 ( .A1(n8705), .A2(n4538), .ZN(n4537) );
  NAND2_X1 U5338 ( .A1(n4335), .A2(n4417), .ZN(n4538) );
  NAND2_X1 U5339 ( .A1(n5927), .A2(n5926), .ZN(n8900) );
  OR3_X1 U5340 ( .A1(n6683), .A2(n6176), .A3(n9886), .ZN(n9821) );
  OAI21_X1 U5341 ( .B1(n6096), .B2(n8862), .A(n6095), .ZN(n6182) );
  NOR2_X1 U5342 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  NOR2_X1 U5343 ( .A1(n8291), .A2(n8864), .ZN(n6093) );
  INV_X1 U5344 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9024) );
  AOI21_X1 U5345 ( .B1(n4319), .B2(n4589), .A(n4381), .ZN(n4587) );
  XNOR2_X1 U5346 ( .A(n6209), .B(n6210), .ZN(n7032) );
  NAND2_X1 U5347 ( .A1(n5289), .A2(n5288), .ZN(n9625) );
  AND2_X1 U5348 ( .A1(n6403), .A2(n9754), .ZN(n10096) );
  NAND2_X1 U5349 ( .A1(n4945), .A2(n4944), .ZN(n9269) );
  OR2_X1 U5350 ( .A1(n4920), .A2(n4943), .ZN(n4944) );
  AND3_X1 U5351 ( .A1(n4942), .A2(n4941), .A3(n4940), .ZN(n4945) );
  INV_X1 U5352 ( .A(n4473), .ZN(n6930) );
  OR2_X1 U5353 ( .A1(n6924), .A2(n6925), .ZN(n4544) );
  NAND2_X1 U5354 ( .A1(n6893), .A2(n4540), .ZN(n6896) );
  NAND2_X1 U5355 ( .A1(n4542), .A2(n4541), .ZN(n4540) );
  NOR2_X1 U5356 ( .A1(n7382), .A2(n7381), .ZN(n7702) );
  XNOR2_X1 U5357 ( .A(n7729), .B(n7732), .ZN(n7704) );
  NAND2_X1 U5358 ( .A1(n4545), .A2(n4414), .ZN(n9339) );
  NAND2_X1 U5359 ( .A1(n7898), .A2(n4546), .ZN(n4545) );
  INV_X1 U5360 ( .A(n7899), .ZN(n4546) );
  INV_X1 U5361 ( .A(n9356), .ZN(n9354) );
  NAND2_X1 U5362 ( .A1(n4582), .A2(n4581), .ZN(n5008) );
  AOI21_X1 U5363 ( .B1(n4584), .B2(n4862), .A(n4862), .ZN(n4581) );
  NAND2_X1 U5364 ( .A1(n5498), .A2(n5497), .ZN(n9370) );
  AOI21_X1 U5365 ( .B1(n8120), .B2(n8106), .A(n9096), .ZN(n9378) );
  OR2_X1 U5366 ( .A1(n9778), .A2(n5619), .ZN(n9760) );
  AND2_X1 U5367 ( .A1(n9372), .A2(n9367), .ZN(n9591) );
  AND2_X1 U5368 ( .A1(n4797), .A2(n4795), .ZN(n8140) );
  NOR2_X1 U5369 ( .A1(n8136), .A2(n4796), .ZN(n4795) );
  INV_X1 U5370 ( .A(n8125), .ZN(n4796) );
  NAND2_X1 U5371 ( .A1(n5425), .A2(n5424), .ZN(n6525) );
  NAND2_X1 U5372 ( .A1(n5404), .A2(n5403), .ZN(n9669) );
  NAND2_X1 U5373 ( .A1(n5251), .A2(n5250), .ZN(n9697) );
  NAND2_X1 U5374 ( .A1(n9713), .A2(n9801), .ZN(n9711) );
  INV_X1 U5375 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5376 ( .A1(n4815), .A2(n4816), .ZN(n5051) );
  INV_X1 U5377 ( .A(n5077), .ZN(n4426) );
  NAND2_X1 U5378 ( .A1(n8768), .A2(n8492), .ZN(n4564) );
  INV_X1 U5379 ( .A(n7091), .ZN(n5519) );
  INV_X1 U5380 ( .A(n4642), .ZN(n4639) );
  INV_X1 U5381 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5680) );
  INV_X1 U5382 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4768) );
  AND2_X1 U5383 ( .A1(n9484), .A2(n4511), .ZN(n9422) );
  NOR2_X1 U5384 ( .A1(n9678), .A2(n4513), .ZN(n4511) );
  INV_X1 U5385 ( .A(n4726), .ZN(n4725) );
  OAI21_X1 U5386 ( .B1(n5347), .B2(n4727), .A(n5383), .ZN(n4726) );
  INV_X1 U5387 ( .A(n5364), .ZN(n4727) );
  INV_X1 U5388 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5002) );
  INV_X1 U5389 ( .A(SI_19_), .ZN(n5268) );
  INV_X1 U5390 ( .A(n5193), .ZN(n5179) );
  AND2_X1 U5391 ( .A1(n4739), .A2(n5154), .ZN(n4731) );
  INV_X1 U5392 ( .A(n5106), .ZN(n4460) );
  INV_X1 U5393 ( .A(n4834), .ZN(n4764) );
  INV_X1 U5394 ( .A(n4747), .ZN(n4746) );
  OAI21_X1 U5395 ( .B1(n4750), .B2(n8247), .A(n8197), .ZN(n4747) );
  AND2_X1 U5396 ( .A1(n8537), .A2(n8302), .ZN(n8525) );
  NAND2_X1 U5397 ( .A1(n4690), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U5398 ( .A1(n4695), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4694) );
  NOR2_X1 U5399 ( .A1(n8685), .A2(n8686), .ZN(n8688) );
  INV_X1 U5400 ( .A(n8687), .ZN(n4672) );
  AND2_X1 U5401 ( .A1(n8691), .A2(n4532), .ZN(n8695) );
  NAND2_X1 U5402 ( .A1(n8693), .A2(n8692), .ZN(n4532) );
  NAND2_X1 U5403 ( .A1(n4730), .A2(n4728), .ZN(n8355) );
  AND2_X1 U5404 ( .A1(n4729), .A2(n6542), .ZN(n4728) );
  INV_X1 U5405 ( .A(n8225), .ZN(n4729) );
  NAND2_X1 U5406 ( .A1(n5752), .A2(n4646), .ZN(n7160) );
  AND2_X1 U5407 ( .A1(n4348), .A2(n5751), .ZN(n4646) );
  NAND2_X1 U5408 ( .A1(n9030), .A2(n8303), .ZN(n4730) );
  OR2_X1 U5409 ( .A1(n8533), .A2(n8524), .ZN(n6540) );
  OR2_X1 U5410 ( .A1(n8839), .A2(n5986), .ZN(n8817) );
  INV_X1 U5411 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U5412 ( .A1(n4445), .A2(n5449), .ZN(n4444) );
  OR2_X1 U5413 ( .A1(n5440), .A2(n5439), .ZN(n5458) );
  INV_X1 U5414 ( .A(n9418), .ZN(n4809) );
  OR2_X1 U5415 ( .A1(n9678), .A2(n5378), .ZN(n6515) );
  INV_X1 U5416 ( .A(n6510), .ZN(n4790) );
  INV_X1 U5417 ( .A(n4793), .ZN(n4792) );
  OAI21_X1 U5418 ( .B1(n9510), .B2(n4794), .A(n9475), .ZN(n4793) );
  INV_X1 U5419 ( .A(n5652), .ZN(n4794) );
  NOR2_X1 U5420 ( .A1(n9614), .A2(n9618), .ZN(n4515) );
  NOR2_X1 U5421 ( .A1(n9697), .A2(n9639), .ZN(n4518) );
  NAND2_X1 U5422 ( .A1(n9271), .A2(n10097), .ZN(n5627) );
  INV_X1 U5423 ( .A(n9251), .ZN(n6494) );
  XNOR2_X1 U5424 ( .A(n5474), .B(n5473), .ZN(n5477) );
  NAND2_X1 U5425 ( .A1(n4714), .A2(n4712), .ZN(n5451) );
  AOI21_X1 U5426 ( .B1(n4716), .B2(n4718), .A(n4713), .ZN(n4712) );
  INV_X1 U5427 ( .A(n5435), .ZN(n4713) );
  INV_X1 U5428 ( .A(n5416), .ZN(n4718) );
  AND2_X1 U5429 ( .A1(n5416), .A2(n5402), .ZN(n5414) );
  AND2_X1 U5430 ( .A1(n5397), .A2(n5389), .ZN(n5395) );
  INV_X1 U5431 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U5432 ( .A1(n5000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5433 ( .A1(n5003), .A2(n5002), .ZN(n5663) );
  INV_X1 U5434 ( .A(SI_20_), .ZN(n5284) );
  INV_X1 U5435 ( .A(n4736), .ZN(n4735) );
  OAI21_X1 U5436 ( .B1(n5141), .B2(n4737), .A(n5140), .ZN(n4736) );
  NAND2_X1 U5437 ( .A1(n5119), .A2(n5118), .ZN(n4737) );
  NOR2_X1 U5438 ( .A1(n5141), .A2(n4740), .ZN(n4739) );
  INV_X1 U5439 ( .A(n5118), .ZN(n4740) );
  XNOR2_X1 U5440 ( .A(n4970), .B(SI_4_), .ZN(n4967) );
  OAI21_X1 U5441 ( .B1(n4907), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n4565), .ZN(
        n4929) );
  NAND2_X1 U5442 ( .A1(n4907), .A2(n4566), .ZN(n4565) );
  NAND2_X1 U5443 ( .A1(n4898), .A2(n4885), .ZN(n4908) );
  AND2_X1 U5444 ( .A1(n8076), .A2(n4777), .ZN(n4776) );
  OR2_X1 U5445 ( .A1(n8002), .A2(n4778), .ZN(n4777) );
  INV_X1 U5446 ( .A(n8051), .ZN(n4778) );
  INV_X1 U5447 ( .A(n8220), .ZN(n4766) );
  INV_X1 U5448 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10034) );
  OAI21_X1 U5449 ( .B1(n8256), .B2(n8255), .A(n8254), .ZN(n8253) );
  INV_X1 U5450 ( .A(n6017), .ZN(n6016) );
  NAND2_X1 U5451 ( .A1(n8003), .A2(n8002), .ZN(n8052) );
  OR2_X1 U5452 ( .A1(n6675), .A2(n6159), .ZN(n6694) );
  INV_X1 U5453 ( .A(n8879), .ZN(n8036) );
  NOR2_X1 U5454 ( .A1(n8530), .A2(n4569), .ZN(n4568) );
  NOR2_X1 U5455 ( .A1(n8535), .A2(n8534), .ZN(n4569) );
  INV_X1 U5456 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5679) );
  AND2_X1 U5457 ( .A1(n8313), .A2(n8312), .ZN(n8555) );
  AND2_X1 U5458 ( .A1(n6038), .A2(n6037), .ZN(n8193) );
  OR2_X1 U5459 ( .A1(n6652), .A2(n7060), .ZN(n6714) );
  NAND2_X1 U5460 ( .A1(n8575), .A2(n6726), .ZN(n4676) );
  NAND2_X1 U5461 ( .A1(n4688), .A2(n6742), .ZN(n6746) );
  INV_X1 U5462 ( .A(n4689), .ZN(n4688) );
  AND2_X1 U5463 ( .A1(n4701), .A2(n4705), .ZN(n7213) );
  NOR2_X1 U5464 ( .A1(n7213), .A2(n7212), .ZN(n7485) );
  NAND2_X1 U5465 ( .A1(n7210), .A2(n7209), .ZN(n7488) );
  OAI21_X1 U5466 ( .B1(n7486), .B2(n4698), .A(n4697), .ZN(n7607) );
  NAND2_X1 U5467 ( .A1(n4699), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U5468 ( .A1(n7547), .A2(n4699), .ZN(n4697) );
  INV_X1 U5469 ( .A(n7608), .ZN(n4699) );
  NOR2_X1 U5470 ( .A1(n5858), .A2(n7550), .ZN(n7818) );
  INV_X1 U5471 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U5472 ( .A1(n7955), .A2(n4664), .ZN(n4663) );
  NOR2_X1 U5473 ( .A1(n7955), .A2(n4664), .ZN(n4662) );
  AND2_X1 U5474 ( .A1(n7941), .A2(n7940), .ZN(n8584) );
  OAI21_X1 U5475 ( .B1(n8623), .B2(n4686), .A(n4685), .ZN(n8669) );
  NAND2_X1 U5476 ( .A1(n4687), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U5477 ( .A1(n8647), .A2(n4687), .ZN(n4685) );
  INV_X1 U5478 ( .A(n8650), .ZN(n4687) );
  NOR2_X1 U5479 ( .A1(n8623), .A2(n8624), .ZN(n8648) );
  NOR2_X1 U5480 ( .A1(n5868), .A2(n4784), .ZN(n5924) );
  NAND2_X1 U5481 ( .A1(n4785), .A2(n5920), .ZN(n4784) );
  INV_X1 U5482 ( .A(n4786), .ZN(n4785) );
  INV_X1 U5483 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U5484 ( .A1(n5924), .A2(n5923), .ZN(n5936) );
  NAND2_X1 U5485 ( .A1(n8695), .A2(n8694), .ZN(n8712) );
  OR2_X1 U5486 ( .A1(n5997), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6004) );
  OR2_X1 U5487 ( .A1(n6004), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U5488 ( .A1(n5990), .A2(n10034), .ZN(n5997) );
  INV_X1 U5489 ( .A(n5991), .ZN(n5990) );
  OR2_X1 U5490 ( .A1(n5979), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5991) );
  AND2_X1 U5491 ( .A1(n8484), .A2(n8475), .ZN(n8860) );
  OR2_X1 U5492 ( .A1(n8859), .A2(n8860), .ZN(n8857) );
  NAND2_X1 U5493 ( .A1(n5942), .A2(n5941), .ZN(n5955) );
  INV_X1 U5494 ( .A(n5943), .ZN(n5942) );
  NAND2_X1 U5495 ( .A1(n5910), .A2(n5909), .ZN(n5928) );
  INV_X1 U5496 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5909) );
  INV_X1 U5497 ( .A(n5911), .ZN(n5910) );
  OR2_X1 U5498 ( .A1(n5928), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5943) );
  OR2_X1 U5499 ( .A1(n5899), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5911) );
  INV_X1 U5500 ( .A(n5875), .ZN(n5874) );
  CLKBUF_X1 U5501 ( .A(n7442), .Z(n7443) );
  NAND2_X1 U5502 ( .A1(n5830), .A2(n5829), .ZN(n5841) );
  INV_X1 U5503 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5829) );
  INV_X1 U5504 ( .A(n5831), .ZN(n5830) );
  NAND2_X1 U5505 ( .A1(n7160), .A2(n5816), .ZN(n7190) );
  INV_X1 U5506 ( .A(n5787), .ZN(n5786) );
  NAND2_X1 U5507 ( .A1(n8395), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5508 ( .A1(n6136), .A2(n8395), .ZN(n4624) );
  NAND2_X1 U5509 ( .A1(n5725), .A2(n5724), .ZN(n4606) );
  INV_X1 U5510 ( .A(n8328), .ZN(n9827) );
  AND2_X1 U5511 ( .A1(n6161), .A2(n8522), .ZN(n6178) );
  NAND2_X1 U5512 ( .A1(n4730), .A2(n6542), .ZN(n6543) );
  INV_X1 U5513 ( .A(n4634), .ZN(n6554) );
  OAI21_X1 U5514 ( .B1(n8757), .B2(n4387), .A(n4635), .ZN(n4634) );
  INV_X1 U5515 ( .A(n4637), .ZN(n4635) );
  NAND2_X1 U5516 ( .A1(n4645), .A2(n4644), .ZN(n4466) );
  OR2_X1 U5517 ( .A1(n8360), .A2(n8361), .ZN(n8750) );
  NAND2_X1 U5518 ( .A1(n6028), .A2(n6027), .ZN(n8244) );
  AND2_X1 U5519 ( .A1(n6149), .A2(n8502), .ZN(n8365) );
  AND2_X1 U5520 ( .A1(n8502), .A2(n8364), .ZN(n8771) );
  AOI21_X1 U5521 ( .B1(n4608), .B2(n4613), .A(n4384), .ZN(n4467) );
  INV_X1 U5522 ( .A(n8496), .ZN(n4657) );
  AND2_X1 U5523 ( .A1(n4619), .A2(n4617), .ZN(n8822) );
  INV_X1 U5524 ( .A(n4620), .ZN(n4617) );
  INV_X1 U5525 ( .A(n8860), .ZN(n8853) );
  OR2_X1 U5526 ( .A1(n8900), .A2(n8036), .ZN(n8469) );
  INV_X1 U5527 ( .A(n8418), .ZN(n9864) );
  OR2_X1 U5528 ( .A1(n6682), .A2(n6683), .ZN(n6695) );
  INV_X1 U5529 ( .A(n6694), .ZN(n6690) );
  XNOR2_X1 U5530 ( .A(n6105), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U5531 ( .A(n6083), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8370) );
  NOR2_X1 U5532 ( .A1(n5868), .A2(n4786), .ZN(n5921) );
  INV_X1 U5533 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U5534 ( .A1(n9092), .A2(n6943), .ZN(n6199) );
  OR2_X1 U5535 ( .A1(n6268), .A2(n9206), .ZN(n6271) );
  OAI22_X1 U5536 ( .A1(n6234), .A2(n10097), .B1(n7305), .B2(n6214), .ZN(n6217)
         );
  OAI21_X1 U5537 ( .B1(n4320), .B2(n4364), .A(n4317), .ZN(n4599) );
  NAND2_X1 U5538 ( .A1(n4602), .A2(n4317), .ZN(n4601) );
  NAND2_X1 U5539 ( .A1(n4603), .A2(n4366), .ZN(n4600) );
  AOI21_X1 U5540 ( .B1(n6943), .B2(n6205), .A(n6204), .ZN(n6206) );
  NOR2_X1 U5541 ( .A1(n6624), .A2(n6203), .ZN(n6204) );
  NAND2_X1 U5542 ( .A1(n6940), .A2(n6941), .ZN(n6939) );
  INV_X1 U5543 ( .A(n6266), .ZN(n9205) );
  AND2_X1 U5544 ( .A1(n4592), .A2(n6310), .ZN(n4591) );
  NAND2_X1 U5545 ( .A1(n4594), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U5546 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  XNOR2_X1 U5547 ( .A(n6293), .B(n6291), .ZN(n9232) );
  NAND2_X1 U5548 ( .A1(n9232), .A2(n9233), .ZN(n9231) );
  OAI21_X1 U5549 ( .B1(n5657), .B2(n5620), .A(n7582), .ZN(n5611) );
  AND2_X1 U5550 ( .A1(n6508), .A2(n5545), .ZN(n6627) );
  OAI211_X1 U5551 ( .C1(n5579), .C2(n4833), .A(n8119), .B(n5578), .ZN(n5580)
         );
  AND2_X1 U5552 ( .A1(n5433), .A2(n5432), .ZN(n8105) );
  INV_X1 U5553 ( .A(n4979), .ZN(n5465) );
  AND4_X1 U5554 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n9109)
         );
  AND4_X1 U5555 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n9195)
         );
  AND4_X1 U5556 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n9223)
         );
  AND4_X1 U5557 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n9137)
         );
  AND4_X1 U5558 ( .A1(n5062), .A2(n5061), .A3(n5060), .A4(n5059), .ZN(n7518)
         );
  AND4_X1 U5559 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n7651)
         );
  OR2_X1 U5560 ( .A1(n4979), .A2(n7337), .ZN(n4940) );
  OR2_X1 U5561 ( .A1(n6910), .A2(n6909), .ZN(n4475) );
  OR2_X1 U5562 ( .A1(n6932), .A2(n6931), .ZN(n4473) );
  AND2_X1 U5563 ( .A1(n4544), .A2(n4543), .ZN(n6772) );
  NAND2_X1 U5564 ( .A1(n6935), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4543) );
  NAND2_X1 U5565 ( .A1(n6772), .A2(n6773), .ZN(n6893) );
  NOR2_X1 U5566 ( .A1(n7012), .A2(n4477), .ZN(n7013) );
  NOR2_X1 U5567 ( .A1(n4478), .A2(n7724), .ZN(n4477) );
  INV_X1 U5568 ( .A(n7017), .ZN(n4478) );
  NOR2_X1 U5569 ( .A1(n7016), .A2(n4396), .ZN(n7020) );
  NAND2_X1 U5570 ( .A1(n7013), .A2(n7014), .ZN(n7232) );
  NAND2_X1 U5571 ( .A1(n7020), .A2(n7019), .ZN(n7236) );
  NOR2_X1 U5572 ( .A1(n7698), .A2(n4480), .ZN(n7733) );
  AND2_X1 U5573 ( .A1(n7703), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U5574 ( .A1(n7701), .A2(n9583), .ZN(n7734) );
  AND2_X1 U5575 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  INV_X1 U5576 ( .A(n4585), .ZN(n4584) );
  OAI21_X1 U5577 ( .B1(n5232), .B2(n4862), .A(n5247), .ZN(n4585) );
  NAND2_X1 U5578 ( .A1(n4521), .A2(n9373), .ZN(n4520) );
  OR2_X1 U5579 ( .A1(n9380), .A2(n9090), .ZN(n8119) );
  NOR2_X1 U5580 ( .A1(n9409), .A2(n4519), .ZN(n8155) );
  INV_X1 U5581 ( .A(n4521), .ZN(n4519) );
  OR2_X1 U5582 ( .A1(n9409), .A2(n4522), .ZN(n8126) );
  OAI21_X1 U5583 ( .B1(n9419), .B2(n4810), .A(n4807), .ZN(n6518) );
  INV_X1 U5584 ( .A(n4811), .ZN(n4810) );
  AOI21_X1 U5585 ( .B1(n4811), .B2(n4809), .A(n4808), .ZN(n4807) );
  NOR2_X1 U5586 ( .A1(n9403), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5587 ( .A1(n6518), .A2(n6519), .ZN(n8100) );
  OR2_X1 U5588 ( .A1(n9431), .A2(n9430), .ZN(n9433) );
  OR2_X1 U5589 ( .A1(n5353), .A2(n5352), .ZN(n5374) );
  NAND2_X1 U5590 ( .A1(n9484), .A2(n4515), .ZN(n9460) );
  NAND2_X1 U5591 ( .A1(n9484), .A2(n9486), .ZN(n9485) );
  OR2_X1 U5592 ( .A1(n5303), .A2(n9178), .ZN(n5291) );
  OR2_X1 U5593 ( .A1(n5291), .A2(n5278), .ZN(n5334) );
  OR2_X1 U5594 ( .A1(n9625), .A2(n6317), .ZN(n9475) );
  OR2_X1 U5595 ( .A1(n5301), .A2(n5300), .ZN(n5303) );
  AND2_X1 U5596 ( .A1(n5596), .A2(n4803), .ZN(n4802) );
  AND2_X1 U5597 ( .A1(n9555), .A2(n4516), .ZN(n9504) );
  NOR2_X1 U5598 ( .A1(n4517), .A2(n9630), .ZN(n4516) );
  INV_X1 U5599 ( .A(n4518), .ZN(n4517) );
  NAND2_X1 U5600 ( .A1(n9555), .A2(n4518), .ZN(n9528) );
  AOI21_X1 U5601 ( .B1(n7247), .B2(n5495), .A(n5299), .ZN(n9505) );
  NAND2_X1 U5602 ( .A1(n5252), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5301) );
  INV_X1 U5603 ( .A(n5254), .ZN(n5252) );
  NAND2_X1 U5604 ( .A1(n9543), .A2(n5595), .ZN(n9542) );
  NAND2_X1 U5605 ( .A1(n5188), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U5606 ( .A1(n5593), .A2(n5592), .ZN(n9562) );
  NOR2_X1 U5607 ( .A1(n4510), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5608 ( .A1(n9718), .A2(n8049), .ZN(n4508) );
  INV_X1 U5609 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5163) );
  OR2_X1 U5610 ( .A1(n5164), .A2(n5163), .ZN(n5203) );
  NOR3_X1 U5611 ( .A1(n7526), .A2(n4510), .A3(n9190), .ZN(n8071) );
  NAND2_X1 U5612 ( .A1(n5127), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5147) );
  INV_X1 U5613 ( .A(n5129), .ZN(n5127) );
  INV_X1 U5614 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9993) );
  OR2_X1 U5615 ( .A1(n5095), .A2(n9993), .ZN(n5129) );
  OR2_X1 U5616 ( .A1(n5057), .A2(n5056), .ZN(n5082) );
  NAND2_X1 U5617 ( .A1(n7453), .A2(n5581), .ZN(n7515) );
  NOR2_X1 U5618 ( .A1(n7762), .A2(n7639), .ZN(n7653) );
  NAND2_X1 U5619 ( .A1(n4420), .A2(n6466), .ZN(n7754) );
  NAND2_X1 U5620 ( .A1(n4388), .A2(n4418), .ZN(n4420) );
  NAND2_X1 U5621 ( .A1(n4418), .A2(n4419), .ZN(n7453) );
  INV_X1 U5622 ( .A(n4506), .ZN(n4505) );
  NOR2_X1 U5623 ( .A1(n7338), .A2(n7458), .ZN(n4504) );
  OR2_X1 U5624 ( .A1(n7302), .A2(n7369), .ZN(n7338) );
  NOR2_X1 U5625 ( .A1(n7338), .A2(n9787), .ZN(n7428) );
  NAND2_X1 U5626 ( .A1(n4503), .A2(n7334), .ZN(n7328) );
  INV_X1 U5627 ( .A(n7326), .ZN(n4503) );
  XNOR2_X1 U5628 ( .A(n9269), .B(n7340), .ZN(n7334) );
  NAND2_X1 U5629 ( .A1(n5518), .A2(n5627), .ZN(n7251) );
  INV_X1 U5630 ( .A(n4787), .ZN(n7094) );
  NAND2_X1 U5631 ( .A1(n5483), .A2(n5482), .ZN(n5540) );
  AND2_X1 U5632 ( .A1(n5647), .A2(n5652), .ZN(n9510) );
  OAI21_X1 U5633 ( .B1(n7871), .B2(n6483), .A(n4827), .ZN(n8064) );
  AOI22_X1 U5634 ( .A1(n7713), .A2(n6478), .B1(n7723), .B2(n6477), .ZN(n7771)
         );
  OR2_X1 U5635 ( .A1(n7117), .A2(n6399), .ZN(n9804) );
  NAND2_X1 U5636 ( .A1(n7582), .A2(n7419), .ZN(n7117) );
  NAND2_X1 U5637 ( .A1(n6381), .A2(n6383), .ZN(n7107) );
  XNOR2_X1 U5638 ( .A(n5477), .B(SI_29_), .ZN(n9030) );
  XNOR2_X1 U5639 ( .A(n5451), .B(n5450), .ZN(n8088) );
  AND2_X1 U5640 ( .A1(n4325), .A2(n4350), .ZN(n4523) );
  NAND2_X1 U5641 ( .A1(n4352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U5642 ( .B1(n5342), .B2(n5341), .A(n5340), .ZN(n5348) );
  NAND2_X1 U5643 ( .A1(n4742), .A2(n4741), .ZN(n5321) );
  INV_X1 U5644 ( .A(n5006), .ZN(n5005) );
  OR2_X1 U5645 ( .A1(n5143), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U5646 ( .A1(n4734), .A2(n5118), .ZN(n5142) );
  INV_X1 U5647 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4817) );
  NAND2_X1 U5648 ( .A1(n4721), .A2(n4719), .ZN(n5064) );
  INV_X1 U5649 ( .A(n4971), .ZN(n4456) );
  NOR2_X1 U5650 ( .A1(n4952), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U5651 ( .A1(n4972), .A2(n4971), .ZN(n4991) );
  NAND2_X1 U5652 ( .A1(n6833), .A2(n6832), .ZN(n6836) );
  NOR2_X1 U5653 ( .A1(n8255), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U5654 ( .A1(n6996), .A2(n6995), .ZN(n7003) );
  NAND2_X1 U5655 ( .A1(n7390), .A2(n7409), .ZN(n4780) );
  NAND2_X1 U5656 ( .A1(n4782), .A2(n7409), .ZN(n4779) );
  AND3_X1 U5657 ( .A1(n5976), .A2(n5975), .A3(n5974), .ZN(n8865) );
  NAND2_X1 U5658 ( .A1(n8235), .A2(n8182), .ZN(n8274) );
  INV_X1 U5659 ( .A(n8290), .ZN(n8266) );
  NAND2_X1 U5660 ( .A1(n8052), .A2(n8051), .ZN(n8077) );
  NAND2_X1 U5661 ( .A1(n7271), .A2(n7270), .ZN(n7274) );
  INV_X1 U5662 ( .A(n8223), .ZN(n8293) );
  OR2_X1 U5663 ( .A1(n5696), .A2(n6078), .ZN(n4539) );
  NAND2_X1 U5664 ( .A1(n6061), .A2(n6060), .ZN(n8751) );
  INV_X1 U5665 ( .A(n8193), .ZN(n8774) );
  INV_X1 U5666 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6619) );
  AND4_X1 U5667 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n7794)
         );
  AND4_X1 U5668 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n8426)
         );
  AND4_X1 U5669 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n7292)
         );
  OR2_X1 U5670 ( .A1(n6646), .A2(n6645), .ZN(n6723) );
  NAND2_X1 U5671 ( .A1(n4673), .A2(n4675), .ZN(n6729) );
  NAND2_X1 U5672 ( .A1(n4690), .A2(n6742), .ZN(n6719) );
  NAND2_X1 U5673 ( .A1(n4679), .A2(n6971), .ZN(n6973) );
  INV_X1 U5674 ( .A(n4680), .ZN(n4679) );
  NAND2_X1 U5675 ( .A1(n4681), .A2(n6971), .ZN(n6863) );
  NAND2_X1 U5676 ( .A1(n6846), .A2(n4525), .ZN(n6852) );
  OR2_X1 U5677 ( .A1(n6847), .A2(n6848), .ZN(n4525) );
  NAND2_X1 U5678 ( .A1(n6852), .A2(n6851), .ZN(n6964) );
  NAND2_X1 U5679 ( .A1(n4695), .A2(n6977), .ZN(n6857) );
  NAND2_X1 U5680 ( .A1(n4702), .A2(n4705), .ZN(n7073) );
  INV_X1 U5681 ( .A(n4701), .ZN(n4700) );
  NOR2_X1 U5682 ( .A1(n7067), .A2(n4524), .ZN(n7208) );
  AND2_X1 U5683 ( .A1(n7068), .A2(n7069), .ZN(n4524) );
  XNOR2_X1 U5684 ( .A(n7544), .B(n7545), .ZN(n7486) );
  NOR2_X1 U5685 ( .A1(n7486), .A2(n5833), .ZN(n7546) );
  OR2_X1 U5686 ( .A1(n7823), .A2(n7822), .ZN(n7941) );
  XNOR2_X1 U5687 ( .A(n8584), .B(n8598), .ZN(n7942) );
  NOR2_X1 U5688 ( .A1(n7942), .A2(n7750), .ZN(n8585) );
  OAI21_X1 U5689 ( .B1(n7942), .B2(n4710), .A(n4709), .ZN(n8610) );
  NAND2_X1 U5690 ( .A1(n4711), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5691 ( .A1(n8586), .A2(n4711), .ZN(n4709) );
  INV_X1 U5692 ( .A(n8588), .ZN(n4711) );
  NOR2_X1 U5693 ( .A1(n8611), .A2(n7971), .ZN(n8631) );
  NAND2_X1 U5694 ( .A1(n4708), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5695 ( .A1(n8632), .A2(n4708), .ZN(n4706) );
  INV_X1 U5696 ( .A(n8634), .ZN(n4708) );
  NAND2_X1 U5697 ( .A1(n8685), .A2(n4413), .ZN(n4667) );
  OAI21_X1 U5698 ( .B1(n4671), .B2(n4410), .A(n4666), .ZN(n4670) );
  AND2_X1 U5699 ( .A1(n6648), .A2(n6091), .ZN(n8727) );
  INV_X1 U5700 ( .A(n8167), .ZN(n4658) );
  NAND2_X1 U5701 ( .A1(n4610), .A2(n4611), .ZN(n8793) );
  OR2_X1 U5702 ( .A1(n8814), .A2(n4613), .ZN(n4610) );
  NAND2_X1 U5703 ( .A1(n5996), .A2(n5995), .ZN(n8923) );
  NAND2_X1 U5704 ( .A1(n5954), .A2(n5953), .ZN(n8935) );
  NAND2_X1 U5705 ( .A1(n4629), .A2(n4630), .ZN(n7805) );
  NAND2_X1 U5706 ( .A1(n7476), .A2(n4631), .ZN(n4629) );
  AND2_X1 U5707 ( .A1(n4651), .A2(n8407), .ZN(n7354) );
  INV_X1 U5708 ( .A(n7398), .ZN(n9870) );
  INV_X1 U5709 ( .A(n9839), .ZN(n8894) );
  NAND2_X1 U5710 ( .A1(n7150), .A2(n8389), .ZN(n7171) );
  OR2_X1 U5711 ( .A1(n6168), .A2(n9823), .ZN(n8738) );
  INV_X1 U5712 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7184) );
  INV_X1 U5713 ( .A(n8903), .ZN(n7811) );
  OR2_X1 U5714 ( .A1(n5827), .A2(n6580), .ZN(n5701) );
  INV_X1 U5715 ( .A(n9821), .ZN(n8898) );
  INV_X1 U5716 ( .A(n8738), .ZN(n8899) );
  INV_X1 U5717 ( .A(n8319), .ZN(n8905) );
  NAND2_X1 U5718 ( .A1(n6182), .A2(n9915), .ZN(n6184) );
  NAND2_X1 U5719 ( .A1(n8298), .A2(n8303), .ZN(n8301) );
  NAND2_X1 U5720 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NAND2_X1 U5721 ( .A1(n6052), .A2(n6051), .ZN(n8958) );
  NAND2_X1 U5722 ( .A1(n4636), .A2(n4336), .ZN(n8741) );
  NAND2_X1 U5723 ( .A1(n4645), .A2(n4642), .ZN(n4636) );
  NAND2_X1 U5724 ( .A1(n6040), .A2(n6039), .ZN(n8964) );
  AOI21_X1 U5725 ( .B1(n4465), .B2(n9829), .A(n4462), .ZN(n8962) );
  NAND2_X1 U5726 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  XNOR2_X1 U5727 ( .A(n4466), .B(n8750), .ZN(n4465) );
  NAND2_X1 U5728 ( .A1(n8774), .A2(n9826), .ZN(n4463) );
  NAND2_X1 U5729 ( .A1(n6014), .A2(n6013), .ZN(n8975) );
  NAND2_X1 U5730 ( .A1(n6003), .A2(n6002), .ZN(n8981) );
  NAND2_X1 U5731 ( .A1(n4619), .A2(n4618), .ZN(n8805) );
  NAND2_X1 U5732 ( .A1(n7247), .A2(n8303), .ZN(n4457) );
  NAND2_X1 U5733 ( .A1(n5939), .A2(n5938), .ZN(n9011) );
  AND2_X1 U5734 ( .A1(n8881), .A2(n8880), .ZN(n9009) );
  NAND2_X1 U5735 ( .A1(n5908), .A2(n5907), .ZN(n8025) );
  AND2_X1 U5736 ( .A1(n7967), .A2(n7966), .ZN(n7975) );
  NAND2_X1 U5737 ( .A1(n5898), .A2(n5897), .ZN(n7918) );
  NAND2_X1 U5738 ( .A1(n5885), .A2(n5884), .ZN(n8451) );
  INV_X1 U5739 ( .A(n9016), .ZN(n9010) );
  AND2_X1 U5740 ( .A1(n6654), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6687) );
  NAND2_X1 U5741 ( .A1(n6600), .A2(n6110), .ZN(n6611) );
  INV_X1 U5742 ( .A(n6107), .ZN(n7981) );
  INV_X1 U5743 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U5744 ( .A1(n6102), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  INV_X1 U5745 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7693) );
  INV_X1 U5746 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7586) );
  INV_X1 U5747 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U5748 ( .A1(n6081), .A2(n6082), .ZN(n8539) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7248) );
  INV_X1 U5750 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7090) );
  INV_X1 U5751 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7028) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6921) );
  INV_X1 U5753 ( .A(n8654), .ZN(n8670) );
  INV_X1 U5754 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6618) );
  INV_X1 U5755 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6608) );
  INV_X1 U5756 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6606) );
  XNOR2_X1 U5757 ( .A(n5812), .B(n4770), .ZN(n7497) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4887) );
  AND2_X1 U5759 ( .A1(n6246), .A2(n4826), .ZN(n7574) );
  AOI21_X1 U5760 ( .B1(n4578), .B2(n4580), .A(n4386), .ZN(n4575) );
  INV_X1 U5761 ( .A(n9505), .ZN(n9630) );
  NAND2_X1 U5762 ( .A1(n6434), .A2(n6433), .ZN(n9105) );
  AOI21_X1 U5763 ( .B1(n4603), .B2(n4602), .A(n4320), .ZN(n4604) );
  NAND2_X1 U5764 ( .A1(n4598), .A2(n4602), .ZN(n4605) );
  INV_X1 U5765 ( .A(n6246), .ZN(n4598) );
  NAND2_X1 U5766 ( .A1(n5187), .A2(n5186), .ZN(n9644) );
  NAND2_X1 U5767 ( .A1(n4597), .A2(n6302), .ZN(n9146) );
  INV_X1 U5768 ( .A(n10098), .ZN(n9224) );
  INV_X1 U5769 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U5770 ( .A1(n4577), .A2(n6278), .ZN(n9183) );
  NAND2_X1 U5771 ( .A1(n9116), .A2(n9117), .ZN(n4577) );
  CLKBUF_X1 U5772 ( .A(n9048), .Z(n9049) );
  AND2_X1 U5773 ( .A1(n5202), .A2(n5201), .ZN(n9648) );
  NAND2_X1 U5774 ( .A1(n6411), .A2(n6410), .ZN(n9242) );
  NAND2_X1 U5775 ( .A1(n5413), .A2(n5412), .ZN(n9249) );
  OAI211_X1 U5776 ( .C1(n4979), .C2(n9439), .A(n5377), .B(n5376), .ZN(n9250)
         );
  AND4_X1 U5777 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n9236)
         );
  NAND2_X1 U5778 ( .A1(n4938), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4925) );
  OR2_X1 U5779 ( .A1(n4920), .A2(n4921), .ZN(n4923) );
  OR2_X2 U5780 ( .A1(n6568), .A2(n6624), .ZN(n9272) );
  OAI21_X1 U5781 ( .B1(n9276), .B2(n4865), .A(n4470), .ZN(n9278) );
  NAND2_X1 U5782 ( .A1(n9276), .A2(n4865), .ZN(n4470) );
  NAND2_X1 U5783 ( .A1(n9305), .A2(n6784), .ZN(n9323) );
  NAND2_X1 U5784 ( .A1(n9323), .A2(n9324), .ZN(n9322) );
  AND2_X1 U5785 ( .A1(n9322), .A2(n4476), .ZN(n6883) );
  NAND2_X1 U5786 ( .A1(n9318), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4476) );
  INV_X1 U5787 ( .A(n4551), .ZN(n6884) );
  INV_X1 U5788 ( .A(n4553), .ZN(n6886) );
  NAND2_X1 U5789 ( .A1(n6887), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4550) );
  INV_X1 U5790 ( .A(n4475), .ZN(n6908) );
  AND2_X1 U5791 ( .A1(n4473), .A2(n4472), .ZN(n6786) );
  NAND2_X1 U5792 ( .A1(n6935), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4472) );
  NOR2_X1 U5793 ( .A1(n6951), .A2(n6950), .ZN(n7012) );
  NOR2_X1 U5794 ( .A1(n6948), .A2(n4479), .ZN(n6951) );
  NOR2_X1 U5795 ( .A1(n6609), .A2(n7525), .ZN(n4479) );
  NOR2_X1 U5796 ( .A1(n6952), .A2(n4399), .ZN(n6956) );
  NOR2_X1 U5797 ( .A1(n6956), .A2(n6955), .ZN(n7016) );
  NOR2_X1 U5798 ( .A1(n7379), .A2(n4548), .ZN(n7382) );
  AND2_X1 U5799 ( .A1(n7380), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4548) );
  XNOR2_X1 U5800 ( .A(n7733), .B(n7732), .ZN(n7701) );
  OR2_X1 U5801 ( .A1(n7737), .A2(n7736), .ZN(n7903) );
  NOR2_X1 U5802 ( .A1(n7730), .A2(n7731), .ZN(n7898) );
  AOI21_X1 U5803 ( .B1(n9339), .B2(n9338), .A(n4409), .ZN(n9343) );
  INV_X1 U5804 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5805 ( .A1(n9417), .A2(n6516), .ZN(n9404) );
  AND2_X1 U5806 ( .A1(n5391), .A2(n5390), .ZN(n9427) );
  AND2_X1 U5807 ( .A1(n5331), .A2(n5330), .ZN(n9463) );
  OAI21_X1 U5808 ( .B1(n9491), .B2(n4494), .A(n4491), .ZN(n9459) );
  AND2_X1 U5809 ( .A1(n4495), .A2(n4345), .ZN(n9480) );
  INV_X1 U5810 ( .A(n9648), .ZN(n9585) );
  NAND2_X1 U5811 ( .A1(n4805), .A2(n5635), .ZN(n8058) );
  NAND2_X1 U5812 ( .A1(n5162), .A2(n5161), .ZN(n9045) );
  NAND2_X1 U5813 ( .A1(n7772), .A2(n5589), .ZN(n7868) );
  NAND2_X1 U5814 ( .A1(n5094), .A2(n5093), .ZN(n9067) );
  NOR2_X1 U5815 ( .A1(n4483), .A2(n4829), .ZN(n4485) );
  INV_X1 U5816 ( .A(n4484), .ZN(n4483) );
  AND2_X1 U5817 ( .A1(n4800), .A2(n5624), .ZN(n7424) );
  INV_X1 U5818 ( .A(n9769), .ZN(n9556) );
  INV_X1 U5819 ( .A(n9760), .ZN(n9772) );
  INV_X1 U5820 ( .A(n5540), .ZN(n9373) );
  OR2_X1 U5821 ( .A1(n9395), .A2(n9389), .ZN(n6526) );
  NAND2_X1 U5822 ( .A1(n4499), .A2(n4497), .ZN(n9571) );
  INV_X1 U5823 ( .A(n4500), .ZN(n4497) );
  NAND2_X1 U5824 ( .A1(n7871), .A2(n4324), .ZN(n4499) );
  INV_X1 U5825 ( .A(n9067), .ZN(n6475) );
  NAND2_X1 U5826 ( .A1(n4926), .A2(n5700), .ZN(n4890) );
  NAND2_X1 U5827 ( .A1(n7108), .A2(n7107), .ZN(n9780) );
  INV_X1 U5828 ( .A(n4866), .ZN(n8092) );
  NAND2_X1 U5829 ( .A1(n4879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4863) );
  INV_X1 U5830 ( .A(n6378), .ZN(n7923) );
  INV_X1 U5831 ( .A(n6379), .ZN(n7814) );
  INV_X1 U5832 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10051) );
  INV_X1 U5833 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7583) );
  INV_X1 U5834 ( .A(n6508), .ZN(n7582) );
  INV_X1 U5835 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7421) );
  INV_X1 U5836 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8145) );
  INV_X1 U5837 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U5838 ( .A1(n4583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U5839 ( .A1(n5233), .A2(n5232), .ZN(n4583) );
  INV_X1 U5840 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7030) );
  INV_X1 U5841 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6922) );
  INV_X1 U5842 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6633) );
  INV_X1 U5843 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6621) );
  OR2_X1 U5844 ( .A1(n5070), .A2(n5069), .ZN(n4573) );
  OAI21_X1 U5845 ( .B1(n5041), .B2(n4452), .A(n4450), .ZN(n5070) );
  INV_X1 U5846 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9977) );
  INV_X1 U5847 ( .A(n4915), .ZN(n4913) );
  XNOR2_X1 U5848 ( .A(n4471), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U5849 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4471) );
  NAND2_X1 U5850 ( .A1(n4759), .A2(n8285), .ZN(n4756) );
  INV_X1 U5851 ( .A(n4684), .ZN(n7826) );
  NAND2_X1 U5852 ( .A1(n8701), .A2(n8700), .ZN(n4533) );
  NAND2_X1 U5853 ( .A1(n4535), .A2(n8713), .ZN(n4534) );
  OR2_X1 U5854 ( .A1(n8706), .A2(n8731), .ZN(n4536) );
  NAND2_X1 U5855 ( .A1(n6182), .A2(n9899), .ZN(n6158) );
  OAI21_X1 U5856 ( .B1(n9410), .B2(n10096), .A(n6417), .ZN(n6418) );
  NAND2_X1 U5857 ( .A1(n5618), .A2(n4412), .ZN(n4427) );
  INV_X1 U5858 ( .A(n4544), .ZN(n6938) );
  NAND2_X1 U5859 ( .A1(n4797), .A2(n8125), .ZN(n8137) );
  MUX2_X1 U5860 ( .A(n9591), .B(n9590), .S(n9816), .Z(n9592) );
  NAND2_X1 U5861 ( .A1(n4799), .A2(n4798), .ZN(n8139) );
  NAND2_X1 U5862 ( .A1(n9816), .A2(n8138), .ZN(n4798) );
  NAND2_X1 U5863 ( .A1(n8140), .A2(n9818), .ZN(n4799) );
  NOR2_X1 U5864 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  MUX2_X1 U5865 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n8112), .S(n9818), .Z(n8110)
         );
  OR2_X1 U5866 ( .A1(n9593), .A2(n9717), .ZN(n4831) );
  MUX2_X1 U5867 ( .A(n8141), .B(n8140), .S(n9794), .Z(n8142) );
  NOR2_X1 U5868 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  MUX2_X1 U5869 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n8112), .S(n9794), .Z(n8114)
         );
  INV_X1 U5870 ( .A(n6196), .ZN(n9088) );
  NAND2_X2 U5871 ( .A1(n6624), .A2(n6191), .ZN(n6196) );
  OR2_X1 U5872 ( .A1(n7631), .A2(n7630), .ZN(n4317) );
  NAND2_X1 U5873 ( .A1(n4876), .A2(n4375), .ZN(n4433) );
  AOI21_X1 U5874 ( .B1(n7027), .B2(n5495), .A(n5234), .ZN(n9537) );
  INV_X1 U5875 ( .A(n9537), .ZN(n9639) );
  OR2_X1 U5876 ( .A1(n8991), .A2(n8825), .ZN(n4318) );
  AND2_X1 U5877 ( .A1(n6377), .A2(n4588), .ZN(n4319) );
  NOR2_X1 U5878 ( .A1(n6251), .A2(n6250), .ZN(n4320) );
  INV_X1 U5879 ( .A(n4815), .ZN(n4952) );
  NAND2_X1 U5880 ( .A1(n8301), .A2(n8300), .ZN(n8318) );
  OAI21_X1 U5881 ( .B1(n5107), .B2(n4461), .A(n4385), .ZN(n5174) );
  NAND2_X1 U5882 ( .A1(n7454), .A2(n9758), .ZN(n4323) );
  AND2_X1 U5883 ( .A1(n4347), .A2(n4827), .ZN(n4324) );
  OAI21_X1 U5884 ( .B1(n8254), .B2(n4753), .A(n4751), .ZN(n4750) );
  INV_X1 U5885 ( .A(n4750), .ZN(n4748) );
  AND2_X1 U5886 ( .A1(n4351), .A2(n4860), .ZN(n4325) );
  NAND2_X1 U5887 ( .A1(n5371), .A2(n5370), .ZN(n9678) );
  INV_X1 U5888 ( .A(n8247), .ZN(n4753) );
  OAI21_X1 U5889 ( .B1(n6062), .B2(n4638), .A(n4382), .ZN(n4637) );
  OR2_X1 U5890 ( .A1(n4498), .A2(n6485), .ZN(n4326) );
  AND2_X1 U5891 ( .A1(n6142), .A2(n8469), .ZN(n4327) );
  AND2_X1 U5892 ( .A1(n8183), .A2(n8182), .ZN(n4328) );
  NAND2_X1 U5893 ( .A1(n4748), .A2(n8795), .ZN(n4329) );
  NAND3_X1 U5894 ( .A1(n5608), .A2(n5620), .A3(n5607), .ZN(n4330) );
  AND4_X1 U5895 ( .A1(n4771), .A2(n5793), .A3(n5745), .A4(n4770), .ZN(n4331)
         );
  OAI21_X1 U5896 ( .B1(n7288), .B2(n4783), .A(n4781), .ZN(n7410) );
  OR2_X1 U5897 ( .A1(n5868), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4332) );
  NOR2_X1 U5898 ( .A1(n7526), .A2(n9662), .ZN(n4333) );
  AND2_X1 U5899 ( .A1(n4505), .A2(n4504), .ZN(n4334) );
  OR2_X1 U5900 ( .A1(n8704), .A2(n8703), .ZN(n4335) );
  INV_X4 U5901 ( .A(n6214), .ZN(n6205) );
  NAND2_X1 U5902 ( .A1(n4791), .A2(n5652), .ZN(n6509) );
  OR2_X1 U5903 ( .A1(n8297), .A2(n8199), .ZN(n4336) );
  OR2_X1 U5904 ( .A1(n9269), .A2(n7340), .ZN(n4337) );
  OR2_X1 U5905 ( .A1(n9409), .A2(n4520), .ZN(n4338) );
  OR2_X1 U5906 ( .A1(n5936), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U5907 ( .A1(n8092), .A2(n9726), .ZN(n4920) );
  AND3_X1 U5908 ( .A1(n5920), .A2(n5950), .A3(n5676), .ZN(n4340) );
  INV_X1 U5909 ( .A(n7755), .ZN(n4482) );
  NAND2_X1 U5910 ( .A1(n5989), .A2(n5988), .ZN(n8991) );
  OR2_X1 U5911 ( .A1(n8202), .A2(n8201), .ZN(n4341) );
  NAND2_X1 U5912 ( .A1(n9479), .A2(n4345), .ZN(n4494) );
  NAND2_X1 U5913 ( .A1(n6080), .A2(n4656), .ZN(n6097) );
  NAND2_X1 U5914 ( .A1(n8473), .A2(n8852), .ZN(n8875) );
  AND2_X1 U5915 ( .A1(n4992), .A2(SI_5_), .ZN(n4342) );
  OR4_X1 U5916 ( .A1(n8358), .A2(n8542), .A3(n8357), .A4(n8527), .ZN(n4343) );
  NAND2_X1 U5917 ( .A1(n5457), .A2(n5456), .ZN(n5463) );
  OR2_X1 U5918 ( .A1(n7825), .A2(n7824), .ZN(n4344) );
  OR2_X1 U5919 ( .A1(n9625), .A2(n9254), .ZN(n4345) );
  AND2_X1 U5920 ( .A1(n4527), .A2(n4531), .ZN(n6080) );
  NAND2_X1 U5921 ( .A1(n6496), .A2(n6495), .ZN(n9435) );
  NAND2_X1 U5922 ( .A1(n6150), .A2(n8365), .ZN(n8756) );
  AND2_X1 U5923 ( .A1(n8407), .A2(n8432), .ZN(n4346) );
  OR2_X1 U5924 ( .A1(n9045), .A2(n9259), .ZN(n4347) );
  INV_X1 U5925 ( .A(n8450), .ZN(n4632) );
  INV_X1 U5926 ( .A(n6517), .ZN(n4808) );
  INV_X1 U5927 ( .A(n8804), .ZN(n4615) );
  NAND2_X1 U5928 ( .A1(n8305), .A2(n8304), .ZN(n8319) );
  OR2_X1 U5929 ( .A1(n8563), .A2(n7048), .ZN(n4348) );
  INV_X1 U5930 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5697) );
  AND4_X1 U5931 ( .A1(n5678), .A2(n5677), .A3(n5865), .A4(n5850), .ZN(n4349)
         );
  AND2_X1 U5932 ( .A1(n4858), .A2(n5547), .ZN(n4350) );
  AND2_X1 U5933 ( .A1(n4838), .A2(n4859), .ZN(n4351) );
  AOI21_X1 U5934 ( .B1(n4990), .B2(n4456), .A(n4342), .ZN(n4455) );
  NAND2_X1 U5935 ( .A1(n5438), .A2(n5437), .ZN(n9380) );
  NAND2_X1 U5936 ( .A1(n4997), .A2(n4351), .ZN(n4352) );
  NAND2_X1 U5937 ( .A1(n6080), .A2(n5679), .ZN(n4353) );
  NAND2_X1 U5938 ( .A1(n4721), .A2(n5043), .ZN(n5048) );
  INV_X1 U5939 ( .A(n8532), .ZN(n4572) );
  INV_X1 U5940 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5777) );
  AND2_X1 U5941 ( .A1(n4551), .A2(n4550), .ZN(n4355) );
  NOR2_X1 U5942 ( .A1(n7498), .A2(n5828), .ZN(n4356) );
  AND2_X1 U5943 ( .A1(n8451), .A2(n8558), .ZN(n4357) );
  NAND2_X1 U5944 ( .A1(n4815), .A2(n4813), .ZN(n4358) );
  OR2_X1 U5945 ( .A1(n9600), .A2(n9159), .ZN(n6516) );
  INV_X1 U5946 ( .A(n6516), .ZN(n4812) );
  NAND2_X1 U5947 ( .A1(n5005), .A2(n4858), .ZN(n5546) );
  NAND2_X1 U5948 ( .A1(n4574), .A2(n4912), .ZN(n4953) );
  AND2_X1 U5949 ( .A1(n8078), .A2(n8842), .ZN(n4359) );
  AND2_X1 U5950 ( .A1(n8792), .A2(n8497), .ZN(n4360) );
  NAND2_X1 U5951 ( .A1(n5276), .A2(n5275), .ZN(n9618) );
  NOR2_X1 U5952 ( .A1(n8631), .A2(n8632), .ZN(n4361) );
  NOR2_X1 U5953 ( .A1(n8648), .A2(n8647), .ZN(n4362) );
  NOR2_X1 U5954 ( .A1(n5590), .A2(n4806), .ZN(n4363) );
  AND2_X1 U5955 ( .A1(n7631), .A2(n7630), .ZN(n4364) );
  AND3_X1 U5956 ( .A1(n5222), .A2(n9258), .A3(n9545), .ZN(n4365) );
  AND2_X1 U5957 ( .A1(n4602), .A2(n4317), .ZN(n4366) );
  NAND2_X1 U5958 ( .A1(n7918), .A2(n8557), .ZN(n4367) );
  OR3_X1 U5959 ( .A1(n6244), .A2(n7505), .A3(n7561), .ZN(n4368) );
  AND2_X1 U5960 ( .A1(n7272), .A2(n7270), .ZN(n4369) );
  NOR2_X1 U5961 ( .A1(n9678), .A2(n9250), .ZN(n4370) );
  NOR2_X1 U5962 ( .A1(n8830), .A2(n8806), .ZN(n4371) );
  NOR2_X1 U5963 ( .A1(n8220), .A2(n4834), .ZN(n4372) );
  AND2_X1 U5964 ( .A1(n7954), .A2(n7953), .ZN(n4373) );
  AND2_X1 U5965 ( .A1(n4426), .A2(n4482), .ZN(n4374) );
  NAND2_X1 U5966 ( .A1(n9267), .A2(n7568), .ZN(n6465) );
  AND2_X1 U5967 ( .A1(n4861), .A2(n4431), .ZN(n4375) );
  NAND2_X1 U5968 ( .A1(n5625), .A2(n5624), .ZN(n4376) );
  AND2_X1 U5969 ( .A1(n9618), .A2(n9253), .ZN(n4377) );
  NAND2_X1 U5970 ( .A1(n9175), .A2(n9174), .ZN(n4378) );
  OR2_X1 U5971 ( .A1(n9463), .A2(n9109), .ZN(n4379) );
  AND2_X1 U5972 ( .A1(n5595), .A2(n5592), .ZN(n4380) );
  AND2_X1 U5973 ( .A1(n8510), .A2(n8511), .ZN(n8758) );
  NAND2_X1 U5974 ( .A1(n4597), .A2(n4594), .ZN(n9071) );
  AND2_X1 U5975 ( .A1(n6424), .A2(n6423), .ZN(n4381) );
  NAND2_X1 U5976 ( .A1(n6063), .A2(n8291), .ZN(n4382) );
  NAND2_X1 U5977 ( .A1(n4997), .A2(n4838), .ZN(n4383) );
  INV_X1 U5978 ( .A(n4513), .ZN(n4512) );
  NAND2_X1 U5979 ( .A1(n4515), .A2(n4514), .ZN(n4513) );
  NOR2_X1 U5980 ( .A1(n8923), .A2(n8807), .ZN(n4384) );
  NOR2_X1 U5981 ( .A1(n4620), .A2(n4371), .ZN(n4618) );
  AND2_X1 U5982 ( .A1(n4732), .A2(n4459), .ZN(n4385) );
  AND2_X1 U5983 ( .A1(n6285), .A2(n6284), .ZN(n4386) );
  INV_X1 U5984 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5985 ( .A1(n4630), .A2(n4367), .ZN(n4628) );
  OR2_X1 U5986 ( .A1(n4640), .A2(n8758), .ZN(n4387) );
  AND2_X1 U5987 ( .A1(n8319), .A2(n8555), .ZN(n8542) );
  INV_X1 U5988 ( .A(n4782), .ZN(n4781) );
  OAI21_X1 U5989 ( .B1(n7287), .B2(n4783), .A(n7392), .ZN(n4782) );
  AND2_X1 U5990 ( .A1(n4419), .A2(n6465), .ZN(n4388) );
  INV_X1 U5991 ( .A(n4494), .ZN(n4493) );
  NAND2_X1 U5992 ( .A1(n4495), .A2(n4493), .ZN(n9481) );
  OR2_X1 U5993 ( .A1(n8688), .A2(n8687), .ZN(n4389) );
  AND2_X1 U5994 ( .A1(n5103), .A2(n5089), .ZN(n4390) );
  INV_X1 U5995 ( .A(n6943), .ZN(n7125) );
  NOR2_X1 U5996 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4391) );
  AND2_X1 U5997 ( .A1(n8493), .A2(n8492), .ZN(n8792) );
  INV_X1 U5998 ( .A(n8792), .ZN(n4609) );
  NAND2_X1 U5999 ( .A1(n6649), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U6000 ( .A1(n9419), .A2(n9418), .ZN(n9417) );
  AND2_X1 U6001 ( .A1(n4502), .A2(n4324), .ZN(n4393) );
  OR2_X1 U6002 ( .A1(n8244), .A2(n8193), .ZN(n8510) );
  INV_X1 U6003 ( .A(n4595), .ZN(n4594) );
  OR2_X1 U6004 ( .A1(n9145), .A2(n4596), .ZN(n4595) );
  INV_X1 U6005 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4770) );
  INV_X1 U6006 ( .A(n6963), .ZN(n4682) );
  INV_X1 U6007 ( .A(n6727), .ZN(n4691) );
  NAND2_X1 U6008 ( .A1(n9562), .A2(n9563), .ZN(n9543) );
  NAND2_X1 U6009 ( .A1(n5351), .A2(n5350), .ZN(n9609) );
  INV_X1 U6010 ( .A(n9609), .ZN(n4514) );
  AND2_X1 U6011 ( .A1(n9504), .A2(n9493), .ZN(n9484) );
  AND2_X1 U6012 ( .A1(n9555), .A2(n9537), .ZN(n4394) );
  AND2_X1 U6013 ( .A1(n9484), .A2(n4512), .ZN(n4395) );
  AND2_X1 U6014 ( .A1(n7017), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4396) );
  AND2_X1 U6015 ( .A1(n7549), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4397) );
  OR2_X1 U6016 ( .A1(n7206), .A2(n7205), .ZN(n4398) );
  AND2_X1 U6017 ( .A1(n6953), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4399) );
  INV_X1 U6018 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4566) );
  OAI22_X1 U6019 ( .A1(n7355), .A2(n4653), .B1(n4652), .B2(n8426), .ZN(n7437)
         );
  NAND2_X1 U6020 ( .A1(n4576), .A2(n4575), .ZN(n9037) );
  OAI21_X1 U6021 ( .B1(n7476), .B2(n5882), .A(n5881), .ZN(n7745) );
  NAND2_X1 U6022 ( .A1(n5146), .A2(n5145), .ZN(n9190) );
  NAND2_X1 U6023 ( .A1(n5116), .A2(n5115), .ZN(n9662) );
  NAND2_X1 U6024 ( .A1(n4633), .A2(n8469), .ZN(n8873) );
  AND3_X1 U6025 ( .A1(n5029), .A2(n5028), .A3(n5027), .ZN(n7767) );
  NAND2_X1 U6026 ( .A1(n5720), .A2(n5699), .ZN(n6704) );
  NOR2_X1 U6027 ( .A1(n8585), .A2(n8586), .ZN(n4400) );
  NOR2_X1 U6028 ( .A1(n9648), .A2(n9137), .ZN(n4401) );
  AND3_X1 U6029 ( .A1(n4958), .A2(n4957), .A3(n4956), .ZN(n7340) );
  INV_X1 U6030 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4862) );
  AND4_X1 U6031 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n7720)
         );
  INV_X1 U6032 ( .A(n6485), .ZN(n4502) );
  NOR2_X1 U6033 ( .A1(n9585), .A2(n9258), .ZN(n6485) );
  NOR2_X1 U6034 ( .A1(n7918), .A2(n8557), .ZN(n4402) );
  AND2_X1 U6035 ( .A1(n5825), .A2(n5824), .ZN(n7545) );
  NAND2_X1 U6036 ( .A1(n6010), .A2(n6009), .ZN(n8773) );
  AND3_X1 U6037 ( .A1(n6649), .A2(n4769), .A3(n9983), .ZN(n4403) );
  AND2_X1 U6038 ( .A1(n5642), .A2(n9572), .ZN(n4404) );
  XNOR2_X1 U6039 ( .A(n6942), .B(n7103), .ZN(n7091) );
  NAND2_X1 U6040 ( .A1(n7288), .A2(n7287), .ZN(n7391) );
  NAND2_X1 U6041 ( .A1(n4509), .A2(n4507), .ZN(n8070) );
  INV_X1 U6042 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U6043 ( .A1(n5752), .A2(n5751), .ZN(n7169) );
  INV_X1 U6044 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4590) );
  OR2_X1 U6045 ( .A1(n7526), .A2(n4510), .ZN(n4405) );
  NOR2_X1 U6046 ( .A1(n7546), .A2(n7547), .ZN(n4406) );
  AND2_X1 U6047 ( .A1(n4849), .A2(n4741), .ZN(n4407) );
  OR2_X1 U6048 ( .A1(n7344), .A2(n8340), .ZN(n4651) );
  INV_X1 U6049 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5869) );
  XNOR2_X1 U6050 ( .A(n4875), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U6051 ( .A(n5008), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5619) );
  NAND4_X1 U6052 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n6942)
         );
  OR2_X1 U6053 ( .A1(n4506), .A2(n7338), .ZN(n4408) );
  AND2_X2 U6054 ( .A1(n6181), .A2(n6180), .ZN(n9915) );
  AND2_X1 U6055 ( .A1(n9337), .A2(n9640), .ZN(n4409) );
  XOR2_X1 U6056 ( .A(n4316), .B(P2_REG1_REG_19__SCAN_IN), .Z(n4410) );
  INV_X1 U6057 ( .A(n7390), .ZN(n4783) );
  INV_X2 U6058 ( .A(n9816), .ZN(n9818) );
  NAND2_X1 U6059 ( .A1(n6532), .A2(n6531), .ZN(n9816) );
  AND2_X1 U6060 ( .A1(n6802), .A2(n6820), .ZN(n6805) );
  INV_X1 U6061 ( .A(n8331), .ZN(n6135) );
  NOR2_X1 U6062 ( .A1(n5675), .A2(n5674), .ZN(n4411) );
  AND2_X1 U6063 ( .A1(n5666), .A2(n5617), .ZN(n4412) );
  AND2_X1 U6064 ( .A1(n4410), .A2(n4672), .ZN(n4413) );
  OR2_X1 U6065 ( .A1(n7901), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4414) );
  AND2_X1 U6066 ( .A1(n4700), .A2(n4705), .ZN(n4415) );
  OR2_X1 U6067 ( .A1(n4410), .A2(n4672), .ZN(n4416) );
  INV_X1 U6068 ( .A(n6898), .ZN(n4542) );
  INV_X1 U6069 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7145) );
  OR2_X1 U6070 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8702), .ZN(n4417) );
  XNOR2_X1 U6071 ( .A(n7824), .B(n7825), .ZN(n7535) );
  NOR2_X1 U6072 ( .A1(n7598), .A2(n7597), .ZN(n7596) );
  XNOR2_X1 U6073 ( .A(n7532), .B(n7545), .ZN(n7498) );
  NOR2_X1 U6074 ( .A1(n7217), .A2(n7216), .ZN(n7220) );
  NOR2_X1 U6075 ( .A1(n8599), .A2(n8600), .ZN(n8603) );
  XNOR2_X1 U6076 ( .A(n8645), .B(n8646), .ZN(n8623) );
  NAND2_X1 U6077 ( .A1(n7072), .A2(n7205), .ZN(n4705) );
  INV_X1 U6078 ( .A(n7205), .ZN(n4703) );
  XNOR2_X1 U6079 ( .A(n8630), .B(n8646), .ZN(n8611) );
  NAND3_X1 U6080 ( .A1(n4421), .A2(n4337), .A3(n4323), .ZN(n4418) );
  OAI211_X1 U6081 ( .C1(n4430), .C2(n4429), .A(n4428), .B(n4427), .ZN(P1_U3242) );
  AOI21_X1 U6082 ( .B1(n5662), .B2(n5666), .A(n4411), .ZN(n4428) );
  NAND2_X1 U6083 ( .A1(n4330), .A2(n5666), .ZN(n4429) );
  INV_X1 U6084 ( .A(n5609), .ZN(n4430) );
  XNOR2_X2 U6085 ( .A(n4432), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4866) );
  NAND3_X1 U6086 ( .A1(n4436), .A2(n5221), .A3(n9545), .ZN(n4435) );
  NAND3_X1 U6087 ( .A1(n5217), .A2(n5643), .A3(n4404), .ZN(n4436) );
  NAND3_X1 U6088 ( .A1(n4322), .A2(n4894), .A3(n6943), .ZN(n4787) );
  NAND4_X1 U6089 ( .A1(n4813), .A2(n4590), .A3(n4815), .A4(n4837), .ZN(n5006)
         );
  AND3_X2 U6090 ( .A1(n4912), .A2(n4574), .A3(n4852), .ZN(n4815) );
  NAND2_X1 U6091 ( .A1(n4444), .A2(n4440), .ZN(n5487) );
  NAND2_X1 U6092 ( .A1(n4441), .A2(n5614), .ZN(n4440) );
  NAND2_X1 U6093 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  OAI21_X1 U6094 ( .B1(n5434), .B2(n5554), .A(n8099), .ZN(n4443) );
  NAND2_X1 U6095 ( .A1(n4446), .A2(n5553), .ZN(n4445) );
  NAND3_X1 U6096 ( .A1(n4454), .A2(n5018), .A3(n4453), .ZN(n4555) );
  NAND2_X1 U6097 ( .A1(n4972), .A2(n4455), .ZN(n4454) );
  OAI21_X1 U6098 ( .B1(n4972), .B2(n4989), .A(n4455), .ZN(n5019) );
  NAND2_X1 U6099 ( .A1(n4607), .A2(n4467), .ZN(n8784) );
  NAND3_X1 U6100 ( .A1(n4469), .A2(n4468), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4886) );
  OAI21_X2 U6101 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4880), .ZN(n4468) );
  NOR2_X1 U6102 ( .A1(n4829), .A2(n4482), .ZN(n4481) );
  OAI21_X1 U6103 ( .B1(n4485), .B2(n7755), .A(n7753), .ZN(n9751) );
  OAI21_X1 U6104 ( .B1(n9491), .B2(n4490), .A(n4487), .ZN(n4486) );
  NAND2_X1 U6105 ( .A1(n7871), .A2(n4393), .ZN(n4496) );
  NAND2_X1 U6106 ( .A1(n4496), .A2(n4326), .ZN(n9554) );
  NAND3_X1 U6107 ( .A1(n4347), .A2(n4827), .A3(n6483), .ZN(n4501) );
  AND2_X2 U6108 ( .A1(n4997), .A2(n4818), .ZN(n4876) );
  AND2_X2 U6109 ( .A1(n5005), .A2(n4350), .ZN(n4997) );
  AND2_X2 U6110 ( .A1(n5091), .A2(n6572), .ZN(n4926) );
  NAND2_X2 U6111 ( .A1(n5673), .A2(n5672), .ZN(n5091) );
  INV_X1 U6112 ( .A(n7526), .ZN(n4509) );
  NOR2_X1 U6113 ( .A1(n9409), .A2(n6525), .ZN(n8108) );
  NAND2_X1 U6114 ( .A1(n5005), .A2(n4523), .ZN(n4873) );
  NAND3_X1 U6115 ( .A1(n4527), .A2(n4531), .A3(n4654), .ZN(n6104) );
  NAND3_X1 U6116 ( .A1(n4531), .A2(n4528), .A3(n4340), .ZN(n6076) );
  NAND4_X1 U6117 ( .A1(n4537), .A2(n4536), .A3(n4534), .A4(n4533), .ZN(
        P2_U3200) );
  NAND3_X1 U6118 ( .A1(n4560), .A2(n8475), .A3(n4556), .ZN(n8478) );
  NAND3_X1 U6119 ( .A1(n8472), .A2(n8471), .A3(n6142), .ZN(n4559) );
  OR2_X1 U6120 ( .A1(n8521), .A2(n4570), .ZN(n4567) );
  NAND2_X1 U6121 ( .A1(n9116), .A2(n4578), .ZN(n4576) );
  NAND2_X1 U6122 ( .A1(n5233), .A2(n4584), .ZN(n4582) );
  NAND2_X1 U6123 ( .A1(n4586), .A2(n4587), .ZN(n6431) );
  NAND2_X1 U6124 ( .A1(n9156), .A2(n4319), .ZN(n4586) );
  NAND2_X1 U6125 ( .A1(n9156), .A2(n6365), .ZN(n9128) );
  NAND3_X1 U6126 ( .A1(n4815), .A2(n4813), .A3(n4837), .ZN(n5183) );
  OAI21_X1 U6127 ( .B1(n9135), .B2(n4595), .A(n4591), .ZN(n9070) );
  NAND2_X1 U6128 ( .A1(n9135), .A2(n9136), .ZN(n4597) );
  INV_X1 U6129 ( .A(n7573), .ZN(n4602) );
  INV_X1 U6130 ( .A(n4826), .ZN(n4603) );
  NAND2_X1 U6131 ( .A1(n4605), .A2(n4604), .ZN(n7633) );
  OAI22_X1 U6132 ( .A1(n7178), .A2(n7177), .B1(n6135), .B2(n4606), .ZN(n7181)
         );
  NAND2_X1 U6133 ( .A1(n4606), .A2(n6134), .ZN(n7178) );
  NAND2_X1 U6134 ( .A1(n8814), .A2(n4608), .ZN(n4607) );
  NAND4_X1 U6135 ( .A1(n7149), .A2(n7148), .A3(n8386), .A4(n8395), .ZN(n4621)
         );
  NAND3_X1 U6136 ( .A1(n7149), .A2(n7148), .A3(n8386), .ZN(n7150) );
  NAND2_X1 U6137 ( .A1(n4648), .A2(n4649), .ZN(n7441) );
  NAND2_X1 U6138 ( .A1(n7344), .A2(n4346), .ZN(n4648) );
  AOI21_X1 U6139 ( .B1(n4346), .B2(n8340), .A(n4650), .ZN(n4649) );
  NAND2_X1 U6140 ( .A1(n6560), .A2(n4658), .ZN(n4819) );
  INV_X1 U6141 ( .A(n6558), .ZN(n6560) );
  NAND2_X1 U6142 ( .A1(n5699), .A2(n4392), .ZN(n4659) );
  OAI21_X1 U6143 ( .B1(n5719), .B2(n4659), .A(n6722), .ZN(n6646) );
  OAI21_X1 U6144 ( .B1(n6704), .B2(n6650), .A(n6713), .ZN(n6652) );
  NAND2_X1 U6145 ( .A1(n7954), .A2(n4662), .ZN(n4661) );
  OAI211_X1 U6146 ( .C1(n7954), .C2(n8598), .A(n4663), .B(n4661), .ZN(n7956)
         );
  NOR2_X1 U6147 ( .A1(n8685), .A2(n4410), .ZN(n4669) );
  NAND2_X1 U6148 ( .A1(n4671), .A2(n4416), .ZN(n4666) );
  NAND3_X1 U6149 ( .A1(n4670), .A2(n4668), .A3(n4667), .ZN(n8728) );
  NAND2_X1 U6150 ( .A1(n4669), .A2(n4671), .ZN(n4668) );
  NAND3_X1 U6151 ( .A1(n4673), .A2(n4675), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n6755) );
  NAND2_X1 U6152 ( .A1(n4674), .A2(n6727), .ZN(n4673) );
  NAND2_X1 U6153 ( .A1(n8575), .A2(n6726), .ZN(n4674) );
  NAND2_X1 U6154 ( .A1(n4677), .A2(n8575), .ZN(n4675) );
  NAND2_X1 U6155 ( .A1(n4676), .A2(n6727), .ZN(n6753) );
  NOR2_X1 U6156 ( .A1(n6727), .A2(n4678), .ZN(n4677) );
  INV_X1 U6157 ( .A(n6726), .ZN(n4678) );
  NAND2_X1 U6158 ( .A1(n4680), .A2(n6971), .ZN(n6969) );
  INV_X1 U6159 ( .A(n6862), .ZN(n4683) );
  NAND2_X1 U6160 ( .A1(n4689), .A2(n6742), .ZN(n6744) );
  NAND2_X1 U6161 ( .A1(n4694), .A2(n6977), .ZN(n6975) );
  INV_X1 U6162 ( .A(n6855), .ZN(n4696) );
  OAI21_X1 U6163 ( .B1(n8611), .B2(n4707), .A(n4706), .ZN(n8657) );
  NAND2_X1 U6164 ( .A1(n5415), .A2(n5414), .ZN(n4715) );
  OAI21_X1 U6165 ( .B1(n5415), .B2(n4718), .A(n4716), .ZN(n5436) );
  NAND2_X1 U6166 ( .A1(n5415), .A2(n4716), .ZN(n4714) );
  INV_X1 U6167 ( .A(n4722), .ZN(n5396) );
  NAND2_X1 U6168 ( .A1(n5348), .A2(n5347), .ZN(n5365) );
  NAND2_X1 U6169 ( .A1(n5090), .A2(n4390), .ZN(n5107) );
  NAND2_X1 U6170 ( .A1(n5287), .A2(n4743), .ZN(n4742) );
  OAI21_X2 U6171 ( .B1(n4745), .B2(n4744), .A(n8283), .ZN(n8282) );
  OAI21_X1 U6172 ( .B1(n8211), .B2(n4329), .A(n4746), .ZN(n4745) );
  NOR2_X2 U6173 ( .A1(n8211), .A2(n8773), .ZN(n8256) );
  AOI21_X1 U6174 ( .B1(n4749), .B2(n4752), .A(n4750), .ZN(n8245) );
  INV_X1 U6175 ( .A(n8256), .ZN(n4749) );
  NAND2_X1 U6176 ( .A1(n8202), .A2(n4755), .ZN(n4754) );
  OAI211_X1 U6177 ( .C1(n8202), .C2(n4756), .A(n4754), .B(n8229), .ZN(P2_U3160) );
  NAND3_X1 U6178 ( .A1(n4331), .A2(n4772), .A3(n4403), .ZN(n5822) );
  INV_X1 U6179 ( .A(n6837), .ZN(n4773) );
  XNOR2_X1 U6180 ( .A(n6993), .B(n8376), .ZN(n6837) );
  NAND2_X1 U6181 ( .A1(n8003), .A2(n4776), .ZN(n4774) );
  NAND2_X1 U6182 ( .A1(n4774), .A2(n4775), .ZN(n8175) );
  OAI21_X2 U6183 ( .B1(n7288), .B2(n4780), .A(n4779), .ZN(n7412) );
  NAND2_X1 U6184 ( .A1(n8235), .A2(n4328), .ZN(n8275) );
  OAI21_X1 U6185 ( .B1(n7091), .B2(n4787), .A(n4900), .ZN(n7249) );
  OAI21_X1 U6186 ( .B1(n7249), .B2(n4919), .A(n5627), .ZN(n7304) );
  NAND2_X1 U6187 ( .A1(n4788), .A2(n4789), .ZN(n6512) );
  NAND2_X1 U6188 ( .A1(n9511), .A2(n4792), .ZN(n4788) );
  NAND2_X1 U6189 ( .A1(n8123), .A2(n9575), .ZN(n4797) );
  NAND2_X1 U6190 ( .A1(n4801), .A2(n4802), .ZN(n5598) );
  NAND2_X1 U6191 ( .A1(n5593), .A2(n4380), .ZN(n4801) );
  NAND2_X1 U6192 ( .A1(n4805), .A2(n4804), .ZN(n8059) );
  AND2_X1 U6193 ( .A1(n9380), .A2(n6528), .ZN(n8113) );
  OR2_X1 U6194 ( .A1(n6796), .A2(n8522), .ZN(n6814) );
  OR2_X1 U6195 ( .A1(n5683), .A2(n6078), .ZN(n5684) );
  INV_X1 U6196 ( .A(n8064), .ZN(n8066) );
  INV_X1 U6197 ( .A(n9270), .ZN(n7201) );
  XNOR2_X1 U6198 ( .A(n8118), .B(n8121), .ZN(n8143) );
  NAND2_X1 U6199 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U6200 ( .A1(n4334), .A2(n7767), .ZN(n7762) );
  AOI21_X2 U6201 ( .B1(n7987), .B2(n7986), .A(n4841), .ZN(n8001) );
  NAND2_X1 U6202 ( .A1(n5670), .A2(n4874), .ZN(n4875) );
  AOI21_X1 U6203 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7549), .A(n7607), .ZN(
        n7817) );
  NAND2_X1 U6204 ( .A1(n7257), .A2(n10097), .ZN(n7302) );
  NAND2_X1 U6205 ( .A1(n4938), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4870) );
  AOI21_X1 U6206 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8670), .A(n8669), .ZN(
        n8684) );
  OAI21_X2 U6207 ( .B1(n7158), .B2(n8339), .A(n8414), .ZN(n7193) );
  AOI21_X1 U6208 ( .B1(n8102), .B2(n8101), .A(n9497), .ZN(n8106) );
  NAND2_X1 U6209 ( .A1(n6800), .A2(n8946), .ZN(n8368) );
  OR2_X1 U6210 ( .A1(n6046), .A2(n6849), .ZN(n5759) );
  NAND2_X1 U6211 ( .A1(n5688), .A2(n5687), .ZN(n5971) );
  AOI21_X1 U6212 ( .B1(n9424), .B2(n5462), .A(n5394), .ZN(n9159) );
  NAND2_X1 U6213 ( .A1(n5517), .A2(n6205), .ZN(n6200) );
  OR2_X1 U6214 ( .A1(n9899), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4820) );
  OR2_X1 U6215 ( .A1(n6624), .A2(n6201), .ZN(n4821) );
  INV_X1 U6216 ( .A(n9794), .ZN(n9809) );
  INV_X1 U6217 ( .A(n10103), .ZN(n6436) );
  INV_X1 U6218 ( .A(n9778), .ZN(n9745) );
  OR2_X1 U6219 ( .A1(n8169), .A2(n9016), .ZN(n4822) );
  AND2_X1 U6220 ( .A1(n8359), .A2(n4343), .ZN(n4823) );
  OR2_X1 U6221 ( .A1(n9899), .A2(n6156), .ZN(n4824) );
  AND4_X1 U6222 ( .A1(n8740), .A2(n8758), .A3(n8771), .A4(n8352), .ZN(n4825)
         );
  INV_X1 U6223 ( .A(n6525), .ZN(n9393) );
  AND2_X1 U6224 ( .A1(n4368), .A2(n6245), .ZN(n4826) );
  OR2_X1 U6225 ( .A1(n9190), .A2(n9260), .ZN(n4827) );
  OR2_X1 U6226 ( .A1(n7117), .A2(n6446), .ZN(n9579) );
  INV_X1 U6227 ( .A(n9579), .ZN(n6447) );
  NOR2_X1 U6228 ( .A1(n6244), .A2(n4843), .ZN(n4828) );
  NOR2_X1 U6229 ( .A1(n6467), .A2(n7452), .ZN(n4829) );
  AND4_X1 U6230 ( .A1(n5581), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n4830)
         );
  OR2_X1 U6231 ( .A1(n8169), .A2(n8942), .ZN(n4832) );
  AND2_X1 U6232 ( .A1(n5577), .A2(n5576), .ZN(n4833) );
  AND2_X1 U6233 ( .A1(n8218), .A2(n8751), .ZN(n4834) );
  NOR2_X1 U6234 ( .A1(n5594), .A2(n5644), .ZN(n4835) );
  OR2_X1 U6235 ( .A1(n9718), .A2(n6484), .ZN(n4836) );
  AND3_X1 U6236 ( .A1(n4999), .A2(n5002), .A3(n5664), .ZN(n4838) );
  OR2_X1 U6237 ( .A1(n9557), .A2(n9236), .ZN(n4839) );
  AND2_X1 U6238 ( .A1(n9639), .A2(n9257), .ZN(n4840) );
  INV_X1 U6239 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5007) );
  INV_X1 U6240 ( .A(n9260), .ZN(n6482) );
  NAND2_X1 U6241 ( .A1(n6049), .A2(n6048), .ZN(n8743) );
  INV_X1 U6242 ( .A(n7518), .ZN(n9264) );
  NOR2_X1 U6243 ( .A1(n7985), .A2(n7984), .ZN(n4841) );
  NAND2_X1 U6244 ( .A1(n9713), .A2(n9788), .ZN(n9717) );
  INV_X1 U6245 ( .A(n9717), .ZN(n6528) );
  INV_X1 U6246 ( .A(n9729), .ZN(n9723) );
  INV_X1 U6247 ( .A(n9659), .ZN(n6535) );
  AND2_X1 U6248 ( .A1(n8172), .A2(n8865), .ZN(n4842) );
  AND2_X1 U6249 ( .A1(n6023), .A2(n6022), .ZN(n8760) );
  INV_X1 U6250 ( .A(n8760), .ZN(n8785) );
  NAND2_X1 U6251 ( .A1(n5619), .A2(n7402), .ZN(n6507) );
  NAND2_X1 U6252 ( .A1(n8550), .A2(n8370), .ZN(n8522) );
  AND2_X1 U6253 ( .A1(n7561), .A2(n7505), .ZN(n4843) );
  AND2_X1 U6254 ( .A1(n6171), .A2(n6170), .ZN(n4844) );
  AND2_X1 U6255 ( .A1(n7306), .A2(n7340), .ZN(n4845) );
  OR2_X1 U6256 ( .A1(n5615), .A2(n5614), .ZN(n4846) );
  AND2_X1 U6257 ( .A1(n6271), .A2(n6270), .ZN(n4847) );
  OR2_X1 U6258 ( .A1(n5323), .A2(SI_21_), .ZN(n4849) );
  INV_X1 U6259 ( .A(n9190), .ZN(n8049) );
  OR2_X1 U6260 ( .A1(n6514), .A2(n5614), .ZN(n4850) );
  NOR2_X1 U6261 ( .A1(n9399), .A2(n6501), .ZN(n4851) );
  AOI21_X1 U6262 ( .B1(n5211), .B2(n4835), .A(n5210), .ZN(n5220) );
  AND2_X1 U6263 ( .A1(n9436), .A2(n4850), .ZN(n5379) );
  NAND2_X1 U6264 ( .A1(n5380), .A2(n5379), .ZN(n5382) );
  NAND2_X1 U6265 ( .A1(n5382), .A2(n5381), .ZN(n5446) );
  AND2_X1 U6266 ( .A1(n8512), .A2(n8353), .ZN(n8513) );
  NOR2_X1 U6267 ( .A1(n5448), .A2(n5614), .ZN(n5449) );
  NAND2_X1 U6268 ( .A1(n8527), .A2(n8536), .ZN(n8528) );
  NAND2_X1 U6269 ( .A1(n8526), .A2(n8522), .ZN(n8529) );
  INV_X1 U6270 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U6271 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U6272 ( .A1(n8356), .A2(n8355), .ZN(n8527) );
  OR2_X1 U6273 ( .A1(n6508), .A2(n5620), .ZN(n5614) );
  INV_X1 U6274 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4859) );
  OR2_X1 U6275 ( .A1(n6797), .A2(n8329), .ZN(n6798) );
  INV_X1 U6276 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4999) );
  INV_X1 U6277 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4881) );
  INV_X1 U6278 ( .A(n8743), .ZN(n8199) );
  OR2_X1 U6279 ( .A1(n6800), .A2(n6801), .ZN(n6802) );
  INV_X1 U6280 ( .A(n7275), .ZN(n7272) );
  OR2_X1 U6281 ( .A1(n5940), .A2(n6810), .ZN(n5690) );
  INV_X1 U6282 ( .A(n7215), .ZN(n7217) );
  INV_X1 U6283 ( .A(n8598), .ZN(n7955) );
  INV_X1 U6284 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5873) );
  INV_X1 U6285 ( .A(n8878), .ZN(n8842) );
  NAND2_X1 U6286 ( .A1(n9770), .A2(n9092), .ZN(n6195) );
  INV_X1 U6287 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5056) );
  OR2_X1 U6288 ( .A1(n7433), .A2(n6234), .ZN(n6238) );
  INV_X1 U6289 ( .A(n5334), .ZN(n5332) );
  INV_X1 U6290 ( .A(n5203), .ZN(n5188) );
  INV_X1 U6291 ( .A(n5082), .ZN(n5080) );
  INV_X1 U6292 ( .A(n5322), .ZN(n5323) );
  INV_X1 U6293 ( .A(SI_17_), .ZN(n5228) );
  INV_X1 U6294 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5785) );
  INV_X1 U6295 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U6296 ( .A1(n5887), .A2(n10009), .ZN(n5899) );
  OR2_X1 U6297 ( .A1(n6067), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6084) );
  INV_X1 U6298 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5694) );
  INV_X1 U6299 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U6300 ( .A1(n5874), .A2(n5873), .ZN(n5888) );
  OR2_X1 U6301 ( .A1(n5770), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5787) );
  OR2_X1 U6302 ( .A1(n6162), .A2(n6178), .ZN(n6164) );
  OR2_X1 U6303 ( .A1(n6110), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6109) );
  INV_X1 U6304 ( .A(n6342), .ZN(n6343) );
  INV_X1 U6305 ( .A(n9085), .ZN(n6372) );
  OR2_X1 U6306 ( .A1(n5406), .A2(n5405), .ZN(n5427) );
  OR2_X1 U6307 ( .A1(n5011), .A2(n5010), .ZN(n5031) );
  INV_X1 U6308 ( .A(n8155), .ZN(n8127) );
  NAND2_X1 U6309 ( .A1(n5332), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5353) );
  OR2_X1 U6310 ( .A1(n5147), .A2(n9186), .ZN(n5164) );
  NAND2_X1 U6311 ( .A1(n5080), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5095) );
  AND2_X1 U6312 ( .A1(n5435), .A2(n5420), .ZN(n5421) );
  AND2_X1 U6313 ( .A1(n5364), .A2(n5346), .ZN(n5347) );
  NAND2_X1 U6314 ( .A1(n6030), .A2(n6029), .ZN(n6041) );
  INV_X1 U6315 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U6316 ( .A1(n6016), .A2(n6015), .ZN(n6031) );
  OR2_X1 U6317 ( .A1(n6123), .A2(n8329), .ZN(n6691) );
  INV_X1 U6318 ( .A(n8751), .ZN(n8291) );
  OR2_X1 U6319 ( .A1(n4848), .A2(n8541), .ZN(n8546) );
  OR2_X1 U6320 ( .A1(n5971), .A2(n10082), .ZN(n5730) );
  AOI21_X1 U6321 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8670), .A(n8657), .ZN(
        n8679) );
  AND2_X1 U6322 ( .A1(n6644), .A2(n8089), .ZN(n6648) );
  OR2_X1 U6323 ( .A1(n6041), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6055) );
  INV_X1 U6324 ( .A(n8773), .ZN(n8795) );
  INV_X1 U6325 ( .A(n8890), .ZN(n8863) );
  AND2_X1 U6326 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  OR2_X1 U6327 ( .A1(n6175), .A2(n6797), .ZN(n6675) );
  INV_X1 U6328 ( .A(n6145), .ZN(n8837) );
  OR2_X1 U6329 ( .A1(n8025), .A2(n7891), .ZN(n8465) );
  NAND2_X1 U6330 ( .A1(n7584), .A2(n7406), .ZN(n9886) );
  OAI22_X1 U6331 ( .A1(n7201), .A2(n9085), .B1(n7321), .B2(n6264), .ZN(n7366)
         );
  INV_X1 U6332 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7635) );
  AND2_X1 U6333 ( .A1(n5458), .A2(n5441), .ZN(n9379) );
  OAI21_X1 U6334 ( .B1(n9448), .B2(n9447), .A(n6514), .ZN(n9431) );
  INV_X1 U6335 ( .A(n9237), .ZN(n9220) );
  NAND2_X1 U6336 ( .A1(n5661), .A2(n5545), .ZN(n7315) );
  INV_X1 U6337 ( .A(n9235), .ZN(n9196) );
  INV_X1 U6338 ( .A(n9575), .ZN(n9497) );
  NAND2_X1 U6339 ( .A1(n6624), .A2(n6567), .ZN(n7110) );
  MUX2_X1 U6340 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5668), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5669) );
  AND2_X1 U6341 ( .A1(n5089), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6342 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  AND2_X1 U6343 ( .A1(n7890), .A2(n7984), .ZN(n8027) );
  INV_X1 U6344 ( .A(n8268), .ZN(n8288) );
  INV_X1 U6345 ( .A(n8272), .ZN(n8285) );
  AND2_X1 U6346 ( .A1(n6074), .A2(n6073), .ZN(n8524) );
  AND3_X1 U6347 ( .A1(n5983), .A2(n5982), .A3(n5981), .ZN(n8843) );
  AND4_X1 U6348 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n7886)
         );
  NOR2_X1 U6349 ( .A1(n7533), .A2(n4356), .ZN(n7598) );
  INV_X1 U6350 ( .A(n8724), .ZN(n8676) );
  AOI21_X1 U6351 ( .B1(n4389), .B2(n8690), .A(n8689), .ZN(n8705) );
  OAI211_X1 U6352 ( .C1(n8738), .C2(n8169), .A(n8168), .B(n4819), .ZN(n8170)
         );
  INV_X1 U6353 ( .A(n8864), .ZN(n9826) );
  NAND2_X1 U6354 ( .A1(n6180), .A2(n6165), .ZN(n6168) );
  INV_X1 U6355 ( .A(n8942), .ZN(n8939) );
  AND3_X1 U6356 ( .A1(n6675), .A2(n6160), .A3(n6678), .ZN(n6180) );
  AND2_X1 U6357 ( .A1(n8846), .A2(n8845), .ZN(n9000) );
  OR2_X1 U6358 ( .A1(n8450), .A2(n4357), .ZN(n8346) );
  INV_X1 U6359 ( .A(n9886), .ZN(n9892) );
  NAND2_X1 U6360 ( .A1(n9833), .A2(n9874), .ZN(n9895) );
  NAND2_X1 U6361 ( .A1(n6680), .A2(n6687), .ZN(n6683) );
  AND2_X1 U6362 ( .A1(n5870), .A2(n4332), .ZN(n7831) );
  OAI21_X1 U6363 ( .B1(n6207), .B2(n9085), .A(n6206), .ZN(n6941) );
  INV_X1 U6364 ( .A(n10096), .ZN(n9228) );
  AND4_X1 U6365 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n9221)
         );
  INV_X1 U6366 ( .A(n9360), .ZN(n7376) );
  INV_X1 U6367 ( .A(n9778), .ZN(n9568) );
  INV_X1 U6368 ( .A(n9589), .ZN(n9763) );
  OR2_X1 U6369 ( .A1(n7110), .A2(n6450), .ZN(n9754) );
  AND2_X1 U6370 ( .A1(n9380), .A2(n6535), .ZN(n8109) );
  AND2_X1 U6371 ( .A1(n6384), .A2(n9721), .ZN(n6531) );
  INV_X1 U6372 ( .A(n9804), .ZN(n9788) );
  NAND2_X1 U6373 ( .A1(n8063), .A2(n9781), .ZN(n9801) );
  INV_X1 U6374 ( .A(n9809), .ZN(n9713) );
  XNOR2_X1 U6375 ( .A(n5665), .B(n5664), .ZN(n6626) );
  INV_X1 U6376 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5232) );
  INV_X1 U6377 ( .A(n8244), .ZN(n8969) );
  AND2_X1 U6378 ( .A1(n6830), .A2(n8553), .ZN(n8223) );
  AND2_X1 U6379 ( .A1(n6693), .A2(n6692), .ZN(n8272) );
  AND2_X1 U6380 ( .A1(n8313), .A2(n6089), .ZN(n8225) );
  INV_X1 U6381 ( .A(n7886), .ZN(n8558) );
  OR2_X1 U6382 ( .A1(n6680), .A2(n6571), .ZN(n8697) );
  OR2_X1 U6383 ( .A1(P2_U3150), .A2(n6655), .ZN(n8704) );
  INV_X1 U6384 ( .A(n8727), .ZN(n8689) );
  OR2_X1 U6385 ( .A1(n6665), .A2(n6091), .ZN(n8731) );
  NAND2_X1 U6386 ( .A1(n6168), .A2(n9821), .ZN(n9837) );
  NAND2_X1 U6387 ( .A1(n8894), .A2(n6167), .ZN(n8903) );
  NAND2_X1 U6388 ( .A1(n9915), .A2(n9895), .ZN(n8943) );
  INV_X1 U6389 ( .A(n9915), .ZN(n9913) );
  NAND2_X1 U6390 ( .A1(n9899), .A2(n9895), .ZN(n9018) );
  AND2_X1 U6391 ( .A1(n6130), .A2(n6129), .ZN(n9901) );
  INV_X2 U6392 ( .A(n9901), .ZN(n9899) );
  INV_X1 U6393 ( .A(n6683), .ZN(n6600) );
  INV_X1 U6394 ( .A(n8370), .ZN(n7406) );
  INV_X1 U6395 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6631) );
  OR2_X1 U6396 ( .A1(n5765), .A2(n5778), .ZN(n6963) );
  INV_X1 U6397 ( .A(n9366), .ZN(n9739) );
  INV_X1 U6398 ( .A(n9242), .ZN(n9226) );
  NAND2_X1 U6399 ( .A1(n6415), .A2(n6400), .ZN(n10103) );
  OR2_X1 U6400 ( .A1(n5358), .A2(n5357), .ZN(n9251) );
  INV_X1 U6401 ( .A(n9137), .ZN(n9258) );
  INV_X1 U6402 ( .A(n7651), .ZN(n9265) );
  OR2_X1 U6403 ( .A1(n9741), .A2(n9735), .ZN(n9356) );
  NAND2_X1 U6404 ( .A1(n6775), .A2(n6774), .ZN(n9366) );
  AND2_X1 U6405 ( .A1(n7777), .A2(n9122), .ZN(n7855) );
  OR2_X1 U6406 ( .A1(n9778), .A2(n7316), .ZN(n9589) );
  AND2_X2 U6407 ( .A1(n7114), .A2(n9754), .ZN(n9778) );
  NAND2_X1 U6408 ( .A1(n9818), .A2(n9788), .ZN(n9659) );
  NAND2_X1 U6409 ( .A1(n9818), .A2(n9801), .ZN(n9653) );
  INV_X1 U6410 ( .A(n9045), .ZN(n9718) );
  AND2_X1 U6411 ( .A1(n6532), .A2(n7113), .ZN(n9794) );
  INV_X1 U6412 ( .A(n9780), .ZN(n9779) );
  INV_X1 U6413 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7925) );
  INV_X1 U6414 ( .A(n7705), .ZN(n7732) );
  INV_X1 U6415 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6604) );
  INV_X1 U6416 ( .A(n7694), .ZN(n9728) );
  INV_X2 U6417 ( .A(n8697), .ZN(P2_U3893) );
  OAI21_X1 U6418 ( .B1(n6174), .B2(n9839), .A(n6173), .ZN(P2_U3205) );
  INV_X1 U6419 ( .A(n9272), .ZN(P1_U3973) );
  INV_X1 U6420 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4860) );
  INV_X1 U6421 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4865) );
  OR2_X1 U6422 ( .A1(n4979), .A2(n4865), .ZN(n4872) );
  NAND2_X1 U6423 ( .A1(n5462), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4871) );
  AND2_X4 U6424 ( .A1(n8092), .A2(n4867), .ZN(n4938) );
  INV_X1 U6425 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4868) );
  OR2_X1 U6426 ( .A1(n4920), .A2(n4868), .ZN(n4869) );
  NAND2_X1 U6427 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4874) );
  OR2_X1 U6428 ( .A1(n4876), .A2(n4862), .ZN(n4877) );
  NAND2_X2 U6429 ( .A1(n4879), .A2(n4878), .ZN(n5672) );
  NAND2_X1 U6430 ( .A1(n4881), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4882) );
  INV_X1 U6431 ( .A(n5038), .ZN(n4883) );
  NAND2_X1 U6432 ( .A1(n4883), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4891) );
  AND2_X1 U6433 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U6434 ( .A1(n4973), .A2(n4884), .ZN(n4898) );
  NAND3_X1 U6435 ( .A1(n4907), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4885) );
  XNOR2_X1 U6436 ( .A(n4908), .B(SI_1_), .ZN(n4888) );
  XNOR2_X1 U6437 ( .A(n4888), .B(n4909), .ZN(n5700) );
  INV_X2 U6438 ( .A(n5091), .ZN(n5160) );
  NAND2_X1 U6439 ( .A1(n5160), .A2(n9276), .ZN(n4889) );
  INV_X1 U6440 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4892) );
  OR2_X1 U6441 ( .A1(n4979), .A2(n4892), .ZN(n4895) );
  INV_X1 U6442 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7121) );
  OR2_X1 U6443 ( .A1(n4939), .A2(n7121), .ZN(n4894) );
  INV_X1 U6444 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4893) );
  INV_X1 U6445 ( .A(SI_0_), .ZN(n4897) );
  INV_X1 U6446 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4896) );
  OAI21_X1 U6447 ( .B1(n4907), .B2(n4897), .A(n4896), .ZN(n4899) );
  AND2_X1 U6448 ( .A1(n4899), .A2(n4898), .ZN(n9733) );
  MUX2_X1 U6449 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9733), .S(n5091), .Z(n6943) );
  INV_X1 U6450 ( .A(n6942), .ZN(n6198) );
  NAND2_X1 U6451 ( .A1(n6198), .A2(n9770), .ZN(n4900) );
  NAND2_X1 U6452 ( .A1(n4938), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4906) );
  INV_X1 U6453 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9288) );
  OR2_X1 U6454 ( .A1(n4939), .A2(n9288), .ZN(n4905) );
  INV_X1 U6455 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n4901) );
  OR2_X1 U6456 ( .A1(n4979), .A2(n4901), .ZN(n4904) );
  INV_X1 U6457 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4902) );
  OR2_X1 U6458 ( .A1(n4920), .A2(n4902), .ZN(n4903) );
  XNOR2_X1 U6459 ( .A(n4929), .B(SI_2_), .ZN(n4927) );
  OAI21_X1 U6460 ( .B1(n4909), .B2(SI_1_), .A(n4908), .ZN(n4911) );
  NAND2_X1 U6461 ( .A1(n4909), .A2(SI_1_), .ZN(n4910) );
  NAND2_X1 U6462 ( .A1(n4911), .A2(n4910), .ZN(n4928) );
  XNOR2_X1 U6463 ( .A(n4927), .B(n4928), .ZN(n6590) );
  NAND2_X1 U6464 ( .A1(n4883), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6465 ( .A1(n4913), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n4916) );
  INV_X1 U6466 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6467 ( .A1(n4915), .A2(n4914), .ZN(n4933) );
  AND2_X1 U6468 ( .A1(n4916), .A2(n4933), .ZN(n9291) );
  NAND2_X1 U6469 ( .A1(n5160), .A2(n9291), .ZN(n4917) );
  NAND2_X1 U6470 ( .A1(n7305), .A2(n7259), .ZN(n5518) );
  INV_X1 U6471 ( .A(n5518), .ZN(n4919) );
  INV_X1 U6472 ( .A(n7305), .ZN(n9271) );
  OR2_X1 U6473 ( .A1(n4939), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4924) );
  INV_X1 U6474 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4921) );
  INV_X1 U6475 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6783) );
  OR2_X1 U6476 ( .A1(n4979), .A2(n6783), .ZN(n4922) );
  INV_X4 U6477 ( .A(n5038), .ZN(n5496) );
  NAND2_X1 U6478 ( .A1(n5496), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6479 ( .A1(n4928), .A2(n4927), .ZN(n4932) );
  INV_X1 U6480 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6481 ( .A1(n4930), .A2(SI_2_), .ZN(n4931) );
  NAND2_X1 U6482 ( .A1(n4932), .A2(n4931), .ZN(n4948) );
  MUX2_X1 U6483 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4973), .Z(n4949) );
  XNOR2_X1 U6484 ( .A(n4949), .B(SI_3_), .ZN(n4946) );
  XNOR2_X1 U6485 ( .A(n4948), .B(n4946), .ZN(n5735) );
  NAND2_X1 U6486 ( .A1(n4926), .A2(n5735), .ZN(n4936) );
  NAND2_X1 U6487 ( .A1(n4933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4934) );
  XNOR2_X1 U6488 ( .A(n4934), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U6489 ( .A1(n5160), .A2(n9304), .ZN(n4935) );
  AND2_X1 U6490 ( .A1(n9270), .A2(n7321), .ZN(n5621) );
  OAI22_X1 U6491 ( .A1(n7304), .A2(n5621), .B1(n7321), .B2(n9270), .ZN(n7333)
         );
  NAND2_X1 U6492 ( .A1(n4938), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6493 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n4960) );
  OAI21_X1 U6494 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n4960), .ZN(n7339) );
  OR2_X1 U6495 ( .A1(n4305), .A2(n7339), .ZN(n4941) );
  INV_X1 U6496 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7337) );
  INV_X1 U6497 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6498 ( .A1(n5496), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4958) );
  MUX2_X1 U6499 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4973), .Z(n4970) );
  INV_X1 U6500 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6501 ( .A1(n4948), .A2(n4947), .ZN(n4951) );
  NAND2_X1 U6502 ( .A1(n4949), .A2(SI_3_), .ZN(n4950) );
  NAND2_X1 U6503 ( .A1(n4951), .A2(n4950), .ZN(n4968) );
  XNOR2_X1 U6504 ( .A(n4967), .B(n4968), .ZN(n5747) );
  NAND2_X1 U6505 ( .A1(n4926), .A2(n5747), .ZN(n4957) );
  NAND2_X1 U6506 ( .A1(n4953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4954) );
  MUX2_X1 U6507 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4954), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n4955) );
  AND2_X1 U6508 ( .A1(n4952), .A2(n4955), .ZN(n9318) );
  NAND2_X1 U6509 ( .A1(n5160), .A2(n9318), .ZN(n4956) );
  NAND2_X1 U6510 ( .A1(n9269), .A2(n7340), .ZN(n5624) );
  NAND2_X1 U6511 ( .A1(n4938), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4966) );
  INV_X1 U6512 ( .A(n4960), .ZN(n4959) );
  NAND2_X1 U6513 ( .A1(n4959), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n4982) );
  INV_X1 U6514 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U6515 ( .A1(n4960), .A2(n7509), .ZN(n4961) );
  NAND2_X1 U6516 ( .A1(n4982), .A2(n4961), .ZN(n9755) );
  OR2_X1 U6517 ( .A1(n4305), .A2(n9755), .ZN(n4965) );
  INV_X1 U6518 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n4962) );
  OR2_X1 U6519 ( .A1(n4920), .A2(n4962), .ZN(n4964) );
  INV_X1 U6520 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9756) );
  OR2_X1 U6521 ( .A1(n4979), .A2(n9756), .ZN(n4963) );
  NAND4_X1 U6522 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n9268)
         );
  INV_X1 U6523 ( .A(n4967), .ZN(n4969) );
  NAND2_X1 U6524 ( .A1(n4969), .A2(n4968), .ZN(n4972) );
  NAND2_X1 U6525 ( .A1(n4970), .A2(SI_4_), .ZN(n4971) );
  MUX2_X1 U6526 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4973), .Z(n4992) );
  XNOR2_X1 U6527 ( .A(n4992), .B(SI_5_), .ZN(n4989) );
  XNOR2_X1 U6528 ( .A(n4991), .B(n4989), .ZN(n5766) );
  NAND2_X1 U6529 ( .A1(n5495), .A2(n5766), .ZN(n4977) );
  NAND2_X1 U6530 ( .A1(n5496), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6531 ( .A1(n4952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  XNOR2_X1 U6532 ( .A(n4974), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U6533 ( .A1(n5160), .A2(n6887), .ZN(n4975) );
  NAND2_X1 U6534 ( .A1(n9268), .A2(n7433), .ZN(n5625) );
  INV_X1 U6535 ( .A(n9268), .ZN(n7454) );
  INV_X1 U6536 ( .A(n7433), .ZN(n9758) );
  NAND2_X1 U6537 ( .A1(n4938), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4988) );
  INV_X1 U6538 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4978) );
  OR2_X1 U6539 ( .A1(n4979), .A2(n4978), .ZN(n4987) );
  INV_X1 U6540 ( .A(n4982), .ZN(n4980) );
  NAND2_X1 U6541 ( .A1(n4980), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5011) );
  INV_X1 U6542 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6543 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NAND2_X1 U6544 ( .A1(n5011), .A2(n4983), .ZN(n7459) );
  OR2_X1 U6545 ( .A1(n4939), .A2(n7459), .ZN(n4986) );
  INV_X1 U6546 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n4984) );
  OR2_X1 U6547 ( .A1(n4920), .A2(n4984), .ZN(n4985) );
  INV_X1 U6548 ( .A(n4989), .ZN(n4990) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6575) );
  INV_X1 U6550 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6615) );
  BUF_X4 U6551 ( .A(n4973), .Z(n6572) );
  MUX2_X1 U6552 ( .A(n6575), .B(n6615), .S(n6572), .Z(n5020) );
  XNOR2_X1 U6553 ( .A(n5020), .B(SI_6_), .ZN(n5018) );
  XNOR2_X1 U6554 ( .A(n5019), .B(n5018), .ZN(n6588) );
  NAND2_X1 U6555 ( .A1(n5496), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4995) );
  OR2_X1 U6556 ( .A1(n4993), .A2(n4862), .ZN(n5024) );
  XNOR2_X1 U6557 ( .A(n5024), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U6558 ( .A1(n5160), .A2(n6874), .ZN(n4994) );
  OAI211_X1 U6559 ( .C1(n6588), .C2(n5074), .A(n4995), .B(n4994), .ZN(n7458)
         );
  NAND2_X1 U6560 ( .A1(n7575), .A2(n7458), .ZN(n6466) );
  NAND2_X1 U6561 ( .A1(n7453), .A2(n6466), .ZN(n4996) );
  INV_X1 U6562 ( .A(n7575), .ZN(n9267) );
  NAND2_X1 U6563 ( .A1(n4996), .A2(n6465), .ZN(n5009) );
  NAND2_X1 U6564 ( .A1(n5507), .A2(n4999), .ZN(n5000) );
  INV_X1 U6565 ( .A(n5003), .ZN(n5001) );
  NAND2_X1 U6566 ( .A1(n5001), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n5004) );
  INV_X1 U6567 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5247) );
  MUX2_X1 U6568 ( .A(n5009), .B(n7754), .S(n5614), .Z(n5030) );
  NAND2_X1 U6569 ( .A1(n4938), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6570 ( .A1(n5011), .A2(n5010), .ZN(n5012) );
  NAND2_X1 U6571 ( .A1(n5031), .A2(n5012), .ZN(n9743) );
  OR2_X1 U6572 ( .A1(n4939), .A2(n9743), .ZN(n5016) );
  INV_X1 U6573 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9744) );
  OR2_X1 U6574 ( .A1(n4979), .A2(n9744), .ZN(n5015) );
  INV_X1 U6575 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5013) );
  OR2_X1 U6576 ( .A1(n5472), .A2(n5013), .ZN(n5014) );
  NAND4_X1 U6577 ( .A1(n5017), .A2(n5016), .A3(n5015), .A4(n5014), .ZN(n9266)
         );
  INV_X1 U6578 ( .A(n5020), .ZN(n5021) );
  NAND2_X1 U6579 ( .A1(n5021), .A2(SI_6_), .ZN(n5022) );
  MUX2_X1 U6580 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6572), .Z(n5042) );
  XNOR2_X1 U6581 ( .A(n5042), .B(SI_7_), .ZN(n5039) );
  XNOR2_X1 U6582 ( .A(n5041), .B(n5039), .ZN(n6577) );
  NAND2_X1 U6583 ( .A1(n5495), .A2(n6577), .ZN(n5029) );
  NAND2_X1 U6584 ( .A1(n5496), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U6585 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6586 ( .A1(n5024), .A2(n5023), .ZN(n5025) );
  NAND2_X1 U6587 ( .A1(n5025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5026) );
  XNOR2_X1 U6588 ( .A(n5026), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U6589 ( .A1(n5160), .A2(n6914), .ZN(n5027) );
  XNOR2_X1 U6590 ( .A(n9266), .B(n7767), .ZN(n7755) );
  NAND2_X1 U6591 ( .A1(n4938), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5037) );
  INV_X1 U6592 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7624) );
  OR2_X1 U6593 ( .A1(n4979), .A2(n7624), .ZN(n5036) );
  NAND2_X1 U6594 ( .A1(n5031), .A2(n7635), .ZN(n5032) );
  NAND2_X1 U6595 ( .A1(n5057), .A2(n5032), .ZN(n7634) );
  OR2_X1 U6596 ( .A1(n4305), .A2(n7634), .ZN(n5035) );
  INV_X1 U6597 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5033) );
  OR2_X1 U6598 ( .A1(n5472), .A2(n5033), .ZN(n5034) );
  INV_X1 U6599 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6600 ( .A1(n5042), .A2(SI_7_), .ZN(n5043) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6599) );
  MUX2_X1 U6602 ( .A(n6599), .B(n9977), .S(n6572), .Z(n5045) );
  INV_X1 U6603 ( .A(SI_8_), .ZN(n5044) );
  NAND2_X1 U6604 ( .A1(n5045), .A2(n5044), .ZN(n5063) );
  INV_X1 U6605 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6606 ( .A1(n5046), .A2(SI_8_), .ZN(n5047) );
  NAND2_X1 U6607 ( .A1(n5063), .A2(n5047), .ZN(n5049) );
  NAND2_X1 U6608 ( .A1(n5048), .A2(n5049), .ZN(n5050) );
  NAND2_X1 U6609 ( .A1(n5064), .A2(n5050), .ZN(n6596) );
  NAND2_X1 U6610 ( .A1(n5495), .A2(n6596), .ZN(n5054) );
  NAND2_X1 U6611 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6612 ( .A(n5052), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U6613 ( .A1(n5160), .A2(n6935), .ZN(n5053) );
  OAI211_X1 U6614 ( .C1(n5298), .C2(n9977), .A(n5054), .B(n5053), .ZN(n7639)
         );
  INV_X1 U6615 ( .A(n7639), .ZN(n9796) );
  NAND2_X1 U6616 ( .A1(n9265), .A2(n9796), .ZN(n7646) );
  NAND2_X1 U6617 ( .A1(n9266), .A2(n7767), .ZN(n5055) );
  AND2_X1 U6618 ( .A1(n7646), .A2(n5055), .ZN(n5516) );
  NAND2_X1 U6619 ( .A1(n7651), .A2(n7639), .ZN(n6470) );
  INV_X1 U6620 ( .A(n9266), .ZN(n7455) );
  INV_X1 U6621 ( .A(n7767), .ZN(n9747) );
  NAND2_X1 U6622 ( .A1(n7455), .A2(n9747), .ZN(n7615) );
  NAND2_X1 U6623 ( .A1(n6470), .A2(n7615), .ZN(n5513) );
  INV_X1 U6624 ( .A(n5513), .ZN(n7645) );
  MUX2_X1 U6625 ( .A(n5516), .B(n7645), .S(n5614), .Z(n5078) );
  INV_X1 U6626 ( .A(n6470), .ZN(n5076) );
  NAND2_X1 U6627 ( .A1(n5466), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5062) );
  OR2_X1 U6628 ( .A1(n5469), .A2(n4541), .ZN(n5061) );
  NAND2_X1 U6629 ( .A1(n5057), .A2(n5056), .ZN(n5058) );
  NAND2_X1 U6630 ( .A1(n5082), .A2(n5058), .ZN(n7863) );
  OR2_X1 U6631 ( .A1(n4939), .A2(n7863), .ZN(n5060) );
  INV_X1 U6632 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7655) );
  OR2_X1 U6633 ( .A1(n4979), .A2(n7655), .ZN(n5059) );
  MUX2_X1 U6634 ( .A(n6606), .B(n6604), .S(n6572), .Z(n5066) );
  INV_X1 U6635 ( .A(SI_9_), .ZN(n5065) );
  NAND2_X1 U6636 ( .A1(n5066), .A2(n5065), .ZN(n5089) );
  INV_X1 U6637 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6638 ( .A1(n5067), .A2(SI_9_), .ZN(n5068) );
  NAND2_X1 U6639 ( .A1(n5496), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6640 ( .A1(n4358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5071) );
  XNOR2_X1 U6641 ( .A(n5071), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U6642 ( .A1(n5160), .A2(n6898), .ZN(n5072) );
  OAI211_X1 U6643 ( .C1(n6605), .C2(n5074), .A(n5073), .B(n5072), .ZN(n7657)
         );
  INV_X1 U6644 ( .A(n7657), .ZN(n9805) );
  NAND2_X1 U6645 ( .A1(n9264), .A2(n9805), .ZN(n6472) );
  NAND2_X1 U6646 ( .A1(n6472), .A2(n7646), .ZN(n5075) );
  MUX2_X1 U6647 ( .A(n5076), .B(n5075), .S(n5614), .Z(n5077) );
  NAND2_X1 U6648 ( .A1(n7518), .A2(n7657), .ZN(n6473) );
  INV_X1 U6649 ( .A(n6472), .ZN(n5079) );
  AOI21_X1 U6650 ( .B1(n5213), .B2(n6473), .A(n5079), .ZN(n5117) );
  NAND2_X1 U6651 ( .A1(n4938), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5088) );
  INV_X1 U6652 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7525) );
  OR2_X1 U6653 ( .A1(n4979), .A2(n7525), .ZN(n5087) );
  INV_X1 U6654 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6655 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  NAND2_X1 U6656 ( .A1(n5095), .A2(n5083), .ZN(n9065) );
  OR2_X1 U6657 ( .A1(n4305), .A2(n9065), .ZN(n5086) );
  INV_X1 U6658 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6659 ( .A1(n5472), .A2(n5084), .ZN(n5085) );
  MUX2_X1 U6660 ( .A(n6608), .B(n6621), .S(n6572), .Z(n5104) );
  XNOR2_X1 U6661 ( .A(n5104), .B(SI_10_), .ZN(n5103) );
  XNOR2_X1 U6662 ( .A(n5102), .B(n5103), .ZN(n6607) );
  NAND2_X1 U6663 ( .A1(n6607), .A2(n5495), .ZN(n5094) );
  NOR2_X1 U6664 ( .A1(n4358), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6665 ( .A1(n5122), .A2(n4862), .ZN(n5112) );
  XNOR2_X1 U6666 ( .A(n5112), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6953) );
  INV_X1 U6667 ( .A(n6953), .ZN(n6609) );
  OAI22_X1 U6668 ( .A1(n5298), .A2(n6621), .B1(n6629), .B2(n6609), .ZN(n5092)
         );
  INV_X1 U6669 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6670 ( .A1(n7720), .A2(n9067), .ZN(n7716) );
  INV_X1 U6671 ( .A(n7716), .ZN(n5586) );
  INV_X1 U6672 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6954) );
  OR2_X1 U6673 ( .A1(n5469), .A2(n6954), .ZN(n5101) );
  NAND2_X1 U6674 ( .A1(n5095), .A2(n9993), .ZN(n5096) );
  NAND2_X1 U6675 ( .A1(n5129), .A2(n5096), .ZN(n9212) );
  OR2_X1 U6676 ( .A1(n4939), .A2(n9212), .ZN(n5100) );
  INV_X1 U6677 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5097) );
  OR2_X1 U6678 ( .A1(n5472), .A2(n5097), .ZN(n5099) );
  INV_X1 U6679 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7724) );
  OR2_X1 U6680 ( .A1(n4979), .A2(n7724), .ZN(n5098) );
  NAND4_X1 U6681 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n9262)
         );
  INV_X1 U6682 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6683 ( .A1(n5105), .A2(SI_10_), .ZN(n5106) );
  MUX2_X1 U6684 ( .A(n6618), .B(n6619), .S(n6572), .Z(n5109) );
  INV_X1 U6685 ( .A(SI_11_), .ZN(n5108) );
  NAND2_X1 U6686 ( .A1(n5109), .A2(n5108), .ZN(n5118) );
  INV_X1 U6687 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6688 ( .A1(n5110), .A2(SI_11_), .ZN(n5111) );
  NAND2_X1 U6689 ( .A1(n5118), .A2(n5111), .ZN(n5119) );
  XNOR2_X1 U6690 ( .A(n5120), .B(n5119), .ZN(n6613) );
  NAND2_X1 U6691 ( .A1(n6613), .A2(n5495), .ZN(n5116) );
  INV_X1 U6692 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U6693 ( .A1(n5112), .A2(n10062), .ZN(n5113) );
  NAND2_X1 U6694 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6695 ( .A(n5114), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7017) );
  AOI22_X1 U6696 ( .A1(n5496), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5160), .B2(
        n7017), .ZN(n5115) );
  OR2_X1 U6697 ( .A1(n6477), .A2(n9662), .ZN(n5588) );
  INV_X1 U6698 ( .A(n7720), .ZN(n9263) );
  NAND2_X1 U6699 ( .A1(n9263), .A2(n6475), .ZN(n5630) );
  OAI211_X1 U6700 ( .C1(n5117), .C2(n5586), .A(n5588), .B(n5630), .ZN(n5135)
         );
  NAND2_X1 U6701 ( .A1(n9662), .A2(n6477), .ZN(n5525) );
  MUX2_X1 U6702 ( .A(n6631), .B(n6633), .S(n6572), .Z(n5138) );
  XNOR2_X1 U6703 ( .A(n5138), .B(SI_12_), .ZN(n5137) );
  XNOR2_X1 U6704 ( .A(n5142), .B(n5137), .ZN(n6630) );
  NAND2_X1 U6705 ( .A1(n6630), .A2(n5495), .ZN(n5126) );
  NOR2_X1 U6706 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5121) );
  NAND2_X1 U6707 ( .A1(n5122), .A2(n5121), .ZN(n5143) );
  NAND2_X1 U6708 ( .A1(n5143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U6709 ( .A(n5123), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7237) );
  INV_X1 U6710 ( .A(n7237), .ZN(n7022) );
  OAI22_X1 U6711 ( .A1(n5298), .A2(n6633), .B1(n6629), .B2(n7022), .ZN(n5124)
         );
  INV_X1 U6712 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6713 ( .A1(n5466), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5134) );
  INV_X1 U6714 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7018) );
  OR2_X1 U6715 ( .A1(n5469), .A2(n7018), .ZN(n5133) );
  INV_X1 U6716 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6717 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  NAND2_X1 U6718 ( .A1(n5147), .A2(n5130), .ZN(n9118) );
  OR2_X1 U6719 ( .A1(n4939), .A2(n9118), .ZN(n5132) );
  INV_X1 U6720 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7849) );
  OR2_X1 U6721 ( .A1(n4979), .A2(n7849), .ZN(n5131) );
  NAND4_X1 U6722 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n9261)
         );
  NAND2_X1 U6723 ( .A1(n9124), .A2(n7721), .ZN(n5526) );
  NAND3_X1 U6724 ( .A1(n5135), .A2(n5525), .A3(n5526), .ZN(n5136) );
  NAND2_X1 U6725 ( .A1(n5136), .A2(n5589), .ZN(n5170) );
  INV_X1 U6726 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6727 ( .A1(n5139), .A2(SI_12_), .ZN(n5140) );
  MUX2_X1 U6728 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6572), .Z(n5156) );
  XNOR2_X1 U6729 ( .A(n5156), .B(SI_13_), .ZN(n5153) );
  XNOR2_X1 U6730 ( .A(n5155), .B(n5153), .ZN(n6634) );
  NAND2_X1 U6731 ( .A1(n6634), .A2(n5495), .ZN(n5146) );
  NAND2_X1 U6732 ( .A1(n5158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  XNOR2_X1 U6733 ( .A(n5144), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7380) );
  AOI22_X1 U6734 ( .A1(n5496), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5160), .B2(
        n7380), .ZN(n5145) );
  NAND2_X1 U6735 ( .A1(n4938), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6736 ( .A1(n5147), .A2(n9186), .ZN(n5148) );
  NAND2_X1 U6737 ( .A1(n5164), .A2(n5148), .ZN(n9185) );
  OR2_X1 U6738 ( .A1(n4305), .A2(n9185), .ZN(n5151) );
  INV_X1 U6739 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7872) );
  OR2_X1 U6740 ( .A1(n4979), .A2(n7872), .ZN(n5150) );
  INV_X1 U6741 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10004) );
  OR2_X1 U6742 ( .A1(n5472), .A2(n10004), .ZN(n5149) );
  NAND4_X1 U6743 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n9260)
         );
  NAND2_X1 U6744 ( .A1(n9190), .A2(n6482), .ZN(n5635) );
  NOR2_X1 U6745 ( .A1(n9190), .A2(n6482), .ZN(n5639) );
  INV_X1 U6746 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6747 ( .A1(n5156), .A2(SI_13_), .ZN(n5157) );
  MUX2_X1 U6748 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6572), .Z(n5175) );
  XNOR2_X1 U6749 ( .A(n5175), .B(SI_14_), .ZN(n5172) );
  XNOR2_X1 U6750 ( .A(n5174), .B(n5172), .ZN(n6701) );
  NAND2_X1 U6751 ( .A1(n6701), .A2(n5495), .ZN(n5162) );
  NAND2_X1 U6752 ( .A1(n5159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5197) );
  XNOR2_X1 U6753 ( .A(n5197), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7703) );
  AOI22_X1 U6754 ( .A1(n5496), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5160), .B2(
        n7703), .ZN(n5161) );
  INV_X1 U6755 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10041) );
  OR2_X1 U6756 ( .A1(n5469), .A2(n10041), .ZN(n5169) );
  NAND2_X1 U6757 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U6758 ( .A1(n5203), .A2(n5165), .ZN(n9043) );
  OR2_X1 U6759 ( .A1(n4305), .A2(n9043), .ZN(n5168) );
  INV_X1 U6760 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9715) );
  OR2_X1 U6761 ( .A1(n5472), .A2(n9715), .ZN(n5167) );
  INV_X1 U6762 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8069) );
  OR2_X1 U6763 ( .A1(n4979), .A2(n8069), .ZN(n5166) );
  NAND4_X1 U6764 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n9259)
         );
  INV_X1 U6765 ( .A(n9259), .ZN(n6484) );
  OR2_X1 U6766 ( .A1(n9045), .A2(n6484), .ZN(n9572) );
  NAND2_X1 U6767 ( .A1(n9045), .A2(n6484), .ZN(n5209) );
  NAND2_X1 U6768 ( .A1(n9572), .A2(n5209), .ZN(n8065) );
  AOI211_X1 U6769 ( .C1(n5170), .C2(n5635), .A(n5639), .B(n8065), .ZN(n5171)
         );
  INV_X1 U6770 ( .A(n5171), .ZN(n5211) );
  INV_X1 U6771 ( .A(n5172), .ZN(n5173) );
  NAND2_X1 U6772 ( .A1(n5175), .A2(SI_14_), .ZN(n5176) );
  NAND2_X1 U6773 ( .A1(n5177), .A2(n5176), .ZN(n5195) );
  MUX2_X1 U6774 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6572), .Z(n5193) );
  NOR2_X1 U6775 ( .A1(n5179), .A2(n5178), .ZN(n5181) );
  NAND2_X1 U6776 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  OAI21_X1 U6777 ( .B1(n5195), .B2(n5181), .A(n5180), .ZN(n5225) );
  MUX2_X1 U6778 ( .A(n6921), .B(n6922), .S(n6572), .Z(n5223) );
  XNOR2_X1 U6779 ( .A(n5223), .B(SI_16_), .ZN(n5182) );
  XNOR2_X1 U6780 ( .A(n5225), .B(n5182), .ZN(n6920) );
  NAND2_X1 U6781 ( .A1(n6920), .A2(n5495), .ZN(n5187) );
  NAND2_X1 U6782 ( .A1(n5183), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6783 ( .A(n5184), .B(n4590), .ZN(n7739) );
  OAI22_X1 U6784 ( .A1(n5298), .A2(n6922), .B1(n6629), .B2(n7739), .ZN(n5185)
         );
  INV_X1 U6785 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6786 ( .A1(n5466), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5192) );
  INV_X1 U6787 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9645) );
  OR2_X1 U6788 ( .A1(n5469), .A2(n9645), .ZN(n5191) );
  INV_X1 U6789 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5236) );
  XNOR2_X1 U6790 ( .A(n5238), .B(n5236), .ZN(n9558) );
  OR2_X1 U6791 ( .A1(n4939), .A2(n9558), .ZN(n5190) );
  INV_X1 U6792 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9559) );
  OR2_X1 U6793 ( .A1(n4979), .A2(n9559), .ZN(n5189) );
  NAND2_X1 U6794 ( .A1(n9644), .A2(n9236), .ZN(n9545) );
  INV_X1 U6795 ( .A(n9545), .ZN(n5594) );
  XNOR2_X1 U6796 ( .A(n5193), .B(SI_15_), .ZN(n5194) );
  XNOR2_X1 U6797 ( .A(n5195), .B(n5194), .ZN(n6764) );
  NAND2_X1 U6798 ( .A1(n6764), .A2(n5495), .ZN(n5202) );
  INV_X1 U6799 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6812) );
  INV_X1 U6800 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6801 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  NAND2_X1 U6802 ( .A1(n5198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5199) );
  XNOR2_X1 U6803 ( .A(n5199), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7705) );
  OAI22_X1 U6804 ( .A1(n5298), .A2(n6812), .B1(n6629), .B2(n7732), .ZN(n5200)
         );
  INV_X1 U6805 ( .A(n5200), .ZN(n5201) );
  NAND2_X1 U6806 ( .A1(n5466), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5208) );
  INV_X1 U6807 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9651) );
  OR2_X1 U6808 ( .A1(n5469), .A2(n9651), .ZN(n5207) );
  INV_X1 U6809 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U6810 ( .A1(n5203), .A2(n9240), .ZN(n5204) );
  NAND2_X1 U6811 ( .A1(n5238), .A2(n5204), .ZN(n9582) );
  OR2_X1 U6812 ( .A1(n4939), .A2(n9582), .ZN(n5206) );
  INV_X1 U6813 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9583) );
  OR2_X1 U6814 ( .A1(n4979), .A2(n9583), .ZN(n5205) );
  NAND2_X1 U6815 ( .A1(n9585), .A2(n9137), .ZN(n5592) );
  NAND2_X1 U6816 ( .A1(n5592), .A2(n5209), .ZN(n5644) );
  INV_X1 U6817 ( .A(n5643), .ZN(n5210) );
  INV_X1 U6818 ( .A(n6473), .ZN(n5212) );
  AND2_X1 U6819 ( .A1(n5525), .A2(n7716), .ZN(n5633) );
  NAND2_X1 U6820 ( .A1(n5589), .A2(n5588), .ZN(n5632) );
  INV_X1 U6821 ( .A(n5526), .ZN(n5636) );
  NOR2_X1 U6822 ( .A1(n5214), .A2(n5636), .ZN(n5216) );
  INV_X1 U6823 ( .A(n8065), .ZN(n5215) );
  OAI211_X1 U6824 ( .C1(n5216), .C2(n5639), .A(n5215), .B(n5635), .ZN(n5217)
         );
  OR2_X1 U6825 ( .A1(n9585), .A2(n9137), .ZN(n5642) );
  INV_X1 U6826 ( .A(n5592), .ZN(n5219) );
  INV_X1 U6827 ( .A(n5614), .ZN(n5549) );
  AND2_X1 U6828 ( .A1(n9648), .A2(n5549), .ZN(n5218) );
  AOI21_X1 U6829 ( .B1(n5643), .B2(n5219), .A(n5218), .ZN(n5221) );
  INV_X1 U6830 ( .A(n5221), .ZN(n5222) );
  NOR2_X1 U6831 ( .A1(n5226), .A2(SI_16_), .ZN(n5224) );
  NAND2_X1 U6832 ( .A1(n5226), .A2(SI_16_), .ZN(n5227) );
  MUX2_X1 U6833 ( .A(n7028), .B(n7030), .S(n6572), .Z(n5229) );
  NAND2_X1 U6834 ( .A1(n5229), .A2(n5228), .ZN(n5246) );
  INV_X1 U6835 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6836 ( .A1(n5230), .A2(SI_17_), .ZN(n5231) );
  NAND2_X1 U6837 ( .A1(n5246), .A2(n5231), .ZN(n5244) );
  XNOR2_X1 U6838 ( .A(n5245), .B(n5244), .ZN(n7027) );
  XNOR2_X1 U6839 ( .A(n5233), .B(n5232), .ZN(n9337) );
  OAI22_X1 U6840 ( .A1(n5298), .A2(n7030), .B1(n6629), .B2(n9337), .ZN(n5234)
         );
  NAND2_X1 U6841 ( .A1(n5466), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5243) );
  INV_X1 U6842 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9640) );
  OR2_X1 U6843 ( .A1(n5469), .A2(n9640), .ZN(n5242) );
  INV_X1 U6844 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5235) );
  OAI21_X1 U6845 ( .B1(n5238), .B2(n5236), .A(n5235), .ZN(n5239) );
  NAND2_X1 U6846 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n5237) );
  NAND2_X1 U6847 ( .A1(n5239), .A2(n5254), .ZN(n9538) );
  OR2_X1 U6848 ( .A1(n4939), .A2(n9538), .ZN(n5241) );
  INV_X1 U6849 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9539) );
  OR2_X1 U6850 ( .A1(n4979), .A2(n9539), .ZN(n5240) );
  OR2_X1 U6851 ( .A1(n9639), .A2(n9221), .ZN(n9518) );
  NAND2_X1 U6852 ( .A1(n9639), .A2(n9221), .ZN(n5308) );
  NAND2_X1 U6853 ( .A1(n9518), .A2(n5308), .ZN(n9534) );
  INV_X1 U6854 ( .A(n9518), .ZN(n5262) );
  MUX2_X1 U6855 ( .A(n7090), .B(n7065), .S(n6572), .Z(n5264) );
  XNOR2_X1 U6856 ( .A(n5264), .B(SI_18_), .ZN(n5263) );
  XNOR2_X1 U6857 ( .A(n5267), .B(n5263), .ZN(n7064) );
  NAND2_X1 U6858 ( .A1(n7064), .A2(n5495), .ZN(n5251) );
  XNOR2_X1 U6859 ( .A(n5248), .B(n5247), .ZN(n9341) );
  OAI22_X1 U6860 ( .A1(n5298), .A2(n7065), .B1(n6629), .B2(n9341), .ZN(n5249)
         );
  INV_X1 U6861 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6862 ( .A1(n4938), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5260) );
  INV_X1 U6863 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6864 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  NAND2_X1 U6865 ( .A1(n5301), .A2(n5255), .ZN(n9526) );
  OR2_X1 U6866 ( .A1(n4305), .A2(n9526), .ZN(n5259) );
  INV_X1 U6867 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6868 ( .A1(n5472), .A2(n5256), .ZN(n5258) );
  INV_X1 U6869 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9527) );
  OR2_X1 U6870 ( .A1(n4979), .A2(n9527), .ZN(n5257) );
  NAND4_X1 U6871 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n9256)
         );
  INV_X1 U6872 ( .A(n9256), .ZN(n6311) );
  OR2_X1 U6873 ( .A1(n9697), .A2(n6311), .ZN(n5648) );
  INV_X1 U6874 ( .A(n5648), .ZN(n5261) );
  INV_X1 U6875 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6876 ( .A1(n5265), .A2(SI_18_), .ZN(n5266) );
  MUX2_X1 U6877 ( .A(n7248), .B(n8145), .S(n6572), .Z(n5269) );
  NAND2_X1 U6878 ( .A1(n5269), .A2(n5268), .ZN(n5272) );
  INV_X1 U6879 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6880 ( .A1(n5270), .A2(SI_19_), .ZN(n5271) );
  NAND2_X1 U6881 ( .A1(n5272), .A2(n5271), .ZN(n5296) );
  MUX2_X1 U6882 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6572), .Z(n5285) );
  INV_X1 U6883 ( .A(n5285), .ZN(n5273) );
  MUX2_X1 U6884 ( .A(n10074), .B(n7421), .S(n6572), .Z(n5322) );
  XNOR2_X1 U6885 ( .A(n5322), .B(SI_21_), .ZN(n5274) );
  XNOR2_X1 U6886 ( .A(n5321), .B(n5274), .ZN(n7405) );
  NAND2_X1 U6887 ( .A1(n7405), .A2(n5495), .ZN(n5276) );
  NAND2_X1 U6888 ( .A1(n5496), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6889 ( .A1(n4938), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5283) );
  INV_X1 U6890 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6891 ( .A1(n5472), .A2(n5277), .ZN(n5282) );
  INV_X1 U6892 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5300) );
  INV_X1 U6893 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9178) );
  INV_X1 U6894 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6895 ( .A1(n5291), .A2(n5278), .ZN(n5279) );
  NAND2_X1 U6896 ( .A1(n5334), .A2(n5279), .ZN(n9482) );
  OR2_X1 U6897 ( .A1(n4305), .A2(n9482), .ZN(n5281) );
  INV_X1 U6898 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9483) );
  OR2_X1 U6899 ( .A1(n4979), .A2(n9483), .ZN(n5280) );
  NAND2_X1 U6900 ( .A1(n9618), .A2(n9195), .ZN(n5511) );
  XNOR2_X1 U6901 ( .A(n5285), .B(n5284), .ZN(n5286) );
  XNOR2_X1 U6902 ( .A(n5287), .B(n5286), .ZN(n7353) );
  NAND2_X1 U6903 ( .A1(n7353), .A2(n5495), .ZN(n5289) );
  NAND2_X1 U6904 ( .A1(n5496), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6905 ( .A1(n4938), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6906 ( .A1(n5303), .A2(n9178), .ZN(n5290) );
  NAND2_X1 U6907 ( .A1(n5291), .A2(n5290), .ZN(n9499) );
  OR2_X1 U6908 ( .A1(n4939), .A2(n9499), .ZN(n5294) );
  INV_X1 U6909 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9688) );
  OR2_X1 U6910 ( .A1(n5472), .A2(n9688), .ZN(n5293) );
  INV_X1 U6911 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10060) );
  OR2_X1 U6912 ( .A1(n4979), .A2(n10060), .ZN(n5292) );
  NAND4_X1 U6913 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n9254)
         );
  INV_X1 U6914 ( .A(n9254), .ZN(n6317) );
  NAND2_X1 U6915 ( .A1(n9625), .A2(n6317), .ZN(n5512) );
  AND2_X1 U6916 ( .A1(n5511), .A2(n5512), .ZN(n6510) );
  OAI22_X1 U6917 ( .A1(n5298), .A2(n8145), .B1(n5620), .B2(n6629), .ZN(n5299)
         );
  NAND2_X1 U6918 ( .A1(n5466), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5307) );
  INV_X1 U6919 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9631) );
  OR2_X1 U6920 ( .A1(n5469), .A2(n9631), .ZN(n5306) );
  INV_X1 U6921 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9507) );
  OR2_X1 U6922 ( .A1(n4979), .A2(n9507), .ZN(n5305) );
  NAND2_X1 U6923 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NAND2_X1 U6924 ( .A1(n5303), .A2(n5302), .ZN(n9506) );
  OR2_X1 U6925 ( .A1(n4305), .A2(n9506), .ZN(n5304) );
  NAND2_X1 U6926 ( .A1(n9630), .A2(n9223), .ZN(n5652) );
  NAND2_X1 U6927 ( .A1(n9697), .A2(n6311), .ZN(n5597) );
  NAND4_X1 U6928 ( .A1(n6510), .A2(n5549), .A3(n5652), .A4(n5597), .ZN(n5319)
         );
  NAND2_X1 U6929 ( .A1(n5597), .A2(n5308), .ZN(n5649) );
  NAND2_X1 U6930 ( .A1(n6511), .A2(n9475), .ZN(n5574) );
  OR2_X1 U6931 ( .A1(n9630), .A2(n9223), .ZN(n5647) );
  INV_X1 U6932 ( .A(n5647), .ZN(n5309) );
  NOR4_X1 U6933 ( .A1(n5574), .A2(n5261), .A3(n5309), .A4(n5549), .ZN(n5310)
         );
  OAI21_X1 U6934 ( .B1(n5311), .B2(n5649), .A(n5310), .ZN(n5318) );
  INV_X1 U6935 ( .A(n6511), .ZN(n5312) );
  NOR2_X1 U6936 ( .A1(n6510), .A2(n5312), .ZN(n5563) );
  NAND2_X1 U6937 ( .A1(n5563), .A2(n5549), .ZN(n5316) );
  NAND3_X1 U6938 ( .A1(n6510), .A2(n5652), .A3(n5614), .ZN(n5315) );
  NAND4_X1 U6939 ( .A1(n6511), .A2(n5549), .A3(n9475), .A4(n5647), .ZN(n5314)
         );
  NAND3_X1 U6940 ( .A1(n5574), .A2(n5511), .A3(n5614), .ZN(n5313) );
  NAND4_X1 U6941 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n5317)
         );
  OAI211_X1 U6942 ( .C1(n5320), .C2(n5319), .A(n5318), .B(n5317), .ZN(n5360)
         );
  NAND2_X1 U6943 ( .A1(n5323), .A2(SI_21_), .ZN(n5324) );
  MUX2_X1 U6944 ( .A(n7586), .B(n7583), .S(n6572), .Z(n5327) );
  INV_X1 U6945 ( .A(SI_22_), .ZN(n5326) );
  NAND2_X1 U6946 ( .A1(n5327), .A2(n5326), .ZN(n5340) );
  INV_X1 U6947 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6948 ( .A1(n5328), .A2(SI_22_), .ZN(n5329) );
  NAND2_X1 U6949 ( .A1(n5340), .A2(n5329), .ZN(n5341) );
  XNOR2_X1 U6950 ( .A(n5342), .B(n5341), .ZN(n7581) );
  NAND2_X1 U6951 ( .A1(n7581), .A2(n5495), .ZN(n5331) );
  NAND2_X1 U6952 ( .A1(n5496), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6953 ( .A1(n4938), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5339) );
  INV_X1 U6954 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10006) );
  OR2_X1 U6955 ( .A1(n5472), .A2(n10006), .ZN(n5338) );
  INV_X1 U6956 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6957 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U6958 ( .A1(n5353), .A2(n5335), .ZN(n9471) );
  OR2_X1 U6959 ( .A1(n4305), .A2(n9471), .ZN(n5337) );
  INV_X1 U6960 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9462) );
  OR2_X1 U6961 ( .A1(n4979), .A2(n9462), .ZN(n5336) );
  NAND2_X1 U6962 ( .A1(n9614), .A2(n9109), .ZN(n5359) );
  MUX2_X1 U6963 ( .A(n7693), .B(n10051), .S(n6572), .Z(n5344) );
  INV_X1 U6964 ( .A(SI_23_), .ZN(n5343) );
  NAND2_X1 U6965 ( .A1(n5344), .A2(n5343), .ZN(n5364) );
  INV_X1 U6966 ( .A(n5344), .ZN(n5345) );
  NAND2_X1 U6967 ( .A1(n5345), .A2(SI_23_), .ZN(n5346) );
  OR2_X1 U6968 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6969 ( .A1(n5365), .A2(n5349), .ZN(n7695) );
  NAND2_X1 U6970 ( .A1(n7695), .A2(n5495), .ZN(n5351) );
  NAND2_X1 U6971 ( .A1(n5496), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5350) );
  INV_X1 U6972 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6973 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U6974 ( .A1(n5374), .A2(n5354), .ZN(n9453) );
  NAND2_X1 U6975 ( .A1(n5465), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5355) );
  OAI21_X1 U6976 ( .B1(n9453), .B2(n4939), .A(n5355), .ZN(n5358) );
  INV_X1 U6977 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U6978 ( .A1(n5466), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5356) );
  OAI21_X1 U6979 ( .B1(n5469), .B2(n9610), .A(n5356), .ZN(n5357) );
  NAND2_X1 U6980 ( .A1(n9609), .A2(n6494), .ZN(n6514) );
  NAND2_X1 U6981 ( .A1(n6514), .A2(n5359), .ZN(n5562) );
  AOI22_X1 U6982 ( .A1(n5360), .A2(n9466), .B1(n5562), .B2(n5614), .ZN(n5363)
         );
  NOR2_X1 U6983 ( .A1(n9609), .A2(n6494), .ZN(n5557) );
  INV_X1 U6984 ( .A(n6513), .ZN(n5361) );
  NOR2_X1 U6985 ( .A1(n5557), .A2(n5361), .ZN(n5362) );
  OAI22_X1 U6986 ( .A1(n5363), .A2(n5557), .B1(n5362), .B2(n5614), .ZN(n5380)
         );
  INV_X1 U6987 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7802) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7816) );
  MUX2_X1 U6989 ( .A(n7802), .B(n7816), .S(n6572), .Z(n5367) );
  INV_X1 U6990 ( .A(SI_24_), .ZN(n5366) );
  NAND2_X1 U6991 ( .A1(n5367), .A2(n5366), .ZN(n5385) );
  INV_X1 U6992 ( .A(n5367), .ZN(n5368) );
  NAND2_X1 U6993 ( .A1(n5368), .A2(SI_24_), .ZN(n5369) );
  XNOR2_X1 U6994 ( .A(n5384), .B(n5383), .ZN(n7801) );
  NAND2_X1 U6995 ( .A1(n7801), .A2(n5495), .ZN(n5371) );
  NAND2_X1 U6996 ( .A1(n5496), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5370) );
  INV_X1 U6997 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9439) );
  INV_X1 U6998 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6999 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U7000 ( .A1(n5406), .A2(n5375), .ZN(n9438) );
  OR2_X1 U7001 ( .A1(n9438), .A2(n4305), .ZN(n5377) );
  AOI22_X1 U7002 ( .A1(n4938), .A2(P1_REG1_REG_24__SCAN_IN), .B1(n5466), .B2(
        P1_REG0_REG_24__SCAN_IN), .ZN(n5376) );
  INV_X1 U7003 ( .A(n9250), .ZN(n5378) );
  NAND2_X1 U7004 ( .A1(n9678), .A2(n5378), .ZN(n5566) );
  NAND2_X1 U7005 ( .A1(n6515), .A2(n5566), .ZN(n9430) );
  INV_X1 U7006 ( .A(n9430), .ZN(n9436) );
  MUX2_X1 U7007 ( .A(n6515), .B(n5566), .S(n5614), .Z(n5381) );
  MUX2_X1 U7008 ( .A(n9991), .B(n7925), .S(n6572), .Z(n5387) );
  INV_X1 U7009 ( .A(SI_25_), .ZN(n5386) );
  NAND2_X1 U7010 ( .A1(n5387), .A2(n5386), .ZN(n5397) );
  INV_X1 U7011 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U7012 ( .A1(n5388), .A2(SI_25_), .ZN(n5389) );
  XNOR2_X1 U7013 ( .A(n5396), .B(n5395), .ZN(n7878) );
  NAND2_X1 U7014 ( .A1(n7878), .A2(n5495), .ZN(n5391) );
  NAND2_X1 U7015 ( .A1(n5496), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U7016 ( .A(n5406), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9424) );
  INV_X1 U7017 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U7018 ( .A1(n5466), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U7019 ( .A1(n5465), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5392) );
  OAI211_X1 U7020 ( .C1(n5469), .C2(n9601), .A(n5393), .B(n5392), .ZN(n5394)
         );
  NAND2_X1 U7021 ( .A1(n5396), .A2(n5395), .ZN(n5398) );
  NAND2_X1 U7022 ( .A1(n5398), .A2(n5397), .ZN(n5415) );
  INV_X1 U7023 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7980) );
  INV_X1 U7024 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8024) );
  MUX2_X1 U7025 ( .A(n7980), .B(n8024), .S(n6572), .Z(n5400) );
  INV_X1 U7026 ( .A(SI_26_), .ZN(n5399) );
  NAND2_X1 U7027 ( .A1(n5400), .A2(n5399), .ZN(n5416) );
  INV_X1 U7028 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U7029 ( .A1(n5401), .A2(SI_26_), .ZN(n5402) );
  XNOR2_X1 U7030 ( .A(n5415), .B(n5414), .ZN(n7979) );
  NAND2_X1 U7031 ( .A1(n7979), .A2(n5495), .ZN(n5404) );
  NAND2_X1 U7032 ( .A1(n5496), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5403) );
  INV_X1 U7033 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9131) );
  INV_X1 U7034 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10036) );
  OAI21_X1 U7035 ( .B1(n5406), .B2(n9131), .A(n10036), .ZN(n5407) );
  NAND2_X1 U7036 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5405) );
  NAND2_X1 U7037 ( .A1(n9411), .A2(n5462), .ZN(n5413) );
  INV_X1 U7038 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U7039 ( .A1(n5466), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U7040 ( .A1(n4938), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5408) );
  OAI211_X1 U7041 ( .C1(n5410), .C2(n4979), .A(n5409), .B(n5408), .ZN(n5411)
         );
  INV_X1 U7042 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U7043 ( .A1(n9669), .A2(n5509), .ZN(n6517) );
  NAND2_X1 U7044 ( .A1(n9600), .A2(n9159), .ZN(n5510) );
  INV_X1 U7045 ( .A(n5510), .ZN(n5567) );
  AOI211_X1 U7046 ( .C1(n5446), .C2(n6516), .A(n4808), .B(n5567), .ZN(n5434)
         );
  NOR2_X1 U7047 ( .A1(n9669), .A2(n5509), .ZN(n5554) );
  INV_X1 U7048 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8087) );
  INV_X1 U7049 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8162) );
  MUX2_X1 U7050 ( .A(n8087), .B(n8162), .S(n6572), .Z(n5418) );
  INV_X1 U7051 ( .A(SI_27_), .ZN(n5417) );
  NAND2_X1 U7052 ( .A1(n5418), .A2(n5417), .ZN(n5435) );
  INV_X1 U7053 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U7054 ( .A1(n5419), .A2(SI_27_), .ZN(n5420) );
  OR2_X1 U7055 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  NAND2_X1 U7056 ( .A1(n5436), .A2(n5423), .ZN(n8086) );
  NAND2_X1 U7057 ( .A1(n8086), .A2(n5495), .ZN(n5425) );
  NAND2_X1 U7058 ( .A1(n5496), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5424) );
  INV_X1 U7059 ( .A(n5427), .ZN(n5426) );
  NAND2_X1 U7060 ( .A1(n5426), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5440) );
  INV_X1 U7061 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U7062 ( .A1(n5427), .A2(n9978), .ZN(n5428) );
  NAND2_X1 U7063 ( .A1(n5440), .A2(n5428), .ZN(n6438) );
  OR2_X1 U7064 ( .A1(n6438), .A2(n4305), .ZN(n5433) );
  INV_X1 U7065 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7066 ( .A1(n5465), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7067 ( .A1(n5466), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5429) );
  OAI211_X1 U7068 ( .C1(n5469), .C2(n6534), .A(n5430), .B(n5429), .ZN(n5431)
         );
  INV_X1 U7069 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7070 ( .A1(n6525), .A2(n8105), .ZN(n8099) );
  INV_X1 U7071 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6064) );
  INV_X1 U7072 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U7073 ( .A(n6064), .B(n9730), .S(n6572), .Z(n5453) );
  XNOR2_X1 U7074 ( .A(n5453), .B(SI_28_), .ZN(n5450) );
  NAND2_X1 U7075 ( .A1(n8088), .A2(n5495), .ZN(n5438) );
  NAND2_X1 U7076 ( .A1(n5496), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5437) );
  INV_X1 U7077 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7078 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  INV_X1 U7079 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7080 ( .A1(n5465), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7081 ( .A1(n5466), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5442) );
  OAI211_X1 U7082 ( .C1(n5469), .C2(n5444), .A(n5443), .B(n5442), .ZN(n5445)
         );
  AOI21_X1 U7083 ( .B1(n9379), .B2(n5462), .A(n5445), .ZN(n9090) );
  AOI211_X1 U7084 ( .C1(n5446), .C2(n5510), .A(n4812), .B(n5554), .ZN(n5447)
         );
  NAND2_X1 U7085 ( .A1(n9380), .A2(n9090), .ZN(n5508) );
  AND2_X1 U7086 ( .A1(n5508), .A2(n8099), .ZN(n5553) );
  INV_X1 U7087 ( .A(n8119), .ZN(n5448) );
  INV_X1 U7088 ( .A(n5508), .ZN(n5464) );
  NAND2_X1 U7089 ( .A1(n5451), .A2(n5450), .ZN(n5455) );
  INV_X1 U7090 ( .A(SI_28_), .ZN(n5452) );
  NAND2_X1 U7091 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  INV_X1 U7092 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9032) );
  INV_X1 U7093 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10021) );
  MUX2_X1 U7094 ( .A(n9032), .B(n10021), .S(n6572), .Z(n5473) );
  NAND2_X1 U7095 ( .A1(n9030), .A2(n5495), .ZN(n5457) );
  NAND2_X1 U7096 ( .A1(n5496), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5456) );
  INV_X1 U7097 ( .A(n5458), .ZN(n8129) );
  INV_X1 U7098 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U7099 ( .A1(n5466), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7100 ( .A1(n5465), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5459) );
  OAI211_X1 U7101 ( .C1(n5469), .C2(n8138), .A(n5460), .B(n5459), .ZN(n5461)
         );
  AOI21_X1 U7102 ( .B1(n8129), .B2(n5462), .A(n5461), .ZN(n8103) );
  NAND2_X1 U7103 ( .A1(n5463), .A2(n8103), .ZN(n5600) );
  AOI21_X1 U7104 ( .B1(n5464), .B2(n5614), .A(n8121), .ZN(n5486) );
  INV_X1 U7105 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U7106 ( .A1(n5465), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7107 ( .A1(n5466), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U7108 ( .C1(n5469), .C2(n8159), .A(n5468), .B(n5467), .ZN(n9246)
         );
  INV_X1 U7109 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U7110 ( .A1(n4938), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5471) );
  INV_X1 U7111 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9368) );
  OR2_X1 U7112 ( .A1(n4979), .A2(n9368), .ZN(n5470) );
  OAI211_X1 U7113 ( .C1(n5472), .C2(n6457), .A(n5471), .B(n5470), .ZN(n6699)
         );
  AND3_X1 U7114 ( .A1(n9246), .A2(n6699), .A3(n5549), .ZN(n5501) );
  AOI22_X1 U7115 ( .A1(n5578), .A2(n5614), .B1(n5600), .B2(n5501), .ZN(n5485)
         );
  INV_X1 U7116 ( .A(SI_29_), .ZN(n5476) );
  INV_X1 U7117 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10033) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8299) );
  MUX2_X1 U7119 ( .A(n10033), .B(n8299), .S(n4907), .Z(n5479) );
  INV_X1 U7120 ( .A(SI_30_), .ZN(n5478) );
  NAND2_X1 U7121 ( .A1(n5479), .A2(n5478), .ZN(n5488) );
  INV_X1 U7122 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U7123 ( .A1(n5480), .A2(SI_30_), .ZN(n5481) );
  NAND2_X1 U7124 ( .A1(n5488), .A2(n5481), .ZN(n5489) );
  NAND2_X1 U7125 ( .A1(n8298), .A2(n5495), .ZN(n5483) );
  NAND2_X1 U7126 ( .A1(n5496), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5482) );
  NAND3_X1 U7127 ( .A1(n9373), .A2(n5549), .A3(n5600), .ZN(n5484) );
  AOI22_X1 U7128 ( .A1(n5487), .A2(n5486), .B1(n5485), .B2(n5484), .ZN(n5506)
         );
  INV_X1 U7129 ( .A(n9246), .ZN(n5539) );
  INV_X1 U7130 ( .A(n6699), .ZN(n5542) );
  OAI21_X1 U7131 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5494) );
  INV_X1 U7132 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5491) );
  INV_X1 U7133 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9026) );
  MUX2_X1 U7134 ( .A(n5491), .B(n9026), .S(n4907), .Z(n5492) );
  XNOR2_X1 U7135 ( .A(n5492), .B(SI_31_), .ZN(n5493) );
  XNOR2_X1 U7136 ( .A(n5494), .B(n5493), .ZN(n9022) );
  NAND2_X1 U7137 ( .A1(n9022), .A2(n5495), .ZN(n5498) );
  NAND2_X1 U7138 ( .A1(n5496), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5497) );
  OAI21_X1 U7139 ( .B1(n5604), .B2(n5542), .A(n9370), .ZN(n5505) );
  AOI21_X1 U7140 ( .B1(n5540), .B2(n5614), .A(n6699), .ZN(n5503) );
  NAND3_X1 U7141 ( .A1(n5539), .A2(n6699), .A3(n5614), .ZN(n5499) );
  NAND2_X1 U7142 ( .A1(n5540), .A2(n5499), .ZN(n5500) );
  OAI21_X1 U7143 ( .B1(n5540), .B2(n5501), .A(n5500), .ZN(n5502) );
  OAI21_X1 U7144 ( .B1(n9370), .B2(n5503), .A(n5502), .ZN(n5504) );
  AOI21_X1 U7145 ( .B1(n5506), .B2(n5505), .A(n5504), .ZN(n5610) );
  OR2_X1 U7146 ( .A1(n9370), .A2(n5542), .ZN(n5657) );
  NAND2_X1 U7147 ( .A1(n5556), .A2(n8099), .ZN(n8094) );
  NAND2_X1 U7148 ( .A1(n8119), .A2(n5508), .ZN(n8101) );
  XNOR2_X1 U7149 ( .A(n9669), .B(n5509), .ZN(n9403) );
  XNOR2_X1 U7150 ( .A(n9609), .B(n6494), .ZN(n9447) );
  NAND2_X1 U7151 ( .A1(n6511), .A2(n5511), .ZN(n9479) );
  INV_X1 U7152 ( .A(n9479), .ZN(n5534) );
  NAND2_X1 U7153 ( .A1(n9475), .A2(n5512), .ZN(n9495) );
  INV_X1 U7154 ( .A(n9534), .ZN(n9544) );
  NAND2_X1 U7155 ( .A1(n5648), .A2(n5597), .ZN(n9519) );
  INV_X1 U7156 ( .A(n9519), .ZN(n9523) );
  NAND2_X1 U7157 ( .A1(n5642), .A2(n5592), .ZN(n9573) );
  INV_X1 U7158 ( .A(n9573), .ZN(n5529) );
  NAND2_X1 U7159 ( .A1(n5513), .A2(n7646), .ZN(n5514) );
  NAND2_X1 U7160 ( .A1(n5514), .A2(n6473), .ZN(n5515) );
  NAND2_X1 U7161 ( .A1(n5515), .A2(n6472), .ZN(n5583) );
  AND2_X1 U7162 ( .A1(n5583), .A2(n6466), .ZN(n5581) );
  NAND3_X1 U7163 ( .A1(n5516), .A2(n6472), .A3(n6465), .ZN(n5582) );
  INV_X1 U7164 ( .A(n5582), .ZN(n5524) );
  XNOR2_X1 U7165 ( .A(n9268), .B(n7433), .ZN(n7425) );
  NOR2_X1 U7166 ( .A1(n7425), .A2(n7334), .ZN(n5523) );
  AND2_X1 U7167 ( .A1(n5517), .A2(n7125), .ZN(n5622) );
  NOR2_X1 U7168 ( .A1(n7094), .A2(n5622), .ZN(n6990) );
  INV_X1 U7169 ( .A(n7251), .ZN(n5520) );
  NAND4_X1 U7170 ( .A1(n6990), .A2(n5520), .A3(n7419), .A4(n5519), .ZN(n5521)
         );
  NOR2_X1 U7171 ( .A1(n5521), .A2(n7303), .ZN(n5522) );
  NAND2_X1 U7172 ( .A1(n7716), .A2(n5630), .ZN(n7523) );
  INV_X1 U7173 ( .A(n7523), .ZN(n5584) );
  NAND2_X1 U7174 ( .A1(n5588), .A2(n5525), .ZN(n7712) );
  INV_X1 U7175 ( .A(n7712), .ZN(n7715) );
  NAND4_X1 U7176 ( .A1(n4830), .A2(n5584), .A3(n7715), .A4(n7773), .ZN(n5527)
         );
  NOR2_X1 U7177 ( .A1(n5527), .A2(n8065), .ZN(n5528) );
  XNOR2_X1 U7178 ( .A(n9190), .B(n6482), .ZN(n5590) );
  INV_X1 U7179 ( .A(n5590), .ZN(n7870) );
  NAND3_X1 U7180 ( .A1(n5529), .A2(n5528), .A3(n7870), .ZN(n5530) );
  NAND2_X1 U7181 ( .A1(n5643), .A2(n9545), .ZN(n9553) );
  NOR2_X1 U7182 ( .A1(n5530), .A2(n9553), .ZN(n5531) );
  NAND4_X1 U7183 ( .A1(n9510), .A2(n9544), .A3(n9523), .A4(n5531), .ZN(n5532)
         );
  NOR2_X1 U7184 ( .A1(n9495), .A2(n5532), .ZN(n5533) );
  NAND3_X1 U7185 ( .A1(n9466), .A2(n5534), .A3(n5533), .ZN(n5535) );
  NOR2_X1 U7186 ( .A1(n9447), .A2(n5535), .ZN(n5536) );
  NAND3_X1 U7187 ( .A1(n9418), .A2(n9436), .A3(n5536), .ZN(n5537) );
  NOR2_X1 U7188 ( .A1(n8121), .A2(n5538), .ZN(n5541) );
  NAND2_X1 U7189 ( .A1(n5540), .A2(n5539), .ZN(n5601) );
  NAND3_X1 U7190 ( .A1(n5657), .A2(n5541), .A3(n5601), .ZN(n5544) );
  NAND2_X1 U7191 ( .A1(n9370), .A2(n5542), .ZN(n5615) );
  INV_X1 U7192 ( .A(n5604), .ZN(n5543) );
  NAND2_X1 U7193 ( .A1(n5615), .A2(n5543), .ZN(n5658) );
  OAI21_X1 U7194 ( .B1(n5610), .B2(n7419), .A(n5607), .ZN(n5552) );
  NAND2_X1 U7195 ( .A1(n5546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5548) );
  INV_X1 U7196 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5547) );
  AOI21_X1 U7197 ( .B1(n5549), .B2(n5545), .A(n7402), .ZN(n5550) );
  INV_X1 U7198 ( .A(n5550), .ZN(n5551) );
  AOI21_X1 U7199 ( .B1(n5552), .B2(n5619), .A(n5551), .ZN(n5609) );
  INV_X1 U7200 ( .A(n5553), .ZN(n5571) );
  INV_X1 U7201 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7202 ( .A1(n5556), .A2(n5555), .ZN(n5572) );
  INV_X1 U7203 ( .A(n6514), .ZN(n5559) );
  INV_X1 U7204 ( .A(n5557), .ZN(n5558) );
  OAI211_X1 U7205 ( .C1(n5559), .C2(n6513), .A(n6515), .B(n5558), .ZN(n5560)
         );
  NAND2_X1 U7206 ( .A1(n5560), .A2(n5566), .ZN(n5561) );
  AND2_X1 U7207 ( .A1(n5561), .A2(n6516), .ZN(n5573) );
  INV_X1 U7208 ( .A(n5562), .ZN(n5565) );
  INV_X1 U7209 ( .A(n5563), .ZN(n5564) );
  NAND3_X1 U7210 ( .A1(n5566), .A2(n5565), .A3(n5564), .ZN(n5568) );
  AOI21_X1 U7211 ( .B1(n5573), .B2(n5568), .A(n5567), .ZN(n5569) );
  NOR2_X1 U7212 ( .A1(n5572), .A2(n5569), .ZN(n5570) );
  NOR2_X1 U7213 ( .A1(n5571), .A2(n5570), .ZN(n5653) );
  INV_X1 U7214 ( .A(n5653), .ZN(n5579) );
  INV_X1 U7215 ( .A(n5572), .ZN(n5577) );
  INV_X1 U7216 ( .A(n5573), .ZN(n5575) );
  OAI21_X1 U7217 ( .B1(n5575), .B2(n5574), .A(n6517), .ZN(n5576) );
  INV_X1 U7218 ( .A(n5580), .ZN(n5656) );
  NAND2_X1 U7219 ( .A1(n5583), .A2(n5582), .ZN(n7514) );
  AND2_X1 U7220 ( .A1(n7514), .A2(n5584), .ZN(n5585) );
  NAND2_X1 U7221 ( .A1(n7515), .A2(n5585), .ZN(n7717) );
  NOR2_X1 U7222 ( .A1(n7712), .A2(n5586), .ZN(n5587) );
  NAND2_X1 U7223 ( .A1(n7717), .A2(n5587), .ZN(n7714) );
  NAND2_X1 U7224 ( .A1(n7714), .A2(n5588), .ZN(n7774) );
  NAND2_X1 U7225 ( .A1(n7774), .A2(n7773), .ZN(n7772) );
  INV_X1 U7226 ( .A(n9572), .ZN(n5640) );
  NOR2_X1 U7227 ( .A1(n9573), .A2(n5640), .ZN(n5591) );
  NAND2_X1 U7228 ( .A1(n8059), .A2(n5591), .ZN(n5593) );
  INV_X1 U7229 ( .A(n9553), .ZN(n9563) );
  NOR2_X1 U7230 ( .A1(n9534), .A2(n5594), .ZN(n5595) );
  NOR2_X1 U7231 ( .A1(n9519), .A2(n5262), .ZN(n5596) );
  NAND2_X1 U7232 ( .A1(n5598), .A2(n5597), .ZN(n9511) );
  INV_X1 U7233 ( .A(n6509), .ZN(n5599) );
  NAND3_X1 U7234 ( .A1(n5653), .A2(n5599), .A3(n6517), .ZN(n5602) );
  NAND2_X1 U7235 ( .A1(n5601), .A2(n5600), .ZN(n5654) );
  AOI21_X1 U7236 ( .B1(n5656), .B2(n5602), .A(n5654), .ZN(n5603) );
  AOI21_X1 U7237 ( .B1(n5604), .B2(n6699), .A(n5603), .ZN(n5606) );
  OAI21_X1 U7238 ( .B1(n9373), .B2(n6699), .A(n5657), .ZN(n5605) );
  OAI211_X1 U7239 ( .C1(n5606), .C2(n5605), .A(n6627), .B(n5615), .ZN(n5608)
         );
  INV_X1 U7240 ( .A(n5610), .ZN(n5613) );
  INV_X1 U7241 ( .A(n7402), .ZN(n6446) );
  NAND2_X1 U7242 ( .A1(n5545), .A2(n6446), .ZN(n6520) );
  INV_X1 U7243 ( .A(n6520), .ZN(n5617) );
  INV_X1 U7244 ( .A(n6507), .ZN(n5661) );
  INV_X1 U7245 ( .A(n6504), .ZN(n6399) );
  INV_X1 U7246 ( .A(n5621), .ZN(n5626) );
  INV_X1 U7247 ( .A(n5622), .ZN(n5623) );
  NAND4_X1 U7248 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n5629)
         );
  OAI211_X1 U7249 ( .C1(n6198), .C2(n9770), .A(n5545), .B(n5627), .ZN(n5628)
         );
  NOR2_X1 U7250 ( .A1(n5629), .A2(n5628), .ZN(n5631) );
  OAI211_X1 U7251 ( .C1(n7515), .C2(n5631), .A(n5630), .B(n7514), .ZN(n5634)
         );
  AOI21_X1 U7252 ( .B1(n5634), .B2(n5633), .A(n5632), .ZN(n5638) );
  INV_X1 U7253 ( .A(n5635), .ZN(n5637) );
  NOR3_X1 U7254 ( .A1(n5638), .A2(n5637), .A3(n5636), .ZN(n5641) );
  NOR3_X1 U7255 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n5645) );
  OAI211_X1 U7256 ( .C1(n5645), .C2(n5644), .A(n5643), .B(n5642), .ZN(n5646)
         );
  AOI21_X1 U7257 ( .B1(n5646), .B2(n9545), .A(n5262), .ZN(n5650) );
  OAI211_X1 U7258 ( .C1(n5650), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5651)
         );
  NAND4_X1 U7259 ( .A1(n5653), .A2(n6517), .A3(n5652), .A4(n5651), .ZN(n5655)
         );
  AOI21_X1 U7260 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5659) );
  OAI21_X1 U7261 ( .B1(n5659), .B2(n5658), .A(n5657), .ZN(n5660) );
  MUX2_X1 U7262 ( .A(n5661), .B(n6399), .S(n5660), .Z(n5662) );
  OR2_X1 U7263 ( .A1(n6626), .A2(P1_U3086), .ZN(n7696) );
  INV_X1 U7264 ( .A(n7696), .ZN(n5666) );
  XNOR2_X1 U7265 ( .A(n5667), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7266 ( .A1(n4383), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7267 ( .A1(n6508), .A2(n5620), .ZN(n6505) );
  NAND2_X1 U7268 ( .A1(n5545), .A2(n7402), .ZN(n6192) );
  OR2_X1 U7269 ( .A1(n6505), .A2(n6192), .ZN(n7116) );
  NOR4_X1 U7270 ( .A1(n7110), .A2(n5672), .A3(n5673), .A4(n7116), .ZN(n5675)
         );
  OAI21_X1 U7271 ( .B1(n7696), .B2(n6508), .A(P1_B_REG_SCAN_IN), .ZN(n5674) );
  NOR2_X1 U7272 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5678) );
  NOR2_X1 U7273 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5677) );
  NAND2_X1 U7274 ( .A1(n5696), .A2(n5697), .ZN(n5693) );
  INV_X1 U7275 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7276 ( .A1(n5683), .A2(n5681), .ZN(n9023) );
  INV_X1 U7277 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7060) );
  INV_X1 U7278 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5685) );
  INV_X1 U7279 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7280 ( .A1(n4290), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7281 ( .A1(n5693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7282 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5698) );
  MUX2_X1 U7283 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5698), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5699) );
  OR2_X1 U7284 ( .A1(n4313), .A2(n4887), .ZN(n5702) );
  INV_X1 U7285 ( .A(n5700), .ZN(n6580) );
  NAND2_X1 U7286 ( .A1(n8368), .A2(n8366), .ZN(n7054) );
  INV_X1 U7287 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5705) );
  INV_X1 U7288 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5706) );
  OR2_X1 U7289 ( .A1(n5971), .A2(n5706), .ZN(n5709) );
  INV_X1 U7290 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7291 ( .A1(n5940), .A2(n6698), .ZN(n5708) );
  NAND2_X1 U7292 ( .A1(n5726), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5707) );
  NAND4_X1 U7293 ( .A1(n5710), .A2(n5709), .A3(n5708), .A4(n5707), .ZN(n6131)
         );
  NAND2_X1 U7294 ( .A1(n4907), .A2(SI_0_), .ZN(n5712) );
  INV_X1 U7295 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5711) );
  XNOR2_X1 U7296 ( .A(n5712), .B(n5711), .ZN(n9035) );
  MUX2_X1 U7297 ( .A(n6649), .B(n9035), .S(n6642), .Z(n6637) );
  INV_X1 U7298 ( .A(n6637), .ZN(n6813) );
  NAND2_X1 U7299 ( .A1(n8566), .A2(n6813), .ZN(n7056) );
  NAND2_X1 U7300 ( .A1(n7054), .A2(n7056), .ZN(n5714) );
  NAND2_X1 U7301 ( .A1(n6800), .A2(n5703), .ZN(n5713) );
  NAND2_X1 U7302 ( .A1(n5714), .A2(n5713), .ZN(n9828) );
  NAND2_X1 U7303 ( .A1(n4290), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5718) );
  INV_X1 U7304 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9822) );
  OR2_X1 U7305 ( .A1(n5940), .A2(n9822), .ZN(n5717) );
  INV_X1 U7306 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6715) );
  INV_X1 U7307 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5715) );
  OR2_X1 U7308 ( .A1(n4315), .A2(n5715), .ZN(n5716) );
  INV_X1 U7309 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U7310 ( .A1(n5720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5721) );
  OR2_X1 U7311 ( .A1(n4288), .A2(n4566), .ZN(n5723) );
  OR2_X1 U7312 ( .A1(n5827), .A2(n6590), .ZN(n5722) );
  NAND2_X1 U7313 ( .A1(n9828), .A2(n9827), .ZN(n5725) );
  OR2_X1 U7314 ( .A1(n8565), .A2(n8377), .ZN(n5724) );
  NAND2_X1 U7315 ( .A1(n5726), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5731) );
  INV_X1 U7316 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5727) );
  OR2_X1 U7317 ( .A1(n4306), .A2(n5727), .ZN(n5729) );
  OR2_X1 U7318 ( .A1(n5940), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7319 ( .A1(n5719), .A2(n9983), .ZN(n5733) );
  NAND2_X1 U7320 ( .A1(n5733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5732) );
  MUX2_X1 U7321 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5732), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5734) );
  INV_X1 U7322 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6574) );
  INV_X1 U7323 ( .A(n5735), .ZN(n6584) );
  OR2_X1 U7324 ( .A1(n5827), .A2(n6584), .ZN(n5736) );
  NAND2_X1 U7325 ( .A1(n8376), .A2(n6839), .ZN(n7176) );
  NAND2_X1 U7326 ( .A1(n7178), .A2(n7176), .ZN(n7153) );
  NAND2_X1 U7327 ( .A1(n5726), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7328 ( .A1(n7184), .A2(n6748), .ZN(n5755) );
  NAND2_X1 U7329 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5739) );
  AND2_X1 U7330 ( .A1(n5755), .A2(n5739), .ZN(n7152) );
  OR2_X1 U7331 ( .A1(n5940), .A2(n7152), .ZN(n5742) );
  INV_X1 U7332 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5740) );
  OR2_X1 U7333 ( .A1(n4306), .A2(n5740), .ZN(n5741) );
  NAND2_X1 U7334 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5746) );
  INV_X1 U7335 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5745) );
  INV_X1 U7336 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6576) );
  OR2_X1 U7337 ( .A1(n4314), .A2(n6576), .ZN(n5749) );
  INV_X1 U7338 ( .A(n5747), .ZN(n6582) );
  OR2_X1 U7339 ( .A1(n5827), .A2(n6582), .ZN(n5748) );
  OAI211_X1 U7340 ( .C1(n4310), .C2(n6859), .A(n5749), .B(n5748), .ZN(n7005)
         );
  NAND2_X1 U7341 ( .A1(n7153), .A2(n8333), .ZN(n5752) );
  INV_X1 U7342 ( .A(n7005), .ZN(n9849) );
  NAND2_X1 U7343 ( .A1(n5750), .A2(n9849), .ZN(n5751) );
  NAND2_X1 U7344 ( .A1(n6069), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5760) );
  INV_X1 U7345 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6849) );
  INV_X1 U7346 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6850) );
  OR2_X1 U7347 ( .A1(n4307), .A2(n6850), .ZN(n5758) );
  INV_X1 U7348 ( .A(n5755), .ZN(n5754) );
  NAND2_X1 U7349 ( .A1(n5754), .A2(n5753), .ZN(n5770) );
  NAND2_X1 U7350 ( .A1(n5755), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5756) );
  AND2_X1 U7351 ( .A1(n5770), .A2(n5756), .ZN(n7172) );
  OR2_X1 U7352 ( .A1(n5940), .A2(n7172), .ZN(n5757) );
  NOR2_X1 U7353 ( .A1(n5764), .A2(n6078), .ZN(n5762) );
  MUX2_X1 U7354 ( .A(n6078), .B(n5762), .S(P2_IR_REG_5__SCAN_IN), .Z(n5765) );
  INV_X1 U7355 ( .A(n5766), .ZN(n6586) );
  OR2_X1 U7356 ( .A1(n5827), .A2(n6586), .ZN(n5768) );
  INV_X1 U7357 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6573) );
  OR2_X1 U7358 ( .A1(n4313), .A2(n6573), .ZN(n5767) );
  OAI211_X1 U7359 ( .C1(n4309), .C2(n6963), .A(n5768), .B(n5767), .ZN(n7048)
         );
  NAND2_X1 U7360 ( .A1(n8563), .A2(n7048), .ZN(n7159) );
  NAND2_X1 U7361 ( .A1(n5738), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5775) );
  INV_X1 U7362 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5769) );
  OR2_X1 U7363 ( .A1(n4315), .A2(n5769), .ZN(n5774) );
  NAND2_X1 U7364 ( .A1(n5770), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5771) );
  AND2_X1 U7365 ( .A1(n5787), .A2(n5771), .ZN(n7264) );
  OR2_X1 U7366 ( .A1(n5940), .A2(n7264), .ZN(n5773) );
  INV_X1 U7367 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8150) );
  OR2_X1 U7368 ( .A1(n4306), .A2(n8150), .ZN(n5772) );
  NOR2_X1 U7369 ( .A1(n5778), .A2(n6078), .ZN(n5776) );
  MUX2_X1 U7370 ( .A(n6078), .B(n5776), .S(P2_IR_REG_6__SCAN_IN), .Z(n5780) );
  NAND2_X1 U7371 ( .A1(n5778), .A2(n5777), .ZN(n5811) );
  INV_X1 U7372 ( .A(n5811), .ZN(n5779) );
  OR2_X1 U7373 ( .A1(n5827), .A2(n6588), .ZN(n5782) );
  OR2_X1 U7374 ( .A1(n4313), .A2(n6575), .ZN(n5781) );
  OAI211_X1 U7375 ( .C1(n6642), .C2(n7074), .A(n5782), .B(n5781), .ZN(n8152)
         );
  INV_X1 U7376 ( .A(n8152), .ZN(n9861) );
  OR2_X1 U7377 ( .A1(n7292), .A2(n9861), .ZN(n8147) );
  AND2_X1 U7378 ( .A1(n7159), .A2(n8147), .ZN(n5798) );
  NAND2_X1 U7379 ( .A1(n5726), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5792) );
  INV_X1 U7380 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5783) );
  OR2_X1 U7381 ( .A1(n6046), .A2(n5783), .ZN(n5791) );
  INV_X1 U7382 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5784) );
  OR2_X1 U7383 ( .A1(n4307), .A2(n5784), .ZN(n5790) );
  NAND2_X1 U7384 ( .A1(n5786), .A2(n5785), .ZN(n5800) );
  NAND2_X1 U7385 ( .A1(n5787), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5788) );
  AND2_X1 U7386 ( .A1(n5800), .A2(n5788), .ZN(n7289) );
  OR2_X1 U7387 ( .A1(n5940), .A2(n7289), .ZN(n5789) );
  AND2_X1 U7389 ( .A1(n8303), .A2(n6577), .ZN(n5797) );
  NAND2_X1 U7390 ( .A1(n5811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  INV_X1 U7391 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5793) );
  XNOR2_X1 U7392 ( .A(n5794), .B(n5793), .ZN(n7205) );
  NOR2_X1 U7393 ( .A1(n4310), .A2(n7205), .ZN(n5796) );
  INV_X1 U7394 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U7395 ( .A1(n4314), .A2(n6578), .ZN(n5795) );
  OR2_X1 U7396 ( .A1(n8419), .A2(n9864), .ZN(n5806) );
  AND2_X1 U7397 ( .A1(n5798), .A2(n5806), .ZN(n5816) );
  NAND2_X1 U7398 ( .A1(n6069), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5805) );
  INV_X1 U7399 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5799) );
  OR2_X1 U7400 ( .A1(n6046), .A2(n5799), .ZN(n5804) );
  NAND2_X1 U7401 ( .A1(n5800), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5801) );
  AND2_X1 U7402 ( .A1(n5831), .A2(n5801), .ZN(n7401) );
  OR2_X1 U7403 ( .A1(n5940), .A2(n7401), .ZN(n5803) );
  INV_X1 U7404 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7194) );
  OR2_X1 U7405 ( .A1(n4307), .A2(n7194), .ZN(n5802) );
  NAND4_X1 U7406 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n8561)
         );
  INV_X1 U7407 ( .A(n5806), .ZN(n5809) );
  NAND2_X1 U7408 ( .A1(n7292), .A2(n9861), .ZN(n8146) );
  NAND2_X1 U7409 ( .A1(n9864), .A2(n8419), .ZN(n5807) );
  AND2_X1 U7410 ( .A1(n8146), .A2(n5807), .ZN(n5808) );
  OR2_X1 U7411 ( .A1(n5809), .A2(n5808), .ZN(n7189) );
  AND2_X1 U7412 ( .A1(n8561), .A2(n7189), .ZN(n5810) );
  NAND2_X1 U7413 ( .A1(n7190), .A2(n5810), .ZN(n5815) );
  NAND2_X1 U7414 ( .A1(n6596), .A2(n8303), .ZN(n5814) );
  OAI21_X1 U7415 ( .B1(n5811), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  INV_X1 U7416 ( .A(n7497), .ZN(n7225) );
  AOI22_X1 U7417 ( .A1(n5965), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5964), .B2(
        n7225), .ZN(n5813) );
  NAND2_X1 U7418 ( .A1(n5814), .A2(n5813), .ZN(n7398) );
  NAND2_X1 U7419 ( .A1(n5815), .A2(n9870), .ZN(n5821) );
  OR2_X1 U7420 ( .A1(n8561), .A2(n7189), .ZN(n5819) );
  INV_X1 U7421 ( .A(n8561), .ZN(n7407) );
  AND2_X1 U7422 ( .A1(n5816), .A2(n7407), .ZN(n5817) );
  NAND2_X1 U7423 ( .A1(n7160), .A2(n5817), .ZN(n5818) );
  AND2_X1 U7424 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  NAND2_X1 U7425 ( .A1(n5821), .A2(n5820), .ZN(n7346) );
  NAND2_X1 U7426 ( .A1(n5822), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  MUX2_X1 U7427 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5823), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5825) );
  INV_X1 U7428 ( .A(n5851), .ZN(n5824) );
  AOI22_X1 U7429 ( .A1(n5965), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5964), .B2(
        n7545), .ZN(n5826) );
  NAND2_X1 U7430 ( .A1(n6069), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5837) );
  INV_X1 U7431 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7432 ( .A1(n6046), .A2(n5828), .ZN(n5836) );
  NAND2_X1 U7433 ( .A1(n5831), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5832) );
  AND2_X1 U7434 ( .A1(n5841), .A2(n5832), .ZN(n7415) );
  OR2_X1 U7435 ( .A1(n5940), .A2(n7415), .ZN(n5835) );
  INV_X1 U7436 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5833) );
  OR2_X1 U7437 ( .A1(n4307), .A2(n5833), .ZN(n5834) );
  NAND4_X1 U7438 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .ZN(n8560)
         );
  OR2_X1 U7439 ( .A1(n9878), .A2(n8431), .ZN(n8407) );
  NAND2_X1 U7440 ( .A1(n9878), .A2(n8431), .ZN(n8406) );
  NAND2_X1 U7441 ( .A1(n8407), .A2(n8406), .ZN(n8340) );
  NAND2_X1 U7442 ( .A1(n7346), .A2(n8340), .ZN(n5839) );
  OR2_X1 U7443 ( .A1(n9878), .A2(n8560), .ZN(n5838) );
  NAND2_X1 U7444 ( .A1(n5839), .A2(n5838), .ZN(n7355) );
  NAND2_X1 U7445 ( .A1(n5726), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5846) );
  INV_X1 U7446 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5840) );
  OR2_X1 U7447 ( .A1(n6046), .A2(n5840), .ZN(n5845) );
  NAND2_X1 U7448 ( .A1(n5841), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5842) );
  AND2_X1 U7449 ( .A1(n5856), .A2(n5842), .ZN(n7672) );
  OR2_X1 U7450 ( .A1(n5940), .A2(n7672), .ZN(n5844) );
  INV_X1 U7451 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7359) );
  OR2_X1 U7452 ( .A1(n4306), .A2(n7359), .ZN(n5843) );
  NAND2_X1 U7453 ( .A1(n6607), .A2(n8303), .ZN(n5849) );
  OR2_X1 U7454 ( .A1(n5851), .A2(n6078), .ZN(n5847) );
  XNOR2_X1 U7455 ( .A(n5847), .B(n5850), .ZN(n7549) );
  INV_X1 U7456 ( .A(n7549), .ZN(n7612) );
  AOI22_X1 U7457 ( .A1(n5965), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5964), .B2(
        n7612), .ZN(n5848) );
  NAND2_X1 U7458 ( .A1(n5849), .A2(n5848), .ZN(n9884) );
  NAND2_X1 U7459 ( .A1(n6613), .A2(n8303), .ZN(n5854) );
  AND2_X1 U7460 ( .A1(n5851), .A2(n5850), .ZN(n5866) );
  OR2_X1 U7461 ( .A1(n5866), .A2(n6078), .ZN(n5852) );
  XNOR2_X1 U7462 ( .A(n5852), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7825) );
  AOI22_X1 U7463 ( .A1(n5965), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5964), .B2(
        n7825), .ZN(n5853) );
  NAND2_X1 U7464 ( .A1(n5854), .A2(n5853), .ZN(n7687) );
  NAND2_X1 U7465 ( .A1(n6069), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5862) );
  INV_X1 U7466 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7467 ( .A1(n6046), .A2(n5855), .ZN(n5861) );
  NAND2_X1 U7468 ( .A1(n5856), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5857) );
  AND2_X1 U7469 ( .A1(n5875), .A2(n5857), .ZN(n7685) );
  OR2_X1 U7470 ( .A1(n5940), .A2(n7685), .ZN(n5860) );
  INV_X1 U7471 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5858) );
  OR2_X1 U7472 ( .A1(n4306), .A2(n5858), .ZN(n5859) );
  NAND2_X1 U7473 ( .A1(n7687), .A2(n7794), .ZN(n8440) );
  NAND2_X1 U7474 ( .A1(n8434), .A2(n8440), .ZN(n8343) );
  INV_X1 U7475 ( .A(n7794), .ZN(n7792) );
  NAND2_X1 U7476 ( .A1(n7687), .A2(n7792), .ZN(n5863) );
  NAND2_X1 U7477 ( .A1(n5864), .A2(n5863), .ZN(n7476) );
  NAND2_X1 U7478 ( .A1(n6630), .A2(n8303), .ZN(n5872) );
  NAND2_X1 U7479 ( .A1(n5866), .A2(n5865), .ZN(n5868) );
  NAND2_X1 U7480 ( .A1(n5868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  MUX2_X1 U7481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5867), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n5870) );
  AOI22_X1 U7482 ( .A1(n5965), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5964), .B2(
        n7831), .ZN(n5871) );
  NAND2_X1 U7483 ( .A1(n5872), .A2(n5871), .ZN(n9893) );
  NAND2_X1 U7484 ( .A1(n6069), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5880) );
  INV_X1 U7485 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7827) );
  OR2_X1 U7486 ( .A1(n6046), .A2(n7827), .ZN(n5879) );
  NAND2_X1 U7487 ( .A1(n5875), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5876) );
  AND2_X1 U7488 ( .A1(n5888), .A2(n5876), .ZN(n7797) );
  OR2_X1 U7489 ( .A1(n5940), .A2(n7797), .ZN(n5878) );
  INV_X1 U7490 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7820) );
  OR2_X1 U7491 ( .A1(n4306), .A2(n7820), .ZN(n5877) );
  NAND4_X1 U7492 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n8559)
         );
  AND2_X1 U7493 ( .A1(n9893), .A2(n8559), .ZN(n5882) );
  OR2_X1 U7494 ( .A1(n9893), .A2(n8559), .ZN(n5881) );
  NAND2_X1 U7495 ( .A1(n6634), .A2(n8303), .ZN(n5885) );
  NAND2_X1 U7496 ( .A1(n4332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7497 ( .A(n5883), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8598) );
  AOI22_X1 U7498 ( .A1(n5965), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5964), .B2(
        n8598), .ZN(n5884) );
  NAND2_X1 U7499 ( .A1(n5726), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5893) );
  INV_X1 U7500 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7501 ( .A1(n6046), .A2(n5886), .ZN(n5892) );
  NAND2_X1 U7502 ( .A1(n5888), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5889) );
  AND2_X1 U7503 ( .A1(n5899), .A2(n5889), .ZN(n7936) );
  OR2_X1 U7504 ( .A1(n5940), .A2(n7936), .ZN(n5891) );
  INV_X1 U7505 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7750) );
  OR2_X1 U7506 ( .A1(n4307), .A2(n7750), .ZN(n5890) );
  NOR2_X1 U7507 ( .A1(n8451), .A2(n8558), .ZN(n8450) );
  NAND2_X1 U7508 ( .A1(n6701), .A2(n8303), .ZN(n5898) );
  OR2_X1 U7509 ( .A1(n5921), .A2(n6078), .ZN(n5895) );
  INV_X1 U7510 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7511 ( .A1(n5895), .A2(n5894), .ZN(n5905) );
  OR2_X1 U7512 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NAND2_X1 U7513 ( .A1(n5905), .A2(n5896), .ZN(n8622) );
  INV_X1 U7514 ( .A(n8622), .ZN(n8607) );
  AOI22_X1 U7515 ( .A1(n5965), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5964), .B2(
        n8607), .ZN(n5897) );
  INV_X1 U7516 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7913) );
  OR2_X1 U7517 ( .A1(n6046), .A2(n7913), .ZN(n5904) );
  INV_X1 U7518 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10042) );
  OR2_X1 U7519 ( .A1(n4315), .A2(n10042), .ZN(n5903) );
  NAND2_X1 U7520 ( .A1(n5899), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5900) );
  AND2_X1 U7521 ( .A1(n5911), .A2(n5900), .ZN(n7894) );
  OR2_X1 U7522 ( .A1(n5940), .A2(n7894), .ZN(n5902) );
  INV_X1 U7523 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7809) );
  OR2_X1 U7524 ( .A1(n4306), .A2(n7809), .ZN(n5901) );
  NAND4_X1 U7525 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n8557)
         );
  NAND2_X1 U7526 ( .A1(n6764), .A2(n8303), .ZN(n5908) );
  NAND2_X1 U7527 ( .A1(n5905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5906) );
  XNOR2_X1 U7528 ( .A(n5906), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8646) );
  AOI22_X1 U7529 ( .A1(n5965), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5964), .B2(
        n8646), .ZN(n5907) );
  NAND2_X1 U7530 ( .A1(n6069), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5916) );
  INV_X1 U7531 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8624) );
  OR2_X1 U7532 ( .A1(n6046), .A2(n8624), .ZN(n5915) );
  NAND2_X1 U7533 ( .A1(n5911), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5912) );
  AND2_X1 U7534 ( .A1(n5928), .A2(n5912), .ZN(n7972) );
  OR2_X1 U7535 ( .A1(n5940), .A2(n7972), .ZN(n5914) );
  INV_X1 U7536 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7971) );
  OR2_X1 U7537 ( .A1(n4306), .A2(n7971), .ZN(n5913) );
  NAND4_X1 U7538 ( .A1(n5916), .A2(n5915), .A3(n5914), .A4(n5913), .ZN(n8891)
         );
  INV_X1 U7539 ( .A(n8891), .ZN(n7891) );
  NAND2_X1 U7540 ( .A1(n8025), .A2(n7891), .ZN(n8467) );
  INV_X1 U7541 ( .A(n8463), .ZN(n5917) );
  NAND2_X1 U7542 ( .A1(n5918), .A2(n5917), .ZN(n7963) );
  NAND2_X1 U7543 ( .A1(n8025), .A2(n8891), .ZN(n5919) );
  NAND2_X1 U7544 ( .A1(n7963), .A2(n5919), .ZN(n8888) );
  NAND2_X1 U7545 ( .A1(n6920), .A2(n8303), .ZN(n5927) );
  OR2_X1 U7546 ( .A1(n5924), .A2(n6078), .ZN(n5922) );
  MUX2_X1 U7547 ( .A(n5922), .B(P2_IR_REG_31__SCAN_IN), .S(n5923), .Z(n5925)
         );
  AND2_X1 U7548 ( .A1(n5925), .A2(n5936), .ZN(n8654) );
  AOI22_X1 U7549 ( .A1(n5965), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5964), .B2(
        n8654), .ZN(n5926) );
  NAND2_X1 U7550 ( .A1(n5726), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5934) );
  INV_X1 U7551 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8649) );
  OR2_X1 U7552 ( .A1(n6046), .A2(n8649), .ZN(n5933) );
  NAND2_X1 U7553 ( .A1(n5928), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5929) );
  AND2_X1 U7554 ( .A1(n5943), .A2(n5929), .ZN(n8896) );
  OR2_X1 U7555 ( .A1(n5940), .A2(n8896), .ZN(n5932) );
  INV_X1 U7556 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7557 ( .A1(n4307), .A2(n5930), .ZN(n5931) );
  NAND4_X1 U7558 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n8879)
         );
  NAND2_X1 U7559 ( .A1(n8900), .A2(n8036), .ZN(n8471) );
  NAND2_X1 U7560 ( .A1(n8469), .A2(n8471), .ZN(n8889) );
  NAND2_X1 U7561 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  NAND2_X1 U7562 ( .A1(n8900), .A2(n8879), .ZN(n8876) );
  NAND2_X1 U7563 ( .A1(n8887), .A2(n8876), .ZN(n5949) );
  NAND2_X1 U7564 ( .A1(n7027), .A2(n8303), .ZN(n5939) );
  NAND2_X1 U7565 ( .A1(n5936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5935) );
  MUX2_X1 U7566 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5935), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5937) );
  AND2_X1 U7567 ( .A1(n5937), .A2(n4339), .ZN(n8692) );
  AOI22_X1 U7568 ( .A1(n5965), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5964), .B2(
        n8692), .ZN(n5938) );
  NAND2_X1 U7569 ( .A1(n5943), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7570 ( .A1(n5955), .A2(n5944), .ZN(n8883) );
  NAND2_X1 U7571 ( .A1(n6085), .A2(n8883), .ZN(n5948) );
  INV_X1 U7572 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8938) );
  OR2_X1 U7573 ( .A1(n6046), .A2(n8938), .ZN(n5947) );
  INV_X1 U7574 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9008) );
  OR2_X1 U7575 ( .A1(n4315), .A2(n9008), .ZN(n5946) );
  INV_X1 U7576 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8882) );
  OR2_X1 U7577 ( .A1(n4306), .A2(n8882), .ZN(n5945) );
  NAND4_X1 U7578 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8890)
         );
  OR2_X1 U7579 ( .A1(n9011), .A2(n8863), .ZN(n8473) );
  NAND2_X1 U7580 ( .A1(n9011), .A2(n8863), .ZN(n8852) );
  NAND2_X1 U7581 ( .A1(n5949), .A2(n8875), .ZN(n8814) );
  NAND2_X1 U7582 ( .A1(n7064), .A2(n8303), .ZN(n5954) );
  OR2_X1 U7583 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  AND2_X1 U7584 ( .A1(n5961), .A2(n5952), .ZN(n8713) );
  AOI22_X1 U7585 ( .A1(n5965), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5964), .B2(
        n8713), .ZN(n5953) );
  NAND2_X1 U7586 ( .A1(n5955), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7587 ( .A1(n5969), .A2(n5956), .ZN(n8867) );
  NAND2_X1 U7588 ( .A1(n6085), .A2(n8867), .ZN(n5960) );
  INV_X1 U7589 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9005) );
  OR2_X1 U7590 ( .A1(n4315), .A2(n9005), .ZN(n5959) );
  INV_X1 U7591 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8936) );
  OR2_X1 U7592 ( .A1(n6046), .A2(n8936), .ZN(n5958) );
  INV_X1 U7593 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8869) );
  OR2_X1 U7594 ( .A1(n4307), .A2(n8869), .ZN(n5957) );
  NAND4_X1 U7595 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8878)
         );
  NAND2_X1 U7596 ( .A1(n8935), .A2(n8842), .ZN(n8475) );
  AOI22_X1 U7597 ( .A1(n5965), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8547), .B2(
        n5964), .ZN(n5966) );
  INV_X1 U7598 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7599 ( .A1(n5969), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7600 ( .A1(n5979), .A2(n5970), .ZN(n8848) );
  NAND2_X1 U7601 ( .A1(n8848), .A2(n6085), .ZN(n5976) );
  INV_X1 U7602 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9982) );
  OR2_X1 U7603 ( .A1(n4315), .A2(n9982), .ZN(n5973) );
  INV_X1 U7604 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8931) );
  OR2_X1 U7605 ( .A1(n6046), .A2(n8931), .ZN(n5972) );
  AND2_X1 U7606 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  INV_X1 U7607 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8847) );
  OR2_X1 U7608 ( .A1(n4306), .A2(n8847), .ZN(n5974) );
  INV_X1 U7609 ( .A(n8865), .ZN(n8824) );
  AND2_X1 U7610 ( .A1(n5985), .A2(n8824), .ZN(n5986) );
  OR2_X1 U7611 ( .A1(n8860), .A2(n5986), .ZN(n8816) );
  NAND2_X1 U7612 ( .A1(n7353), .A2(n8303), .ZN(n5978) );
  INV_X1 U7613 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10068) );
  OR2_X1 U7614 ( .A1(n4314), .A2(n10068), .ZN(n5977) );
  NAND2_X1 U7615 ( .A1(n5979), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7616 ( .A1(n5991), .A2(n5980), .ZN(n8829) );
  NAND2_X1 U7617 ( .A1(n8829), .A2(n6085), .ZN(n5983) );
  AOI22_X1 U7618 ( .A1(n6069), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n5738), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5982) );
  INV_X1 U7619 ( .A(n4307), .ZN(n6043) );
  NAND2_X1 U7620 ( .A1(n6043), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7621 ( .A1(n8830), .A2(n8843), .ZN(n8488) );
  NOR2_X1 U7622 ( .A1(n8816), .A2(n8819), .ZN(n5984) );
  NAND2_X1 U7623 ( .A1(n9011), .A2(n8890), .ZN(n8815) );
  AND2_X1 U7624 ( .A1(n5984), .A2(n8815), .ZN(n5987) );
  XNOR2_X1 U7625 ( .A(n5985), .B(n8865), .ZN(n6145) );
  OR2_X1 U7626 ( .A1(n8935), .A2(n8878), .ZN(n8836) );
  AND2_X1 U7627 ( .A1(n6145), .A2(n8836), .ZN(n8839) );
  INV_X1 U7628 ( .A(n8843), .ZN(n8806) );
  NAND2_X1 U7629 ( .A1(n7405), .A2(n8303), .ZN(n5989) );
  OR2_X1 U7630 ( .A1(n4314), .A2(n10074), .ZN(n5988) );
  INV_X1 U7631 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U7632 ( .A1(n5991), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7633 ( .A1(n5997), .A2(n5992), .ZN(n8810) );
  NAND2_X1 U7634 ( .A1(n8810), .A2(n6085), .ZN(n5994) );
  AOI22_X1 U7635 ( .A1(n5726), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5738), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5993) );
  OAI211_X1 U7636 ( .C1(n4306), .C2(n8809), .A(n5994), .B(n5993), .ZN(n8825)
         );
  NAND2_X1 U7637 ( .A1(n8991), .A2(n8796), .ZN(n8498) );
  INV_X1 U7638 ( .A(n8991), .ZN(n8243) );
  NAND2_X1 U7639 ( .A1(n7581), .A2(n8303), .ZN(n5996) );
  OR2_X1 U7640 ( .A1(n4314), .A2(n7586), .ZN(n5995) );
  NAND2_X1 U7641 ( .A1(n5997), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7642 ( .A1(n6004), .A2(n5998), .ZN(n8797) );
  INV_X1 U7643 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U7644 ( .A1(n6069), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7645 ( .A1(n5738), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7646 ( .C1(n8798), .C2(n4307), .A(n6000), .B(n5999), .ZN(n6001)
         );
  NAND2_X1 U7647 ( .A1(n8923), .A2(n8238), .ZN(n8492) );
  INV_X1 U7648 ( .A(n8238), .ZN(n8807) );
  NAND2_X1 U7649 ( .A1(n7695), .A2(n8303), .ZN(n6003) );
  OR2_X1 U7650 ( .A1(n4313), .A2(n7693), .ZN(n6002) );
  NAND2_X1 U7651 ( .A1(n6004), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7652 ( .A1(n6017), .A2(n6005), .ZN(n8788) );
  NAND2_X1 U7653 ( .A1(n8788), .A2(n6085), .ZN(n6010) );
  INV_X1 U7654 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U7655 ( .A1(n5738), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7656 ( .A1(n5726), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6006) );
  OAI211_X1 U7657 ( .C1(n8787), .C2(n4306), .A(n6007), .B(n6006), .ZN(n6008)
         );
  INV_X1 U7658 ( .A(n6008), .ZN(n6009) );
  NOR2_X1 U7659 ( .A1(n8981), .A2(n8773), .ZN(n6012) );
  INV_X1 U7660 ( .A(n8981), .ZN(n6011) );
  OAI22_X1 U7661 ( .A1(n8784), .A2(n6012), .B1(n6011), .B2(n8795), .ZN(n8772)
         );
  INV_X1 U7662 ( .A(n8772), .ZN(n6026) );
  NAND2_X1 U7663 ( .A1(n7801), .A2(n8303), .ZN(n6014) );
  OR2_X1 U7664 ( .A1(n4314), .A2(n7802), .ZN(n6013) );
  INV_X1 U7665 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7666 ( .A1(n6017), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7667 ( .A1(n6031), .A2(n6018), .ZN(n8776) );
  NAND2_X1 U7668 ( .A1(n8776), .A2(n6085), .ZN(n6023) );
  INV_X1 U7669 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7670 ( .A1(n6069), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7671 ( .A1(n6043), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6019) );
  OAI211_X1 U7672 ( .C1(n6046), .C2(n8916), .A(n6020), .B(n6019), .ZN(n6021)
         );
  INV_X1 U7673 ( .A(n6021), .ZN(n6022) );
  INV_X1 U7674 ( .A(n8975), .ZN(n8778) );
  NAND2_X1 U7675 ( .A1(n7878), .A2(n8303), .ZN(n6028) );
  OR2_X1 U7676 ( .A1(n4313), .A2(n9991), .ZN(n6027) );
  INV_X1 U7677 ( .A(n6031), .ZN(n6030) );
  INV_X1 U7678 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7679 ( .A1(n6031), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7680 ( .A1(n6041), .A2(n6032), .ZN(n8761) );
  NAND2_X1 U7681 ( .A1(n8761), .A2(n6085), .ZN(n6038) );
  INV_X1 U7682 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7683 ( .A1(n5738), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7684 ( .A1(n6069), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6033) );
  OAI211_X1 U7685 ( .C1(n4306), .C2(n6035), .A(n6034), .B(n6033), .ZN(n6036)
         );
  INV_X1 U7686 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7687 ( .A1(n8244), .A2(n8193), .ZN(n8511) );
  NAND2_X1 U7688 ( .A1(n7979), .A2(n8303), .ZN(n6040) );
  OR2_X1 U7689 ( .A1(n4314), .A2(n7980), .ZN(n6039) );
  NAND2_X1 U7690 ( .A1(n6041), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7691 ( .A1(n6055), .A2(n6042), .ZN(n8753) );
  NAND2_X1 U7692 ( .A1(n8753), .A2(n6085), .ZN(n6049) );
  INV_X1 U7693 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U7694 ( .A1(n5726), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7695 ( .A1(n6043), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6044) );
  OAI211_X1 U7696 ( .C1(n6046), .C2(n10077), .A(n6045), .B(n6044), .ZN(n6047)
         );
  INV_X1 U7697 ( .A(n6047), .ZN(n6048) );
  NOR2_X1 U7698 ( .A1(n8964), .A2(n8743), .ZN(n6050) );
  INV_X1 U7699 ( .A(n8964), .ZN(n8297) );
  NAND2_X1 U7700 ( .A1(n8086), .A2(n8303), .ZN(n6052) );
  OR2_X1 U7701 ( .A1(n4314), .A2(n8087), .ZN(n6051) );
  INV_X1 U7702 ( .A(n6055), .ZN(n6054) );
  INV_X1 U7703 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7704 ( .A1(n6054), .A2(n6053), .ZN(n6067) );
  NAND2_X1 U7705 ( .A1(n6055), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7706 ( .A1(n6067), .A2(n6056), .ZN(n8746) );
  NAND2_X1 U7707 ( .A1(n8746), .A2(n6085), .ZN(n6061) );
  INV_X1 U7708 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U7709 ( .A1(n5726), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7710 ( .A1(n5738), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6057) );
  OAI211_X1 U7711 ( .C1(n8745), .C2(n4307), .A(n6058), .B(n6057), .ZN(n6059)
         );
  INV_X1 U7712 ( .A(n6059), .ZN(n6060) );
  INV_X1 U7713 ( .A(n8958), .ZN(n6063) );
  NAND2_X1 U7714 ( .A1(n8088), .A2(n8303), .ZN(n6066) );
  OR2_X1 U7715 ( .A1(n4314), .A2(n6064), .ZN(n6065) );
  NAND2_X1 U7716 ( .A1(n6067), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7717 ( .A1(n6084), .A2(n6068), .ZN(n8222) );
  NAND2_X1 U7718 ( .A1(n8222), .A2(n6085), .ZN(n6074) );
  INV_X1 U7719 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7720 ( .A1(n5738), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7721 ( .A1(n6069), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6070) );
  OAI211_X1 U7722 ( .C1(n6169), .C2(n4307), .A(n6071), .B(n6070), .ZN(n6072)
         );
  INV_X1 U7723 ( .A(n6072), .ZN(n6073) );
  NAND2_X1 U7724 ( .A1(n8533), .A2(n8524), .ZN(n6538) );
  NAND2_X1 U7725 ( .A1(n6540), .A2(n6538), .ZN(n8326) );
  XNOR2_X1 U7726 ( .A(n6554), .B(n8326), .ZN(n6096) );
  NAND2_X1 U7727 ( .A1(n4353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7728 ( .A1(n8547), .A2(n8550), .ZN(n6123) );
  AND2_X1 U7729 ( .A1(n6076), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6077) );
  MUX2_X1 U7730 ( .A(n6078), .B(n6077), .S(P2_IR_REG_20__SCAN_IN), .Z(n6079)
         );
  INV_X1 U7731 ( .A(n6079), .ZN(n6081) );
  INV_X1 U7732 ( .A(n8539), .ZN(n8322) );
  NAND2_X1 U7733 ( .A1(n6082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7734 ( .A1(n8322), .A2(n8370), .ZN(n8320) );
  NAND2_X1 U7735 ( .A1(n8164), .A2(n6085), .ZN(n8313) );
  INV_X1 U7736 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U7737 ( .A1(n5738), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7738 ( .A1(n5726), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6086) );
  OAI211_X1 U7739 ( .C1(n4306), .C2(n8165), .A(n6087), .B(n6086), .ZN(n6088)
         );
  INV_X1 U7740 ( .A(n6088), .ZN(n6089) );
  INV_X1 U7741 ( .A(n6090), .ZN(n6640) );
  NAND2_X1 U7742 ( .A1(n6640), .A2(n8715), .ZN(n6092) );
  NAND2_X1 U7743 ( .A1(n4310), .A2(n6092), .ZN(n6792) );
  NOR2_X1 U7744 ( .A1(n8225), .A2(n8866), .ZN(n6094) );
  NAND2_X1 U7745 ( .A1(n6122), .A2(n4299), .ZN(n6098) );
  NAND2_X1 U7746 ( .A1(n6100), .A2(n4300), .ZN(n6102) );
  XNOR2_X1 U7747 ( .A(n7803), .B(P2_B_REG_SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7748 ( .A1(n7879), .A2(n6103), .ZN(n6106) );
  NAND2_X1 U7749 ( .A1(n6104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7750 ( .A1(n7879), .A2(n7981), .ZN(n6108) );
  NAND2_X1 U7751 ( .A1(n7803), .A2(n7981), .ZN(n6601) );
  NOR2_X1 U7752 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n6114) );
  NOR4_X1 U7753 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6113) );
  NOR4_X1 U7754 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6112) );
  NOR4_X1 U7755 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6111) );
  NAND4_X1 U7756 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n6120)
         );
  NOR4_X1 U7757 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6118) );
  NOR4_X1 U7758 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6117) );
  NOR4_X1 U7759 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6116) );
  NOR4_X1 U7760 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6115) );
  NAND4_X1 U7761 ( .A1(n6118), .A2(n6117), .A3(n6116), .A4(n6115), .ZN(n6119)
         );
  NOR2_X1 U7762 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  NOR2_X1 U7763 ( .A1(n6110), .A2(n6121), .ZN(n6676) );
  INV_X1 U7764 ( .A(n6676), .ZN(n6126) );
  NAND3_X1 U7765 ( .A1(n6175), .A2(n6797), .A3(n6126), .ZN(n6682) );
  XNOR2_X1 U7766 ( .A(n6122), .B(n4299), .ZN(n6654) );
  INV_X1 U7767 ( .A(n6695), .ZN(n6125) );
  OR2_X1 U7768 ( .A1(n8539), .A2(n8370), .ZN(n8329) );
  INV_X1 U7769 ( .A(n8550), .ZN(n7584) );
  AND2_X1 U7770 ( .A1(n8522), .A2(n9886), .ZN(n6124) );
  NAND2_X1 U7771 ( .A1(n6691), .A2(n6124), .ZN(n6688) );
  NAND2_X1 U7772 ( .A1(n6176), .A2(n9892), .ZN(n9823) );
  NAND2_X1 U7773 ( .A1(n6688), .A2(n9823), .ZN(n6674) );
  NAND2_X1 U7774 ( .A1(n6125), .A2(n6674), .ZN(n6130) );
  NAND2_X1 U7775 ( .A1(n6126), .A2(n6600), .ZN(n6159) );
  NAND2_X1 U7776 ( .A1(n6127), .A2(n8539), .ZN(n6796) );
  NAND2_X1 U7777 ( .A1(n6814), .A2(n6691), .ZN(n6128) );
  NAND2_X1 U7778 ( .A1(n6690), .A2(n6128), .ZN(n6129) );
  INV_X1 U7779 ( .A(n6131), .ZN(n6132) );
  OR2_X1 U7780 ( .A1(n8565), .A2(n9841), .ZN(n8379) );
  NAND2_X1 U7781 ( .A1(n8376), .A2(n6835), .ZN(n8380) );
  AND2_X1 U7782 ( .A1(n8379), .A2(n8380), .ZN(n6133) );
  INV_X1 U7783 ( .A(n8380), .ZN(n8397) );
  NAND2_X1 U7784 ( .A1(n6135), .A2(n8380), .ZN(n7148) );
  OR2_X1 U7785 ( .A1(n8563), .A2(n9855), .ZN(n8399) );
  INV_X1 U7786 ( .A(n8399), .ZN(n6136) );
  NAND2_X1 U7787 ( .A1(n8563), .A2(n9855), .ZN(n8395) );
  NOR2_X1 U7788 ( .A1(n7292), .A2(n8152), .ZN(n8401) );
  NAND2_X1 U7789 ( .A1(n7292), .A2(n8152), .ZN(n8400) );
  XNOR2_X1 U7790 ( .A(n8419), .B(n8418), .ZN(n8339) );
  OR2_X1 U7791 ( .A1(n8419), .A2(n8418), .ZN(n8414) );
  AND2_X1 U7792 ( .A1(n9870), .A2(n8561), .ZN(n7188) );
  OR2_X1 U7793 ( .A1(n8561), .A2(n9870), .ZN(n8420) );
  OR2_X1 U7794 ( .A1(n9884), .A2(n8426), .ZN(n8432) );
  NAND2_X1 U7795 ( .A1(n9884), .A2(n8426), .ZN(n8435) );
  INV_X1 U7796 ( .A(n8343), .ZN(n7444) );
  NAND2_X1 U7797 ( .A1(n7441), .A2(n7444), .ZN(n7442) );
  INV_X1 U7798 ( .A(n8559), .ZN(n7682) );
  OR2_X1 U7799 ( .A1(n9893), .A2(n7682), .ZN(n8446) );
  NAND2_X1 U7800 ( .A1(n9893), .A2(n7682), .ZN(n8447) );
  NAND2_X1 U7801 ( .A1(n8446), .A2(n8447), .ZN(n8344) );
  INV_X1 U7802 ( .A(n8440), .ZN(n6137) );
  NOR2_X1 U7803 ( .A1(n8344), .A2(n6137), .ZN(n6138) );
  NOR2_X1 U7804 ( .A1(n8451), .A2(n7886), .ZN(n6140) );
  NAND2_X1 U7805 ( .A1(n8451), .A2(n7886), .ZN(n6139) );
  INV_X1 U7806 ( .A(n8557), .ZN(n7990) );
  AND2_X1 U7807 ( .A1(n7918), .A2(n7990), .ZN(n8460) );
  OR2_X1 U7808 ( .A1(n7918), .A2(n7990), .ZN(n8458) );
  NAND2_X1 U7809 ( .A1(n7962), .A2(n8467), .ZN(n6141) );
  INV_X1 U7810 ( .A(n8875), .ZN(n6142) );
  INV_X1 U7811 ( .A(n8852), .ZN(n6143) );
  NOR2_X1 U7812 ( .A1(n8853), .A2(n6143), .ZN(n6144) );
  NAND2_X1 U7813 ( .A1(n8855), .A2(n8484), .ZN(n8833) );
  OR2_X1 U7814 ( .A1(n5985), .A2(n8865), .ZN(n8479) );
  INV_X1 U7815 ( .A(n8498), .ZN(n6146) );
  NAND2_X1 U7816 ( .A1(n8791), .A2(n8492), .ZN(n6147) );
  NAND2_X1 U7817 ( .A1(n8975), .A2(n8760), .ZN(n8364) );
  NAND2_X1 U7818 ( .A1(n8981), .A2(n8795), .ZN(n8768) );
  INV_X1 U7819 ( .A(n8503), .ZN(n6148) );
  OR2_X1 U7820 ( .A1(n6148), .A2(n8767), .ZN(n6149) );
  NAND2_X1 U7821 ( .A1(n8958), .A2(n8291), .ZN(n8516) );
  NAND2_X1 U7822 ( .A1(n8739), .A2(n8516), .ZN(n6151) );
  NAND2_X1 U7823 ( .A1(n6151), .A2(n8515), .ZN(n6539) );
  XOR2_X1 U7824 ( .A(n8326), .B(n6539), .Z(n6185) );
  OAI21_X1 U7825 ( .B1(n8550), .B2(n8539), .A(n9886), .ZN(n6152) );
  INV_X1 U7826 ( .A(n6152), .ZN(n6153) );
  AND2_X1 U7827 ( .A1(n4316), .A2(n6153), .ZN(n6154) );
  INV_X1 U7828 ( .A(n8533), .ZN(n8523) );
  NAND2_X1 U7829 ( .A1(n9899), .A2(n9892), .ZN(n9016) );
  OAI22_X1 U7830 ( .A1(n6185), .A2(n9018), .B1(n8523), .B2(n9016), .ZN(n6155)
         );
  INV_X1 U7831 ( .A(n6155), .ZN(n6157) );
  INV_X1 U7832 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6156) );
  NAND3_X1 U7833 ( .A1(n6158), .A2(n6157), .A3(n4824), .ZN(P2_U3455) );
  INV_X1 U7834 ( .A(n6182), .ZN(n6174) );
  INV_X1 U7835 ( .A(n6159), .ZN(n6160) );
  NAND2_X1 U7836 ( .A1(n6796), .A2(n8536), .ZN(n6678) );
  INV_X1 U7837 ( .A(n6797), .ZN(n6162) );
  NAND3_X1 U7838 ( .A1(n4316), .A2(n8550), .A3(n8322), .ZN(n6161) );
  NAND2_X1 U7839 ( .A1(n6178), .A2(n6175), .ZN(n6163) );
  NOR2_X1 U7840 ( .A1(n6176), .A2(n7406), .ZN(n9836) );
  INV_X1 U7841 ( .A(n9836), .ZN(n6166) );
  NAND2_X1 U7842 ( .A1(n6166), .A2(n9833), .ZN(n6167) );
  AOI22_X1 U7843 ( .A1(n8533), .A2(n8899), .B1(n8898), .B2(n8222), .ZN(n6171)
         );
  NAND2_X1 U7844 ( .A1(n9839), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7845 ( .B1(n6185), .B2(n8903), .A(n4844), .ZN(n6172) );
  INV_X1 U7846 ( .A(n6172), .ZN(n6173) );
  INV_X1 U7847 ( .A(n6175), .ZN(n6591) );
  INV_X1 U7848 ( .A(n6176), .ZN(n6177) );
  AOI21_X1 U7849 ( .B1(n6177), .B2(n9892), .A(n6797), .ZN(n6179) );
  MUX2_X1 U7850 ( .A(n6591), .B(n6179), .S(n6178), .Z(n6181) );
  NAND2_X1 U7851 ( .A1(n9913), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7852 ( .A1(n6184), .A2(n6183), .ZN(n6187) );
  NAND2_X1 U7853 ( .A1(n9915), .A2(n9892), .ZN(n8942) );
  OAI22_X1 U7854 ( .A1(n6185), .A2(n8943), .B1(n8523), .B2(n8942), .ZN(n6186)
         );
  OR2_X1 U7855 ( .A1(n6187), .A2(n6186), .ZN(P2_U3487) );
  OAI21_X1 U7856 ( .B1(n6508), .B2(n6504), .A(n7315), .ZN(n6188) );
  INV_X1 U7857 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7858 ( .A1(n6505), .A2(n7419), .ZN(n6190) );
  NAND2_X1 U7859 ( .A1(n6190), .A2(n6520), .ZN(n6191) );
  INV_X1 U7860 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7861 ( .A1(n6624), .A2(n6193), .ZN(n6214) );
  NAND2_X1 U7862 ( .A1(n6942), .A2(n6205), .ZN(n6194) );
  NAND2_X1 U7863 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  OAI22_X1 U7864 ( .A1(n6198), .A2(n4312), .B1(n7103), .B2(n6214), .ZN(n6210)
         );
  AND2_X1 U7865 ( .A1(n6200), .A2(n6199), .ZN(n6202) );
  INV_X1 U7866 ( .A(n6202), .ZN(n6208) );
  INV_X1 U7867 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7868 ( .A1(n6202), .A2(n4821), .ZN(n6940) );
  INV_X1 U7869 ( .A(n5517), .ZN(n6207) );
  INV_X1 U7870 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6203) );
  OAI21_X1 U7871 ( .B1(n6208), .B2(n6355), .A(n6939), .ZN(n7031) );
  NAND2_X1 U7872 ( .A1(n9270), .A2(n6205), .ZN(n6212) );
  NAND2_X1 U7873 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  OR2_X1 U7874 ( .A1(n7305), .A2(n9085), .ZN(n6216) );
  NAND2_X1 U7875 ( .A1(n7259), .A2(n6205), .ZN(n6215) );
  NAND2_X1 U7876 ( .A1(n6216), .A2(n6215), .ZN(n10101) );
  AOI22_X1 U7877 ( .A1(n7365), .A2(n7366), .B1(n10101), .B2(n7363), .ZN(n6218)
         );
  NAND2_X1 U7878 ( .A1(n7364), .A2(n6218), .ZN(n6225) );
  INV_X1 U7879 ( .A(n7363), .ZN(n6220) );
  INV_X1 U7880 ( .A(n10101), .ZN(n6219) );
  NAND2_X1 U7881 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  AOI21_X1 U7882 ( .B1(n6221), .B2(n7366), .A(n7365), .ZN(n6223) );
  NOR3_X1 U7883 ( .A1(n7363), .A2(n10101), .A3(n7366), .ZN(n6222) );
  NOR2_X1 U7884 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  NAND2_X1 U7885 ( .A1(n9269), .A2(n6372), .ZN(n6227) );
  OR2_X1 U7886 ( .A1(n7340), .A2(n6214), .ZN(n6226) );
  NAND2_X1 U7887 ( .A1(n6227), .A2(n6226), .ZN(n6232) );
  NAND2_X1 U7888 ( .A1(n9269), .A2(n6205), .ZN(n6229) );
  OR2_X1 U7889 ( .A1(n7340), .A2(n6234), .ZN(n6228) );
  NAND2_X1 U7890 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  XNOR2_X1 U7891 ( .A(n6230), .B(n6355), .ZN(n6231) );
  XOR2_X1 U7892 ( .A(n6232), .B(n6231), .Z(n7199) );
  NAND2_X1 U7893 ( .A1(n7200), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U7894 ( .A1(n6231), .A2(n6232), .ZN(n6233) );
  NAND2_X1 U7895 ( .A1(n7198), .A2(n6233), .ZN(n7504) );
  INV_X1 U7896 ( .A(n7504), .ZN(n6243) );
  OAI22_X1 U7897 ( .A1(n7575), .A2(n6264), .B1(n6234), .B2(n7568), .ZN(n6235)
         );
  XNOR2_X1 U7898 ( .A(n6235), .B(n9088), .ZN(n7563) );
  OR2_X1 U7899 ( .A1(n7575), .A2(n9085), .ZN(n6237) );
  NAND2_X1 U7900 ( .A1(n7458), .A2(n6205), .ZN(n6236) );
  AND2_X1 U7901 ( .A1(n6237), .A2(n6236), .ZN(n7562) );
  NOR2_X1 U7902 ( .A1(n7563), .A2(n7562), .ZN(n6244) );
  NAND2_X1 U7903 ( .A1(n9268), .A2(n6205), .ZN(n6239) );
  NAND2_X1 U7904 ( .A1(n6239), .A2(n6238), .ZN(n6240) );
  XNOR2_X1 U7905 ( .A(n6240), .B(n6355), .ZN(n7561) );
  NAND2_X1 U7906 ( .A1(n9268), .A2(n6372), .ZN(n6242) );
  OR2_X1 U7907 ( .A1(n7433), .A2(n6264), .ZN(n6241) );
  NAND2_X1 U7908 ( .A1(n6242), .A2(n6241), .ZN(n7505) );
  NAND2_X1 U7909 ( .A1(n7563), .A2(n7562), .ZN(n6245) );
  NAND2_X1 U7910 ( .A1(n9266), .A2(n6205), .ZN(n6248) );
  OR2_X1 U7911 ( .A1(n7767), .A2(n6234), .ZN(n6247) );
  NAND2_X1 U7912 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  XNOR2_X1 U7913 ( .A(n6249), .B(n6355), .ZN(n6251) );
  OAI22_X1 U7914 ( .A1(n7455), .A2(n9085), .B1(n7767), .B2(n6264), .ZN(n6250)
         );
  XNOR2_X1 U7915 ( .A(n6251), .B(n6250), .ZN(n7573) );
  AOI22_X1 U7916 ( .A1(n9265), .A2(n6205), .B1(n9092), .B2(n7639), .ZN(n6252)
         );
  XNOR2_X1 U7917 ( .A(n6252), .B(n6355), .ZN(n7631) );
  AOI22_X1 U7918 ( .A1(n9265), .A2(n6372), .B1(n6205), .B2(n7639), .ZN(n7630)
         );
  OAI22_X1 U7919 ( .A1(n7518), .A2(n9085), .B1(n9805), .B2(n6264), .ZN(n6254)
         );
  OAI22_X1 U7920 ( .A1(n7518), .A2(n6264), .B1(n6234), .B2(n9805), .ZN(n6253)
         );
  XNOR2_X1 U7921 ( .A(n6253), .B(n6355), .ZN(n6255) );
  XOR2_X1 U7922 ( .A(n6254), .B(n6255), .Z(n7857) );
  NAND2_X1 U7923 ( .A1(n7856), .A2(n7857), .ZN(n6257) );
  OR2_X1 U7924 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  NAND2_X1 U7925 ( .A1(n6257), .A2(n6256), .ZN(n9060) );
  OR2_X1 U7926 ( .A1(n7720), .A2(n9085), .ZN(n6259) );
  NAND2_X1 U7927 ( .A1(n9067), .A2(n6205), .ZN(n6258) );
  NAND2_X1 U7928 ( .A1(n6259), .A2(n6258), .ZN(n9061) );
  OAI22_X1 U7929 ( .A1(n7720), .A2(n6264), .B1(n6475), .B2(n6234), .ZN(n6260)
         );
  XNOR2_X1 U7930 ( .A(n6260), .B(n6355), .ZN(n6266) );
  NAND2_X1 U7931 ( .A1(n9662), .A2(n9092), .ZN(n6262) );
  NAND2_X1 U7932 ( .A1(n9262), .A2(n6205), .ZN(n6261) );
  NAND2_X1 U7933 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  XNOR2_X1 U7934 ( .A(n6263), .B(n6355), .ZN(n9206) );
  INV_X1 U7935 ( .A(n9662), .ZN(n7723) );
  OAI22_X1 U7936 ( .A1(n7723), .A2(n6264), .B1(n6477), .B2(n9085), .ZN(n6267)
         );
  AOI22_X1 U7937 ( .A1(n9061), .A2(n6266), .B1(n9206), .B2(n6267), .ZN(n6265)
         );
  NAND2_X1 U7938 ( .A1(n9060), .A2(n6265), .ZN(n6272) );
  INV_X1 U7939 ( .A(n9061), .ZN(n6269) );
  INV_X1 U7940 ( .A(n6267), .ZN(n9207) );
  AOI21_X1 U7941 ( .B1(n9205), .B2(n6269), .A(n9207), .ZN(n6268) );
  NAND3_X1 U7942 ( .A1(n9205), .A2(n6269), .A3(n9207), .ZN(n6270) );
  NAND2_X1 U7943 ( .A1(n6272), .A2(n4847), .ZN(n9116) );
  INV_X1 U7944 ( .A(n9124), .ZN(n7778) );
  OAI22_X1 U7945 ( .A1(n7778), .A2(n6264), .B1(n7721), .B2(n9085), .ZN(n6276)
         );
  NAND2_X1 U7946 ( .A1(n9124), .A2(n9092), .ZN(n6274) );
  NAND2_X1 U7947 ( .A1(n9261), .A2(n6205), .ZN(n6273) );
  NAND2_X1 U7948 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  XNOR2_X1 U7949 ( .A(n6275), .B(n6355), .ZN(n6277) );
  XOR2_X1 U7950 ( .A(n6276), .B(n6277), .Z(n9117) );
  OAI22_X1 U7951 ( .A1(n8049), .A2(n6264), .B1(n6482), .B2(n9085), .ZN(n6283)
         );
  NAND2_X1 U7952 ( .A1(n9190), .A2(n9092), .ZN(n6280) );
  NAND2_X1 U7953 ( .A1(n9260), .A2(n6205), .ZN(n6279) );
  NAND2_X1 U7954 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  XNOR2_X1 U7955 ( .A(n6281), .B(n6355), .ZN(n6282) );
  XOR2_X1 U7956 ( .A(n6283), .B(n6282), .Z(n9184) );
  INV_X1 U7957 ( .A(n6282), .ZN(n6285) );
  INV_X1 U7958 ( .A(n6283), .ZN(n6284) );
  INV_X1 U7959 ( .A(n9037), .ZN(n6289) );
  AOI22_X1 U7960 ( .A1(n9045), .A2(n9092), .B1(n6205), .B2(n9259), .ZN(n6286)
         );
  XNOR2_X1 U7961 ( .A(n6286), .B(n6355), .ZN(n9039) );
  INV_X1 U7962 ( .A(n9039), .ZN(n6288) );
  AOI22_X1 U7963 ( .A1(n9045), .A2(n6205), .B1(n6372), .B2(n9259), .ZN(n9038)
         );
  OAI21_X2 U7964 ( .B1(n6289), .B2(n6288), .A(n6287), .ZN(n6293) );
  OAI22_X1 U7965 ( .A1(n9648), .A2(n6234), .B1(n9137), .B2(n6264), .ZN(n6290)
         );
  XNOR2_X1 U7966 ( .A(n6290), .B(n6355), .ZN(n6291) );
  AOI22_X1 U7967 ( .A1(n9585), .A2(n6205), .B1(n6372), .B2(n9258), .ZN(n9233)
         );
  INV_X1 U7968 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U7969 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  NAND2_X1 U7970 ( .A1(n9231), .A2(n6294), .ZN(n9135) );
  INV_X1 U7971 ( .A(n9644), .ZN(n9557) );
  OAI22_X1 U7972 ( .A1(n9557), .A2(n6264), .B1(n9236), .B2(n9085), .ZN(n6299)
         );
  NAND2_X1 U7973 ( .A1(n9644), .A2(n9092), .ZN(n6296) );
  OR2_X1 U7974 ( .A1(n9236), .A2(n6214), .ZN(n6295) );
  NAND2_X1 U7975 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  XNOR2_X1 U7976 ( .A(n6297), .B(n6355), .ZN(n6298) );
  XOR2_X1 U7977 ( .A(n6299), .B(n6298), .Z(n9136) );
  INV_X1 U7978 ( .A(n6298), .ZN(n6301) );
  INV_X1 U7979 ( .A(n6299), .ZN(n6300) );
  NAND2_X1 U7980 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  OAI22_X1 U7981 ( .A1(n9537), .A2(n6234), .B1(n9221), .B2(n6264), .ZN(n6303)
         );
  XNOR2_X1 U7982 ( .A(n6303), .B(n6355), .ZN(n6308) );
  OR2_X1 U7983 ( .A1(n9537), .A2(n6264), .ZN(n6305) );
  OR2_X1 U7984 ( .A1(n9221), .A2(n9085), .ZN(n6304) );
  NAND2_X1 U7985 ( .A1(n6305), .A2(n6304), .ZN(n6307) );
  XNOR2_X1 U7986 ( .A(n6308), .B(n6307), .ZN(n9145) );
  AOI22_X1 U7987 ( .A1(n9697), .A2(n9092), .B1(n6205), .B2(n9256), .ZN(n6306)
         );
  XOR2_X1 U7988 ( .A(n6355), .B(n6306), .Z(n9073) );
  NAND2_X1 U7989 ( .A1(n6308), .A2(n6307), .ZN(n9072) );
  INV_X1 U7990 ( .A(n9072), .ZN(n6309) );
  NOR2_X1 U7991 ( .A1(n9073), .A2(n6309), .ZN(n6310) );
  INV_X1 U7992 ( .A(n9697), .ZN(n9529) );
  OAI22_X1 U7993 ( .A1(n9529), .A2(n6264), .B1(n6311), .B2(n9085), .ZN(n9219)
         );
  NAND2_X1 U7994 ( .A1(n9070), .A2(n9219), .ZN(n9167) );
  OAI22_X1 U7995 ( .A1(n9505), .A2(n6234), .B1(n9223), .B2(n6264), .ZN(n6312)
         );
  XNOR2_X1 U7996 ( .A(n6312), .B(n9088), .ZN(n6326) );
  INV_X1 U7997 ( .A(n6326), .ZN(n6316) );
  OR2_X1 U7998 ( .A1(n9505), .A2(n6264), .ZN(n6314) );
  OR2_X1 U7999 ( .A1(n9223), .A2(n9085), .ZN(n6313) );
  AND2_X1 U8000 ( .A1(n6314), .A2(n6313), .ZN(n6325) );
  INV_X1 U8001 ( .A(n6325), .ZN(n6315) );
  NAND2_X1 U8002 ( .A1(n6316), .A2(n6315), .ZN(n9076) );
  AND2_X1 U8003 ( .A1(n9072), .A2(n9076), .ZN(n9168) );
  INV_X1 U8004 ( .A(n9625), .ZN(n9493) );
  OAI22_X1 U8005 ( .A1(n9493), .A2(n6264), .B1(n6317), .B2(n9085), .ZN(n6327)
         );
  AOI22_X1 U8006 ( .A1(n9625), .A2(n9092), .B1(n6205), .B2(n9254), .ZN(n6318)
         );
  XNOR2_X1 U8007 ( .A(n6318), .B(n6355), .ZN(n6329) );
  XOR2_X1 U8008 ( .A(n6327), .B(n6329), .Z(n9177) );
  INV_X1 U8009 ( .A(n9177), .ZN(n6319) );
  AND2_X1 U8010 ( .A1(n9168), .A2(n6319), .ZN(n6320) );
  NAND2_X1 U8011 ( .A1(n9071), .A2(n6320), .ZN(n6323) );
  INV_X1 U8012 ( .A(n9076), .ZN(n6321) );
  OR2_X1 U8013 ( .A1(n6321), .A2(n9073), .ZN(n9169) );
  OR2_X1 U8014 ( .A1(n9177), .A2(n9169), .ZN(n6322) );
  NAND2_X1 U8015 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U8016 ( .A1(n9167), .A2(n6324), .ZN(n9175) );
  NAND2_X1 U8017 ( .A1(n6326), .A2(n6325), .ZN(n9172) );
  OR2_X1 U8018 ( .A1(n9177), .A2(n9172), .ZN(n9174) );
  INV_X1 U8019 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U8020 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  AND2_X1 U8021 ( .A1(n9174), .A2(n6330), .ZN(n6331) );
  NAND2_X1 U8022 ( .A1(n9175), .A2(n6331), .ZN(n9107) );
  INV_X1 U8023 ( .A(n9618), .ZN(n9486) );
  OAI22_X1 U8024 ( .A1(n9486), .A2(n6264), .B1(n9195), .B2(n9085), .ZN(n6336)
         );
  NAND2_X1 U8025 ( .A1(n9618), .A2(n9092), .ZN(n6333) );
  OR2_X1 U8026 ( .A1(n9195), .A2(n6264), .ZN(n6332) );
  NAND2_X1 U8027 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  XNOR2_X1 U8028 ( .A(n6334), .B(n6355), .ZN(n6335) );
  XOR2_X1 U8029 ( .A(n6336), .B(n6335), .Z(n9108) );
  NAND2_X1 U8030 ( .A1(n9107), .A2(n9108), .ZN(n6340) );
  INV_X1 U8031 ( .A(n6335), .ZN(n6338) );
  INV_X1 U8032 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U8033 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  NAND2_X1 U8034 ( .A1(n6340), .A2(n6339), .ZN(n6344) );
  OAI22_X1 U8035 ( .A1(n9463), .A2(n6234), .B1(n9109), .B2(n6264), .ZN(n6341)
         );
  XNOR2_X1 U8036 ( .A(n6341), .B(n6196), .ZN(n6342) );
  XNOR2_X1 U8037 ( .A(n6344), .B(n6342), .ZN(n9193) );
  INV_X1 U8038 ( .A(n9109), .ZN(n9252) );
  AOI22_X1 U8039 ( .A1(n9614), .A2(n6205), .B1(n6372), .B2(n9252), .ZN(n9194)
         );
  NAND2_X1 U8040 ( .A1(n9193), .A2(n9194), .ZN(n9048) );
  NAND2_X1 U8041 ( .A1(n6344), .A2(n6343), .ZN(n9050) );
  NAND2_X1 U8042 ( .A1(n9609), .A2(n9092), .ZN(n6346) );
  NAND2_X1 U8043 ( .A1(n9251), .A2(n6205), .ZN(n6345) );
  NAND2_X1 U8044 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U8045 ( .A(n6347), .B(n6196), .ZN(n6362) );
  INV_X1 U8046 ( .A(n6362), .ZN(n6351) );
  NAND2_X1 U8047 ( .A1(n9609), .A2(n6205), .ZN(n6349) );
  NAND2_X1 U8048 ( .A1(n9251), .A2(n6372), .ZN(n6348) );
  NAND2_X1 U8049 ( .A1(n6349), .A2(n6348), .ZN(n6361) );
  INV_X1 U8050 ( .A(n6361), .ZN(n6350) );
  NAND2_X1 U8051 ( .A1(n6351), .A2(n6350), .ZN(n9051) );
  AND2_X1 U8052 ( .A1(n9050), .A2(n9051), .ZN(n6352) );
  NAND2_X1 U8053 ( .A1(n9048), .A2(n6352), .ZN(n9155) );
  NAND2_X1 U8054 ( .A1(n9678), .A2(n9092), .ZN(n6354) );
  NAND2_X1 U8055 ( .A1(n9250), .A2(n6205), .ZN(n6353) );
  NAND2_X1 U8056 ( .A1(n6354), .A2(n6353), .ZN(n6356) );
  XNOR2_X1 U8057 ( .A(n6356), .B(n6355), .ZN(n6360) );
  NAND2_X1 U8058 ( .A1(n9678), .A2(n6205), .ZN(n6358) );
  NAND2_X1 U8059 ( .A1(n9250), .A2(n6372), .ZN(n6357) );
  NAND2_X1 U8060 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NOR2_X1 U8061 ( .A1(n6360), .A2(n6359), .ZN(n6364) );
  AOI21_X1 U8062 ( .B1(n6360), .B2(n6359), .A(n6364), .ZN(n9158) );
  NAND2_X1 U8063 ( .A1(n6362), .A2(n6361), .ZN(n9154) );
  AND2_X1 U8064 ( .A1(n9158), .A2(n9154), .ZN(n6363) );
  NAND2_X1 U8065 ( .A1(n9155), .A2(n6363), .ZN(n9156) );
  INV_X1 U8066 ( .A(n6364), .ZN(n6365) );
  OAI22_X1 U8067 ( .A1(n9427), .A2(n6214), .B1(n9159), .B2(n4312), .ZN(n6367)
         );
  OAI22_X1 U8068 ( .A1(n9427), .A2(n6234), .B1(n9159), .B2(n6264), .ZN(n6366)
         );
  XNOR2_X1 U8069 ( .A(n6366), .B(n6196), .ZN(n6368) );
  XOR2_X1 U8070 ( .A(n6367), .B(n6368), .Z(n9129) );
  INV_X1 U8071 ( .A(n9127), .ZN(n6374) );
  NOR2_X1 U8072 ( .A1(n6368), .A2(n6367), .ZN(n6375) );
  NAND2_X1 U8073 ( .A1(n9669), .A2(n9092), .ZN(n6370) );
  NAND2_X1 U8074 ( .A1(n9249), .A2(n6205), .ZN(n6369) );
  NAND2_X1 U8075 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  XNOR2_X1 U8076 ( .A(n6371), .B(n9088), .ZN(n6421) );
  AND2_X1 U8077 ( .A1(n9249), .A2(n6372), .ZN(n6373) );
  AOI21_X1 U8078 ( .B1(n9669), .B2(n6205), .A(n6373), .ZN(n6422) );
  XNOR2_X1 U8079 ( .A(n6421), .B(n6422), .ZN(n6376) );
  OAI21_X1 U8080 ( .B1(n6374), .B2(n6375), .A(n6376), .ZN(n6401) );
  NOR2_X1 U8081 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  NAND2_X1 U8082 ( .A1(n7923), .A2(P1_B_REG_SCAN_IN), .ZN(n6380) );
  MUX2_X1 U8083 ( .A(P1_B_REG_SCAN_IN), .B(n6380), .S(n7814), .Z(n6381) );
  INV_X1 U8084 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8085 ( .A1(n6453), .A2(n6382), .ZN(n6384) );
  INV_X1 U8086 ( .A(n6383), .ZN(n8022) );
  NAND2_X1 U8087 ( .A1(n8022), .A2(n7814), .ZN(n9721) );
  NOR4_X1 U8088 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6388) );
  NOR4_X1 U8089 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6387) );
  NOR4_X1 U8090 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6386) );
  NOR4_X1 U8091 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6385) );
  AND4_X1 U8092 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n6394)
         );
  NOR2_X1 U8093 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .ZN(
        n6392) );
  NOR4_X1 U8094 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6391) );
  NOR4_X1 U8095 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6390) );
  NOR4_X1 U8096 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6389) );
  AND4_X1 U8097 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .ZN(n6393)
         );
  NAND2_X1 U8098 ( .A1(n6394), .A2(n6393), .ZN(n6452) );
  INV_X1 U8099 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6395) );
  OR2_X1 U8100 ( .A1(n6452), .A2(n6395), .ZN(n7109) );
  INV_X1 U8101 ( .A(n7109), .ZN(n6396) );
  NAND2_X1 U8102 ( .A1(n8022), .A2(n7923), .ZN(n9720) );
  OAI21_X1 U8103 ( .B1(n7107), .B2(n6396), .A(n9720), .ZN(n6397) );
  INV_X1 U8104 ( .A(n6397), .ZN(n6398) );
  INV_X1 U8105 ( .A(n6627), .ZN(n6412) );
  NAND2_X1 U8106 ( .A1(n6412), .A2(n9804), .ZN(n6404) );
  NOR2_X1 U8107 ( .A1(n7110), .A2(n6404), .ZN(n6400) );
  NAND3_X1 U8108 ( .A1(n6401), .A2(n6434), .A3(n6436), .ZN(n6420) );
  INV_X1 U8109 ( .A(n9669), .ZN(n9410) );
  OR2_X1 U8110 ( .A1(n7117), .A2(n7402), .ZN(n7115) );
  NOR2_X1 U8111 ( .A1(n7110), .A2(n7115), .ZN(n6402) );
  NAND2_X1 U8112 ( .A1(n6415), .A2(n6402), .ZN(n6403) );
  OR2_X1 U8113 ( .A1(n7117), .A2(n6507), .ZN(n6450) );
  INV_X1 U8114 ( .A(n6415), .ZN(n6409) );
  NAND2_X1 U8115 ( .A1(n6404), .A2(n7115), .ZN(n6405) );
  NAND2_X1 U8116 ( .A1(n6409), .A2(n6405), .ZN(n6406) );
  NAND2_X1 U8117 ( .A1(n6627), .A2(n6504), .ZN(n7111) );
  NAND4_X1 U8118 ( .A1(n6406), .A2(n6624), .A3(n6626), .A4(n7111), .ZN(n6407)
         );
  NAND2_X1 U8119 ( .A1(n6407), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6411) );
  INV_X1 U8120 ( .A(n7116), .ZN(n6408) );
  NAND3_X1 U8121 ( .A1(n6409), .A2(n7108), .A3(n6408), .ZN(n6410) );
  INV_X1 U8122 ( .A(n8105), .ZN(n9248) );
  NAND2_X1 U8123 ( .A1(n5672), .A2(n6627), .ZN(n9235) );
  NOR2_X2 U8124 ( .A1(n5672), .A2(n6412), .ZN(n9237) );
  NOR2_X1 U8125 ( .A1(n9159), .A2(n9220), .ZN(n6413) );
  AOI21_X1 U8126 ( .B1(n9248), .B2(n9196), .A(n6413), .ZN(n9405) );
  NOR2_X1 U8127 ( .A1(n7110), .A2(n6504), .ZN(n6414) );
  NAND2_X1 U8128 ( .A1(n6415), .A2(n6414), .ZN(n10098) );
  OAI22_X1 U8129 ( .A1(n9405), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10036), .ZN(n6416) );
  AOI21_X1 U8130 ( .B1(n9411), .B2(n9242), .A(n6416), .ZN(n6417) );
  INV_X1 U8131 ( .A(n6418), .ZN(n6419) );
  NAND2_X1 U8132 ( .A1(n6420), .A2(n6419), .ZN(P1_U3240) );
  INV_X1 U8133 ( .A(n6421), .ZN(n6424) );
  INV_X1 U8134 ( .A(n6422), .ZN(n6423) );
  NAND2_X1 U8135 ( .A1(n6525), .A2(n9092), .ZN(n6426) );
  NAND2_X1 U8136 ( .A1(n9248), .A2(n6205), .ZN(n6425) );
  NAND2_X1 U8137 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  XNOR2_X1 U8138 ( .A(n6427), .B(n9088), .ZN(n6430) );
  NOR2_X1 U8139 ( .A1(n8105), .A2(n9085), .ZN(n6428) );
  AOI21_X1 U8140 ( .B1(n6525), .B2(n6205), .A(n6428), .ZN(n6429) );
  NAND2_X1 U8141 ( .A1(n6430), .A2(n6429), .ZN(n9099) );
  OAI21_X1 U8142 ( .B1(n6430), .B2(n6429), .A(n9099), .ZN(n6432) );
  NAND2_X1 U8143 ( .A1(n6431), .A2(n6432), .ZN(n6435) );
  NOR2_X1 U8144 ( .A1(n6432), .A2(n4381), .ZN(n6433) );
  NAND2_X1 U8145 ( .A1(n6435), .A2(n9105), .ZN(n6437) );
  NAND2_X1 U8146 ( .A1(n6437), .A2(n6436), .ZN(n6445) );
  INV_X1 U8147 ( .A(n6438), .ZN(n9390) );
  OR2_X1 U8148 ( .A1(n9090), .A2(n9235), .ZN(n6440) );
  NAND2_X1 U8149 ( .A1(n9249), .A2(n9237), .ZN(n6439) );
  AND2_X1 U8150 ( .A1(n6440), .A2(n6439), .ZN(n6523) );
  OAI22_X1 U8151 ( .A1(n6523), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9978), .ZN(n6441) );
  AOI21_X1 U8152 ( .B1(n9390), .B2(n9242), .A(n6441), .ZN(n6442) );
  OAI21_X1 U8153 ( .B1(n9393), .B2(n10096), .A(n6442), .ZN(n6443) );
  INV_X1 U8154 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8155 ( .A1(n6445), .A2(n6444), .ZN(P1_U3214) );
  INV_X1 U8156 ( .A(n7321), .ZN(n7369) );
  INV_X1 U8157 ( .A(n7340), .ZN(n9787) );
  NAND2_X1 U8158 ( .A1(n7527), .A2(n6475), .ZN(n7526) );
  INV_X1 U8159 ( .A(n9678), .ZN(n9441) );
  NAND2_X1 U8160 ( .A1(n9422), .A2(n9427), .ZN(n9408) );
  INV_X1 U8161 ( .A(n9380), .ZN(n8107) );
  XOR2_X1 U8162 ( .A(n4338), .B(n9370), .Z(n6448) );
  NAND2_X1 U8163 ( .A1(n6448), .A2(n6447), .ZN(n9372) );
  INV_X1 U8164 ( .A(n5673), .ZN(n9735) );
  AND2_X1 U8165 ( .A1(n9735), .A2(P1_B_REG_SCAN_IN), .ZN(n6449) );
  NOR2_X1 U8166 ( .A1(n9235), .A2(n6449), .ZN(n8124) );
  NAND2_X1 U8167 ( .A1(n6699), .A2(n8124), .ZN(n9367) );
  NAND2_X1 U8168 ( .A1(n7111), .A2(n6450), .ZN(n6451) );
  NOR2_X1 U8169 ( .A1(n7110), .A2(n6451), .ZN(n6456) );
  OAI21_X1 U8170 ( .B1(n7107), .B2(P1_D_REG_1__SCAN_IN), .A(n9720), .ZN(n6455)
         );
  NAND2_X1 U8171 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  MUX2_X1 U8172 ( .A(n9591), .B(n6457), .S(n9809), .Z(n6458) );
  INV_X1 U8173 ( .A(n9370), .ZN(n9593) );
  NAND2_X1 U8174 ( .A1(n6458), .A2(n4831), .ZN(P1_U3521) );
  INV_X1 U8175 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6527) );
  INV_X1 U8176 ( .A(n9269), .ZN(n7306) );
  NAND2_X1 U8177 ( .A1(n7201), .A2(n7321), .ZN(n7326) );
  INV_X1 U8178 ( .A(n7328), .ZN(n6459) );
  NOR2_X1 U8179 ( .A1(n4845), .A2(n6459), .ZN(n6463) );
  NAND2_X1 U8180 ( .A1(n5517), .A2(n6943), .ZN(n7093) );
  NAND2_X1 U8181 ( .A1(n7091), .A2(n7093), .ZN(n7092) );
  NAND2_X1 U8182 ( .A1(n6198), .A2(n7103), .ZN(n6460) );
  NAND2_X1 U8183 ( .A1(n7092), .A2(n6460), .ZN(n7252) );
  NAND2_X1 U8184 ( .A1(n7252), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U8185 ( .A1(n7305), .A2(n10097), .ZN(n6461) );
  NAND2_X1 U8186 ( .A1(n7250), .A2(n6461), .ZN(n7300) );
  AND2_X1 U8187 ( .A1(n7334), .A2(n7303), .ZN(n6462) );
  NAND2_X1 U8188 ( .A1(n7300), .A2(n6462), .ZN(n7329) );
  NAND2_X1 U8189 ( .A1(n6463), .A2(n7329), .ZN(n7423) );
  NAND2_X1 U8190 ( .A1(n7423), .A2(n7425), .ZN(n7422) );
  NAND2_X1 U8191 ( .A1(n7454), .A2(n7433), .ZN(n7449) );
  NAND2_X1 U8192 ( .A1(n7575), .A2(n7568), .ZN(n6464) );
  AND2_X1 U8193 ( .A1(n7449), .A2(n6464), .ZN(n6468) );
  INV_X1 U8194 ( .A(n6464), .ZN(n6467) );
  NAND2_X1 U8195 ( .A1(n6466), .A2(n6465), .ZN(n7452) );
  NAND2_X1 U8196 ( .A1(n7455), .A2(n7767), .ZN(n6469) );
  NAND2_X1 U8197 ( .A1(n7753), .A2(n6469), .ZN(n7619) );
  NAND2_X1 U8198 ( .A1(n6470), .A2(n7646), .ZN(n7618) );
  NAND2_X1 U8199 ( .A1(n7619), .A2(n7618), .ZN(n7617) );
  NAND2_X1 U8200 ( .A1(n7651), .A2(n9796), .ZN(n6471) );
  NAND2_X1 U8201 ( .A1(n7617), .A2(n6471), .ZN(n7642) );
  NAND2_X1 U8202 ( .A1(n6473), .A2(n6472), .ZN(n7648) );
  NAND2_X1 U8203 ( .A1(n7642), .A2(n7648), .ZN(n7644) );
  NAND2_X1 U8204 ( .A1(n7518), .A2(n9805), .ZN(n6474) );
  NAND2_X1 U8205 ( .A1(n7644), .A2(n6474), .ZN(n7524) );
  NAND2_X1 U8206 ( .A1(n7524), .A2(n7523), .ZN(n7522) );
  NAND2_X1 U8207 ( .A1(n7720), .A2(n6475), .ZN(n6476) );
  NAND2_X1 U8208 ( .A1(n7522), .A2(n6476), .ZN(n7713) );
  NAND2_X1 U8209 ( .A1(n9262), .A2(n9662), .ZN(n6478) );
  OR2_X1 U8210 ( .A1(n9124), .A2(n9261), .ZN(n6479) );
  NAND2_X1 U8211 ( .A1(n7771), .A2(n6479), .ZN(n6481) );
  OR2_X1 U8212 ( .A1(n7778), .A2(n7721), .ZN(n6480) );
  NAND2_X1 U8213 ( .A1(n9554), .A2(n9553), .ZN(n9552) );
  NAND2_X1 U8214 ( .A1(n9552), .A2(n4839), .ZN(n9535) );
  NAND2_X1 U8215 ( .A1(n9537), .A2(n9221), .ZN(n6486) );
  INV_X1 U8216 ( .A(n9221), .ZN(n9257) );
  NAND2_X1 U8217 ( .A1(n9697), .A2(n9256), .ZN(n6488) );
  NOR2_X1 U8218 ( .A1(n9697), .A2(n9256), .ZN(n6487) );
  NAND2_X1 U8219 ( .A1(n9505), .A2(n9223), .ZN(n6490) );
  NOR2_X1 U8220 ( .A1(n9505), .A2(n9223), .ZN(n6489) );
  NAND2_X1 U8221 ( .A1(n9625), .A2(n9254), .ZN(n6491) );
  INV_X1 U8222 ( .A(n9195), .ZN(n9253) );
  NAND2_X1 U8223 ( .A1(n9463), .A2(n9109), .ZN(n6492) );
  NAND2_X1 U8224 ( .A1(n9609), .A2(n9251), .ZN(n6493) );
  NAND2_X1 U8225 ( .A1(n9446), .A2(n6493), .ZN(n6496) );
  NAND2_X1 U8226 ( .A1(n4514), .A2(n6494), .ZN(n6495) );
  NAND2_X1 U8227 ( .A1(n9678), .A2(n9250), .ZN(n6497) );
  INV_X1 U8228 ( .A(n9398), .ZN(n6498) );
  NOR2_X1 U8229 ( .A1(n9427), .A2(n9159), .ZN(n9399) );
  AND2_X1 U8230 ( .A1(n9669), .A2(n9249), .ZN(n6501) );
  NAND2_X1 U8231 ( .A1(n6498), .A2(n4851), .ZN(n6503) );
  OR2_X1 U8232 ( .A1(n9669), .A2(n9249), .ZN(n6499) );
  NAND2_X1 U8233 ( .A1(n9427), .A2(n9159), .ZN(n9400) );
  AND2_X1 U8234 ( .A1(n6499), .A2(n9400), .ZN(n6500) );
  XNOR2_X1 U8235 ( .A(n8095), .B(n8094), .ZN(n9388) );
  NAND2_X1 U8236 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  NAND3_X1 U8237 ( .A1(n7116), .A2(n7117), .A3(n6506), .ZN(n8063) );
  OR2_X1 U8238 ( .A1(n6508), .A2(n6507), .ZN(n9781) );
  INV_X1 U8239 ( .A(n8094), .ZN(n6519) );
  NAND2_X1 U8240 ( .A1(n6512), .A2(n6511), .ZN(n9467) );
  NAND2_X1 U8241 ( .A1(n9467), .A2(n9466), .ZN(n9465) );
  NAND2_X1 U8242 ( .A1(n9465), .A2(n6513), .ZN(n9448) );
  OAI21_X1 U8243 ( .B1(n6519), .B2(n6518), .A(n8100), .ZN(n6522) );
  OR2_X1 U8244 ( .A1(n7582), .A2(n5620), .ZN(n6521) );
  NAND2_X1 U8245 ( .A1(n6522), .A2(n9575), .ZN(n6524) );
  NAND2_X1 U8246 ( .A1(n6524), .A2(n6523), .ZN(n9395) );
  AOI211_X1 U8247 ( .C1(n6525), .C2(n9409), .A(n9579), .B(n8108), .ZN(n9389)
         );
  AOI21_X1 U8248 ( .B1(n9388), .B2(n9801), .A(n6526), .ZN(n6533) );
  MUX2_X1 U8249 ( .A(n6527), .B(n6533), .S(n9713), .Z(n6530) );
  NAND2_X1 U8250 ( .A1(n6525), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8251 ( .A1(n6530), .A2(n6529), .ZN(P1_U3517) );
  MUX2_X1 U8252 ( .A(n6534), .B(n6533), .S(n9818), .Z(n6537) );
  NAND2_X1 U8253 ( .A1(n6525), .A2(n6535), .ZN(n6536) );
  NAND2_X1 U8254 ( .A1(n6537), .A2(n6536), .ZN(P1_U3549) );
  NAND2_X1 U8255 ( .A1(n6539), .A2(n6538), .ZN(n6541) );
  NAND2_X1 U8256 ( .A1(n6541), .A2(n6540), .ZN(n8316) );
  OR2_X1 U8257 ( .A1(n4314), .A2(n9032), .ZN(n6542) );
  NAND2_X1 U8258 ( .A1(n6543), .A2(n8225), .ZN(n8302) );
  NAND2_X1 U8259 ( .A1(n8355), .A2(n8302), .ZN(n8532) );
  AND2_X1 U8260 ( .A1(n4310), .A2(P2_B_REG_SCAN_IN), .ZN(n6544) );
  NOR2_X1 U8261 ( .A1(n8866), .A2(n6544), .ZN(n8732) );
  INV_X1 U8262 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U8263 ( .A1(n5738), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6547) );
  INV_X1 U8264 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6545) );
  OR2_X1 U8265 ( .A1(n4315), .A2(n6545), .ZN(n6546) );
  OAI211_X1 U8266 ( .C1(n6548), .C2(n4307), .A(n6547), .B(n6546), .ZN(n6549)
         );
  INV_X1 U8267 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8268 ( .A1(n8313), .A2(n6550), .ZN(n8556) );
  AOI22_X1 U8269 ( .A1(n8742), .A2(n9826), .B1(n8732), .B2(n8556), .ZN(n6551)
         );
  NAND2_X1 U8270 ( .A1(n8523), .A2(n8524), .ZN(n6553) );
  AOI21_X1 U8271 ( .B1(n6554), .B2(n6553), .A(n6552), .ZN(n6555) );
  XNOR2_X1 U8272 ( .A(n6555), .B(n8532), .ZN(n6556) );
  NAND2_X1 U8273 ( .A1(n6556), .A2(n9829), .ZN(n6557) );
  INV_X1 U8274 ( .A(n9874), .ZN(n6559) );
  NAND2_X1 U8275 ( .A1(n8163), .A2(n6561), .ZN(n6565) );
  INV_X1 U8276 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8277 ( .A1(n9913), .A2(n6562), .ZN(n6563) );
  OAI21_X1 U8278 ( .B1(n6565), .B2(n9913), .A(n6563), .ZN(n6564) );
  NAND2_X1 U8279 ( .A1(n6564), .A2(n4832), .ZN(P2_U3488) );
  OAI21_X1 U8280 ( .B1(n6565), .B2(n9901), .A(n4820), .ZN(n6566) );
  NAND2_X1 U8281 ( .A1(n6566), .A2(n4822), .ZN(P2_U3456) );
  INV_X1 U8282 ( .A(n6567), .ZN(n6568) );
  NAND2_X1 U8283 ( .A1(n6680), .A2(n8522), .ZN(n6569) );
  NAND2_X1 U8284 ( .A1(n6569), .A2(n6654), .ZN(n6644) );
  NAND2_X1 U8285 ( .A1(n6644), .A2(n6642), .ZN(n6570) );
  NAND2_X1 U8286 ( .A1(n6570), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8287 ( .A(n6687), .ZN(n6571) );
  NAND2_X1 U8288 ( .A1(n6572), .A2(P2_U3151), .ZN(n9031) );
  AND2_X1 U8289 ( .A1(n4907), .A2(P2_U3151), .ZN(n7691) );
  INV_X2 U8290 ( .A(n7691), .ZN(n9034) );
  OAI222_X1 U8291 ( .A1(n9031), .A2(n4887), .B1(n9034), .B2(n6580), .C1(
        P2_U3151), .C2(n6704), .ZN(P2_U3294) );
  INV_X1 U8292 ( .A(n9031), .ZN(n8090) );
  INV_X1 U8293 ( .A(n8090), .ZN(n9025) );
  OAI222_X1 U8294 ( .A1(n9025), .A2(n6573), .B1(n9034), .B2(n6586), .C1(
        P2_U3151), .C2(n6963), .ZN(P2_U3290) );
  OAI222_X1 U8295 ( .A1(n9025), .A2(n4566), .B1(n9034), .B2(n6590), .C1(
        P2_U3151), .C2(n4289), .ZN(P2_U3293) );
  OAI222_X1 U8296 ( .A1(n9025), .A2(n6574), .B1(n9034), .B2(n6584), .C1(
        P2_U3151), .C2(n6727), .ZN(P2_U3292) );
  OAI222_X1 U8297 ( .A1(n9025), .A2(n6575), .B1(n9034), .B2(n6588), .C1(
        P2_U3151), .C2(n7074), .ZN(P2_U3289) );
  OAI222_X1 U8298 ( .A1(n9025), .A2(n6576), .B1(n9034), .B2(n6582), .C1(
        P2_U3151), .C2(n6859), .ZN(P2_U3291) );
  INV_X1 U8299 ( .A(n6577), .ZN(n6595) );
  OAI222_X1 U8300 ( .A1(n9025), .A2(n6578), .B1(n9034), .B2(n6595), .C1(
        P2_U3151), .C2(n7205), .ZN(P2_U3288) );
  NAND2_X1 U8301 ( .A1(n6572), .A2(P1_U3086), .ZN(n9732) );
  NAND2_X1 U8302 ( .A1(n4907), .A2(P1_U3086), .ZN(n9729) );
  AOI22_X1 U8303 ( .A1(n9723), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9276), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6579) );
  OAI21_X1 U8304 ( .B1(n6580), .B2(n9732), .A(n6579), .ZN(P1_U3354) );
  INV_X1 U8305 ( .A(n9732), .ZN(n7694) );
  AOI22_X1 U8306 ( .A1(n9318), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9723), .ZN(n6581) );
  OAI21_X1 U8307 ( .B1(n6582), .B2(n9728), .A(n6581), .ZN(P1_U3351) );
  AOI22_X1 U8308 ( .A1(n9304), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9723), .ZN(n6583) );
  OAI21_X1 U8309 ( .B1(n6584), .B2(n9728), .A(n6583), .ZN(P1_U3352) );
  AOI22_X1 U8310 ( .A1(n6887), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9723), .ZN(n6585) );
  OAI21_X1 U8311 ( .B1(n6586), .B2(n9728), .A(n6585), .ZN(P1_U3350) );
  AOI22_X1 U8312 ( .A1(n6874), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9723), .ZN(n6587) );
  OAI21_X1 U8313 ( .B1(n6588), .B2(n9732), .A(n6587), .ZN(P1_U3349) );
  AOI22_X1 U8314 ( .A1(n9291), .A2(P1_STATE_REG_SCAN_IN), .B1(n9723), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n6589) );
  OAI21_X1 U8315 ( .B1(n6590), .B2(n9728), .A(n6589), .ZN(P1_U3353) );
  INV_X1 U8316 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8317 ( .A1(n6591), .A2(n6600), .ZN(n6592) );
  OAI21_X1 U8318 ( .B1(n6600), .B2(n6593), .A(n6592), .ZN(P2_U3377) );
  AOI22_X1 U8319 ( .A1(n6914), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9723), .ZN(n6594) );
  OAI21_X1 U8320 ( .B1(n6595), .B2(n9732), .A(n6594), .ZN(P1_U3348) );
  INV_X1 U8321 ( .A(n6596), .ZN(n6598) );
  INV_X1 U8322 ( .A(n6935), .ZN(n6597) );
  OAI222_X1 U8323 ( .A1(n9729), .A2(n9977), .B1(n9728), .B2(n6598), .C1(
        P1_U3086), .C2(n6597), .ZN(P1_U3347) );
  OAI222_X1 U8324 ( .A1(n9031), .A2(n6599), .B1(n9034), .B2(n6598), .C1(
        P2_U3151), .C2(n7497), .ZN(P2_U3287) );
  INV_X1 U8325 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6603) );
  INV_X1 U8326 ( .A(n6601), .ZN(n6602) );
  AOI22_X1 U8327 ( .A1(n6611), .A2(n6603), .B1(n6602), .B2(n6687), .ZN(
        P2_U3376) );
  OAI222_X1 U8328 ( .A1(n9729), .A2(n6604), .B1(n9728), .B2(n6605), .C1(
        P1_U3086), .C2(n4542), .ZN(P1_U3346) );
  INV_X1 U8329 ( .A(n7545), .ZN(n7537) );
  OAI222_X1 U8330 ( .A1(n9031), .A2(n6606), .B1(n9034), .B2(n6605), .C1(
        P2_U3151), .C2(n7537), .ZN(P2_U3286) );
  INV_X1 U8331 ( .A(n6607), .ZN(n6610) );
  OAI222_X1 U8332 ( .A1(n9034), .A2(n6610), .B1(n7549), .B2(P2_U3151), .C1(
        n6608), .C2(n9031), .ZN(P2_U3285) );
  AND2_X1 U8333 ( .A1(n6611), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8334 ( .A1(n6611), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8335 ( .A1(n6611), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8336 ( .A1(n6611), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8337 ( .A1(n6611), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8338 ( .A1(n6611), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8339 ( .A1(n6611), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8340 ( .A1(n6611), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8341 ( .A1(n6611), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8342 ( .A1(n6611), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8343 ( .A1(n6611), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8344 ( .A1(n6611), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8345 ( .A1(n6611), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8346 ( .A1(n6611), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8347 ( .A1(n6611), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8348 ( .A1(n6611), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8349 ( .A1(n6611), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8350 ( .A1(n6611), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8351 ( .A1(n6611), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8352 ( .A1(n6611), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8353 ( .A1(n6611), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8354 ( .A1(n6611), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8355 ( .A1(n6611), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8356 ( .A1(n6611), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8357 ( .A1(n6611), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8358 ( .A1(n6611), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8359 ( .A1(n6611), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8360 ( .A1(n6611), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  OAI222_X1 U8361 ( .A1(n9729), .A2(n6621), .B1(n9728), .B2(n6610), .C1(n6609), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8362 ( .A(n6611), .ZN(n6612) );
  INV_X1 U8363 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U8364 ( .A1(n6612), .A2(n10083), .ZN(P2_U3252) );
  INV_X1 U8365 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U8366 ( .A1(n6612), .A2(n10048), .ZN(P2_U3263) );
  INV_X1 U8367 ( .A(n6613), .ZN(n6617) );
  AOI22_X1 U8368 ( .A1(n7017), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9723), .ZN(n6614) );
  OAI21_X1 U8369 ( .B1(n6617), .B2(n9728), .A(n6614), .ZN(P1_U3344) );
  MUX2_X1 U8370 ( .A(n6615), .B(n7292), .S(P2_U3893), .Z(n6616) );
  INV_X1 U8371 ( .A(n6616), .ZN(P2_U3497) );
  INV_X1 U8372 ( .A(n7825), .ZN(n7832) );
  OAI222_X1 U8373 ( .A1(n9031), .A2(n6618), .B1(n9034), .B2(n6617), .C1(
        P2_U3151), .C2(n7832), .ZN(P2_U3284) );
  MUX2_X1 U8374 ( .A(n6619), .B(n7794), .S(P2_U3893), .Z(n6620) );
  INV_X1 U8375 ( .A(n6620), .ZN(P2_U3502) );
  MUX2_X1 U8376 ( .A(n6621), .B(n8426), .S(P2_U3893), .Z(n6622) );
  INV_X1 U8377 ( .A(n6622), .ZN(P2_U3501) );
  INV_X1 U8378 ( .A(n6626), .ZN(n6623) );
  OR2_X1 U8379 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  AND2_X1 U8380 ( .A1(n6625), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6775) );
  NAND2_X1 U8381 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  NAND2_X1 U8382 ( .A1(n6629), .A2(n6628), .ZN(n6774) );
  NOR2_X1 U8383 ( .A1(n9739), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8384 ( .A(n6630), .ZN(n6632) );
  INV_X1 U8385 ( .A(n7831), .ZN(n7952) );
  OAI222_X1 U8386 ( .A1(n9034), .A2(n6632), .B1(n7952), .B2(P2_U3151), .C1(
        n6631), .C2(n9031), .ZN(P2_U3283) );
  OAI222_X1 U8387 ( .A1(n9729), .A2(n6633), .B1(n9728), .B2(n6632), .C1(n7022), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8388 ( .A(n6634), .ZN(n6673) );
  AOI22_X1 U8389 ( .A1(n7380), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9723), .ZN(n6635) );
  OAI21_X1 U8390 ( .B1(n6673), .B2(n9728), .A(n6635), .ZN(P1_U3342) );
  INV_X1 U8391 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8392 ( .A1(n8566), .A2(n6637), .ZN(n8371) );
  NAND2_X1 U8393 ( .A1(n7055), .A2(n8371), .ZN(n8332) );
  OAI21_X1 U8394 ( .B1(n9829), .B2(n9895), .A(n8332), .ZN(n6636) );
  NAND2_X1 U8395 ( .A1(n5704), .A2(n9824), .ZN(n6815) );
  OAI211_X1 U8396 ( .C1(n6637), .C2(n9886), .A(n6636), .B(n6815), .ZN(n6663)
         );
  NAND2_X1 U8397 ( .A1(n6663), .A2(n9899), .ZN(n6638) );
  OAI21_X1 U8398 ( .B1(n6639), .B2(n9899), .A(n6638), .ZN(P2_U3390) );
  AND2_X1 U8399 ( .A1(n6644), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6641) );
  MUX2_X1 U8400 ( .A(n6641), .B(P2_U3893), .S(n6640), .Z(n6643) );
  NAND2_X1 U8401 ( .A1(n6643), .A2(n4309), .ZN(n8724) );
  NOR2_X1 U8402 ( .A1(n6090), .A2(P2_U3151), .ZN(n8089) );
  NAND2_X1 U8403 ( .A1(n5719), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6722) );
  INV_X1 U8404 ( .A(n6646), .ZN(n6647) );
  INV_X1 U8405 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6645) );
  OAI21_X1 U8406 ( .B1(n6647), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6723), .ZN(
        n6658) );
  INV_X1 U8407 ( .A(n6648), .ZN(n6665) );
  AND2_X1 U8408 ( .A1(n6649), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8409 ( .A1(n5719), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6713) );
  INV_X1 U8410 ( .A(n6714), .ZN(n6651) );
  AOI21_X1 U8411 ( .B1(n7060), .B2(n6652), .A(n6651), .ZN(n6653) );
  OAI22_X1 U8412 ( .A1(n8731), .A2(n6653), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6810), .ZN(n6657) );
  INV_X1 U8413 ( .A(n6654), .ZN(n6829) );
  NOR2_X1 U8414 ( .A1(n6680), .A2(n6829), .ZN(n6655) );
  INV_X1 U8415 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U8416 ( .A1(n8704), .A2(n9920), .ZN(n6656) );
  AOI211_X1 U8417 ( .C1(n8727), .C2(n6658), .A(n6657), .B(n6656), .ZN(n6662)
         );
  MUX2_X1 U8418 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6091), .Z(n6705) );
  XOR2_X1 U8419 ( .A(n6704), .B(n6705), .Z(n6660) );
  MUX2_X1 U8420 ( .A(n5705), .B(n5706), .S(n6091), .Z(n6667) );
  NAND2_X1 U8421 ( .A1(n6667), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8422 ( .A1(n6660), .A2(n6666), .ZN(n6706) );
  NAND2_X1 U8423 ( .A1(P2_U3893), .A2(n6090), .ZN(n8719) );
  OAI211_X1 U8424 ( .C1(n6660), .C2(n6666), .A(n6706), .B(n8664), .ZN(n6661)
         );
  OAI211_X1 U8425 ( .C1(n8724), .C2(n6704), .A(n6662), .B(n6661), .ZN(P2_U3183) );
  NAND2_X1 U8426 ( .A1(n6663), .A2(n9915), .ZN(n6664) );
  OAI21_X1 U8427 ( .B1(n9915), .B2(n5706), .A(n6664), .ZN(P2_U3459) );
  INV_X1 U8428 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8429 ( .A1(n8676), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8430 ( .A1(n6665), .A2(n8719), .ZN(n6669) );
  OAI21_X1 U8431 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6667), .A(n6666), .ZN(n6668) );
  AOI22_X1 U8432 ( .A1(n6669), .A2(n6668), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6670) );
  OAI211_X1 U8433 ( .C1(n8704), .C2(n6672), .A(n6671), .B(n6670), .ZN(P2_U3182) );
  INV_X1 U8434 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10008) );
  OAI222_X1 U8435 ( .A1(n9031), .A2(n10008), .B1(n9034), .B2(n6673), .C1(
        P2_U3151), .C2(n7955), .ZN(P2_U3282) );
  OAI21_X1 U8436 ( .B1(n6676), .B2(n6675), .A(n6674), .ZN(n6681) );
  INV_X1 U8437 ( .A(n6691), .ZN(n6677) );
  NAND2_X1 U8438 ( .A1(n6682), .A2(n6677), .ZN(n6679) );
  NAND4_X1 U8439 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6686)
         );
  INV_X1 U8440 ( .A(n6682), .ZN(n6684) );
  OR2_X1 U8441 ( .A1(n6814), .A2(n6683), .ZN(n8549) );
  NOR2_X1 U8442 ( .A1(n6684), .A2(n8549), .ZN(n6685) );
  AOI21_X1 U8443 ( .B1(n6686), .B2(P2_STATE_REG_SCAN_IN), .A(n6685), .ZN(n6830) );
  AND2_X1 U8444 ( .A1(n6830), .A2(n6687), .ZN(n6828) );
  INV_X1 U8445 ( .A(n6688), .ZN(n6689) );
  NAND2_X1 U8446 ( .A1(n6690), .A2(n6689), .ZN(n6693) );
  OR2_X1 U8447 ( .A1(n6695), .A2(n6691), .ZN(n6692) );
  OAI21_X2 U8448 ( .B1(n6694), .B2(n9886), .A(n9821), .ZN(n8228) );
  AOI22_X1 U8449 ( .A1(n8285), .A2(n8332), .B1(n6813), .B2(n8228), .ZN(n6697)
         );
  NOR2_X1 U8450 ( .A1(n6695), .A2(n6814), .ZN(n6794) );
  NAND2_X1 U8451 ( .A1(n6794), .A2(n6792), .ZN(n8290) );
  NAND2_X1 U8452 ( .A1(n8266), .A2(n5704), .ZN(n6696) );
  OAI211_X1 U8453 ( .C1(n6828), .C2(n6698), .A(n6697), .B(n6696), .ZN(P2_U3172) );
  NAND2_X1 U8454 ( .A1(n6699), .A2(P1_U3973), .ZN(n6700) );
  OAI21_X1 U8455 ( .B1(P1_U3973), .B2(n9026), .A(n6700), .ZN(P1_U3585) );
  INV_X1 U8456 ( .A(n6701), .ZN(n6762) );
  AOI22_X1 U8457 ( .A1(n7703), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9723), .ZN(n6702) );
  OAI21_X1 U8458 ( .B1(n6762), .B2(n9732), .A(n6702), .ZN(P1_U3341) );
  NAND2_X1 U8459 ( .A1(n5517), .A2(P1_U3973), .ZN(n6703) );
  OAI21_X1 U8460 ( .B1(P1_U3973), .B2(n5711), .A(n6703), .ZN(P1_U3554) );
  MUX2_X1 U8461 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6091), .Z(n6736) );
  XNOR2_X1 U8462 ( .A(n6736), .B(n6727), .ZN(n6712) );
  INV_X1 U8463 ( .A(n4289), .ZN(n8579) );
  MUX2_X1 U8464 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6091), .Z(n6709) );
  INV_X1 U8465 ( .A(n6709), .ZN(n6710) );
  INV_X1 U8466 ( .A(n6704), .ZN(n6708) );
  INV_X1 U8467 ( .A(n6705), .ZN(n6707) );
  OAI21_X1 U8468 ( .B1(n6708), .B2(n6707), .A(n6706), .ZN(n8569) );
  XOR2_X1 U8469 ( .A(n4289), .B(n6709), .Z(n8568) );
  NAND2_X1 U8470 ( .A1(n8569), .A2(n8568), .ZN(n8567) );
  OAI21_X1 U8471 ( .B1(n8579), .B2(n6710), .A(n8567), .ZN(n6711) );
  NOR2_X1 U8472 ( .A1(n6711), .A2(n6712), .ZN(n6737) );
  AOI21_X1 U8473 ( .B1(n6712), .B2(n6711), .A(n6737), .ZN(n6735) );
  NAND2_X1 U8474 ( .A1(n6714), .A2(n6713), .ZN(n8571) );
  XNOR2_X1 U8475 ( .A(n4289), .B(n6715), .ZN(n8572) );
  NAND2_X1 U8476 ( .A1(n8571), .A2(n8572), .ZN(n8570) );
  NAND2_X1 U8477 ( .A1(n4289), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8478 ( .A1(n8570), .A2(n6716), .ZN(n6717) );
  INV_X1 U8479 ( .A(n6746), .ZN(n6718) );
  AOI21_X1 U8480 ( .B1(n5727), .B2(n6719), .A(n6718), .ZN(n6721) );
  NOR2_X1 U8481 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7184), .ZN(n6840) );
  INV_X1 U8482 ( .A(n6840), .ZN(n6720) );
  OAI21_X1 U8483 ( .B1(n8731), .B2(n6721), .A(n6720), .ZN(n6733) );
  INV_X1 U8484 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U8485 ( .A1(n6723), .A2(n6722), .ZN(n8576) );
  INV_X1 U8486 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6724) );
  XNOR2_X1 U8487 ( .A(n6725), .B(n6724), .ZN(n8577) );
  NAND2_X1 U8488 ( .A1(n8576), .A2(n8577), .ZN(n8575) );
  NAND2_X1 U8489 ( .A1(n4289), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6726) );
  INV_X1 U8490 ( .A(n6755), .ZN(n6728) );
  AOI21_X1 U8491 ( .B1(n10082), .B2(n6729), .A(n6728), .ZN(n6731) );
  INV_X1 U8492 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6730) );
  OAI22_X1 U8493 ( .A1(n8689), .A2(n6731), .B1(n8704), .B2(n6730), .ZN(n6732)
         );
  AOI211_X1 U8494 ( .C1(n4691), .C2(n8676), .A(n6733), .B(n6732), .ZN(n6734)
         );
  OAI21_X1 U8495 ( .B1(n6735), .B2(n8719), .A(n6734), .ZN(P2_U3185) );
  INV_X1 U8496 ( .A(n6736), .ZN(n6738) );
  MUX2_X1 U8497 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6091), .Z(n6845) );
  XOR2_X1 U8498 ( .A(n6859), .B(n6845), .Z(n6739) );
  OAI211_X1 U8499 ( .C1(n6740), .C2(n6739), .A(n6846), .B(n8664), .ZN(n6760)
         );
  INV_X1 U8500 ( .A(n8704), .ZN(n8721) );
  INV_X1 U8501 ( .A(n6742), .ZN(n6741) );
  MUX2_X1 U8502 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5740), .S(n6859), .Z(n6743)
         );
  NOR2_X1 U8503 ( .A1(n6741), .A2(n6743), .ZN(n6747) );
  NAND2_X1 U8504 ( .A1(n6744), .A2(n6743), .ZN(n6854) );
  INV_X1 U8505 ( .A(n6854), .ZN(n6745) );
  AOI21_X1 U8506 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(n6750) );
  NOR2_X1 U8507 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6748), .ZN(n7004) );
  INV_X1 U8508 ( .A(n7004), .ZN(n6749) );
  OAI21_X1 U8509 ( .B1(n8731), .B2(n6750), .A(n6749), .ZN(n6758) );
  NAND2_X1 U8510 ( .A1(n6755), .A2(n6753), .ZN(n6751) );
  INV_X1 U8511 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9904) );
  MUX2_X1 U8512 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9904), .S(n6859), .Z(n6752)
         );
  NAND2_X1 U8513 ( .A1(n6751), .A2(n6752), .ZN(n6861) );
  INV_X1 U8514 ( .A(n6752), .ZN(n6754) );
  NAND3_X1 U8515 ( .A1(n6755), .A2(n6754), .A3(n6753), .ZN(n6756) );
  AOI21_X1 U8516 ( .B1(n6861), .B2(n6756), .A(n8689), .ZN(n6757) );
  AOI211_X1 U8517 ( .C1(n8721), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6758), .B(
        n6757), .ZN(n6759) );
  OAI211_X1 U8518 ( .C1(n8724), .C2(n6859), .A(n6760), .B(n6759), .ZN(P2_U3186) );
  NAND2_X1 U8519 ( .A1(n9272), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6761) );
  OAI21_X1 U8520 ( .B1(n9236), .B2(n9272), .A(n6761), .ZN(P1_U3570) );
  INV_X1 U8521 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6763) );
  OAI222_X1 U8522 ( .A1(n9031), .A2(n6763), .B1(n9034), .B2(n6762), .C1(
        P2_U3151), .C2(n8622), .ZN(P2_U3281) );
  INV_X1 U8523 ( .A(n6764), .ZN(n6811) );
  AOI22_X1 U8524 ( .A1(n8646), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8090), .ZN(n6765) );
  OAI21_X1 U8525 ( .B1(n6811), .B2(n9034), .A(n6765), .ZN(P2_U3280) );
  NOR2_X1 U8526 ( .A1(n6898), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6766) );
  AOI21_X1 U8527 ( .B1(n6898), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6766), .ZN(
        n6773) );
  INV_X1 U8528 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9811) );
  MUX2_X1 U8529 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9811), .S(n9291), .Z(n9297)
         );
  INV_X1 U8530 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7102) );
  MUX2_X1 U8531 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7102), .S(n9276), .Z(n9275)
         );
  AND2_X1 U8532 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9274) );
  NAND2_X1 U8533 ( .A1(n9275), .A2(n9274), .ZN(n9273) );
  NAND2_X1 U8534 ( .A1(n9276), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U8535 ( .A1(n9273), .A2(n6767), .ZN(n9296) );
  NAND2_X1 U8536 ( .A1(n9297), .A2(n9296), .ZN(n9295) );
  NAND2_X1 U8537 ( .A1(n9291), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8538 ( .A1(n9295), .A2(n6768), .ZN(n9309) );
  INV_X1 U8539 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6769) );
  XNOR2_X1 U8540 ( .A(n9304), .B(n6769), .ZN(n9310) );
  NAND2_X1 U8541 ( .A1(n9309), .A2(n9310), .ZN(n9308) );
  NAND2_X1 U8542 ( .A1(n9304), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U8543 ( .A1(n9308), .A2(n6770), .ZN(n9320) );
  INV_X1 U8544 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9990) );
  MUX2_X1 U8545 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9990), .S(n9318), .Z(n9321)
         );
  NAND2_X1 U8546 ( .A1(n9320), .A2(n9321), .ZN(n9319) );
  XNOR2_X1 U8547 ( .A(n6887), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6885) );
  XNOR2_X1 U8548 ( .A(n6874), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U8549 ( .A1(n4355), .A2(n6873), .ZN(n6872) );
  AOI21_X1 U8550 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6874), .A(n6872), .ZN(
        n6913) );
  NAND2_X1 U8551 ( .A1(n6914), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6771) );
  OAI21_X1 U8552 ( .B1(n6914), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6771), .ZN(
        n6912) );
  NOR2_X1 U8553 ( .A1(n6913), .A2(n6912), .ZN(n6911) );
  AOI21_X1 U8554 ( .B1(n6914), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6911), .ZN(
        n6924) );
  XNOR2_X1 U8555 ( .A(n6935), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6925) );
  OAI21_X1 U8556 ( .B1(n6773), .B2(n6772), .A(n6893), .ZN(n6779) );
  INV_X1 U8557 ( .A(n6774), .ZN(n6776) );
  NAND2_X1 U8558 ( .A1(n6776), .A2(n6775), .ZN(n9741) );
  INV_X1 U8559 ( .A(n5672), .ZN(n9285) );
  NOR2_X2 U8560 ( .A1(n9741), .A2(n9285), .ZN(n9359) );
  INV_X1 U8561 ( .A(n9359), .ZN(n7907) );
  NAND2_X1 U8562 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U8563 ( .A1(n9739), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6777) );
  OAI211_X1 U8564 ( .C1(n7907), .C2(n4542), .A(n7861), .B(n6777), .ZN(n6778)
         );
  AOI21_X1 U8565 ( .B1(n6779), .B2(n9354), .A(n6778), .ZN(n6791) );
  NOR2_X1 U8566 ( .A1(n6898), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6780) );
  AOI21_X1 U8567 ( .B1(n6898), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6780), .ZN(
        n6787) );
  MUX2_X1 U8568 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n4901), .S(n9291), .Z(n9294)
         );
  AND2_X1 U8569 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9284) );
  NAND2_X1 U8570 ( .A1(n9278), .A2(n9284), .ZN(n9277) );
  NAND2_X1 U8571 ( .A1(n9276), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U8572 ( .A1(n9277), .A2(n6781), .ZN(n9293) );
  NAND2_X1 U8573 ( .A1(n9294), .A2(n9293), .ZN(n9292) );
  NAND2_X1 U8574 ( .A1(n9291), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8575 ( .A1(n9292), .A2(n6782), .ZN(n9306) );
  XNOR2_X1 U8576 ( .A(n9304), .B(n6783), .ZN(n9307) );
  NAND2_X1 U8577 ( .A1(n9306), .A2(n9307), .ZN(n9305) );
  NAND2_X1 U8578 ( .A1(n9304), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6784) );
  MUX2_X1 U8579 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7337), .S(n9318), .Z(n9324)
         );
  XNOR2_X1 U8580 ( .A(n6887), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6882) );
  NOR2_X1 U8581 ( .A1(n6883), .A2(n6882), .ZN(n6881) );
  AOI21_X1 U8582 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6887), .A(n6881), .ZN(
        n6871) );
  XNOR2_X1 U8583 ( .A(n6874), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6870) );
  NOR2_X1 U8584 ( .A1(n6871), .A2(n6870), .ZN(n6869) );
  AOI21_X1 U8585 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6874), .A(n6869), .ZN(
        n6910) );
  NAND2_X1 U8586 ( .A1(n6914), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6785) );
  OAI21_X1 U8587 ( .B1(n6914), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6785), .ZN(
        n6909) );
  XNOR2_X1 U8588 ( .A(n6935), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8589 ( .A1(n6786), .A2(n6787), .ZN(n6897) );
  OAI21_X1 U8590 ( .B1(n6787), .B2(n6786), .A(n6897), .ZN(n6789) );
  NAND2_X1 U8591 ( .A1(n9285), .A2(n9735), .ZN(n6788) );
  NOR2_X2 U8592 ( .A1(n9741), .A2(n6788), .ZN(n9360) );
  NAND2_X1 U8593 ( .A1(n6789), .A2(n9360), .ZN(n6790) );
  NAND2_X1 U8594 ( .A1(n6791), .A2(n6790), .ZN(P1_U3252) );
  INV_X1 U8595 ( .A(n8228), .ZN(n8296) );
  INV_X1 U8596 ( .A(n6792), .ZN(n6793) );
  NAND2_X1 U8597 ( .A1(n6794), .A2(n6793), .ZN(n8268) );
  OAI22_X1 U8598 ( .A1(n5703), .A2(n8296), .B1(n8268), .B2(n6132), .ZN(n6795)
         );
  AOI21_X1 U8599 ( .B1(n8266), .B2(n8565), .A(n6795), .ZN(n6809) );
  NAND2_X1 U8600 ( .A1(n8539), .A2(n8370), .ZN(n8543) );
  AND2_X1 U8601 ( .A1(n6796), .A2(n8543), .ZN(n6799) );
  XNOR2_X1 U8602 ( .A(n8946), .B(n6803), .ZN(n6801) );
  NAND2_X1 U8603 ( .A1(n6801), .A2(n6800), .ZN(n6820) );
  INV_X1 U8604 ( .A(n6803), .ZN(n6834) );
  OR2_X1 U8605 ( .A1(n6803), .A2(n6813), .ZN(n6804) );
  NAND2_X1 U8606 ( .A1(n7055), .A2(n6804), .ZN(n6806) );
  OAI21_X1 U8607 ( .B1(n6805), .B2(n6806), .A(n6821), .ZN(n6807) );
  NAND2_X1 U8608 ( .A1(n6807), .A2(n8285), .ZN(n6808) );
  OAI211_X1 U8609 ( .C1(n6828), .C2(n6810), .A(n6809), .B(n6808), .ZN(P2_U3162) );
  OAI222_X1 U8610 ( .A1(n9729), .A2(n6812), .B1(n9728), .B2(n6811), .C1(
        P1_U3086), .C2(n7732), .ZN(P1_U3340) );
  AOI22_X1 U8611 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n9839), .B1(n8899), .B2(
        n6813), .ZN(n6819) );
  NAND3_X1 U8612 ( .A1(n8332), .A2(n9886), .A3(n6814), .ZN(n6816) );
  OAI211_X1 U8613 ( .C1(n6698), .C2(n9821), .A(n6816), .B(n6815), .ZN(n6817)
         );
  NAND2_X1 U8614 ( .A1(n6817), .A2(n9837), .ZN(n6818) );
  NAND2_X1 U8615 ( .A1(n6819), .A2(n6818), .ZN(P2_U3233) );
  XNOR2_X1 U8616 ( .A(n6803), .B(n8377), .ZN(n6831) );
  XNOR2_X1 U8617 ( .A(n6831), .B(n8565), .ZN(n6823) );
  NAND2_X1 U8618 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  NAND2_X1 U8619 ( .A1(n6822), .A2(n6823), .ZN(n6833) );
  OAI21_X1 U8620 ( .B1(n6823), .B2(n6822), .A(n6833), .ZN(n6824) );
  NAND2_X1 U8621 ( .A1(n6824), .A2(n8285), .ZN(n6827) );
  INV_X1 U8622 ( .A(n8376), .ZN(n9825) );
  OAI22_X1 U8623 ( .A1(n9841), .A2(n8296), .B1(n8268), .B2(n6800), .ZN(n6825)
         );
  AOI21_X1 U8624 ( .B1(n8266), .B2(n9825), .A(n6825), .ZN(n6826) );
  OAI211_X1 U8625 ( .C1(n6828), .C2(n9822), .A(n6827), .B(n6826), .ZN(P2_U3177) );
  NAND2_X1 U8626 ( .A1(n6829), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8553) );
  INV_X1 U8627 ( .A(n8565), .ZN(n8378) );
  NAND2_X1 U8628 ( .A1(n6831), .A2(n8378), .ZN(n6832) );
  INV_X2 U8629 ( .A(n6834), .ZN(n8219) );
  XNOR2_X1 U8630 ( .A(n6835), .B(n8219), .ZN(n6993) );
  AOI21_X1 U8631 ( .B1(n6836), .B2(n6837), .A(n8272), .ZN(n6838) );
  NAND2_X1 U8632 ( .A1(n6838), .A2(n6996), .ZN(n6844) );
  AOI21_X1 U8633 ( .B1(n8228), .B2(n6835), .A(n6840), .ZN(n6841) );
  OAI21_X1 U8634 ( .B1(n8290), .B2(n5750), .A(n6841), .ZN(n6842) );
  AOI21_X1 U8635 ( .B1(n8288), .B2(n8565), .A(n6842), .ZN(n6843) );
  OAI211_X1 U8636 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8223), .A(n6844), .B(
        n6843), .ZN(P2_U3158) );
  INV_X1 U8637 ( .A(n6859), .ZN(n6848) );
  INV_X1 U8638 ( .A(n6845), .ZN(n6847) );
  MUX2_X1 U8639 ( .A(n6850), .B(n6849), .S(n6091), .Z(n6965) );
  XNOR2_X1 U8640 ( .A(n6965), .B(n6963), .ZN(n6851) );
  OAI211_X1 U8641 ( .C1(n6852), .C2(n6851), .A(n6964), .B(n8664), .ZN(n6868)
         );
  NAND2_X1 U8642 ( .A1(n6859), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8643 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  INV_X1 U8644 ( .A(n6979), .ZN(n6856) );
  AOI21_X1 U8645 ( .B1(n6850), .B2(n6857), .A(n6856), .ZN(n6858) );
  NAND2_X1 U8646 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7046) );
  OAI21_X1 U8647 ( .B1(n6858), .B2(n8731), .A(n7046), .ZN(n6866) );
  NAND2_X1 U8648 ( .A1(n6859), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8649 ( .A1(n6861), .A2(n6860), .ZN(n6862) );
  NAND2_X1 U8650 ( .A1(n6863), .A2(n6849), .ZN(n6864) );
  AOI21_X1 U8651 ( .B1(n6973), .B2(n6864), .A(n8689), .ZN(n6865) );
  AOI211_X1 U8652 ( .C1(n8721), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6866), .B(
        n6865), .ZN(n6867) );
  OAI211_X1 U8653 ( .C1(n8724), .C2(n6963), .A(n6868), .B(n6867), .ZN(P2_U3187) );
  AOI211_X1 U8654 ( .C1(n6871), .C2(n6870), .A(n6869), .B(n7376), .ZN(n6880)
         );
  AOI211_X1 U8655 ( .C1(n4355), .C2(n6873), .A(n6872), .B(n9356), .ZN(n6879)
         );
  INV_X1 U8656 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U8657 ( .A1(n9359), .A2(n6874), .ZN(n6876) );
  NAND2_X1 U8658 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6875) );
  OAI211_X1 U8659 ( .C1(n6877), .C2(n9366), .A(n6876), .B(n6875), .ZN(n6878)
         );
  OR3_X1 U8660 ( .A1(n6880), .A2(n6879), .A3(n6878), .ZN(P1_U3249) );
  AOI211_X1 U8661 ( .C1(n6883), .C2(n6882), .A(n6881), .B(n7376), .ZN(n6892)
         );
  AOI211_X1 U8662 ( .C1(n6886), .C2(n6885), .A(n6884), .B(n9356), .ZN(n6891)
         );
  INV_X1 U8663 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U8664 ( .A1(n9359), .A2(n6887), .ZN(n6889) );
  NAND2_X1 U8665 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n6888) );
  OAI211_X1 U8666 ( .C1(n10019), .C2(n9366), .A(n6889), .B(n6888), .ZN(n6890)
         );
  OR3_X1 U8667 ( .A1(n6892), .A2(n6891), .A3(n6890), .ZN(P1_U3248) );
  INV_X1 U8668 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6894) );
  MUX2_X1 U8669 ( .A(n6894), .B(P1_REG1_REG_10__SCAN_IN), .S(n6953), .Z(n6895)
         );
  NOR2_X1 U8670 ( .A1(n6895), .A2(n6896), .ZN(n6952) );
  AOI211_X1 U8671 ( .C1(n6896), .C2(n6895), .A(n6952), .B(n9356), .ZN(n6907)
         );
  OAI21_X1 U8672 ( .B1(n6898), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6897), .ZN(
        n6901) );
  NAND2_X1 U8673 ( .A1(n6953), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6899) );
  OAI21_X1 U8674 ( .B1(n6953), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6899), .ZN(
        n6900) );
  NOR2_X1 U8675 ( .A1(n6900), .A2(n6901), .ZN(n6948) );
  AOI211_X1 U8676 ( .C1(n6901), .C2(n6900), .A(n6948), .B(n7376), .ZN(n6906)
         );
  INV_X1 U8677 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8678 ( .A1(n9359), .A2(n6953), .ZN(n6903) );
  NAND2_X1 U8679 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n6902) );
  OAI211_X1 U8680 ( .C1(n6904), .C2(n9366), .A(n6903), .B(n6902), .ZN(n6905)
         );
  OR3_X1 U8681 ( .A1(n6907), .A2(n6906), .A3(n6905), .ZN(P1_U3253) );
  AOI211_X1 U8682 ( .C1(n6910), .C2(n6909), .A(n7376), .B(n6908), .ZN(n6919)
         );
  AOI211_X1 U8683 ( .C1(n6913), .C2(n6912), .A(n9356), .B(n6911), .ZN(n6918)
         );
  INV_X1 U8684 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U8685 ( .A1(n9359), .A2(n6914), .ZN(n6916) );
  NAND2_X1 U8686 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6915) );
  OAI211_X1 U8687 ( .C1(n10069), .C2(n9366), .A(n6916), .B(n6915), .ZN(n6917)
         );
  OR3_X1 U8688 ( .A1(n6919), .A2(n6918), .A3(n6917), .ZN(P1_U3250) );
  INV_X1 U8689 ( .A(n6920), .ZN(n6923) );
  OAI222_X1 U8690 ( .A1(n9034), .A2(n6923), .B1(n8670), .B2(P2_U3151), .C1(
        n6921), .C2(n9025), .ZN(P2_U3279) );
  OAI222_X1 U8691 ( .A1(P1_U3086), .A2(n7739), .B1(n9732), .B2(n6923), .C1(
        n6922), .C2(n9729), .ZN(P1_U3339) );
  INV_X1 U8692 ( .A(n6924), .ZN(n6927) );
  INV_X1 U8693 ( .A(n6925), .ZN(n6926) );
  OAI21_X1 U8694 ( .B1(n6927), .B2(n6926), .A(n9354), .ZN(n6937) );
  INV_X1 U8695 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8696 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n6928) );
  OAI21_X1 U8697 ( .B1(n9366), .B2(n6929), .A(n6928), .ZN(n6934) );
  AOI211_X1 U8698 ( .C1(n6932), .C2(n6931), .A(n7376), .B(n6930), .ZN(n6933)
         );
  AOI211_X1 U8699 ( .C1(n9359), .C2(n6935), .A(n6934), .B(n6933), .ZN(n6936)
         );
  OAI21_X1 U8700 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(P1_U3251) );
  OAI21_X1 U8701 ( .B1(n6941), .B2(n6940), .A(n6939), .ZN(n9283) );
  NAND2_X1 U8702 ( .A1(n6942), .A2(n9196), .ZN(n7119) );
  NAND2_X1 U8703 ( .A1(n9228), .A2(n6943), .ZN(n6944) );
  NAND2_X1 U8704 ( .A1(P1_U3086), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9737) );
  OAI211_X1 U8705 ( .C1(n10098), .C2(n7119), .A(n6944), .B(n9737), .ZN(n6945)
         );
  AOI21_X1 U8706 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9242), .A(n6945), .ZN(
        n6946) );
  OAI21_X1 U8707 ( .B1(n9283), .B2(n10103), .A(n6946), .ZN(P1_U3232) );
  NAND2_X1 U8708 ( .A1(n9272), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6947) );
  OAI21_X1 U8709 ( .B1(n9159), .B2(n9272), .A(n6947), .ZN(P1_U3579) );
  NAND2_X1 U8710 ( .A1(n7017), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6949) );
  OAI21_X1 U8711 ( .B1(n7017), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6949), .ZN(
        n6950) );
  AOI211_X1 U8712 ( .C1(n6951), .C2(n6950), .A(n7012), .B(n7376), .ZN(n6962)
         );
  MUX2_X1 U8713 ( .A(n6954), .B(P1_REG1_REG_11__SCAN_IN), .S(n7017), .Z(n6955)
         );
  AOI211_X1 U8714 ( .C1(n6956), .C2(n6955), .A(n7016), .B(n9356), .ZN(n6961)
         );
  INV_X1 U8715 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U8716 ( .A1(n9359), .A2(n7017), .ZN(n6958) );
  NAND2_X1 U8717 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n6957) );
  OAI211_X1 U8718 ( .C1(n6959), .C2(n9366), .A(n6958), .B(n6957), .ZN(n6960)
         );
  OR3_X1 U8719 ( .A1(n6962), .A2(n6961), .A3(n6960), .ZN(P1_U3254) );
  MUX2_X1 U8720 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6091), .Z(n7066) );
  XNOR2_X1 U8721 ( .A(n7066), .B(n7074), .ZN(n6967) );
  OAI21_X1 U8722 ( .B1(n4682), .B2(n6965), .A(n6964), .ZN(n6966) );
  NOR2_X1 U8723 ( .A1(n6966), .A2(n6967), .ZN(n7067) );
  AOI21_X1 U8724 ( .B1(n6967), .B2(n6966), .A(n7067), .ZN(n6989) );
  INV_X1 U8725 ( .A(n7074), .ZN(n7069) );
  INV_X1 U8726 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6986) );
  INV_X1 U8727 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6968) );
  XNOR2_X1 U8728 ( .A(n7074), .B(n6968), .ZN(n6970) );
  NAND2_X1 U8729 ( .A1(n6969), .A2(n6970), .ZN(n7076) );
  INV_X1 U8730 ( .A(n6970), .ZN(n6972) );
  NAND3_X1 U8731 ( .A1(n6973), .A2(n6972), .A3(n6971), .ZN(n6974) );
  AOI21_X1 U8732 ( .B1(n7076), .B2(n6974), .A(n8689), .ZN(n6982) );
  XNOR2_X1 U8733 ( .A(n7074), .B(n8150), .ZN(n6976) );
  NAND2_X1 U8734 ( .A1(n6975), .A2(n6976), .ZN(n7071) );
  INV_X1 U8735 ( .A(n6976), .ZN(n6978) );
  NAND3_X1 U8736 ( .A1(n6979), .A2(n6978), .A3(n6977), .ZN(n6980) );
  AOI21_X1 U8737 ( .B1(n7071), .B2(n6980), .A(n8731), .ZN(n6981) );
  NOR2_X1 U8738 ( .A1(n6982), .A2(n6981), .ZN(n6985) );
  INV_X1 U8739 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U8740 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6983), .ZN(n7265) );
  INV_X1 U8741 ( .A(n7265), .ZN(n6984) );
  OAI211_X1 U8742 ( .C1(n8704), .C2(n6986), .A(n6985), .B(n6984), .ZN(n6987)
         );
  AOI21_X1 U8743 ( .B1(n7069), .B2(n8676), .A(n6987), .ZN(n6988) );
  OAI21_X1 U8744 ( .B1(n6989), .B2(n8719), .A(n6988), .ZN(P2_U3188) );
  INV_X1 U8745 ( .A(n6990), .ZN(n7118) );
  OAI21_X1 U8746 ( .B1(n9575), .B2(n9801), .A(n7118), .ZN(n6991) );
  OAI211_X1 U8747 ( .C1(n7117), .C2(n7125), .A(n6991), .B(n7119), .ZN(n9666)
         );
  NAND2_X1 U8748 ( .A1(n9666), .A2(n9713), .ZN(n6992) );
  OAI21_X1 U8749 ( .B1(n9794), .B2(n4893), .A(n6992), .ZN(P1_U3453) );
  INV_X1 U8750 ( .A(n6993), .ZN(n6994) );
  NAND2_X1 U8751 ( .A1(n6994), .A2(n9825), .ZN(n6995) );
  INV_X1 U8752 ( .A(n6803), .ZN(n8079) );
  XNOR2_X1 U8753 ( .A(n8219), .B(n7005), .ZN(n6997) );
  NAND2_X1 U8754 ( .A1(n6997), .A2(n5750), .ZN(n7040) );
  INV_X1 U8755 ( .A(n6997), .ZN(n6998) );
  INV_X1 U8756 ( .A(n5750), .ZN(n8564) );
  NAND2_X1 U8757 ( .A1(n6998), .A2(n8564), .ZN(n6999) );
  NAND2_X1 U8758 ( .A1(n7040), .A2(n6999), .ZN(n7002) );
  INV_X1 U8759 ( .A(n7003), .ZN(n7001) );
  NAND2_X1 U8760 ( .A1(n7001), .A2(n7000), .ZN(n7041) );
  INV_X1 U8761 ( .A(n7041), .ZN(n7039) );
  AOI21_X1 U8762 ( .B1(n7003), .B2(n7002), .A(n7039), .ZN(n7010) );
  INV_X1 U8763 ( .A(n8563), .ZN(n7268) );
  AOI21_X1 U8764 ( .B1(n8228), .B2(n7005), .A(n7004), .ZN(n7006) );
  OAI21_X1 U8765 ( .B1(n8290), .B2(n7268), .A(n7006), .ZN(n7008) );
  NOR2_X1 U8766 ( .A1(n8223), .A2(n7152), .ZN(n7007) );
  AOI211_X1 U8767 ( .C1(n8288), .C2(n9825), .A(n7008), .B(n7007), .ZN(n7009)
         );
  OAI21_X1 U8768 ( .B1(n7010), .B2(n8272), .A(n7009), .ZN(P2_U3170) );
  NOR2_X1 U8769 ( .A1(n7237), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7011) );
  AOI21_X1 U8770 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7237), .A(n7011), .ZN(
        n7014) );
  OAI21_X1 U8771 ( .B1(n7014), .B2(n7013), .A(n7232), .ZN(n7015) );
  NAND2_X1 U8772 ( .A1(n7015), .A2(n9360), .ZN(n7026) );
  AOI22_X1 U8773 ( .A1(n7237), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n7018), .B2(
        n7022), .ZN(n7019) );
  OAI21_X1 U8774 ( .B1(n7020), .B2(n7019), .A(n7236), .ZN(n7024) );
  NAND2_X1 U8775 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U8776 ( .A1(n9739), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7021) );
  OAI211_X1 U8777 ( .C1(n7907), .C2(n7022), .A(n9120), .B(n7021), .ZN(n7023)
         );
  AOI21_X1 U8778 ( .B1(n7024), .B2(n9354), .A(n7023), .ZN(n7025) );
  NAND2_X1 U8779 ( .A1(n7026), .A2(n7025), .ZN(P1_U3255) );
  INV_X1 U8780 ( .A(n7027), .ZN(n7029) );
  INV_X1 U8781 ( .A(n8692), .ZN(n8671) );
  OAI222_X1 U8782 ( .A1(n9031), .A2(n7028), .B1(n9034), .B2(n7029), .C1(
        P2_U3151), .C2(n8671), .ZN(P2_U3278) );
  OAI222_X1 U8783 ( .A1(n9729), .A2(n7030), .B1(n9732), .B2(n7029), .C1(
        P1_U3086), .C2(n9337), .ZN(P1_U3338) );
  XOR2_X1 U8784 ( .A(n7032), .B(n7031), .Z(n7037) );
  OR2_X1 U8785 ( .A1(n7305), .A2(n9235), .ZN(n7034) );
  NAND2_X1 U8786 ( .A1(n5517), .A2(n9237), .ZN(n7033) );
  NAND2_X1 U8787 ( .A1(n7034), .A2(n7033), .ZN(n7097) );
  AOI22_X1 U8788 ( .A1(n7097), .A2(n9224), .B1(n9770), .B2(n9228), .ZN(n7036)
         );
  NAND2_X1 U8789 ( .A1(n9226), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10107) );
  NAND2_X1 U8790 ( .A1(n10107), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7035) );
  OAI211_X1 U8791 ( .C1(n7037), .C2(n10103), .A(n7036), .B(n7035), .ZN(
        P1_U3222) );
  INV_X1 U8792 ( .A(n7040), .ZN(n7038) );
  XNOR2_X1 U8793 ( .A(n8219), .B(n7048), .ZN(n7269) );
  XNOR2_X1 U8794 ( .A(n7269), .B(n8563), .ZN(n7042) );
  NOR3_X1 U8795 ( .A1(n7039), .A2(n7038), .A3(n7042), .ZN(n7045) );
  NAND2_X1 U8796 ( .A1(n7041), .A2(n7040), .ZN(n7043) );
  INV_X1 U8797 ( .A(n7271), .ZN(n7044) );
  OAI21_X1 U8798 ( .B1(n7045), .B2(n7044), .A(n8285), .ZN(n7052) );
  INV_X1 U8799 ( .A(n7046), .ZN(n7047) );
  AOI21_X1 U8800 ( .B1(n8228), .B2(n7048), .A(n7047), .ZN(n7049) );
  OAI21_X1 U8801 ( .B1(n8290), .B2(n7292), .A(n7049), .ZN(n7050) );
  AOI21_X1 U8802 ( .B1(n8288), .B2(n8564), .A(n7050), .ZN(n7051) );
  OAI211_X1 U8803 ( .C1(n7172), .C2(n8223), .A(n7052), .B(n7051), .ZN(P2_U3167) );
  NAND2_X1 U8804 ( .A1(n9272), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7053) );
  OAI21_X1 U8805 ( .B1(n8103), .B2(n9272), .A(n7053), .ZN(P1_U3583) );
  XNOR2_X1 U8806 ( .A(n7055), .B(n7054), .ZN(n8947) );
  INV_X1 U8807 ( .A(n8947), .ZN(n7063) );
  XNOR2_X1 U8808 ( .A(n7054), .B(n7056), .ZN(n7057) );
  NAND2_X1 U8809 ( .A1(n7057), .A2(n9829), .ZN(n7059) );
  AOI22_X1 U8810 ( .A1(n9826), .A2(n8566), .B1(n8565), .B2(n9824), .ZN(n7058)
         );
  AND2_X1 U8811 ( .A1(n7059), .A2(n7058), .ZN(n8948) );
  MUX2_X1 U8812 ( .A(n8948), .B(n7060), .S(n9839), .Z(n7062) );
  AOI22_X1 U8813 ( .A1(n8899), .A2(n8946), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8898), .ZN(n7061) );
  OAI211_X1 U8814 ( .C1(n7063), .C2(n8903), .A(n7062), .B(n7061), .ZN(P2_U3232) );
  INV_X1 U8815 ( .A(n7064), .ZN(n7089) );
  OAI222_X1 U8816 ( .A1(P1_U3086), .A2(n9341), .B1(n9732), .B2(n7089), .C1(
        n7065), .C2(n9729), .ZN(P1_U3337) );
  INV_X1 U8817 ( .A(n7066), .ZN(n7068) );
  MUX2_X1 U8818 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6091), .Z(n7206) );
  XNOR2_X1 U8819 ( .A(n7206), .B(n7205), .ZN(n7207) );
  XNOR2_X1 U8820 ( .A(n7208), .B(n7207), .ZN(n7087) );
  NAND2_X1 U8821 ( .A1(n7074), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7070) );
  NAND2_X1 U8822 ( .A1(n7071), .A2(n7070), .ZN(n7072) );
  AOI21_X1 U8823 ( .B1(n7073), .B2(n5784), .A(n4415), .ZN(n7085) );
  NAND2_X1 U8824 ( .A1(n7074), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8825 ( .A1(n7076), .A2(n7075), .ZN(n7078) );
  NAND2_X1 U8826 ( .A1(n7078), .A2(n7205), .ZN(n7215) );
  NAND2_X1 U8827 ( .A1(n7077), .A2(n7215), .ZN(n7079) );
  NOR2_X1 U8828 ( .A1(n5783), .A2(n7079), .ZN(n7216) );
  AOI21_X1 U8829 ( .B1(n7079), .B2(n5783), .A(n7216), .ZN(n7080) );
  OR2_X1 U8830 ( .A1(n7080), .A2(n8689), .ZN(n7084) );
  INV_X1 U8831 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8832 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7290) );
  OAI21_X1 U8833 ( .B1(n8704), .B2(n7081), .A(n7290), .ZN(n7082) );
  AOI21_X1 U8834 ( .B1(n8676), .B2(n4703), .A(n7082), .ZN(n7083) );
  OAI211_X1 U8835 ( .C1(n7085), .C2(n8731), .A(n7084), .B(n7083), .ZN(n7086)
         );
  AOI21_X1 U8836 ( .B1(n7087), .B2(n8664), .A(n7086), .ZN(n7088) );
  INV_X1 U8837 ( .A(n7088), .ZN(P2_U3189) );
  INV_X1 U8838 ( .A(n8713), .ZN(n8700) );
  OAI222_X1 U8839 ( .A1(n9031), .A2(n7090), .B1(n8700), .B2(P2_U3151), .C1(
        n9034), .C2(n7089), .ZN(P2_U3277) );
  OAI21_X1 U8840 ( .B1(n7091), .B2(n7093), .A(n7092), .ZN(n9774) );
  INV_X1 U8841 ( .A(n9774), .ZN(n7099) );
  INV_X1 U8842 ( .A(n8063), .ZN(n7761) );
  XNOR2_X1 U8843 ( .A(n7091), .B(n7094), .ZN(n7095) );
  NOR2_X1 U8844 ( .A1(n7095), .A2(n9497), .ZN(n7096) );
  AOI211_X1 U8845 ( .C1(n7761), .C2(n9774), .A(n7097), .B(n7096), .ZN(n9777)
         );
  INV_X1 U8846 ( .A(n7257), .ZN(n7098) );
  OAI211_X1 U8847 ( .C1(n7103), .C2(n7125), .A(n7098), .B(n6447), .ZN(n9768)
         );
  OAI211_X1 U8848 ( .C1(n7099), .C2(n9781), .A(n9777), .B(n9768), .ZN(n7105)
         );
  OAI22_X1 U8849 ( .A1(n9717), .A2(n7103), .B1(n9713), .B2(n4868), .ZN(n7100)
         );
  AOI21_X1 U8850 ( .B1(n7105), .B2(n9713), .A(n7100), .ZN(n7101) );
  INV_X1 U8851 ( .A(n7101), .ZN(P1_U3456) );
  OAI22_X1 U8852 ( .A1(n9659), .A2(n7103), .B1(n9818), .B2(n7102), .ZN(n7104)
         );
  AOI21_X1 U8853 ( .B1(n7105), .B2(n9818), .A(n7104), .ZN(n7106) );
  INV_X1 U8854 ( .A(n7106), .ZN(P1_U3523) );
  OAI21_X1 U8855 ( .B1(n7110), .B2(n7109), .A(n9780), .ZN(n7112) );
  NAND4_X1 U8856 ( .A1(n7113), .A2(n9720), .A3(n7112), .A4(n7111), .ZN(n7114)
         );
  NOR2_X2 U8857 ( .A1(n9778), .A2(n7115), .ZN(n9769) );
  AOI21_X1 U8858 ( .B1(n9772), .B2(n6447), .A(n9769), .ZN(n7126) );
  NAND3_X1 U8859 ( .A1(n7118), .A2(n7117), .A3(n7116), .ZN(n7120) );
  OAI211_X1 U8860 ( .C1(n9754), .C2(n7121), .A(n7120), .B(n7119), .ZN(n7123)
         );
  NOR2_X1 U8861 ( .A1(n9745), .A2(n4892), .ZN(n7122) );
  AOI21_X1 U8862 ( .B1(n7123), .B2(n9745), .A(n7122), .ZN(n7124) );
  OAI21_X1 U8863 ( .B1(n7126), .B2(n7125), .A(n7124), .ZN(P1_U3293) );
  INV_X1 U8864 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9922) );
  NOR2_X1 U8865 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7127) );
  AOI21_X1 U8866 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7127), .ZN(n9927) );
  NOR2_X1 U8867 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7128) );
  AOI21_X1 U8868 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7128), .ZN(n9930) );
  NOR2_X1 U8869 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7129) );
  AOI21_X1 U8870 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7129), .ZN(n9933) );
  NOR2_X1 U8871 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7130) );
  AOI21_X1 U8872 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7130), .ZN(n9936) );
  NOR2_X1 U8873 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7131) );
  AOI21_X1 U8874 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7131), .ZN(n9939) );
  NOR2_X1 U8875 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7132) );
  AOI21_X1 U8876 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7132), .ZN(n9942) );
  NOR2_X1 U8877 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7133) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7133), .ZN(n9945) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7134) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7134), .ZN(n9948) );
  NOR2_X1 U8881 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7135) );
  AOI21_X1 U8882 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7135), .ZN(n10118) );
  NOR2_X1 U8883 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7136) );
  AOI21_X1 U8884 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7136), .ZN(n10124) );
  NOR2_X1 U8885 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7137) );
  AOI21_X1 U8886 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7137), .ZN(n10121) );
  NOR2_X1 U8887 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7138) );
  AOI21_X1 U8888 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7138), .ZN(n10112) );
  NOR2_X1 U8889 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7139) );
  AOI21_X1 U8890 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7139), .ZN(n10115) );
  AND2_X1 U8891 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7140) );
  NOR2_X1 U8892 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7140), .ZN(n9917) );
  INV_X1 U8893 ( .A(n9917), .ZN(n9918) );
  NAND3_X1 U8894 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U8895 ( .A1(n9920), .A2(n9919), .ZN(n9916) );
  NAND2_X1 U8896 ( .A1(n9918), .A2(n9916), .ZN(n10127) );
  NAND2_X1 U8897 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7141) );
  OAI21_X1 U8898 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7141), .ZN(n10126) );
  NOR2_X1 U8899 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  AOI21_X1 U8900 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10125), .ZN(n10130) );
  NAND2_X1 U8901 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7142) );
  OAI21_X1 U8902 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7142), .ZN(n10129) );
  NOR2_X1 U8903 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  AOI21_X1 U8904 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10128), .ZN(n10133) );
  NOR2_X1 U8905 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7143) );
  AOI21_X1 U8906 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7143), .ZN(n10132) );
  NAND2_X1 U8907 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  OAI21_X1 U8908 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10131), .ZN(n10114) );
  NAND2_X1 U8909 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  OAI21_X1 U8910 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10113), .ZN(n10111) );
  NAND2_X1 U8911 ( .A1(n10112), .A2(n10111), .ZN(n10110) );
  OAI21_X1 U8912 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10110), .ZN(n10120) );
  NAND2_X1 U8913 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  OAI21_X1 U8914 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10119), .ZN(n10123) );
  NAND2_X1 U8915 ( .A1(n10124), .A2(n10123), .ZN(n10122) );
  OAI21_X1 U8916 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10122), .ZN(n10117) );
  NAND2_X1 U8917 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OAI21_X1 U8918 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10116), .ZN(n9947) );
  NAND2_X1 U8919 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  OAI21_X1 U8920 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9946), .ZN(n9944) );
  NAND2_X1 U8921 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U8922 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9943), .ZN(n9941) );
  NAND2_X1 U8923 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  OAI21_X1 U8924 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9940), .ZN(n9938) );
  NAND2_X1 U8925 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  OAI21_X1 U8926 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9937), .ZN(n9935) );
  NAND2_X1 U8927 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  OAI21_X1 U8928 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9934), .ZN(n9932) );
  NAND2_X1 U8929 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  OAI21_X1 U8930 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9931), .ZN(n9929) );
  NAND2_X1 U8931 ( .A1(n9930), .A2(n9929), .ZN(n9928) );
  OAI21_X1 U8932 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9928), .ZN(n9926) );
  NAND2_X1 U8933 ( .A1(n9927), .A2(n9926), .ZN(n9925) );
  OAI21_X1 U8934 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9925), .ZN(n9923) );
  NOR2_X1 U8935 ( .A1(n9922), .A2(n9923), .ZN(n7144) );
  NAND2_X1 U8936 ( .A1(n9922), .A2(n9923), .ZN(n9921) );
  OAI21_X1 U8937 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7144), .A(n9921), .ZN(
        n7147) );
  XNOR2_X1 U8938 ( .A(n7145), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7146) );
  XNOR2_X1 U8939 ( .A(n7147), .B(n7146), .ZN(ADD_1068_U4) );
  AND2_X1 U8940 ( .A1(n7149), .A2(n7148), .ZN(n7151) );
  OAI21_X1 U8941 ( .B1(n7151), .B2(n8386), .A(n7150), .ZN(n9852) );
  OAI22_X1 U8942 ( .A1(n8738), .A2(n9849), .B1(n7152), .B2(n9821), .ZN(n7156)
         );
  XNOR2_X1 U8943 ( .A(n7153), .B(n8386), .ZN(n7154) );
  OAI222_X1 U8944 ( .A1(n8866), .A2(n7268), .B1(n8864), .B2(n8376), .C1(n8862), 
        .C2(n7154), .ZN(n9850) );
  MUX2_X1 U8945 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9850), .S(n9837), .Z(n7155)
         );
  AOI211_X1 U8946 ( .C1(n7811), .C2(n9852), .A(n7156), .B(n7155), .ZN(n7157)
         );
  INV_X1 U8947 ( .A(n7157), .ZN(P2_U3229) );
  XNOR2_X1 U8948 ( .A(n7158), .B(n8339), .ZN(n9865) );
  NAND2_X1 U8949 ( .A1(n8894), .A2(n9836), .ZN(n8167) );
  NAND2_X1 U8950 ( .A1(n7160), .A2(n7159), .ZN(n8148) );
  NAND2_X1 U8951 ( .A1(n8148), .A2(n8146), .ZN(n7161) );
  NAND2_X1 U8952 ( .A1(n7161), .A2(n8147), .ZN(n7162) );
  INV_X1 U8953 ( .A(n8339), .ZN(n8410) );
  XNOR2_X1 U8954 ( .A(n7162), .B(n8410), .ZN(n7164) );
  OAI22_X1 U8955 ( .A1(n7407), .A2(n8866), .B1(n7292), .B2(n8864), .ZN(n7163)
         );
  AOI21_X1 U8956 ( .B1(n7164), .B2(n9829), .A(n7163), .ZN(n7165) );
  OAI21_X1 U8957 ( .B1(n9865), .B2(n9833), .A(n7165), .ZN(n9867) );
  NAND2_X1 U8958 ( .A1(n9867), .A2(n9837), .ZN(n7168) );
  OAI22_X1 U8959 ( .A1(n8894), .A2(n5784), .B1(n7289), .B2(n9821), .ZN(n7166)
         );
  AOI21_X1 U8960 ( .B1(n8899), .B2(n8418), .A(n7166), .ZN(n7167) );
  OAI211_X1 U8961 ( .C1(n9865), .C2(n8167), .A(n7168), .B(n7167), .ZN(P2_U3226) );
  AND2_X1 U8962 ( .A1(n8399), .A2(n8395), .ZN(n8337) );
  XOR2_X1 U8963 ( .A(n7169), .B(n8337), .Z(n7170) );
  INV_X1 U8964 ( .A(n7292), .ZN(n7280) );
  AOI222_X1 U8965 ( .A1(n9829), .A2(n7170), .B1(n7280), .B2(n9824), .C1(n8564), 
        .C2(n9826), .ZN(n9854) );
  XNOR2_X1 U8966 ( .A(n7171), .B(n8337), .ZN(n9857) );
  NOR2_X1 U8967 ( .A1(n9837), .A2(n6850), .ZN(n7174) );
  OAI22_X1 U8968 ( .A1(n8738), .A2(n9855), .B1(n7172), .B2(n9821), .ZN(n7173)
         );
  AOI211_X1 U8969 ( .C1(n9857), .C2(n7811), .A(n7174), .B(n7173), .ZN(n7175)
         );
  OAI21_X1 U8970 ( .B1(n9854), .B2(n9839), .A(n7175), .ZN(P2_U3228) );
  INV_X1 U8971 ( .A(n7176), .ZN(n7177) );
  NAND2_X1 U8972 ( .A1(n8565), .A2(n9826), .ZN(n7179) );
  OAI21_X1 U8973 ( .B1(n5750), .B2(n8866), .A(n7179), .ZN(n7180) );
  AOI21_X1 U8974 ( .B1(n7181), .B2(n9829), .A(n7180), .ZN(n9845) );
  NAND2_X1 U8975 ( .A1(n7182), .A2(n8379), .ZN(n7183) );
  XNOR2_X1 U8976 ( .A(n8331), .B(n7183), .ZN(n9847) );
  AOI22_X1 U8977 ( .A1(n8899), .A2(n6835), .B1(n8898), .B2(n7184), .ZN(n7185)
         );
  OAI21_X1 U8978 ( .B1(n5727), .B2(n9837), .A(n7185), .ZN(n7186) );
  AOI21_X1 U8979 ( .B1(n9847), .B2(n7811), .A(n7186), .ZN(n7187) );
  OAI21_X1 U8980 ( .B1(n9845), .B2(n9839), .A(n7187), .ZN(P2_U3230) );
  INV_X1 U8981 ( .A(n7188), .ZN(n8415) );
  NAND2_X1 U8982 ( .A1(n8415), .A2(n8420), .ZN(n8338) );
  AND2_X1 U8983 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  XOR2_X1 U8984 ( .A(n8338), .B(n7191), .Z(n7192) );
  INV_X1 U8985 ( .A(n8419), .ZN(n8562) );
  AOI222_X1 U8986 ( .A1(n9829), .A2(n7192), .B1(n8560), .B2(n9824), .C1(n8562), 
        .C2(n9826), .ZN(n9869) );
  XNOR2_X1 U8987 ( .A(n7193), .B(n8338), .ZN(n9872) );
  NOR2_X1 U8988 ( .A1(n8738), .A2(n9870), .ZN(n7196) );
  OAI22_X1 U8989 ( .A1(n8894), .A2(n7194), .B1(n7401), .B2(n9821), .ZN(n7195)
         );
  AOI211_X1 U8990 ( .C1(n9872), .C2(n7811), .A(n7196), .B(n7195), .ZN(n7197)
         );
  OAI21_X1 U8991 ( .B1(n9869), .B2(n9839), .A(n7197), .ZN(P2_U3225) );
  OAI211_X1 U8992 ( .C1(n7200), .C2(n7199), .A(n7198), .B(n6436), .ZN(n7204)
         );
  OAI22_X1 U8993 ( .A1(n7454), .A2(n9235), .B1(n7201), .B2(n9220), .ZN(n7335)
         );
  AND2_X1 U8994 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9314) );
  NOR2_X1 U8995 ( .A1(n10096), .A2(n7340), .ZN(n7202) );
  AOI211_X1 U8996 ( .C1(n7335), .C2(n9224), .A(n9314), .B(n7202), .ZN(n7203)
         );
  OAI211_X1 U8997 ( .C1(n9226), .C2(n7339), .A(n7204), .B(n7203), .ZN(P1_U3230) );
  MUX2_X1 U8998 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6091), .Z(n7487) );
  XNOR2_X1 U8999 ( .A(n7487), .B(n7225), .ZN(n7209) );
  OAI21_X1 U9000 ( .B1(n7210), .B2(n7209), .A(n7488), .ZN(n7230) );
  NAND2_X1 U9001 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7497), .ZN(n7211) );
  OAI21_X1 U9002 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7497), .A(n7211), .ZN(
        n7212) );
  AOI21_X1 U9003 ( .B1(n7213), .B2(n7212), .A(n7485), .ZN(n7214) );
  NOR2_X1 U9004 ( .A1(n7214), .A2(n8731), .ZN(n7229) );
  NAND2_X1 U9005 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7497), .ZN(n7218) );
  OAI21_X1 U9006 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7497), .A(n7218), .ZN(
        n7219) );
  AOI21_X1 U9007 ( .B1(n7220), .B2(n7219), .A(n7496), .ZN(n7227) );
  INV_X1 U9008 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7223) );
  INV_X1 U9009 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7221) );
  NOR2_X1 U9010 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7221), .ZN(n7395) );
  INV_X1 U9011 ( .A(n7395), .ZN(n7222) );
  OAI21_X1 U9012 ( .B1(n8704), .B2(n7223), .A(n7222), .ZN(n7224) );
  AOI21_X1 U9013 ( .B1(n8676), .B2(n7225), .A(n7224), .ZN(n7226) );
  OAI21_X1 U9014 ( .B1(n7227), .B2(n8689), .A(n7226), .ZN(n7228) );
  AOI211_X1 U9015 ( .C1(n7230), .C2(n8664), .A(n7229), .B(n7228), .ZN(n7231)
         );
  INV_X1 U9016 ( .A(n7231), .ZN(P2_U3190) );
  OAI21_X1 U9017 ( .B1(n7237), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7232), .ZN(
        n7235) );
  NAND2_X1 U9018 ( .A1(n7380), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7233) );
  OAI21_X1 U9019 ( .B1(n7380), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7233), .ZN(
        n7234) );
  NOR2_X1 U9020 ( .A1(n7234), .A2(n7235), .ZN(n7375) );
  AOI211_X1 U9021 ( .C1(n7235), .C2(n7234), .A(n7375), .B(n7376), .ZN(n7245)
         );
  OAI21_X1 U9022 ( .B1(n7237), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7236), .ZN(
        n7239) );
  XNOR2_X1 U9023 ( .A(n7380), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7238) );
  NOR2_X1 U9024 ( .A1(n7238), .A2(n7239), .ZN(n7379) );
  AOI211_X1 U9025 ( .C1(n7239), .C2(n7238), .A(n7379), .B(n9356), .ZN(n7244)
         );
  INV_X1 U9026 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U9027 ( .A1(n9359), .A2(n7380), .ZN(n7241) );
  NAND2_X1 U9028 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7240) );
  OAI211_X1 U9029 ( .C1(n7242), .C2(n9366), .A(n7241), .B(n7240), .ZN(n7243)
         );
  OR3_X1 U9030 ( .A1(n7245), .A2(n7244), .A3(n7243), .ZN(P1_U3256) );
  NAND2_X1 U9031 ( .A1(n8697), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7246) );
  OAI21_X1 U9032 ( .B1(n8225), .B2(n8697), .A(n7246), .ZN(P2_U3520) );
  INV_X1 U9033 ( .A(n7247), .ZN(n8144) );
  OAI222_X1 U9034 ( .A1(n9031), .A2(n7248), .B1(n9034), .B2(n8144), .C1(n4316), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XNOR2_X1 U9035 ( .A(n7249), .B(n7251), .ZN(n7256) );
  OAI21_X1 U9036 ( .B1(n7252), .B2(n7251), .A(n7250), .ZN(n9785) );
  NAND2_X1 U9037 ( .A1(n9785), .A2(n7761), .ZN(n7255) );
  NAND2_X1 U9038 ( .A1(n6942), .A2(n9237), .ZN(n7254) );
  NAND2_X1 U9039 ( .A1(n9270), .A2(n9196), .ZN(n7253) );
  AND2_X1 U9040 ( .A1(n7254), .A2(n7253), .ZN(n10099) );
  OAI211_X1 U9041 ( .C1(n9497), .C2(n7256), .A(n7255), .B(n10099), .ZN(n9783)
         );
  INV_X1 U9042 ( .A(n9783), .ZN(n7263) );
  NOR2_X1 U9043 ( .A1(n9778), .A2(n7315), .ZN(n9773) );
  OAI211_X1 U9044 ( .C1(n7257), .C2(n10097), .A(n7302), .B(n6447), .ZN(n9782)
         );
  OAI22_X1 U9045 ( .A1(n9745), .A2(n4901), .B1(n9288), .B2(n9754), .ZN(n7258)
         );
  AOI21_X1 U9046 ( .B1(n9769), .B2(n7259), .A(n7258), .ZN(n7260) );
  OAI21_X1 U9047 ( .B1(n9760), .B2(n9782), .A(n7260), .ZN(n7261) );
  AOI21_X1 U9048 ( .B1(n9785), .B2(n9773), .A(n7261), .ZN(n7262) );
  OAI21_X1 U9049 ( .B1(n7263), .B2(n9778), .A(n7262), .ZN(P1_U3291) );
  INV_X1 U9050 ( .A(n7264), .ZN(n8151) );
  OR2_X1 U9051 ( .A1(n8268), .A2(n7268), .ZN(n7267) );
  AOI21_X1 U9052 ( .B1(n8228), .B2(n8152), .A(n7265), .ZN(n7266) );
  OAI211_X1 U9053 ( .C1(n8290), .C2(n8419), .A(n7267), .B(n7266), .ZN(n7277)
         );
  XNOR2_X1 U9054 ( .A(n6803), .B(n8152), .ZN(n7279) );
  XNOR2_X1 U9055 ( .A(n7279), .B(n7292), .ZN(n7275) );
  NAND2_X1 U9056 ( .A1(n7269), .A2(n7268), .ZN(n7270) );
  INV_X1 U9057 ( .A(n7283), .ZN(n7273) );
  AOI211_X1 U9058 ( .C1(n7275), .C2(n7274), .A(n8272), .B(n7273), .ZN(n7276)
         );
  AOI211_X1 U9059 ( .C1(n8151), .C2(n8293), .A(n7277), .B(n7276), .ZN(n7278)
         );
  INV_X1 U9060 ( .A(n7278), .ZN(P2_U3179) );
  INV_X1 U9061 ( .A(n7279), .ZN(n7281) );
  NAND2_X1 U9062 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  AND2_X2 U9063 ( .A1(n7283), .A2(n7282), .ZN(n7288) );
  XNOR2_X1 U9064 ( .A(n6803), .B(n8418), .ZN(n7284) );
  NAND2_X1 U9065 ( .A1(n7284), .A2(n8419), .ZN(n7390) );
  INV_X1 U9066 ( .A(n7284), .ZN(n7285) );
  NAND2_X1 U9067 ( .A1(n7285), .A2(n8562), .ZN(n7286) );
  AND2_X1 U9068 ( .A1(n7390), .A2(n7286), .ZN(n7287) );
  OAI21_X1 U9069 ( .B1(n7288), .B2(n7287), .A(n7391), .ZN(n7298) );
  OR2_X1 U9070 ( .A1(n8223), .A2(n7289), .ZN(n7296) );
  INV_X1 U9071 ( .A(n7290), .ZN(n7291) );
  AOI21_X1 U9072 ( .B1(n8266), .B2(n8561), .A(n7291), .ZN(n7295) );
  NAND2_X1 U9073 ( .A1(n8228), .A2(n8418), .ZN(n7294) );
  OR2_X1 U9074 ( .A1(n8268), .A2(n7292), .ZN(n7293) );
  NAND4_X1 U9075 ( .A1(n7296), .A2(n7295), .A3(n7294), .A4(n7293), .ZN(n7297)
         );
  AOI21_X1 U9076 ( .B1(n7298), .B2(n8285), .A(n7297), .ZN(n7299) );
  INV_X1 U9077 ( .A(n7299), .ZN(P2_U3153) );
  NAND2_X1 U9078 ( .A1(n7300), .A2(n7303), .ZN(n7327) );
  OAI21_X1 U9079 ( .B1(n7300), .B2(n7303), .A(n7327), .ZN(n7323) );
  INV_X1 U9080 ( .A(n7338), .ZN(n7301) );
  AOI211_X1 U9081 ( .C1(n7369), .C2(n7302), .A(n9579), .B(n7301), .ZN(n7317)
         );
  XOR2_X1 U9082 ( .A(n7304), .B(n7303), .Z(n7308) );
  OAI22_X1 U9083 ( .A1(n7306), .A2(n9235), .B1(n7305), .B2(n9220), .ZN(n7370)
         );
  INV_X1 U9084 ( .A(n7370), .ZN(n7307) );
  OAI21_X1 U9085 ( .B1(n7308), .B2(n9497), .A(n7307), .ZN(n7314) );
  AOI211_X1 U9086 ( .C1(n9801), .C2(n7323), .A(n7317), .B(n7314), .ZN(n7313)
         );
  OAI22_X1 U9087 ( .A1(n9659), .A2(n7321), .B1(n9818), .B2(n6769), .ZN(n7309)
         );
  INV_X1 U9088 ( .A(n7309), .ZN(n7310) );
  OAI21_X1 U9089 ( .B1(n7313), .B2(n9816), .A(n7310), .ZN(P1_U3525) );
  OAI22_X1 U9090 ( .A1(n9717), .A2(n7321), .B1(n9794), .B2(n4921), .ZN(n7311)
         );
  INV_X1 U9091 ( .A(n7311), .ZN(n7312) );
  OAI21_X1 U9092 ( .B1(n7313), .B2(n9809), .A(n7312), .ZN(P1_U3462) );
  INV_X1 U9093 ( .A(n7314), .ZN(n7325) );
  AND2_X1 U9094 ( .A1(n8063), .A2(n7315), .ZN(n7316) );
  NAND2_X1 U9095 ( .A1(n7317), .A2(n9772), .ZN(n7320) );
  INV_X1 U9096 ( .A(n9754), .ZN(n9767) );
  INV_X1 U9097 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7318) );
  AOI22_X1 U9098 ( .A1(n9778), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9767), .B2(
        n7318), .ZN(n7319) );
  OAI211_X1 U9099 ( .C1(n7321), .C2(n9556), .A(n7320), .B(n7319), .ZN(n7322)
         );
  AOI21_X1 U9100 ( .B1(n9763), .B2(n7323), .A(n7322), .ZN(n7324) );
  OAI21_X1 U9101 ( .B1(n9778), .B2(n7325), .A(n7324), .ZN(P1_U3290) );
  NAND2_X1 U9102 ( .A1(n7327), .A2(n7326), .ZN(n7331) );
  AND2_X1 U9103 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  OAI21_X1 U9104 ( .B1(n7331), .B2(n7334), .A(n7330), .ZN(n7332) );
  INV_X1 U9105 ( .A(n7332), .ZN(n9791) );
  XOR2_X1 U9106 ( .A(n7334), .B(n7333), .Z(n7336) );
  AOI21_X1 U9107 ( .B1(n7336), .B2(n9575), .A(n7335), .ZN(n9790) );
  MUX2_X1 U9108 ( .A(n9790), .B(n7337), .S(n9778), .Z(n7343) );
  AOI211_X1 U9109 ( .C1(n9787), .C2(n7338), .A(n9579), .B(n7428), .ZN(n9786)
         );
  OAI22_X1 U9110 ( .A1(n9556), .A2(n7340), .B1(n9754), .B2(n7339), .ZN(n7341)
         );
  AOI21_X1 U9111 ( .B1(n9786), .B2(n9772), .A(n7341), .ZN(n7342) );
  OAI211_X1 U9112 ( .C1(n9791), .C2(n9589), .A(n7343), .B(n7342), .ZN(P1_U3289) );
  NAND2_X1 U9113 ( .A1(n7344), .A2(n8340), .ZN(n7345) );
  NAND2_X1 U9114 ( .A1(n4651), .A2(n7345), .ZN(n9875) );
  INV_X1 U9115 ( .A(n8426), .ZN(n7681) );
  AOI22_X1 U9116 ( .A1(n7681), .A2(n9824), .B1(n9826), .B2(n8561), .ZN(n7349)
         );
  XNOR2_X1 U9117 ( .A(n7346), .B(n8340), .ZN(n7347) );
  NAND2_X1 U9118 ( .A1(n7347), .A2(n9829), .ZN(n7348) );
  OAI211_X1 U9119 ( .C1(n9875), .C2(n9833), .A(n7349), .B(n7348), .ZN(n9876)
         );
  NAND2_X1 U9120 ( .A1(n9876), .A2(n9837), .ZN(n7352) );
  OAI22_X1 U9121 ( .A1(n8894), .A2(n5833), .B1(n7415), .B2(n9821), .ZN(n7350)
         );
  AOI21_X1 U9122 ( .B1(n8899), .B2(n9878), .A(n7350), .ZN(n7351) );
  OAI211_X1 U9123 ( .C1(n9875), .C2(n8167), .A(n7352), .B(n7351), .ZN(P2_U3224) );
  INV_X1 U9124 ( .A(n7353), .ZN(n7403) );
  OAI222_X1 U9125 ( .A1(n9034), .A2(n7403), .B1(P2_U3151), .B2(n8539), .C1(
        n10068), .C2(n9031), .ZN(P2_U3275) );
  NAND2_X1 U9126 ( .A1(n8432), .A2(n8435), .ZN(n8342) );
  XNOR2_X1 U9127 ( .A(n7354), .B(n8342), .ZN(n9881) );
  XNOR2_X1 U9128 ( .A(n7355), .B(n8342), .ZN(n7356) );
  NAND2_X1 U9129 ( .A1(n7356), .A2(n9829), .ZN(n7358) );
  AOI22_X1 U9130 ( .A1(n7792), .A2(n9824), .B1(n9826), .B2(n8560), .ZN(n7357)
         );
  NAND2_X1 U9131 ( .A1(n7358), .A2(n7357), .ZN(n9883) );
  NAND2_X1 U9132 ( .A1(n9883), .A2(n9837), .ZN(n7362) );
  OAI22_X1 U9133 ( .A1(n8894), .A2(n7359), .B1(n7672), .B2(n9821), .ZN(n7360)
         );
  AOI21_X1 U9134 ( .B1(n8899), .B2(n9884), .A(n7360), .ZN(n7361) );
  OAI211_X1 U9135 ( .C1(n9881), .C2(n8903), .A(n7362), .B(n7361), .ZN(P2_U3223) );
  XNOR2_X1 U9136 ( .A(n7364), .B(n6220), .ZN(n10102) );
  NOR2_X1 U9137 ( .A1(n10102), .A2(n10101), .ZN(n10100) );
  AOI21_X1 U9138 ( .B1(n6220), .B2(n7364), .A(n10100), .ZN(n7368) );
  XOR2_X1 U9139 ( .A(n7366), .B(n7365), .Z(n7367) );
  XNOR2_X1 U9140 ( .A(n7368), .B(n7367), .ZN(n7373) );
  AOI22_X1 U9141 ( .A1(n7370), .A2(n9224), .B1(n7369), .B2(n9228), .ZN(n7372)
         );
  MUX2_X1 U9142 ( .A(n9226), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7371) );
  OAI211_X1 U9143 ( .C1(n7373), .C2(n10103), .A(n7372), .B(n7371), .ZN(
        P1_U3218) );
  NAND2_X1 U9144 ( .A1(n7703), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7374) );
  OAI21_X1 U9145 ( .B1(n7703), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7374), .ZN(
        n7378) );
  AOI21_X1 U9146 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7380), .A(n7375), .ZN(
        n7377) );
  NOR2_X1 U9147 ( .A1(n7377), .A2(n7378), .ZN(n7698) );
  AOI211_X1 U9148 ( .C1(n7378), .C2(n7377), .A(n7698), .B(n7376), .ZN(n7388)
         );
  XNOR2_X1 U9149 ( .A(n7703), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7381) );
  AOI211_X1 U9150 ( .C1(n7382), .C2(n7381), .A(n7702), .B(n9356), .ZN(n7387)
         );
  INV_X1 U9151 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U9152 ( .A1(n9359), .A2(n7703), .ZN(n7384) );
  NAND2_X1 U9153 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n7383) );
  OAI211_X1 U9154 ( .C1(n7385), .C2(n9366), .A(n7384), .B(n7383), .ZN(n7386)
         );
  OR3_X1 U9155 ( .A1(n7388), .A2(n7387), .A3(n7386), .ZN(P1_U3257) );
  INV_X1 U9156 ( .A(n7391), .ZN(n7389) );
  XNOR2_X1 U9157 ( .A(n7398), .B(n6803), .ZN(n7408) );
  XNOR2_X1 U9158 ( .A(n7408), .B(n8561), .ZN(n7392) );
  NOR3_X1 U9159 ( .A1(n7389), .A2(n4783), .A3(n7392), .ZN(n7394) );
  INV_X1 U9160 ( .A(n7410), .ZN(n7393) );
  OAI21_X1 U9161 ( .B1(n7394), .B2(n7393), .A(n8285), .ZN(n7400) );
  AOI21_X1 U9162 ( .B1(n8266), .B2(n8560), .A(n7395), .ZN(n7396) );
  OAI21_X1 U9163 ( .B1(n8419), .B2(n8268), .A(n7396), .ZN(n7397) );
  AOI21_X1 U9164 ( .B1(n7398), .B2(n8228), .A(n7397), .ZN(n7399) );
  OAI211_X1 U9165 ( .C1(n7401), .C2(n8223), .A(n7400), .B(n7399), .ZN(P2_U3161) );
  INV_X1 U9166 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7404) );
  OAI222_X1 U9167 ( .A1(n9729), .A2(n7404), .B1(n9732), .B2(n7403), .C1(n7402), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U9168 ( .A(n7405), .ZN(n7420) );
  OAI222_X1 U9169 ( .A1(n9034), .A2(n7420), .B1(P2_U3151), .B2(n7406), .C1(
        n10074), .C2(n9025), .ZN(P2_U3274) );
  NAND2_X1 U9170 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  XNOR2_X1 U9171 ( .A(n9878), .B(n6803), .ZN(n7662) );
  XNOR2_X1 U9172 ( .A(n7662), .B(n8560), .ZN(n7411) );
  NAND2_X1 U9173 ( .A1(n7412), .A2(n7411), .ZN(n7665) );
  OAI211_X1 U9174 ( .C1(n7412), .C2(n7411), .A(n7665), .B(n8285), .ZN(n7418)
         );
  AND2_X1 U9175 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7493) );
  AOI21_X1 U9176 ( .B1(n8288), .B2(n8561), .A(n7493), .ZN(n7414) );
  OR2_X1 U9177 ( .A1(n8290), .A2(n8426), .ZN(n7413) );
  OAI211_X1 U9178 ( .C1(n8223), .C2(n7415), .A(n7414), .B(n7413), .ZN(n7416)
         );
  AOI21_X1 U9179 ( .B1(n9878), .B2(n8228), .A(n7416), .ZN(n7417) );
  NAND2_X1 U9180 ( .A1(n7418), .A2(n7417), .ZN(P2_U3171) );
  OAI222_X1 U9181 ( .A1(n9729), .A2(n7421), .B1(n9732), .B2(n7420), .C1(n7419), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9182 ( .A(n9801), .ZN(n9792) );
  OAI21_X1 U9183 ( .B1(n7423), .B2(n7425), .A(n7422), .ZN(n9764) );
  INV_X1 U9184 ( .A(n9764), .ZN(n7429) );
  XOR2_X1 U9185 ( .A(n7425), .B(n7424), .Z(n7427) );
  AOI22_X1 U9186 ( .A1(n9267), .A2(n9196), .B1(n9237), .B2(n9269), .ZN(n7510)
         );
  INV_X1 U9187 ( .A(n7510), .ZN(n7426) );
  AOI21_X1 U9188 ( .B1(n7427), .B2(n9575), .A(n7426), .ZN(n9766) );
  OAI211_X1 U9189 ( .C1(n7433), .C2(n7428), .A(n4408), .B(n6447), .ZN(n9761)
         );
  OAI211_X1 U9190 ( .C1(n9792), .C2(n7429), .A(n9766), .B(n9761), .ZN(n7435)
         );
  OAI22_X1 U9191 ( .A1(n9717), .A2(n7433), .B1(n9713), .B2(n4962), .ZN(n7430)
         );
  AOI21_X1 U9192 ( .B1(n7435), .B2(n9713), .A(n7430), .ZN(n7431) );
  INV_X1 U9193 ( .A(n7431), .ZN(P1_U3468) );
  INV_X1 U9194 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7432) );
  OAI22_X1 U9195 ( .A1(n9659), .A2(n7433), .B1(n9818), .B2(n7432), .ZN(n7434)
         );
  AOI21_X1 U9196 ( .B1(n7435), .B2(n9818), .A(n7434), .ZN(n7436) );
  INV_X1 U9197 ( .A(n7436), .ZN(P1_U3527) );
  XNOR2_X1 U9198 ( .A(n7437), .B(n7444), .ZN(n7438) );
  NAND2_X1 U9199 ( .A1(n7438), .A2(n9829), .ZN(n7440) );
  AOI22_X1 U9200 ( .A1(n7681), .A2(n9826), .B1(n9824), .B2(n8559), .ZN(n7439)
         );
  NAND2_X1 U9201 ( .A1(n7440), .A2(n7439), .ZN(n9888) );
  INV_X1 U9202 ( .A(n9888), .ZN(n7448) );
  OAI21_X1 U9203 ( .B1(n7441), .B2(n7444), .A(n7443), .ZN(n9890) );
  INV_X1 U9204 ( .A(n7687), .ZN(n9887) );
  NOR2_X1 U9205 ( .A1(n9887), .A2(n8738), .ZN(n7446) );
  OAI22_X1 U9206 ( .A1(n8894), .A2(n5858), .B1(n7685), .B2(n9821), .ZN(n7445)
         );
  AOI211_X1 U9207 ( .C1(n9890), .C2(n7811), .A(n7446), .B(n7445), .ZN(n7447)
         );
  OAI21_X1 U9208 ( .B1(n7448), .B2(n9839), .A(n7447), .ZN(P2_U3222) );
  NAND2_X1 U9209 ( .A1(n7422), .A2(n7449), .ZN(n7451) );
  NAND2_X1 U9210 ( .A1(n7451), .A2(n7452), .ZN(n7450) );
  OAI21_X1 U9211 ( .B1(n7451), .B2(n7452), .A(n7450), .ZN(n7473) );
  INV_X1 U9212 ( .A(n7473), .ZN(n7464) );
  XOR2_X1 U9213 ( .A(n7453), .B(n7452), .Z(n7457) );
  OAI22_X1 U9214 ( .A1(n7455), .A2(n9235), .B1(n7454), .B2(n9220), .ZN(n7566)
         );
  INV_X1 U9215 ( .A(n7566), .ZN(n7456) );
  OAI21_X1 U9216 ( .B1(n7457), .B2(n9497), .A(n7456), .ZN(n7466) );
  NAND2_X1 U9217 ( .A1(n7466), .A2(n9568), .ZN(n7463) );
  AOI211_X1 U9218 ( .C1(n7458), .C2(n4408), .A(n9579), .B(n4334), .ZN(n7465)
         );
  INV_X1 U9219 ( .A(n7459), .ZN(n7570) );
  AOI22_X1 U9220 ( .A1(n9778), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7570), .B2(
        n9767), .ZN(n7460) );
  OAI21_X1 U9221 ( .B1(n9556), .B2(n7568), .A(n7460), .ZN(n7461) );
  AOI21_X1 U9222 ( .B1(n7465), .B2(n9772), .A(n7461), .ZN(n7462) );
  OAI211_X1 U9223 ( .C1(n7464), .C2(n9589), .A(n7463), .B(n7462), .ZN(P1_U3287) );
  NOR2_X1 U9224 ( .A1(n7466), .A2(n7465), .ZN(n7475) );
  INV_X1 U9225 ( .A(n9653), .ZN(n7469) );
  INV_X1 U9226 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7467) );
  OAI22_X1 U9227 ( .A1(n9659), .A2(n7568), .B1(n9818), .B2(n7467), .ZN(n7468)
         );
  AOI21_X1 U9228 ( .B1(n7473), .B2(n7469), .A(n7468), .ZN(n7470) );
  OAI21_X1 U9229 ( .B1(n7475), .B2(n9816), .A(n7470), .ZN(P1_U3528) );
  INV_X1 U9230 ( .A(n9711), .ZN(n7472) );
  OAI22_X1 U9231 ( .A1(n9717), .A2(n7568), .B1(n9713), .B2(n4984), .ZN(n7471)
         );
  AOI21_X1 U9232 ( .B1(n7473), .B2(n7472), .A(n7471), .ZN(n7474) );
  OAI21_X1 U9233 ( .B1(n7475), .B2(n9809), .A(n7474), .ZN(P1_U3471) );
  INV_X1 U9234 ( .A(n8344), .ZN(n8444) );
  XNOR2_X1 U9235 ( .A(n7476), .B(n8444), .ZN(n7478) );
  OAI22_X1 U9236 ( .A1(n7794), .A2(n8864), .B1(n7886), .B2(n8866), .ZN(n7477)
         );
  AOI21_X1 U9237 ( .B1(n7478), .B2(n9829), .A(n7477), .ZN(n9898) );
  OAI22_X1 U9238 ( .A1(n8894), .A2(n7820), .B1(n7797), .B2(n9821), .ZN(n7479)
         );
  AOI21_X1 U9239 ( .B1(n9893), .B2(n8899), .A(n7479), .ZN(n7484) );
  NAND2_X1 U9240 ( .A1(n7443), .A2(n8440), .ZN(n7480) );
  NAND2_X1 U9241 ( .A1(n7480), .A2(n8344), .ZN(n7481) );
  AND2_X1 U9242 ( .A1(n7482), .A2(n7481), .ZN(n9896) );
  NAND2_X1 U9243 ( .A1(n9896), .A2(n7811), .ZN(n7483) );
  OAI211_X1 U9244 ( .C1(n9898), .C2(n9839), .A(n7484), .B(n7483), .ZN(P2_U3221) );
  AOI21_X1 U9245 ( .B1(n7486), .B2(n5833), .A(n7546), .ZN(n7503) );
  INV_X1 U9246 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U9247 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6091), .Z(n7538) );
  XNOR2_X1 U9248 ( .A(n7538), .B(n7545), .ZN(n7491) );
  OR2_X1 U9249 ( .A1(n7487), .A2(n7497), .ZN(n7489) );
  NAND2_X1 U9250 ( .A1(n7491), .A2(n7490), .ZN(n7539) );
  OAI21_X1 U9251 ( .B1(n7491), .B2(n7490), .A(n7539), .ZN(n7492) );
  NAND2_X1 U9252 ( .A1(n7492), .A2(n8664), .ZN(n7495) );
  INV_X1 U9253 ( .A(n7493), .ZN(n7494) );
  OAI211_X1 U9254 ( .C1(n10061), .C2(n8704), .A(n7495), .B(n7494), .ZN(n7501)
         );
  AOI21_X1 U9255 ( .B1(n5828), .B2(n7498), .A(n4356), .ZN(n7499) );
  NOR2_X1 U9256 ( .A1(n7499), .A2(n8689), .ZN(n7500) );
  AOI211_X1 U9257 ( .C1(n8676), .C2(n7545), .A(n7501), .B(n7500), .ZN(n7502)
         );
  OAI21_X1 U9258 ( .B1(n7503), .B2(n8731), .A(n7502), .ZN(P2_U3191) );
  XOR2_X1 U9259 ( .A(n7504), .B(n7561), .Z(n7507) );
  INV_X1 U9260 ( .A(n7505), .ZN(n7506) );
  NAND2_X1 U9261 ( .A1(n7507), .A2(n7506), .ZN(n7560) );
  OAI21_X1 U9262 ( .B1(n7507), .B2(n7506), .A(n7560), .ZN(n7508) );
  NAND2_X1 U9263 ( .A1(n7508), .A2(n6436), .ZN(n7513) );
  OAI22_X1 U9264 ( .A1(n7510), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7509), .ZN(n7511) );
  AOI21_X1 U9265 ( .B1(n9758), .B2(n9228), .A(n7511), .ZN(n7512) );
  OAI211_X1 U9266 ( .C1(n9226), .C2(n9755), .A(n7513), .B(n7512), .ZN(P1_U3227) );
  NAND2_X1 U9267 ( .A1(n7515), .A2(n7514), .ZN(n7516) );
  NAND2_X1 U9268 ( .A1(n7516), .A2(n7523), .ZN(n7517) );
  NAND2_X1 U9269 ( .A1(n7517), .A2(n7717), .ZN(n7521) );
  OR2_X1 U9270 ( .A1(n7518), .A2(n9220), .ZN(n7520) );
  NAND2_X1 U9271 ( .A1(n9262), .A2(n9196), .ZN(n7519) );
  NAND2_X1 U9272 ( .A1(n7520), .A2(n7519), .ZN(n9063) );
  AOI21_X1 U9273 ( .B1(n7521), .B2(n9575), .A(n9063), .ZN(n7589) );
  OAI21_X1 U9274 ( .B1(n7524), .B2(n7523), .A(n7522), .ZN(n7587) );
  NAND2_X1 U9275 ( .A1(n7587), .A2(n9763), .ZN(n7531) );
  OAI22_X1 U9276 ( .A1(n9568), .A2(n7525), .B1(n9065), .B2(n9754), .ZN(n7529)
         );
  OAI211_X1 U9277 ( .C1(n7527), .C2(n6475), .A(n6447), .B(n7526), .ZN(n7588)
         );
  NOR2_X1 U9278 ( .A1(n7588), .A2(n9760), .ZN(n7528) );
  AOI211_X1 U9279 ( .C1(n9769), .C2(n9067), .A(n7529), .B(n7528), .ZN(n7530)
         );
  OAI211_X1 U9280 ( .C1(n9778), .C2(n7589), .A(n7531), .B(n7530), .ZN(P1_U3283) );
  NOR2_X1 U9281 ( .A1(n7545), .A2(n7532), .ZN(n7533) );
  NAND2_X1 U9282 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7549), .ZN(n7534) );
  OAI21_X1 U9283 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7549), .A(n7534), .ZN(
        n7597) );
  AOI21_X1 U9284 ( .B1(n5855), .B2(n7535), .A(n7826), .ZN(n7559) );
  MUX2_X1 U9285 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6091), .Z(n7833) );
  XNOR2_X1 U9286 ( .A(n7833), .B(n7825), .ZN(n7543) );
  MUX2_X1 U9287 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6091), .Z(n7536) );
  OR2_X1 U9288 ( .A1(n7536), .A2(n7549), .ZN(n7541) );
  XNOR2_X1 U9289 ( .A(n7536), .B(n7612), .ZN(n7601) );
  OR2_X1 U9290 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  NAND2_X1 U9291 ( .A1(n7540), .A2(n7539), .ZN(n7600) );
  NAND2_X1 U9292 ( .A1(n7601), .A2(n7600), .ZN(n7599) );
  NAND2_X1 U9293 ( .A1(n7541), .A2(n7599), .ZN(n7542) );
  NAND2_X1 U9294 ( .A1(n7543), .A2(n7542), .ZN(n7834) );
  OAI21_X1 U9295 ( .B1(n7543), .B2(n7542), .A(n7834), .ZN(n7557) );
  INV_X1 U9296 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7554) );
  NOR2_X1 U9297 ( .A1(n7545), .A2(n7544), .ZN(n7547) );
  NAND2_X1 U9298 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7549), .ZN(n7548) );
  OAI21_X1 U9299 ( .B1(n7549), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7548), .ZN(
        n7608) );
  XNOR2_X1 U9300 ( .A(n7825), .B(n7817), .ZN(n7550) );
  AOI21_X1 U9301 ( .B1(n7550), .B2(n5858), .A(n7818), .ZN(n7551) );
  OR2_X1 U9302 ( .A1(n8731), .A2(n7551), .ZN(n7553) );
  AND2_X1 U9303 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7680) );
  INV_X1 U9304 ( .A(n7680), .ZN(n7552) );
  OAI211_X1 U9305 ( .C1(n8704), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7556)
         );
  NOR2_X1 U9306 ( .A1(n8724), .A2(n7832), .ZN(n7555) );
  AOI211_X1 U9307 ( .C1(n8664), .C2(n7557), .A(n7556), .B(n7555), .ZN(n7558)
         );
  OAI21_X1 U9308 ( .B1(n7559), .B2(n8689), .A(n7558), .ZN(P2_U3193) );
  OAI21_X1 U9309 ( .B1(n7561), .B2(n7504), .A(n7560), .ZN(n7565) );
  XNOR2_X1 U9310 ( .A(n7563), .B(n7562), .ZN(n7564) );
  XNOR2_X1 U9311 ( .A(n7565), .B(n7564), .ZN(n7572) );
  AOI22_X1 U9312 ( .A1(n7566), .A2(n9224), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7567) );
  OAI21_X1 U9313 ( .B1(n7568), .B2(n10096), .A(n7567), .ZN(n7569) );
  AOI21_X1 U9314 ( .B1(n7570), .B2(n9242), .A(n7569), .ZN(n7571) );
  OAI21_X1 U9315 ( .B1(n7572), .B2(n10103), .A(n7571), .ZN(P1_U3239) );
  XOR2_X1 U9316 ( .A(n7574), .B(n7573), .Z(n7580) );
  INV_X1 U9317 ( .A(n9743), .ZN(n7578) );
  OAI22_X1 U9318 ( .A1(n7575), .A2(n9220), .B1(n7651), .B2(n9235), .ZN(n7760)
         );
  AOI22_X1 U9319 ( .A1(n7760), .A2(n9224), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7576) );
  OAI21_X1 U9320 ( .B1(n7767), .B2(n10096), .A(n7576), .ZN(n7577) );
  AOI21_X1 U9321 ( .B1(n7578), .B2(n9242), .A(n7577), .ZN(n7579) );
  OAI21_X1 U9322 ( .B1(n7580), .B2(n10103), .A(n7579), .ZN(P1_U3213) );
  INV_X1 U9323 ( .A(n7581), .ZN(n7585) );
  OAI222_X1 U9324 ( .A1(n9729), .A2(n7583), .B1(n9732), .B2(n7585), .C1(
        P1_U3086), .C2(n7582), .ZN(P1_U3333) );
  OAI222_X1 U9325 ( .A1(n9025), .A2(n7586), .B1(n9034), .B2(n7585), .C1(n7584), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U9326 ( .A(n7587), .ZN(n7595) );
  NAND2_X1 U9327 ( .A1(n7589), .A2(n7588), .ZN(n7593) );
  OAI22_X1 U9328 ( .A1(n9717), .A2(n6475), .B1(n9794), .B2(n5084), .ZN(n7590)
         );
  AOI21_X1 U9329 ( .B1(n7593), .B2(n9713), .A(n7590), .ZN(n7591) );
  OAI21_X1 U9330 ( .B1(n7595), .B2(n9711), .A(n7591), .ZN(P1_U3483) );
  OAI22_X1 U9331 ( .A1(n9659), .A2(n6475), .B1(n9818), .B2(n6894), .ZN(n7592)
         );
  AOI21_X1 U9332 ( .B1(n7593), .B2(n9818), .A(n7592), .ZN(n7594) );
  OAI21_X1 U9333 ( .B1(n7595), .B2(n9653), .A(n7594), .ZN(P1_U3532) );
  AOI21_X1 U9334 ( .B1(n7598), .B2(n7597), .A(n7596), .ZN(n7614) );
  INV_X1 U9335 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7606) );
  OAI21_X1 U9336 ( .B1(n7601), .B2(n7600), .A(n7599), .ZN(n7602) );
  NAND2_X1 U9337 ( .A1(n7602), .A2(n8664), .ZN(n7605) );
  INV_X1 U9338 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7603) );
  NOR2_X1 U9339 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7603), .ZN(n7669) );
  INV_X1 U9340 ( .A(n7669), .ZN(n7604) );
  OAI211_X1 U9341 ( .C1(n7606), .C2(n8704), .A(n7605), .B(n7604), .ZN(n7611)
         );
  AOI21_X1 U9342 ( .B1(n4406), .B2(n7608), .A(n7607), .ZN(n7609) );
  NOR2_X1 U9343 ( .A1(n7609), .A2(n8731), .ZN(n7610) );
  AOI211_X1 U9344 ( .C1(n8676), .C2(n7612), .A(n7611), .B(n7610), .ZN(n7613)
         );
  OAI21_X1 U9345 ( .B1(n7614), .B2(n8689), .A(n7613), .ZN(P2_U3192) );
  NAND2_X1 U9346 ( .A1(n7754), .A2(n4482), .ZN(n7757) );
  NAND2_X1 U9347 ( .A1(n7757), .A2(n7615), .ZN(n7616) );
  XNOR2_X1 U9348 ( .A(n7616), .B(n7618), .ZN(n7621) );
  AOI22_X1 U9349 ( .A1(n9264), .A2(n9196), .B1(n9237), .B2(n9266), .ZN(n7636)
         );
  OAI21_X1 U9350 ( .B1(n7619), .B2(n7618), .A(n7617), .ZN(n9799) );
  NAND2_X1 U9351 ( .A1(n9799), .A2(n7761), .ZN(n7620) );
  OAI211_X1 U9352 ( .C1(n7621), .C2(n9497), .A(n7636), .B(n7620), .ZN(n9797)
         );
  INV_X1 U9353 ( .A(n9797), .ZN(n7629) );
  INV_X1 U9354 ( .A(n7762), .ZN(n7623) );
  INV_X1 U9355 ( .A(n7653), .ZN(n7622) );
  OAI211_X1 U9356 ( .C1(n9796), .C2(n7623), .A(n7622), .B(n6447), .ZN(n9795)
         );
  OAI22_X1 U9357 ( .A1(n9745), .A2(n7624), .B1(n7634), .B2(n9754), .ZN(n7625)
         );
  AOI21_X1 U9358 ( .B1(n9769), .B2(n7639), .A(n7625), .ZN(n7626) );
  OAI21_X1 U9359 ( .B1(n9795), .B2(n9760), .A(n7626), .ZN(n7627) );
  AOI21_X1 U9360 ( .B1(n9799), .B2(n9773), .A(n7627), .ZN(n7628) );
  OAI21_X1 U9361 ( .B1(n7629), .B2(n9778), .A(n7628), .ZN(P1_U3285) );
  XNOR2_X1 U9362 ( .A(n7631), .B(n7630), .ZN(n7632) );
  XNOR2_X1 U9363 ( .A(n7633), .B(n7632), .ZN(n7641) );
  NOR2_X1 U9364 ( .A1(n9226), .A2(n7634), .ZN(n7638) );
  OAI22_X1 U9365 ( .A1(n7636), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7635), .ZN(n7637) );
  AOI211_X1 U9366 ( .C1(n7639), .C2(n9228), .A(n7638), .B(n7637), .ZN(n7640)
         );
  OAI21_X1 U9367 ( .B1(n7641), .B2(n10103), .A(n7640), .ZN(P1_U3221) );
  OR2_X1 U9368 ( .A1(n7642), .A2(n7648), .ZN(n7643) );
  NAND2_X1 U9369 ( .A1(n7644), .A2(n7643), .ZN(n9802) );
  INV_X1 U9370 ( .A(n9802), .ZN(n7661) );
  NAND2_X1 U9371 ( .A1(n7757), .A2(n7645), .ZN(n7647) );
  NAND2_X1 U9372 ( .A1(n7647), .A2(n7646), .ZN(n7649) );
  XNOR2_X1 U9373 ( .A(n7649), .B(n7648), .ZN(n7650) );
  NAND2_X1 U9374 ( .A1(n7650), .A2(n9575), .ZN(n7652) );
  OR2_X1 U9375 ( .A1(n7651), .A2(n9220), .ZN(n7858) );
  NAND2_X1 U9376 ( .A1(n7652), .A2(n7858), .ZN(n9807) );
  XNOR2_X1 U9377 ( .A(n7653), .B(n7657), .ZN(n7654) );
  NOR2_X1 U9378 ( .A1(n7720), .A2(n9235), .ZN(n7860) );
  AOI21_X1 U9379 ( .B1(n7654), .B2(n6447), .A(n7860), .ZN(n9803) );
  OAI22_X1 U9380 ( .A1(n9745), .A2(n7655), .B1(n7863), .B2(n9754), .ZN(n7656)
         );
  AOI21_X1 U9381 ( .B1(n9769), .B2(n7657), .A(n7656), .ZN(n7658) );
  OAI21_X1 U9382 ( .B1(n9803), .B2(n9760), .A(n7658), .ZN(n7659) );
  AOI21_X1 U9383 ( .B1(n9807), .B2(n9745), .A(n7659), .ZN(n7660) );
  OAI21_X1 U9384 ( .B1(n7661), .B2(n9589), .A(n7660), .ZN(P1_U3284) );
  INV_X1 U9385 ( .A(n7662), .ZN(n7663) );
  NAND2_X1 U9386 ( .A1(n7663), .A2(n8560), .ZN(n7664) );
  NAND2_X1 U9387 ( .A1(n7665), .A2(n7664), .ZN(n7676) );
  XNOR2_X1 U9388 ( .A(n7676), .B(n8426), .ZN(n7667) );
  XNOR2_X1 U9389 ( .A(n9884), .B(n8219), .ZN(n7666) );
  OAI21_X1 U9390 ( .B1(n7667), .B2(n7666), .A(n7679), .ZN(n7668) );
  NAND2_X1 U9391 ( .A1(n7668), .A2(n8285), .ZN(n7675) );
  AOI21_X1 U9392 ( .B1(n8288), .B2(n8560), .A(n7669), .ZN(n7671) );
  OR2_X1 U9393 ( .A1(n8290), .A2(n7794), .ZN(n7670) );
  OAI211_X1 U9394 ( .C1(n8223), .C2(n7672), .A(n7671), .B(n7670), .ZN(n7673)
         );
  AOI21_X1 U9395 ( .B1(n9884), .B2(n8228), .A(n7673), .ZN(n7674) );
  NAND2_X1 U9396 ( .A1(n7675), .A2(n7674), .ZN(P2_U3157) );
  OR2_X1 U9397 ( .A1(n7676), .A2(n7681), .ZN(n7678) );
  XNOR2_X1 U9398 ( .A(n8343), .B(n8079), .ZN(n7791) );
  AND2_X1 U9399 ( .A1(n7678), .A2(n7791), .ZN(n7677) );
  NAND2_X1 U9400 ( .A1(n7679), .A2(n7677), .ZN(n7987) );
  NAND2_X1 U9401 ( .A1(n7987), .A2(n8285), .ZN(n7690) );
  AOI21_X1 U9402 ( .B1(n7679), .B2(n7678), .A(n7791), .ZN(n7689) );
  AOI21_X1 U9403 ( .B1(n8288), .B2(n7681), .A(n7680), .ZN(n7684) );
  OR2_X1 U9404 ( .A1(n8290), .A2(n7682), .ZN(n7683) );
  OAI211_X1 U9405 ( .C1(n8223), .C2(n7685), .A(n7684), .B(n7683), .ZN(n7686)
         );
  AOI21_X1 U9406 ( .B1(n7687), .B2(n8228), .A(n7686), .ZN(n7688) );
  OAI21_X1 U9407 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(P2_U3176) );
  NAND2_X1 U9408 ( .A1(n7695), .A2(n7691), .ZN(n7692) );
  OAI211_X1 U9409 ( .C1(n7693), .C2(n9025), .A(n7692), .B(n8553), .ZN(P2_U3272) );
  NAND2_X1 U9410 ( .A1(n7695), .A2(n7694), .ZN(n7697) );
  OAI211_X1 U9411 ( .C1(n10051), .C2(n9729), .A(n7697), .B(n7696), .ZN(
        P1_U3332) );
  INV_X1 U9412 ( .A(n7734), .ZN(n7699) );
  NAND2_X1 U9413 ( .A1(n9360), .A2(n7699), .ZN(n7700) );
  AOI21_X1 U9414 ( .B1(n7701), .B2(n9583), .A(n7700), .ZN(n7711) );
  NOR2_X1 U9415 ( .A1(n9651), .A2(n7704), .ZN(n7730) );
  AOI211_X1 U9416 ( .C1(n7704), .C2(n9651), .A(n7730), .B(n9356), .ZN(n7710)
         );
  INV_X1 U9417 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U9418 ( .A1(n9359), .A2(n7705), .ZN(n7707) );
  NAND2_X1 U9419 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n7706) );
  OAI211_X1 U9420 ( .C1(n7708), .C2(n9366), .A(n7707), .B(n7706), .ZN(n7709)
         );
  OR3_X1 U9421 ( .A1(n7711), .A2(n7710), .A3(n7709), .ZN(P1_U3258) );
  XNOR2_X1 U9422 ( .A(n7713), .B(n7712), .ZN(n9660) );
  INV_X1 U9423 ( .A(n7714), .ZN(n7719) );
  AOI21_X1 U9424 ( .B1(n7717), .B2(n7716), .A(n7715), .ZN(n7718) );
  NOR3_X1 U9425 ( .A1(n7719), .A2(n7718), .A3(n9497), .ZN(n7722) );
  OAI22_X1 U9426 ( .A1(n7721), .A2(n9235), .B1(n7720), .B2(n9220), .ZN(n9210)
         );
  AOI211_X1 U9427 ( .C1(n9660), .C2(n7761), .A(n7722), .B(n9210), .ZN(n9664)
         );
  AOI211_X1 U9428 ( .C1(n9662), .C2(n7526), .A(n9579), .B(n4333), .ZN(n9661)
         );
  NOR2_X1 U9429 ( .A1(n9556), .A2(n7723), .ZN(n7726) );
  OAI22_X1 U9430 ( .A1(n9568), .A2(n7724), .B1(n9212), .B2(n9754), .ZN(n7725)
         );
  AOI211_X1 U9431 ( .C1(n9661), .C2(n9772), .A(n7726), .B(n7725), .ZN(n7728)
         );
  NAND2_X1 U9432 ( .A1(n9660), .A2(n9773), .ZN(n7727) );
  OAI211_X1 U9433 ( .C1(n9664), .C2(n9778), .A(n7728), .B(n7727), .ZN(P1_U3282) );
  NOR2_X1 U9434 ( .A1(n7729), .A2(n7732), .ZN(n7731) );
  XNOR2_X1 U9435 ( .A(n7739), .B(n9645), .ZN(n7899) );
  XNOR2_X1 U9436 ( .A(n7898), .B(n7899), .ZN(n7744) );
  NOR2_X1 U9437 ( .A1(n7733), .A2(n7732), .ZN(n7735) );
  XNOR2_X1 U9438 ( .A(n7739), .B(n9559), .ZN(n7736) );
  NAND2_X1 U9439 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  NAND3_X1 U9440 ( .A1(n7903), .A2(n9360), .A3(n7738), .ZN(n7743) );
  INV_X1 U9441 ( .A(n7739), .ZN(n7901) );
  INV_X1 U9442 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U9443 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9140) );
  OAI21_X1 U9444 ( .B1(n9366), .B2(n7740), .A(n9140), .ZN(n7741) );
  AOI21_X1 U9445 ( .B1(n9359), .B2(n7901), .A(n7741), .ZN(n7742) );
  OAI211_X1 U9446 ( .C1(n7744), .C2(n9356), .A(n7743), .B(n7742), .ZN(P1_U3259) );
  XOR2_X1 U9447 ( .A(n7745), .B(n8346), .Z(n7746) );
  AOI222_X1 U9448 ( .A1(n9829), .A2(n7746), .B1(n8557), .B2(n9824), .C1(n8559), 
        .C2(n9826), .ZN(n7787) );
  INV_X1 U9449 ( .A(n9823), .ZN(n7807) );
  INV_X1 U9450 ( .A(n7936), .ZN(n7747) );
  AOI22_X1 U9451 ( .A1(n8451), .A2(n7807), .B1(n8898), .B2(n7747), .ZN(n7748)
         );
  AOI21_X1 U9452 ( .B1(n7787), .B2(n7748), .A(n9839), .ZN(n7752) );
  XNOR2_X1 U9453 ( .A(n7749), .B(n8346), .ZN(n7790) );
  OAI22_X1 U9454 ( .A1(n7790), .A2(n8903), .B1(n7750), .B2(n9837), .ZN(n7751)
         );
  OR2_X1 U9455 ( .A1(n7752), .A2(n7751), .ZN(P2_U3220) );
  INV_X1 U9456 ( .A(n9751), .ZN(n7763) );
  INV_X1 U9457 ( .A(n7754), .ZN(n7756) );
  NAND2_X1 U9458 ( .A1(n7756), .A2(n7755), .ZN(n7758) );
  AOI21_X1 U9459 ( .B1(n7758), .B2(n7757), .A(n9497), .ZN(n7759) );
  AOI211_X1 U9460 ( .C1(n7761), .C2(n9751), .A(n7760), .B(n7759), .ZN(n9753)
         );
  OAI211_X1 U9461 ( .C1(n4334), .C2(n7767), .A(n6447), .B(n7762), .ZN(n9749)
         );
  OAI211_X1 U9462 ( .C1(n7763), .C2(n9781), .A(n9753), .B(n9749), .ZN(n7769)
         );
  OAI22_X1 U9463 ( .A1(n9717), .A2(n7767), .B1(n9794), .B2(n5013), .ZN(n7764)
         );
  AOI21_X1 U9464 ( .B1(n7769), .B2(n9713), .A(n7764), .ZN(n7765) );
  INV_X1 U9465 ( .A(n7765), .ZN(P1_U3474) );
  INV_X1 U9466 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7766) );
  OAI22_X1 U9467 ( .A1(n9659), .A2(n7767), .B1(n9818), .B2(n7766), .ZN(n7768)
         );
  AOI21_X1 U9468 ( .B1(n7769), .B2(n9818), .A(n7768), .ZN(n7770) );
  INV_X1 U9469 ( .A(n7770), .ZN(P1_U3529) );
  XOR2_X1 U9470 ( .A(n7771), .B(n7773), .Z(n7847) );
  AOI22_X1 U9471 ( .A1(n9124), .A2(n6528), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n9809), .ZN(n7780) );
  OAI211_X1 U9472 ( .C1(n7774), .C2(n7773), .A(n7772), .B(n9575), .ZN(n7777)
         );
  NAND2_X1 U9473 ( .A1(n9262), .A2(n9237), .ZN(n7776) );
  NAND2_X1 U9474 ( .A1(n9260), .A2(n9196), .ZN(n7775) );
  AND2_X1 U9475 ( .A1(n7776), .A2(n7775), .ZN(n9122) );
  OAI211_X1 U9476 ( .C1(n4333), .C2(n7778), .A(n6447), .B(n4405), .ZN(n7850)
         );
  NAND2_X1 U9477 ( .A1(n7855), .A2(n7850), .ZN(n7781) );
  NAND2_X1 U9478 ( .A1(n7781), .A2(n9713), .ZN(n7779) );
  OAI211_X1 U9479 ( .C1(n7847), .C2(n9711), .A(n7780), .B(n7779), .ZN(P1_U3489) );
  AOI22_X1 U9480 ( .A1(n9124), .A2(n6535), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n9816), .ZN(n7783) );
  NAND2_X1 U9481 ( .A1(n7781), .A2(n9818), .ZN(n7782) );
  OAI211_X1 U9482 ( .C1(n7847), .C2(n9653), .A(n7783), .B(n7782), .ZN(P1_U3534) );
  INV_X1 U9483 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7784) );
  MUX2_X1 U9484 ( .A(n7784), .B(n7787), .S(n9899), .Z(n7786) );
  NAND2_X1 U9485 ( .A1(n8451), .A2(n9010), .ZN(n7785) );
  OAI211_X1 U9486 ( .C1(n7790), .C2(n9018), .A(n7786), .B(n7785), .ZN(P2_U3429) );
  MUX2_X1 U9487 ( .A(n5886), .B(n7787), .S(n9915), .Z(n7789) );
  NAND2_X1 U9488 ( .A1(n8451), .A2(n8939), .ZN(n7788) );
  OAI211_X1 U9489 ( .C1(n8943), .C2(n7790), .A(n7789), .B(n7788), .ZN(P2_U3472) );
  INV_X1 U9490 ( .A(n7791), .ZN(n7793) );
  NAND2_X1 U9491 ( .A1(n7793), .A2(n7792), .ZN(n7883) );
  NAND2_X1 U9492 ( .A1(n7987), .A2(n7883), .ZN(n7929) );
  XNOR2_X1 U9493 ( .A(n9893), .B(n8219), .ZN(n7880) );
  XNOR2_X1 U9494 ( .A(n7880), .B(n8559), .ZN(n7928) );
  XNOR2_X1 U9495 ( .A(n7929), .B(n7928), .ZN(n7800) );
  AND2_X1 U9496 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7840) );
  NOR2_X1 U9497 ( .A1(n8268), .A2(n7794), .ZN(n7795) );
  AOI211_X1 U9498 ( .C1(n8266), .C2(n8558), .A(n7840), .B(n7795), .ZN(n7796)
         );
  OAI21_X1 U9499 ( .B1(n7797), .B2(n8223), .A(n7796), .ZN(n7798) );
  AOI21_X1 U9500 ( .B1(n9893), .B2(n8228), .A(n7798), .ZN(n7799) );
  OAI21_X1 U9501 ( .B1(n7800), .B2(n8272), .A(n7799), .ZN(P2_U3164) );
  INV_X1 U9502 ( .A(n7801), .ZN(n7815) );
  OAI222_X1 U9503 ( .A1(n9034), .A2(n7815), .B1(P2_U3151), .B2(n7803), .C1(
        n7802), .C2(n9025), .ZN(P2_U3271) );
  INV_X1 U9504 ( .A(n8460), .ZN(n7804) );
  INV_X1 U9505 ( .A(n8348), .ZN(n8455) );
  XNOR2_X1 U9506 ( .A(n7805), .B(n8455), .ZN(n7806) );
  OAI222_X1 U9507 ( .A1(n8866), .A2(n7891), .B1(n8864), .B2(n7886), .C1(n7806), 
        .C2(n8862), .ZN(n7912) );
  AOI21_X1 U9508 ( .B1(n7807), .B2(n7918), .A(n7912), .ZN(n7813) );
  XNOR2_X1 U9509 ( .A(n7808), .B(n8348), .ZN(n7920) );
  OAI22_X1 U9510 ( .A1(n8894), .A2(n7809), .B1(n7894), .B2(n9821), .ZN(n7810)
         );
  AOI21_X1 U9511 ( .B1(n7920), .B2(n7811), .A(n7810), .ZN(n7812) );
  OAI21_X1 U9512 ( .B1(n7813), .B2(n9839), .A(n7812), .ZN(P2_U3219) );
  OAI222_X1 U9513 ( .A1(n9729), .A2(n7816), .B1(n9732), .B2(n7815), .C1(n7814), 
        .C2(P1_U3086), .ZN(P1_U3331) );
  NOR2_X1 U9514 ( .A1(n7825), .A2(n7817), .ZN(n7819) );
  NOR2_X1 U9515 ( .A1(n7819), .A2(n7818), .ZN(n7823) );
  MUX2_X1 U9516 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7820), .S(n7831), .Z(n7822)
         );
  INV_X1 U9517 ( .A(n7941), .ZN(n7821) );
  AOI21_X1 U9518 ( .B1(n7823), .B2(n7822), .A(n7821), .ZN(n7846) );
  MUX2_X1 U9519 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7827), .S(n7831), .Z(n7828)
         );
  INV_X1 U9520 ( .A(n7828), .ZN(n7830) );
  OAI21_X1 U9521 ( .B1(n7829), .B2(n7830), .A(n7954), .ZN(n7844) );
  MUX2_X1 U9522 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6091), .Z(n7943) );
  XNOR2_X1 U9523 ( .A(n7943), .B(n7831), .ZN(n7837) );
  OR2_X1 U9524 ( .A1(n7833), .A2(n7832), .ZN(n7835) );
  NAND2_X1 U9525 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NAND2_X1 U9526 ( .A1(n7837), .A2(n7836), .ZN(n7944) );
  OAI21_X1 U9527 ( .B1(n7837), .B2(n7836), .A(n7944), .ZN(n7841) );
  INV_X1 U9528 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7838) );
  NOR2_X1 U9529 ( .A1(n8704), .A2(n7838), .ZN(n7839) );
  AOI211_X1 U9530 ( .C1(n8664), .C2(n7841), .A(n7840), .B(n7839), .ZN(n7842)
         );
  OAI21_X1 U9531 ( .B1(n7952), .B2(n8724), .A(n7842), .ZN(n7843) );
  AOI21_X1 U9532 ( .B1(n7844), .B2(n8727), .A(n7843), .ZN(n7845) );
  OAI21_X1 U9533 ( .B1(n7846), .B2(n8731), .A(n7845), .ZN(P2_U3194) );
  INV_X1 U9534 ( .A(n7847), .ZN(n7848) );
  NAND2_X1 U9535 ( .A1(n7848), .A2(n9763), .ZN(n7854) );
  OAI22_X1 U9536 ( .A1(n9568), .A2(n7849), .B1(n9118), .B2(n9754), .ZN(n7852)
         );
  NOR2_X1 U9537 ( .A1(n7850), .A2(n9760), .ZN(n7851) );
  AOI211_X1 U9538 ( .C1(n9769), .C2(n9124), .A(n7852), .B(n7851), .ZN(n7853)
         );
  OAI211_X1 U9539 ( .C1(n9778), .C2(n7855), .A(n7854), .B(n7853), .ZN(P1_U3281) );
  XNOR2_X1 U9540 ( .A(n7856), .B(n7857), .ZN(n7866) );
  NOR2_X1 U9541 ( .A1(n10096), .A2(n9805), .ZN(n7865) );
  INV_X1 U9542 ( .A(n7858), .ZN(n7859) );
  OAI21_X1 U9543 ( .B1(n7860), .B2(n7859), .A(n9224), .ZN(n7862) );
  OAI211_X1 U9544 ( .C1(n9226), .C2(n7863), .A(n7862), .B(n7861), .ZN(n7864)
         );
  AOI211_X1 U9545 ( .C1(n7866), .C2(n6436), .A(n7865), .B(n7864), .ZN(n7867)
         );
  INV_X1 U9546 ( .A(n7867), .ZN(P1_U3231) );
  XNOR2_X1 U9547 ( .A(n7868), .B(n7870), .ZN(n7869) );
  AOI22_X1 U9548 ( .A1(n9237), .A2(n9261), .B1(n9259), .B2(n9196), .ZN(n9187)
         );
  OAI21_X1 U9549 ( .B1(n7869), .B2(n9497), .A(n9187), .ZN(n8042) );
  INV_X1 U9550 ( .A(n8042), .ZN(n7877) );
  XNOR2_X1 U9551 ( .A(n7871), .B(n7870), .ZN(n8044) );
  NAND2_X1 U9552 ( .A1(n8044), .A2(n9763), .ZN(n7876) );
  AOI211_X1 U9553 ( .C1(n9190), .C2(n4405), .A(n9579), .B(n8071), .ZN(n8043)
         );
  NOR2_X1 U9554 ( .A1(n8049), .A2(n9556), .ZN(n7874) );
  OAI22_X1 U9555 ( .A1(n9568), .A2(n7872), .B1(n9185), .B2(n9754), .ZN(n7873)
         );
  AOI211_X1 U9556 ( .C1(n8043), .C2(n9772), .A(n7874), .B(n7873), .ZN(n7875)
         );
  OAI211_X1 U9557 ( .C1(n9778), .C2(n7877), .A(n7876), .B(n7875), .ZN(P1_U3280) );
  INV_X1 U9558 ( .A(n7878), .ZN(n7924) );
  OAI222_X1 U9559 ( .A1(n9034), .A2(n7924), .B1(P2_U3151), .B2(n7879), .C1(
        n9991), .C2(n9025), .ZN(P2_U3270) );
  XNOR2_X1 U9560 ( .A(n7918), .B(n8079), .ZN(n7989) );
  XNOR2_X1 U9561 ( .A(n7989), .B(n8557), .ZN(n8026) );
  INV_X1 U9562 ( .A(n7880), .ZN(n7881) );
  NAND2_X1 U9563 ( .A1(n7881), .A2(n8559), .ZN(n7930) );
  XNOR2_X1 U9564 ( .A(n8451), .B(n8219), .ZN(n7887) );
  INV_X1 U9565 ( .A(n7887), .ZN(n7882) );
  NAND2_X1 U9566 ( .A1(n7882), .A2(n8558), .ZN(n7927) );
  AND2_X1 U9567 ( .A1(n7930), .A2(n7927), .ZN(n7884) );
  AND2_X1 U9568 ( .A1(n7883), .A2(n7884), .ZN(n7983) );
  NAND2_X1 U9569 ( .A1(n7987), .A2(n7983), .ZN(n7890) );
  INV_X1 U9570 ( .A(n7884), .ZN(n7885) );
  NOR2_X1 U9571 ( .A1(n7885), .A2(n7928), .ZN(n7889) );
  NAND2_X1 U9572 ( .A1(n7887), .A2(n7886), .ZN(n7926) );
  INV_X1 U9573 ( .A(n7926), .ZN(n7888) );
  NOR2_X1 U9574 ( .A1(n7889), .A2(n7888), .ZN(n7984) );
  XOR2_X1 U9575 ( .A(n8026), .B(n8027), .Z(n7897) );
  NAND2_X1 U9576 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8595) );
  OAI21_X1 U9577 ( .B1(n8290), .B2(n7891), .A(n8595), .ZN(n7892) );
  AOI21_X1 U9578 ( .B1(n8288), .B2(n8558), .A(n7892), .ZN(n7893) );
  OAI21_X1 U9579 ( .B1(n7894), .B2(n8223), .A(n7893), .ZN(n7895) );
  AOI21_X1 U9580 ( .B1(n7918), .B2(n8228), .A(n7895), .ZN(n7896) );
  OAI21_X1 U9581 ( .B1(n7897), .B2(n8272), .A(n7896), .ZN(P2_U3155) );
  XNOR2_X1 U9582 ( .A(n9337), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9338) );
  XOR2_X1 U9583 ( .A(n9338), .B(n9339), .Z(n7911) );
  OR2_X1 U9584 ( .A1(n9337), .A2(n9539), .ZN(n7900) );
  NAND2_X1 U9585 ( .A1(n9337), .A2(n9539), .ZN(n9329) );
  AND2_X1 U9586 ( .A1(n7900), .A2(n9329), .ZN(n7905) );
  NAND2_X1 U9587 ( .A1(n7901), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U9588 ( .A1(n7904), .A2(n7905), .ZN(n9330) );
  OAI21_X1 U9589 ( .B1(n7905), .B2(n7904), .A(n9330), .ZN(n7906) );
  NAND2_X1 U9590 ( .A1(n7906), .A2(n9360), .ZN(n7910) );
  AND2_X1 U9591 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9151) );
  NOR2_X1 U9592 ( .A1(n7907), .A2(n9337), .ZN(n7908) );
  AOI211_X1 U9593 ( .C1(n9739), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9151), .B(
        n7908), .ZN(n7909) );
  OAI211_X1 U9594 ( .C1(n7911), .C2(n9356), .A(n7910), .B(n7909), .ZN(P1_U3260) );
  INV_X1 U9595 ( .A(n7912), .ZN(n7917) );
  MUX2_X1 U9596 ( .A(n7913), .B(n7917), .S(n9915), .Z(n7916) );
  INV_X1 U9597 ( .A(n8943), .ZN(n7914) );
  AOI22_X1 U9598 ( .A1(n7920), .A2(n7914), .B1(n8939), .B2(n7918), .ZN(n7915)
         );
  NAND2_X1 U9599 ( .A1(n7916), .A2(n7915), .ZN(P2_U3473) );
  MUX2_X1 U9600 ( .A(n10042), .B(n7917), .S(n9899), .Z(n7922) );
  INV_X1 U9601 ( .A(n9018), .ZN(n7919) );
  AOI22_X1 U9602 ( .A1(n7920), .A2(n7919), .B1(n9010), .B2(n7918), .ZN(n7921)
         );
  NAND2_X1 U9603 ( .A1(n7922), .A2(n7921), .ZN(P2_U3432) );
  OAI222_X1 U9604 ( .A1(n9729), .A2(n7925), .B1(n9728), .B2(n7924), .C1(n7923), 
        .C2(P1_U3086), .ZN(P1_U3330) );
  NAND2_X1 U9605 ( .A1(n7927), .A2(n7926), .ZN(n7933) );
  NAND2_X1 U9606 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  NAND2_X1 U9607 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  XOR2_X1 U9608 ( .A(n7933), .B(n7932), .Z(n7939) );
  OR2_X1 U9609 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10009), .ZN(n7949) );
  OAI21_X1 U9610 ( .B1(n8290), .B2(n7990), .A(n7949), .ZN(n7934) );
  AOI21_X1 U9611 ( .B1(n8288), .B2(n8559), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9612 ( .B1(n7936), .B2(n8223), .A(n7935), .ZN(n7937) );
  AOI21_X1 U9613 ( .B1(n8451), .B2(n8228), .A(n7937), .ZN(n7938) );
  OAI21_X1 U9614 ( .B1(n7939), .B2(n8272), .A(n7938), .ZN(P2_U3174) );
  NAND2_X1 U9615 ( .A1(n7952), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7940) );
  AOI21_X1 U9616 ( .B1(n7942), .B2(n7750), .A(n8585), .ZN(n7961) );
  INV_X1 U9617 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7951) );
  MUX2_X1 U9618 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6091), .Z(n8589) );
  XNOR2_X1 U9619 ( .A(n8589), .B(n8598), .ZN(n7947) );
  OR2_X1 U9620 ( .A1(n7943), .A2(n7952), .ZN(n7945) );
  NAND2_X1 U9621 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U9622 ( .A1(n7947), .A2(n7946), .ZN(n8590) );
  OAI21_X1 U9623 ( .B1(n7947), .B2(n7946), .A(n8590), .ZN(n7948) );
  NAND2_X1 U9624 ( .A1(n7948), .A2(n8664), .ZN(n7950) );
  OAI211_X1 U9625 ( .C1(n7951), .C2(n8704), .A(n7950), .B(n7949), .ZN(n7959)
         );
  NAND2_X1 U9626 ( .A1(n7952), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7953) );
  AOI21_X1 U9627 ( .B1(n5886), .B2(n7956), .A(n8599), .ZN(n7957) );
  NOR2_X1 U9628 ( .A1(n7957), .A2(n8689), .ZN(n7958) );
  AOI211_X1 U9629 ( .C1(n8676), .C2(n8598), .A(n7959), .B(n7958), .ZN(n7960)
         );
  OAI21_X1 U9630 ( .B1(n7961), .B2(n8731), .A(n7960), .ZN(P2_U3195) );
  XNOR2_X1 U9631 ( .A(n7962), .B(n8463), .ZN(n7978) );
  NAND2_X1 U9632 ( .A1(n7964), .A2(n8463), .ZN(n7965) );
  NAND3_X1 U9633 ( .A1(n7963), .A2(n9829), .A3(n7965), .ZN(n7967) );
  AOI22_X1 U9634 ( .A1(n9826), .A2(n8557), .B1(n8879), .B2(n9824), .ZN(n7966)
         );
  INV_X1 U9635 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7968) );
  MUX2_X1 U9636 ( .A(n7975), .B(n7968), .S(n9901), .Z(n7970) );
  NAND2_X1 U9637 ( .A1(n8025), .A2(n9010), .ZN(n7969) );
  OAI211_X1 U9638 ( .C1(n7978), .C2(n9018), .A(n7970), .B(n7969), .ZN(P2_U3435) );
  MUX2_X1 U9639 ( .A(n7975), .B(n7971), .S(n9839), .Z(n7974) );
  INV_X1 U9640 ( .A(n7972), .ZN(n8038) );
  AOI22_X1 U9641 ( .A1(n8025), .A2(n8899), .B1(n8898), .B2(n8038), .ZN(n7973)
         );
  OAI211_X1 U9642 ( .C1(n7978), .C2(n8903), .A(n7974), .B(n7973), .ZN(P2_U3218) );
  MUX2_X1 U9643 ( .A(n8624), .B(n7975), .S(n9915), .Z(n7977) );
  NAND2_X1 U9644 ( .A1(n8025), .A2(n8939), .ZN(n7976) );
  OAI211_X1 U9645 ( .C1(n7978), .C2(n8943), .A(n7977), .B(n7976), .ZN(P2_U3474) );
  INV_X1 U9646 ( .A(n7979), .ZN(n8023) );
  OAI222_X1 U9647 ( .A1(n9034), .A2(n8023), .B1(P2_U3151), .B2(n7981), .C1(
        n7980), .C2(n9025), .ZN(P2_U3269) );
  INV_X1 U9648 ( .A(n9011), .ZN(n8010) );
  XNOR2_X1 U9649 ( .A(n8025), .B(n8079), .ZN(n7988) );
  AND2_X1 U9650 ( .A1(n7988), .A2(n8891), .ZN(n7993) );
  OR2_X1 U9651 ( .A1(n8026), .A2(n7993), .ZN(n8011) );
  XNOR2_X1 U9652 ( .A(n8900), .B(n8219), .ZN(n7995) );
  XNOR2_X1 U9653 ( .A(n7995), .B(n8879), .ZN(n8015) );
  INV_X1 U9654 ( .A(n8015), .ZN(n7994) );
  OR2_X1 U9655 ( .A1(n8011), .A2(n7994), .ZN(n7985) );
  INV_X1 U9656 ( .A(n7985), .ZN(n7982) );
  AND2_X1 U9657 ( .A1(n7983), .A2(n7982), .ZN(n7986) );
  XNOR2_X1 U9658 ( .A(n7988), .B(n8891), .ZN(n8029) );
  INV_X1 U9659 ( .A(n8029), .ZN(n7992) );
  INV_X1 U9660 ( .A(n7989), .ZN(n7991) );
  NAND2_X1 U9661 ( .A1(n7991), .A2(n7990), .ZN(n8028) );
  AND2_X1 U9662 ( .A1(n7992), .A2(n8028), .ZN(n8031) );
  OR2_X1 U9663 ( .A1(n7993), .A2(n8031), .ZN(n8012) );
  OR2_X1 U9664 ( .A1(n7994), .A2(n8012), .ZN(n7999) );
  AND2_X1 U9665 ( .A1(n8001), .A2(n7999), .ZN(n8014) );
  INV_X1 U9666 ( .A(n8014), .ZN(n7997) );
  NAND2_X1 U9667 ( .A1(n7995), .A2(n8036), .ZN(n7998) );
  INV_X1 U9668 ( .A(n7998), .ZN(n7996) );
  XNOR2_X1 U9669 ( .A(n9011), .B(n8219), .ZN(n8050) );
  XNOR2_X1 U9670 ( .A(n8050), .B(n8890), .ZN(n8002) );
  NOR3_X1 U9671 ( .A1(n7997), .A2(n7996), .A3(n8002), .ZN(n8005) );
  AND2_X1 U9672 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  NAND2_X1 U9673 ( .A1(n8001), .A2(n8000), .ZN(n8003) );
  INV_X1 U9674 ( .A(n8052), .ZN(n8004) );
  OAI21_X1 U9675 ( .B1(n8005), .B2(n8004), .A(n8285), .ZN(n8009) );
  NAND2_X1 U9676 ( .A1(n8266), .A2(n8878), .ZN(n8006) );
  NAND2_X1 U9677 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8666) );
  OAI211_X1 U9678 ( .C1(n8036), .C2(n8268), .A(n8006), .B(n8666), .ZN(n8007)
         );
  AOI21_X1 U9679 ( .B1(n8293), .B2(n8883), .A(n8007), .ZN(n8008) );
  OAI211_X1 U9680 ( .C1(n8010), .C2(n8296), .A(n8009), .B(n8008), .ZN(P2_U3168) );
  INV_X1 U9681 ( .A(n8900), .ZN(n9017) );
  OR2_X1 U9682 ( .A1(n8027), .A2(n8011), .ZN(n8013) );
  NAND2_X1 U9683 ( .A1(n8013), .A2(n8012), .ZN(n8016) );
  OAI21_X1 U9684 ( .B1(n8016), .B2(n8015), .A(n8014), .ZN(n8017) );
  NAND2_X1 U9685 ( .A1(n8017), .A2(n8285), .ZN(n8021) );
  NAND2_X1 U9686 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8642) );
  OAI21_X1 U9687 ( .B1(n8290), .B2(n8863), .A(n8642), .ZN(n8019) );
  NOR2_X1 U9688 ( .A1(n8223), .A2(n8896), .ZN(n8018) );
  AOI211_X1 U9689 ( .C1(n8288), .C2(n8891), .A(n8019), .B(n8018), .ZN(n8020)
         );
  OAI211_X1 U9690 ( .C1(n9017), .C2(n8296), .A(n8021), .B(n8020), .ZN(P2_U3166) );
  OAI222_X1 U9691 ( .A1(n9729), .A2(n8024), .B1(n9732), .B2(n8023), .C1(n8022), 
        .C2(P1_U3086), .ZN(P1_U3329) );
  INV_X1 U9692 ( .A(n8025), .ZN(n8041) );
  OR2_X1 U9693 ( .A1(n8027), .A2(n8026), .ZN(n8032) );
  NAND2_X1 U9694 ( .A1(n8032), .A2(n8028), .ZN(n8030) );
  AOI21_X1 U9695 ( .B1(n8030), .B2(n8029), .A(n8272), .ZN(n8034) );
  NAND2_X1 U9696 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U9697 ( .A1(n8034), .A2(n8033), .ZN(n8040) );
  NAND2_X1 U9698 ( .A1(n8288), .A2(n8557), .ZN(n8035) );
  NAND2_X1 U9699 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8618) );
  OAI211_X1 U9700 ( .C1(n8036), .C2(n8290), .A(n8035), .B(n8618), .ZN(n8037)
         );
  AOI21_X1 U9701 ( .B1(n8293), .B2(n8038), .A(n8037), .ZN(n8039) );
  OAI211_X1 U9702 ( .C1(n8041), .C2(n8296), .A(n8040), .B(n8039), .ZN(P2_U3181) );
  AOI211_X1 U9703 ( .C1(n8044), .C2(n9801), .A(n8043), .B(n8042), .ZN(n8046)
         );
  MUX2_X1 U9704 ( .A(n10004), .B(n8046), .S(n9794), .Z(n8045) );
  OAI21_X1 U9705 ( .B1(n8049), .B2(n9717), .A(n8045), .ZN(P1_U3492) );
  INV_X1 U9706 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8047) );
  MUX2_X1 U9707 ( .A(n8047), .B(n8046), .S(n9818), .Z(n8048) );
  OAI21_X1 U9708 ( .B1(n8049), .B2(n9659), .A(n8048), .ZN(P1_U3535) );
  NAND2_X1 U9709 ( .A1(n8050), .A2(n8863), .ZN(n8051) );
  XNOR2_X1 U9710 ( .A(n8935), .B(n8219), .ZN(n8078) );
  XNOR2_X1 U9711 ( .A(n8078), .B(n8878), .ZN(n8076) );
  XOR2_X1 U9712 ( .A(n8077), .B(n8076), .Z(n8057) );
  NAND2_X1 U9713 ( .A1(n8293), .A2(n8867), .ZN(n8054) );
  AOI22_X1 U9714 ( .A1(n8266), .A2(n8824), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8053) );
  OAI211_X1 U9715 ( .C1(n8863), .C2(n8268), .A(n8054), .B(n8053), .ZN(n8055)
         );
  AOI21_X1 U9716 ( .B1(n8935), .B2(n8228), .A(n8055), .ZN(n8056) );
  OAI21_X1 U9717 ( .B1(n8057), .B2(n8272), .A(n8056), .ZN(P2_U3178) );
  AOI21_X1 U9718 ( .B1(n8058), .B2(n8065), .A(n9497), .ZN(n8062) );
  OR2_X1 U9719 ( .A1(n9137), .A2(n9235), .ZN(n8061) );
  NAND2_X1 U9720 ( .A1(n9260), .A2(n9237), .ZN(n8060) );
  NAND2_X1 U9721 ( .A1(n8061), .A2(n8060), .ZN(n9041) );
  AOI21_X1 U9722 ( .B1(n8062), .B2(n8059), .A(n9041), .ZN(n9655) );
  NOR2_X1 U9723 ( .A1(n9778), .A2(n8063), .ZN(n8068) );
  XNOR2_X1 U9724 ( .A(n8066), .B(n8065), .ZN(n9656) );
  INV_X1 U9725 ( .A(n9656), .ZN(n8067) );
  OAI21_X1 U9726 ( .B1(n9773), .B2(n8068), .A(n8067), .ZN(n8075) );
  OAI22_X1 U9727 ( .A1(n9568), .A2(n8069), .B1(n9043), .B2(n9754), .ZN(n8073)
         );
  OAI211_X1 U9728 ( .C1(n8071), .C2(n9718), .A(n8070), .B(n6447), .ZN(n9654)
         );
  NOR2_X1 U9729 ( .A1(n9654), .A2(n9760), .ZN(n8072) );
  AOI211_X1 U9730 ( .C1(n9769), .C2(n9045), .A(n8073), .B(n8072), .ZN(n8074)
         );
  OAI211_X1 U9731 ( .C1(n9778), .C2(n9655), .A(n8075), .B(n8074), .ZN(P1_U3279) );
  XNOR2_X1 U9732 ( .A(n5985), .B(n6803), .ZN(n8172) );
  XNOR2_X1 U9733 ( .A(n8172), .B(n8865), .ZN(n8080) );
  XNOR2_X1 U9734 ( .A(n8175), .B(n8080), .ZN(n8085) );
  NAND2_X1 U9735 ( .A1(n8288), .A2(n8878), .ZN(n8081) );
  NAND2_X1 U9736 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8723) );
  OAI211_X1 U9737 ( .C1(n8843), .C2(n8290), .A(n8081), .B(n8723), .ZN(n8082)
         );
  AOI21_X1 U9738 ( .B1(n8293), .B2(n8848), .A(n8082), .ZN(n8084) );
  NAND2_X1 U9739 ( .A1(n5985), .A2(n8228), .ZN(n8083) );
  OAI211_X1 U9740 ( .C1(n8085), .C2(n8272), .A(n8084), .B(n8083), .ZN(P2_U3159) );
  INV_X1 U9741 ( .A(n8086), .ZN(n8161) );
  OAI222_X1 U9742 ( .A1(n9031), .A2(n8087), .B1(n9034), .B2(n8161), .C1(
        P2_U3151), .C2(n6091), .ZN(P2_U3268) );
  INV_X1 U9743 ( .A(n8088), .ZN(n9731) );
  AOI21_X1 U9744 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8090), .A(n8089), .ZN(
        n8091) );
  OAI21_X1 U9745 ( .B1(n9731), .B2(n9034), .A(n8091), .ZN(P2_U3267) );
  INV_X1 U9746 ( .A(n8298), .ZN(n8093) );
  OAI222_X1 U9747 ( .A1(n9729), .A2(n10033), .B1(n9728), .B2(n8093), .C1(n8092), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U9748 ( .A1(n9025), .A2(n8299), .B1(n9034), .B2(n8093), .C1(
        P2_U3151), .C2(n5688), .ZN(P2_U3265) );
  NAND2_X1 U9749 ( .A1(n8096), .A2(n8101), .ZN(n8117) );
  OAI21_X1 U9750 ( .B1(n8096), .B2(n8101), .A(n8117), .ZN(n9387) );
  INV_X1 U9751 ( .A(n8099), .ZN(n8097) );
  NOR2_X1 U9752 ( .A1(n8101), .A2(n8097), .ZN(n8098) );
  NAND2_X1 U9753 ( .A1(n8100), .A2(n8098), .ZN(n8120) );
  NAND2_X1 U9754 ( .A1(n8100), .A2(n8099), .ZN(n8102) );
  OR2_X1 U9755 ( .A1(n8103), .A2(n9235), .ZN(n8104) );
  OAI21_X1 U9756 ( .B1(n8105), .B2(n9220), .A(n8104), .ZN(n9096) );
  OAI211_X1 U9757 ( .C1(n8108), .C2(n8107), .A(n8126), .B(n6447), .ZN(n9383)
         );
  NAND2_X1 U9758 ( .A1(n9378), .A2(n9383), .ZN(n8112) );
  OAI21_X1 U9759 ( .B1(n9387), .B2(n9653), .A(n8111), .ZN(P1_U3550) );
  OAI21_X1 U9760 ( .B1(n9387), .B2(n9711), .A(n8115), .ZN(P1_U3518) );
  INV_X1 U9761 ( .A(n9090), .ZN(n9247) );
  NAND2_X1 U9762 ( .A1(n9380), .A2(n9247), .ZN(n8116) );
  NAND2_X1 U9763 ( .A1(n8120), .A2(n8119), .ZN(n8122) );
  XNOR2_X1 U9764 ( .A(n8122), .B(n8121), .ZN(n8123) );
  AOI22_X1 U9765 ( .A1(n9247), .A2(n9237), .B1(n8124), .B2(n9246), .ZN(n8125)
         );
  AOI21_X1 U9766 ( .B1(n8126), .B2(n5463), .A(n9579), .ZN(n8128) );
  NAND2_X1 U9767 ( .A1(n8128), .A2(n8127), .ZN(n8134) );
  AOI22_X1 U9768 ( .A1(n8129), .A2(n9767), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9778), .ZN(n8131) );
  NAND2_X1 U9769 ( .A1(n5463), .A2(n9769), .ZN(n8130) );
  OAI211_X1 U9770 ( .C1(n8134), .C2(n9760), .A(n8131), .B(n8130), .ZN(n8132)
         );
  AOI21_X1 U9771 ( .B1(n8137), .B2(n9745), .A(n8132), .ZN(n8133) );
  OAI21_X1 U9772 ( .B1(n8143), .B2(n9589), .A(n8133), .ZN(P1_U3356) );
  INV_X1 U9773 ( .A(n5463), .ZN(n8135) );
  OAI21_X1 U9774 ( .B1(n8135), .B2(n9804), .A(n8134), .ZN(n8136) );
  OAI21_X1 U9775 ( .B1(n8143), .B2(n9653), .A(n8139), .ZN(P1_U3551) );
  INV_X1 U9776 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8141) );
  OAI21_X1 U9777 ( .B1(n8143), .B2(n9711), .A(n8142), .ZN(P1_U3519) );
  OAI222_X1 U9778 ( .A1(n9729), .A2(n8145), .B1(n9732), .B2(n8144), .C1(
        P1_U3086), .C2(n5620), .ZN(P1_U3336) );
  NAND2_X1 U9779 ( .A1(n8147), .A2(n8146), .ZN(n8335) );
  XNOR2_X1 U9780 ( .A(n8148), .B(n8335), .ZN(n8149) );
  AOI222_X1 U9781 ( .A1(n9829), .A2(n8149), .B1(n8562), .B2(n9824), .C1(n8563), 
        .C2(n9826), .ZN(n9860) );
  MUX2_X1 U9782 ( .A(n8150), .B(n9860), .S(n9837), .Z(n8154) );
  AOI22_X1 U9783 ( .A1(n8899), .A2(n8152), .B1(n8898), .B2(n8151), .ZN(n8153)
         );
  OAI211_X1 U9784 ( .C1(n8903), .C2(n9859), .A(n8154), .B(n8153), .ZN(P2_U3227) );
  INV_X1 U9785 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8156) );
  OAI211_X1 U9786 ( .C1(n8155), .C2(n9373), .A(n6447), .B(n4338), .ZN(n9377)
         );
  AND2_X1 U9787 ( .A1(n9377), .A2(n9367), .ZN(n8158) );
  MUX2_X1 U9788 ( .A(n8156), .B(n8158), .S(n9794), .Z(n8157) );
  OAI21_X1 U9789 ( .B1(n9373), .B2(n9717), .A(n8157), .ZN(P1_U3520) );
  MUX2_X1 U9790 ( .A(n8159), .B(n8158), .S(n9818), .Z(n8160) );
  OAI21_X1 U9791 ( .B1(n9373), .B2(n9659), .A(n8160), .ZN(P1_U3552) );
  OAI222_X1 U9792 ( .A1(n8162), .A2(n9729), .B1(P1_U3086), .B2(n5673), .C1(
        n9728), .C2(n8161), .ZN(P1_U3328) );
  INV_X1 U9793 ( .A(n6543), .ZN(n8169) );
  NAND2_X1 U9794 ( .A1(n8164), .A2(n8898), .ZN(n8734) );
  OAI21_X1 U9795 ( .B1(n8894), .B2(n8165), .A(n8734), .ZN(n8166) );
  INV_X1 U9796 ( .A(n8166), .ZN(n8168) );
  INV_X1 U9797 ( .A(n8170), .ZN(n8171) );
  OAI21_X1 U9798 ( .B1(n8163), .B2(n9839), .A(n8171), .ZN(P2_U3204) );
  INV_X1 U9799 ( .A(n8172), .ZN(n8173) );
  NAND2_X1 U9800 ( .A1(n8173), .A2(n8824), .ZN(n8174) );
  OAI21_X1 U9801 ( .B1(n8175), .B2(n4842), .A(n8174), .ZN(n8176) );
  INV_X1 U9802 ( .A(n8176), .ZN(n8263) );
  XNOR2_X1 U9803 ( .A(n8830), .B(n6803), .ZN(n8177) );
  NAND2_X1 U9804 ( .A1(n8177), .A2(n8843), .ZN(n8231) );
  INV_X1 U9805 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U9806 ( .A1(n8178), .A2(n8806), .ZN(n8179) );
  AND2_X1 U9807 ( .A1(n8231), .A2(n8179), .ZN(n8264) );
  NAND2_X1 U9808 ( .A1(n8263), .A2(n8264), .ZN(n8230) );
  NAND2_X1 U9809 ( .A1(n8230), .A2(n8231), .ZN(n8180) );
  XNOR2_X1 U9810 ( .A(n8991), .B(n6803), .ZN(n8181) );
  XNOR2_X1 U9811 ( .A(n8181), .B(n8825), .ZN(n8232) );
  NAND2_X1 U9812 ( .A1(n8181), .A2(n8796), .ZN(n8182) );
  XNOR2_X1 U9813 ( .A(n8923), .B(n6803), .ZN(n8184) );
  XNOR2_X1 U9814 ( .A(n8184), .B(n8238), .ZN(n8273) );
  INV_X1 U9815 ( .A(n8273), .ZN(n8183) );
  INV_X1 U9816 ( .A(n8184), .ZN(n8185) );
  NAND2_X1 U9817 ( .A1(n8185), .A2(n8807), .ZN(n8186) );
  AND2_X2 U9818 ( .A1(n8275), .A2(n8186), .ZN(n8188) );
  XNOR2_X1 U9819 ( .A(n8981), .B(n6803), .ZN(n8187) );
  INV_X1 U9820 ( .A(n8189), .ZN(n8255) );
  XNOR2_X1 U9821 ( .A(n8975), .B(n8219), .ZN(n8190) );
  NAND2_X1 U9822 ( .A1(n8190), .A2(n8760), .ZN(n8247) );
  INV_X1 U9823 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U9824 ( .A1(n8191), .A2(n8785), .ZN(n8192) );
  AND2_X1 U9825 ( .A1(n8247), .A2(n8192), .ZN(n8254) );
  XNOR2_X1 U9826 ( .A(n8244), .B(n8219), .ZN(n8194) );
  NAND2_X1 U9827 ( .A1(n8194), .A2(n8193), .ZN(n8197) );
  INV_X1 U9828 ( .A(n8194), .ZN(n8195) );
  NAND2_X1 U9829 ( .A1(n8195), .A2(n8774), .ZN(n8196) );
  NAND2_X1 U9830 ( .A1(n8197), .A2(n8196), .ZN(n8246) );
  INV_X1 U9831 ( .A(n8197), .ZN(n8284) );
  XNOR2_X1 U9832 ( .A(n8964), .B(n6803), .ZN(n8198) );
  XNOR2_X1 U9833 ( .A(n8198), .B(n8743), .ZN(n8283) );
  NAND2_X1 U9834 ( .A1(n8198), .A2(n8199), .ZN(n8200) );
  NAND2_X1 U9835 ( .A1(n8282), .A2(n8200), .ZN(n8202) );
  XNOR2_X1 U9836 ( .A(n8958), .B(n6803), .ZN(n8217) );
  XOR2_X1 U9837 ( .A(n8751), .B(n8217), .Z(n8201) );
  AOI21_X1 U9838 ( .B1(n8202), .B2(n8201), .A(n8272), .ZN(n8209) );
  AOI22_X1 U9839 ( .A1(n8743), .A2(n8288), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8204) );
  NAND2_X1 U9840 ( .A1(n8746), .A2(n8293), .ZN(n8203) );
  OAI211_X1 U9841 ( .C1(n8524), .C2(n8290), .A(n8204), .B(n8203), .ZN(n8205)
         );
  INV_X1 U9842 ( .A(n8205), .ZN(n8206) );
  INV_X1 U9843 ( .A(n8210), .ZN(P2_U3154) );
  AOI21_X1 U9844 ( .B1(n8773), .B2(n8211), .A(n8256), .ZN(n8216) );
  AOI22_X1 U9845 ( .A1(n8785), .A2(n8266), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8213) );
  NAND2_X1 U9846 ( .A1(n8293), .A2(n8788), .ZN(n8212) );
  OAI211_X1 U9847 ( .C1(n8238), .C2(n8268), .A(n8213), .B(n8212), .ZN(n8214)
         );
  AOI21_X1 U9848 ( .B1(n8981), .B2(n8228), .A(n8214), .ZN(n8215) );
  OAI21_X1 U9849 ( .B1(n8216), .B2(n8272), .A(n8215), .ZN(P2_U3156) );
  INV_X1 U9850 ( .A(n8217), .ZN(n8218) );
  XNOR2_X1 U9851 ( .A(n8326), .B(n8219), .ZN(n8220) );
  INV_X1 U9852 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8221) );
  OAI22_X1 U9853 ( .A1(n8291), .A2(n8268), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8221), .ZN(n8227) );
  INV_X1 U9854 ( .A(n8222), .ZN(n8224) );
  OAI22_X1 U9855 ( .A1(n8225), .A2(n8290), .B1(n8224), .B2(n8223), .ZN(n8226)
         );
  AOI211_X1 U9856 ( .C1(n8533), .C2(n8228), .A(n8227), .B(n8226), .ZN(n8229)
         );
  INV_X1 U9857 ( .A(n8230), .ZN(n8234) );
  INV_X1 U9858 ( .A(n8231), .ZN(n8233) );
  NOR3_X1 U9859 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(n8237) );
  INV_X1 U9860 ( .A(n8235), .ZN(n8236) );
  OAI21_X1 U9861 ( .B1(n8237), .B2(n8236), .A(n8285), .ZN(n8242) );
  NOR2_X1 U9862 ( .A1(n8843), .A2(n8268), .ZN(n8240) );
  OAI22_X1 U9863 ( .A1(n8238), .A2(n8290), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10034), .ZN(n8239) );
  AOI211_X1 U9864 ( .C1(n8810), .C2(n8293), .A(n8240), .B(n8239), .ZN(n8241)
         );
  OAI211_X1 U9865 ( .C1(n8243), .C2(n8296), .A(n8242), .B(n8241), .ZN(P2_U3163) );
  AND3_X1 U9866 ( .A1(n8253), .A2(n8247), .A3(n8246), .ZN(n8248) );
  OAI21_X1 U9867 ( .B1(n8245), .B2(n8248), .A(n8285), .ZN(n8252) );
  AOI22_X1 U9868 ( .A1(n8785), .A2(n8288), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8249) );
  OAI21_X1 U9869 ( .B1(n8199), .B2(n8290), .A(n8249), .ZN(n8250) );
  AOI21_X1 U9870 ( .B1(n8761), .B2(n8293), .A(n8250), .ZN(n8251) );
  OAI211_X1 U9871 ( .C1(n8969), .C2(n8296), .A(n8252), .B(n8251), .ZN(P2_U3165) );
  INV_X1 U9872 ( .A(n8253), .ZN(n8258) );
  NOR3_X1 U9873 ( .A1(n8256), .A2(n8255), .A3(n8254), .ZN(n8257) );
  OAI21_X1 U9874 ( .B1(n8258), .B2(n8257), .A(n8285), .ZN(n8262) );
  AOI22_X1 U9875 ( .A1(n8774), .A2(n8266), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8259) );
  OAI21_X1 U9876 ( .B1(n8795), .B2(n8268), .A(n8259), .ZN(n8260) );
  AOI21_X1 U9877 ( .B1(n8776), .B2(n8293), .A(n8260), .ZN(n8261) );
  OAI211_X1 U9878 ( .C1(n8778), .C2(n8296), .A(n8262), .B(n8261), .ZN(P2_U3169) );
  INV_X1 U9879 ( .A(n8830), .ZN(n8996) );
  OAI21_X1 U9880 ( .B1(n8264), .B2(n8263), .A(n8230), .ZN(n8265) );
  NAND2_X1 U9881 ( .A1(n8265), .A2(n8285), .ZN(n8271) );
  AOI22_X1 U9882 ( .A1(n8825), .A2(n8266), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8267) );
  OAI21_X1 U9883 ( .B1(n8865), .B2(n8268), .A(n8267), .ZN(n8269) );
  AOI21_X1 U9884 ( .B1(n8829), .B2(n8293), .A(n8269), .ZN(n8270) );
  OAI211_X1 U9885 ( .C1(n8996), .C2(n8296), .A(n8271), .B(n8270), .ZN(P2_U3173) );
  INV_X1 U9886 ( .A(n8923), .ZN(n8281) );
  AOI21_X1 U9887 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8276) );
  NAND2_X1 U9888 ( .A1(n8276), .A2(n8275), .ZN(n8280) );
  AOI22_X1 U9889 ( .A1(n8825), .A2(n8288), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8277) );
  OAI21_X1 U9890 ( .B1(n8795), .B2(n8290), .A(n8277), .ZN(n8278) );
  AOI21_X1 U9891 ( .B1(n8797), .B2(n8293), .A(n8278), .ZN(n8279) );
  OAI211_X1 U9892 ( .C1(n8281), .C2(n8296), .A(n8280), .B(n8279), .ZN(P2_U3175) );
  INV_X1 U9893 ( .A(n8282), .ZN(n8287) );
  NOR3_X1 U9894 ( .A1(n8245), .A2(n8284), .A3(n8283), .ZN(n8286) );
  OAI21_X1 U9895 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8295) );
  AOI22_X1 U9896 ( .A1(n8774), .A2(n8288), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8289) );
  OAI21_X1 U9897 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n8292) );
  AOI21_X1 U9898 ( .B1(n8753), .B2(n8293), .A(n8292), .ZN(n8294) );
  OAI211_X1 U9899 ( .C1(n8297), .C2(n8296), .A(n8295), .B(n8294), .ZN(P2_U3180) );
  INV_X1 U9900 ( .A(n8355), .ZN(n8315) );
  OR2_X1 U9901 ( .A1(n4313), .A2(n8299), .ZN(n8300) );
  INV_X1 U9902 ( .A(n8556), .ZN(n8317) );
  NAND2_X1 U9903 ( .A1(n8318), .A2(n8317), .ZN(n8537) );
  NAND2_X1 U9904 ( .A1(n9022), .A2(n8303), .ZN(n8305) );
  OR2_X1 U9905 ( .A1(n4288), .A2(n9026), .ZN(n8304) );
  INV_X1 U9906 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U9907 ( .A1(n5738), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8308) );
  INV_X1 U9908 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8306) );
  OR2_X1 U9909 ( .A1(n4315), .A2(n8306), .ZN(n8307) );
  OAI211_X1 U9910 ( .C1(n8310), .C2(n4306), .A(n8308), .B(n8307), .ZN(n8311)
         );
  INV_X1 U9911 ( .A(n8311), .ZN(n8312) );
  NOR2_X1 U9912 ( .A1(n8319), .A2(n8555), .ZN(n8358) );
  OAI211_X1 U9913 ( .C1(n8316), .C2(n8315), .A(n8525), .B(n8314), .ZN(n8325)
         );
  INV_X1 U9914 ( .A(n8356), .ZN(n8321) );
  AOI211_X1 U9915 ( .C1(n8321), .C2(n8319), .A(n8320), .B(n8542), .ZN(n8324)
         );
  NOR3_X1 U9916 ( .A1(n8319), .A2(n8322), .A3(n8555), .ZN(n8323) );
  AOI21_X1 U9917 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8359) );
  INV_X1 U9918 ( .A(n8326), .ZN(n8354) );
  INV_X1 U9919 ( .A(n8327), .ZN(n8360) );
  INV_X1 U9920 ( .A(n8750), .ZN(n8353) );
  NAND2_X1 U9921 ( .A1(n8767), .A2(n8768), .ZN(n8783) );
  INV_X1 U9922 ( .A(n8329), .ZN(n8330) );
  NAND2_X1 U9923 ( .A1(n8331), .A2(n8330), .ZN(n8334) );
  NOR4_X1 U9924 ( .A1(n7054), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n8336)
         );
  NAND4_X1 U9925 ( .A1(n8328), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n8341)
         );
  OR4_X1 U9926 ( .A1(n8341), .A2(n8340), .A3(n8339), .A4(n8338), .ZN(n8345) );
  NOR4_X1 U9927 ( .A1(n8345), .A2(n8344), .A3(n8343), .A4(n8342), .ZN(n8347)
         );
  NAND4_X1 U9928 ( .A1(n8463), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n8349)
         );
  NOR4_X1 U9929 ( .A1(n8853), .A2(n8875), .A3(n8889), .A4(n8349), .ZN(n8350)
         );
  NAND3_X1 U9930 ( .A1(n8819), .A2(n8350), .A3(n8837), .ZN(n8351) );
  NOR4_X1 U9931 ( .A1(n4609), .A2(n8783), .A3(n8804), .A4(n8351), .ZN(n8352)
         );
  NAND4_X1 U9932 ( .A1(n8525), .A2(n8354), .A3(n8353), .A4(n4825), .ZN(n8357)
         );
  MUX2_X1 U9933 ( .A(n8361), .B(n8360), .S(n8522), .Z(n8363) );
  INV_X1 U9934 ( .A(n8740), .ZN(n8362) );
  NOR2_X1 U9935 ( .A1(n8363), .A2(n8362), .ZN(n8520) );
  MUX2_X1 U9936 ( .A(n8365), .B(n8364), .S(n8522), .Z(n8508) );
  NAND2_X1 U9937 ( .A1(n5985), .A2(n8865), .ZN(n8481) );
  AND2_X1 U9938 ( .A1(n8488), .A2(n8481), .ZN(n8483) );
  INV_X1 U9939 ( .A(n8371), .ZN(n8367) );
  NAND2_X1 U9940 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  AND2_X1 U9941 ( .A1(n8366), .A2(n8369), .ZN(n8375) );
  AND2_X1 U9942 ( .A1(n8371), .A2(n8370), .ZN(n8372) );
  OAI21_X1 U9943 ( .B1(n8373), .B2(n8372), .A(n8366), .ZN(n8374) );
  MUX2_X1 U9944 ( .A(n8375), .B(n8374), .S(n8522), .Z(n8385) );
  OR2_X1 U9945 ( .A1(n8376), .A2(n6835), .ZN(n8388) );
  OAI21_X1 U9946 ( .B1(n8378), .B2(n8377), .A(n8388), .ZN(n8382) );
  NAND2_X1 U9947 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  MUX2_X1 U9948 ( .A(n8382), .B(n8381), .S(n8522), .Z(n8383) );
  INV_X1 U9949 ( .A(n8383), .ZN(n8384) );
  OAI21_X1 U9950 ( .B1(n8385), .B2(n9827), .A(n8384), .ZN(n8387) );
  NAND2_X1 U9951 ( .A1(n8387), .A2(n8386), .ZN(n8398) );
  INV_X1 U9952 ( .A(n8388), .ZN(n8390) );
  OAI211_X1 U9953 ( .C1(n8398), .C2(n8390), .A(n8399), .B(n8389), .ZN(n8394)
         );
  INV_X1 U9954 ( .A(n8395), .ZN(n8391) );
  NOR2_X1 U9955 ( .A1(n8401), .A2(n8391), .ZN(n8393) );
  INV_X1 U9956 ( .A(n8400), .ZN(n8392) );
  AOI21_X1 U9957 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8405) );
  OAI211_X1 U9958 ( .C1(n8398), .C2(n8397), .A(n8396), .B(n8395), .ZN(n8403)
         );
  AND2_X1 U9959 ( .A1(n8400), .A2(n8399), .ZN(n8402) );
  AOI21_X1 U9960 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8404) );
  MUX2_X1 U9961 ( .A(n8405), .B(n8404), .S(n8536), .Z(n8413) );
  AND2_X1 U9962 ( .A1(n8440), .A2(n8435), .ZN(n8430) );
  NAND2_X1 U9963 ( .A1(n8406), .A2(n8420), .ZN(n8409) );
  NAND2_X1 U9964 ( .A1(n8407), .A2(n8415), .ZN(n8408) );
  MUX2_X1 U9965 ( .A(n8409), .B(n8408), .S(n8536), .Z(n8423) );
  NAND2_X1 U9966 ( .A1(n8432), .A2(n8410), .ZN(n8411) );
  NOR2_X1 U9967 ( .A1(n8423), .A2(n8411), .ZN(n8412) );
  OR2_X1 U9968 ( .A1(n8434), .A2(n8522), .ZN(n8437) );
  NAND4_X1 U9969 ( .A1(n8413), .A2(n8430), .A3(n8412), .A4(n8437), .ZN(n8445)
         );
  INV_X1 U9970 ( .A(n8430), .ZN(n8417) );
  AND2_X1 U9971 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  OR3_X1 U9972 ( .A1(n8417), .A2(n8536), .A3(n8416), .ZN(n8425) );
  NAND2_X1 U9973 ( .A1(n8419), .A2(n8418), .ZN(n8421) );
  AOI21_X1 U9974 ( .B1(n8421), .B2(n8420), .A(n8522), .ZN(n8422) );
  NAND3_X1 U9975 ( .A1(n8434), .A2(n8422), .A3(n8432), .ZN(n8424) );
  AOI21_X1 U9976 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8442) );
  OR2_X1 U9977 ( .A1(n8426), .A2(n8536), .ZN(n8428) );
  NAND2_X1 U9978 ( .A1(n8560), .A2(n8522), .ZN(n8427) );
  OAI22_X1 U9979 ( .A1(n9884), .A2(n8428), .B1(n9878), .B2(n8427), .ZN(n8429)
         );
  NAND2_X1 U9980 ( .A1(n8430), .A2(n8429), .ZN(n8439) );
  NAND4_X1 U9981 ( .A1(n8432), .A2(n8431), .A3(n8536), .A4(n9878), .ZN(n8433)
         );
  OAI211_X1 U9982 ( .C1(n8522), .C2(n8435), .A(n8434), .B(n8433), .ZN(n8436)
         );
  NAND2_X1 U9983 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  OAI211_X1 U9984 ( .C1(n8440), .C2(n8522), .A(n8439), .B(n8438), .ZN(n8441)
         );
  NOR2_X1 U9985 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  NAND3_X1 U9986 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8449) );
  MUX2_X1 U9987 ( .A(n8447), .B(n8446), .S(n8536), .Z(n8448) );
  NAND2_X1 U9988 ( .A1(n8449), .A2(n8448), .ZN(n8454) );
  MUX2_X1 U9989 ( .A(n8558), .B(n8451), .S(n8536), .Z(n8452) );
  INV_X1 U9990 ( .A(n8452), .ZN(n8453) );
  OAI21_X1 U9991 ( .B1(n8454), .B2(n4632), .A(n8453), .ZN(n8457) );
  NAND2_X1 U9992 ( .A1(n8454), .A2(n4357), .ZN(n8456) );
  AOI21_X1 U9993 ( .B1(n8457), .B2(n8456), .A(n8455), .ZN(n8462) );
  INV_X1 U9994 ( .A(n8458), .ZN(n8459) );
  MUX2_X1 U9995 ( .A(n8460), .B(n8459), .S(n8536), .Z(n8461) );
  OR2_X1 U9996 ( .A1(n8462), .A2(n8461), .ZN(n8464) );
  NAND2_X1 U9997 ( .A1(n8464), .A2(n8463), .ZN(n8468) );
  NAND3_X1 U9998 ( .A1(n8468), .A2(n8469), .A3(n8465), .ZN(n8466) );
  AOI21_X1 U9999 ( .B1(n8466), .B2(n8471), .A(n8875), .ZN(n8474) );
  NAND2_X1 U10000 ( .A1(n8468), .A2(n8467), .ZN(n8470) );
  NAND2_X1 U10001 ( .A1(n8470), .A2(n8469), .ZN(n8472) );
  NAND2_X1 U10002 ( .A1(n8475), .A2(n8852), .ZN(n8476) );
  NAND2_X1 U10003 ( .A1(n8476), .A2(n8536), .ZN(n8477) );
  NAND2_X1 U10004 ( .A1(n8478), .A2(n8477), .ZN(n8485) );
  NAND2_X1 U10005 ( .A1(n8819), .A2(n8479), .ZN(n8480) );
  AOI21_X1 U10006 ( .B1(n8485), .B2(n8481), .A(n8480), .ZN(n8482) );
  MUX2_X1 U10007 ( .A(n8483), .B(n8482), .S(n8522), .Z(n8487) );
  NAND3_X1 U10008 ( .A1(n8485), .A2(n8484), .A3(n8837), .ZN(n8486) );
  NAND2_X1 U10009 ( .A1(n8487), .A2(n8486), .ZN(n8491) );
  NAND2_X1 U10010 ( .A1(n8498), .A2(n8488), .ZN(n8489) );
  NAND2_X1 U10011 ( .A1(n8489), .A2(n8522), .ZN(n8490) );
  NAND2_X1 U10012 ( .A1(n8491), .A2(n8490), .ZN(n8495) );
  INV_X1 U10013 ( .A(n8493), .ZN(n8494) );
  NAND2_X1 U10014 ( .A1(n8495), .A2(n4615), .ZN(n8501) );
  NAND2_X1 U10015 ( .A1(n8497), .A2(n8496), .ZN(n8499) );
  NAND3_X1 U10016 ( .A1(n8499), .A2(n8536), .A3(n8498), .ZN(n8500) );
  AOI21_X1 U10017 ( .B1(n8501), .B2(n8500), .A(n4609), .ZN(n8506) );
  AND2_X1 U10018 ( .A1(n8502), .A2(n8767), .ZN(n8504) );
  MUX2_X1 U10019 ( .A(n8504), .B(n8503), .S(n8536), .Z(n8505) );
  NAND2_X1 U10020 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  NAND2_X1 U10021 ( .A1(n8509), .A2(n8758), .ZN(n8514) );
  MUX2_X1 U10022 ( .A(n8511), .B(n8510), .S(n8536), .Z(n8512) );
  NAND2_X1 U10023 ( .A1(n8514), .A2(n8513), .ZN(n8519) );
  MUX2_X1 U10024 ( .A(n8516), .B(n8515), .S(n8536), .Z(n8517) );
  INV_X1 U10025 ( .A(n8517), .ZN(n8518) );
  AOI21_X1 U10026 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8521) );
  MUX2_X1 U10027 ( .A(n8524), .B(n8523), .S(n8522), .Z(n8531) );
  INV_X1 U10028 ( .A(n8525), .ZN(n8526) );
  OR2_X1 U10029 ( .A1(n8532), .A2(n8531), .ZN(n8535) );
  MUX2_X1 U10030 ( .A(n8742), .B(n8533), .S(n8536), .Z(n8534) );
  INV_X1 U10031 ( .A(n8542), .ZN(n8540) );
  NAND2_X1 U10032 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  NAND4_X1 U10033 ( .A1(n8540), .A2(n8539), .A3(n8356), .A4(n8538), .ZN(n8541)
         );
  INV_X1 U10034 ( .A(n8543), .ZN(n8544) );
  NAND4_X1 U10035 ( .A1(n4848), .A2(n8540), .A3(n8544), .A4(n8550), .ZN(n8545)
         );
  NAND3_X1 U10036 ( .A1(n4823), .A2(n8546), .A3(n8545), .ZN(n8548) );
  XNOR2_X1 U10037 ( .A(n8548), .B(n8547), .ZN(n8554) );
  NOR3_X1 U10038 ( .A1(n8549), .A2(n8715), .A3(n6090), .ZN(n8552) );
  OAI21_X1 U10039 ( .B1(n8553), .B2(n8550), .A(P2_B_REG_SCAN_IN), .ZN(n8551)
         );
  OAI22_X1 U10040 ( .A1(n8554), .A2(n8553), .B1(n8552), .B2(n8551), .ZN(
        P2_U3296) );
  INV_X1 U10041 ( .A(n8555), .ZN(n8733) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8733), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8556), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8742), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8751), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10046 ( .A(n8743), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8697), .Z(
        P2_U3517) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8774), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8785), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10049 ( .A(n8773), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8697), .Z(
        P2_U3514) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8807), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10051 ( .A(n8825), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8697), .Z(
        P2_U3512) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8806), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8824), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8878), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8890), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10056 ( .A(n8879), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8697), .Z(
        P2_U3507) );
  MUX2_X1 U10057 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8891), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8557), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10059 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8558), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10060 ( .A(n8559), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8697), .Z(
        P2_U3503) );
  MUX2_X1 U10061 ( .A(n8560), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8697), .Z(
        P2_U3500) );
  MUX2_X1 U10062 ( .A(n8561), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8697), .Z(
        P2_U3499) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8562), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10064 ( .A(n8563), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8697), .Z(
        P2_U3496) );
  MUX2_X1 U10065 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8564), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10066 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9825), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10067 ( .A(n8565), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8697), .Z(
        P2_U3493) );
  MUX2_X1 U10068 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5704), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10069 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8566), .S(P2_U3893), .Z(
        P2_U3491) );
  OAI211_X1 U10070 ( .C1(n8569), .C2(n8568), .A(n8567), .B(n8664), .ZN(n8583)
         );
  INV_X1 U10071 ( .A(n8731), .ZN(n8574) );
  OAI21_X1 U10072 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8573) );
  AOI22_X1 U10073 ( .A1(n8574), .A2(n8573), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n8582) );
  OAI21_X1 U10074 ( .B1(n8577), .B2(n8576), .A(n8575), .ZN(n8578) );
  AOI22_X1 U10075 ( .A1(n8721), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8727), .B2(
        n8578), .ZN(n8581) );
  NAND2_X1 U10076 ( .A1(n8676), .A2(n8579), .ZN(n8580) );
  NAND4_X1 U10077 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(
        P2_U3184) );
  NOR2_X1 U10078 ( .A1(n8598), .A2(n8584), .ZN(n8586) );
  NAND2_X1 U10079 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8622), .ZN(n8587) );
  OAI21_X1 U10080 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8622), .A(n8587), .ZN(
        n8588) );
  AOI21_X1 U10081 ( .B1(n4400), .B2(n8588), .A(n8610), .ZN(n8609) );
  INV_X1 U10082 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8597) );
  MUX2_X1 U10083 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6091), .Z(n8612) );
  XNOR2_X1 U10084 ( .A(n8612), .B(n8607), .ZN(n8593) );
  OR2_X1 U10085 ( .A1(n8589), .A2(n7955), .ZN(n8591) );
  NAND2_X1 U10086 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  NAND2_X1 U10087 ( .A1(n8593), .A2(n8592), .ZN(n8613) );
  OAI21_X1 U10088 ( .B1(n8593), .B2(n8592), .A(n8613), .ZN(n8594) );
  NAND2_X1 U10089 ( .A1(n8594), .A2(n8664), .ZN(n8596) );
  OAI211_X1 U10090 ( .C1(n8704), .C2(n8597), .A(n8596), .B(n8595), .ZN(n8606)
         );
  NOR2_X1 U10091 ( .A1(n8598), .A2(n4373), .ZN(n8600) );
  NAND2_X1 U10092 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8622), .ZN(n8601) );
  OAI21_X1 U10093 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8622), .A(n8601), .ZN(
        n8602) );
  NOR2_X1 U10094 ( .A1(n8603), .A2(n8602), .ZN(n8621) );
  AOI21_X1 U10095 ( .B1(n8603), .B2(n8602), .A(n8621), .ZN(n8604) );
  NOR2_X1 U10096 ( .A1(n8604), .A2(n8689), .ZN(n8605) );
  AOI211_X1 U10097 ( .C1(n8676), .C2(n8607), .A(n8606), .B(n8605), .ZN(n8608)
         );
  OAI21_X1 U10098 ( .B1(n8609), .B2(n8731), .A(n8608), .ZN(P2_U3196) );
  AOI21_X1 U10099 ( .B1(n8611), .B2(n7971), .A(n8631), .ZN(n8629) );
  INV_X1 U10100 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8620) );
  MUX2_X1 U10101 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6091), .Z(n8635) );
  XNOR2_X1 U10102 ( .A(n8635), .B(n8646), .ZN(n8616) );
  OR2_X1 U10103 ( .A1(n8612), .A2(n8622), .ZN(n8614) );
  NAND2_X1 U10104 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U10105 ( .A1(n8616), .A2(n8615), .ZN(n8637) );
  OAI21_X1 U10106 ( .B1(n8616), .B2(n8615), .A(n8637), .ZN(n8617) );
  NAND2_X1 U10107 ( .A1(n8617), .A2(n8664), .ZN(n8619) );
  OAI211_X1 U10108 ( .C1(n8620), .C2(n8704), .A(n8619), .B(n8618), .ZN(n8627)
         );
  AOI21_X1 U10109 ( .B1(n8624), .B2(n8623), .A(n8648), .ZN(n8625) );
  NOR2_X1 U10110 ( .A1(n8625), .A2(n8689), .ZN(n8626) );
  AOI211_X1 U10111 ( .C1(n8676), .C2(n8646), .A(n8627), .B(n8626), .ZN(n8628)
         );
  OAI21_X1 U10112 ( .B1(n8629), .B2(n8731), .A(n8628), .ZN(P2_U3197) );
  NOR2_X1 U10113 ( .A1(n8646), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U10114 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8670), .ZN(n8633) );
  OAI21_X1 U10115 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8670), .A(n8633), .ZN(
        n8634) );
  AOI21_X1 U10116 ( .B1(n4361), .B2(n8634), .A(n8657), .ZN(n8656) );
  INV_X1 U10117 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8644) );
  MUX2_X1 U10118 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6091), .Z(n8659) );
  XNOR2_X1 U10119 ( .A(n8659), .B(n8654), .ZN(n8640) );
  INV_X1 U10120 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U10121 ( .A1(n8646), .A2(n8636), .ZN(n8638) );
  NAND2_X1 U10122 ( .A1(n8638), .A2(n8637), .ZN(n8639) );
  NAND2_X1 U10123 ( .A1(n8640), .A2(n8639), .ZN(n8660) );
  OAI21_X1 U10124 ( .B1(n8640), .B2(n8639), .A(n8660), .ZN(n8641) );
  NAND2_X1 U10125 ( .A1(n8641), .A2(n8664), .ZN(n8643) );
  OAI211_X1 U10126 ( .C1(n8704), .C2(n8644), .A(n8643), .B(n8642), .ZN(n8653)
         );
  NOR2_X1 U10127 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  AOI22_X1 U10128 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8654), .B1(n8670), .B2(
        n8649), .ZN(n8650) );
  AOI21_X1 U10129 ( .B1(n4362), .B2(n8650), .A(n8669), .ZN(n8651) );
  NOR2_X1 U10130 ( .A1(n8651), .A2(n8689), .ZN(n8652) );
  AOI211_X1 U10131 ( .C1(n8676), .C2(n8654), .A(n8653), .B(n8652), .ZN(n8655)
         );
  OAI21_X1 U10132 ( .B1(n8656), .B2(n8731), .A(n8655), .ZN(P2_U3198) );
  XOR2_X1 U10133 ( .A(n8679), .B(n8671), .Z(n8658) );
  NOR2_X1 U10134 ( .A1(n8882), .A2(n8658), .ZN(n8680) );
  AOI21_X1 U10135 ( .B1(n8882), .B2(n8658), .A(n8680), .ZN(n8678) );
  INV_X1 U10136 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8668) );
  MUX2_X1 U10137 ( .A(n8882), .B(n8938), .S(n6091), .Z(n8693) );
  XNOR2_X1 U10138 ( .A(n8693), .B(n8671), .ZN(n8663) );
  OR2_X1 U10139 ( .A1(n8659), .A2(n8670), .ZN(n8661) );
  NAND2_X1 U10140 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  NAND2_X1 U10141 ( .A1(n8663), .A2(n8662), .ZN(n8691) );
  OAI21_X1 U10142 ( .B1(n8663), .B2(n8662), .A(n8691), .ZN(n8665) );
  NAND2_X1 U10143 ( .A1(n8665), .A2(n8664), .ZN(n8667) );
  OAI211_X1 U10144 ( .C1(n8704), .C2(n8668), .A(n8667), .B(n8666), .ZN(n8675)
         );
  XNOR2_X1 U10145 ( .A(n8684), .B(n8692), .ZN(n8672) );
  AOI21_X1 U10146 ( .B1(n8938), .B2(n8672), .A(n8685), .ZN(n8673) );
  NOR2_X1 U10147 ( .A1(n8673), .A2(n8689), .ZN(n8674) );
  OAI21_X1 U10148 ( .B1(n8678), .B2(n8731), .A(n8677), .ZN(P2_U3199) );
  NOR2_X1 U10149 ( .A1(n8692), .A2(n8679), .ZN(n8681) );
  NAND2_X1 U10150 ( .A1(n8700), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8707) );
  OAI21_X1 U10151 ( .B1(n8700), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8707), .ZN(
        n8682) );
  NOR2_X1 U10152 ( .A1(n8683), .A2(n8682), .ZN(n8709) );
  AOI21_X1 U10153 ( .B1(n8683), .B2(n8682), .A(n8709), .ZN(n8706) );
  NOR2_X1 U10154 ( .A1(n8692), .A2(n8684), .ZN(n8686) );
  NAND2_X1 U10155 ( .A1(n8700), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8711) );
  OAI21_X1 U10156 ( .B1(n8700), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8711), .ZN(
        n8687) );
  NAND2_X1 U10157 ( .A1(n8688), .A2(n8687), .ZN(n8690) );
  MUX2_X1 U10158 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6091), .Z(n8694) );
  NOR2_X1 U10159 ( .A1(n8695), .A2(n8694), .ZN(n8714) );
  NOR2_X1 U10160 ( .A1(n8714), .A2(n8696), .ZN(n8699) );
  INV_X1 U10161 ( .A(n8699), .ZN(n8698) );
  NOR2_X1 U10162 ( .A1(n8699), .A2(n8719), .ZN(n8701) );
  INV_X1 U10163 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8702) );
  INV_X1 U10164 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8703) );
  INV_X1 U10165 ( .A(n8707), .ZN(n8708) );
  NOR2_X1 U10166 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  MUX2_X1 U10167 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8847), .S(n4316), .Z(n8716) );
  XNOR2_X1 U10168 ( .A(n8710), .B(n8716), .ZN(n8730) );
  OAI21_X1 U10169 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8718) );
  MUX2_X1 U10170 ( .A(n4410), .B(n8716), .S(n8715), .Z(n8717) );
  XNOR2_X1 U10171 ( .A(n8718), .B(n8717), .ZN(n8720) );
  NOR2_X1 U10172 ( .A1(n8720), .A2(n8719), .ZN(n8726) );
  NAND2_X1 U10173 ( .A1(n8721), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U10174 ( .C1(n8724), .C2(n4316), .A(n8723), .B(n8722), .ZN(n8725)
         );
  OAI21_X1 U10175 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(P2_U3201) );
  NAND2_X1 U10176 ( .A1(n8733), .A2(n8732), .ZN(n8951) );
  OAI21_X1 U10177 ( .B1(n8951), .B2(n9839), .A(n8734), .ZN(n8736) );
  AOI21_X1 U10178 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n9839), .A(n8736), .ZN(
        n8735) );
  OAI21_X1 U10179 ( .B1(n8905), .B2(n8738), .A(n8735), .ZN(P2_U3202) );
  INV_X1 U10180 ( .A(n8318), .ZN(n8908) );
  AOI21_X1 U10181 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n9839), .A(n8736), .ZN(
        n8737) );
  OAI21_X1 U10182 ( .B1(n8908), .B2(n8738), .A(n8737), .ZN(P2_U3203) );
  XNOR2_X1 U10183 ( .A(n8739), .B(n8740), .ZN(n8961) );
  XNOR2_X1 U10184 ( .A(n8741), .B(n8740), .ZN(n8744) );
  AOI222_X1 U10185 ( .A1(n9829), .A2(n8744), .B1(n8743), .B2(n9826), .C1(n8742), .C2(n9824), .ZN(n8956) );
  MUX2_X1 U10186 ( .A(n8745), .B(n8956), .S(n9837), .Z(n8748) );
  AOI22_X1 U10187 ( .A1(n8958), .A2(n8899), .B1(n8898), .B2(n8746), .ZN(n8747)
         );
  OAI211_X1 U10188 ( .C1(n8961), .C2(n8903), .A(n8748), .B(n8747), .ZN(
        P2_U3206) );
  XNOR2_X1 U10189 ( .A(n8749), .B(n8750), .ZN(n8967) );
  INV_X1 U10190 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8752) );
  MUX2_X1 U10191 ( .A(n8752), .B(n8962), .S(n9837), .Z(n8755) );
  AOI22_X1 U10192 ( .A1(n8964), .A2(n8899), .B1(n8898), .B2(n8753), .ZN(n8754)
         );
  OAI211_X1 U10193 ( .C1(n8967), .C2(n8903), .A(n8755), .B(n8754), .ZN(
        P2_U3207) );
  XNOR2_X1 U10194 ( .A(n8756), .B(n8758), .ZN(n8970) );
  XOR2_X1 U10195 ( .A(n8758), .B(n8757), .Z(n8759) );
  OAI222_X1 U10196 ( .A1(n8864), .A2(n8760), .B1(n8866), .B2(n8199), .C1(n8862), .C2(n8759), .ZN(n8968) );
  INV_X1 U10197 ( .A(n8761), .ZN(n8762) );
  OAI22_X1 U10198 ( .A1(n8969), .A2(n9823), .B1(n8762), .B2(n9821), .ZN(n8763)
         );
  OAI21_X1 U10199 ( .B1(n8968), .B2(n8763), .A(n9837), .ZN(n8765) );
  NAND2_X1 U10200 ( .A1(n9839), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U10201 ( .C1(n8970), .C2(n8903), .A(n8765), .B(n8764), .ZN(
        P2_U3208) );
  INV_X1 U10202 ( .A(n8767), .ZN(n8769) );
  OAI21_X1 U10203 ( .B1(n8766), .B2(n8769), .A(n8768), .ZN(n8770) );
  XOR2_X1 U10204 ( .A(n8771), .B(n8770), .Z(n8978) );
  XNOR2_X1 U10205 ( .A(n8772), .B(n8771), .ZN(n8775) );
  AOI222_X1 U10206 ( .A1(n9829), .A2(n8775), .B1(n8774), .B2(n9824), .C1(n8773), .C2(n9826), .ZN(n8973) );
  INV_X1 U10207 ( .A(n8973), .ZN(n8780) );
  INV_X1 U10208 ( .A(n8776), .ZN(n8777) );
  OAI22_X1 U10209 ( .A1(n8778), .A2(n9823), .B1(n8777), .B2(n9821), .ZN(n8779)
         );
  OAI21_X1 U10210 ( .B1(n8780), .B2(n8779), .A(n9837), .ZN(n8782) );
  NAND2_X1 U10211 ( .A1(n9839), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8781) );
  OAI211_X1 U10212 ( .C1(n8978), .C2(n8903), .A(n8782), .B(n8781), .ZN(
        P2_U3209) );
  XOR2_X1 U10213 ( .A(n8766), .B(n8783), .Z(n8984) );
  XNOR2_X1 U10214 ( .A(n8784), .B(n8783), .ZN(n8786) );
  AOI222_X1 U10215 ( .A1(n9829), .A2(n8786), .B1(n8785), .B2(n9824), .C1(n8807), .C2(n9826), .ZN(n8979) );
  MUX2_X1 U10216 ( .A(n8787), .B(n8979), .S(n8894), .Z(n8790) );
  AOI22_X1 U10217 ( .A1(n8981), .A2(n8899), .B1(n8898), .B2(n8788), .ZN(n8789)
         );
  OAI211_X1 U10218 ( .C1(n8984), .C2(n8903), .A(n8790), .B(n8789), .ZN(
        P2_U3210) );
  XNOR2_X1 U10219 ( .A(n8791), .B(n8792), .ZN(n8988) );
  XNOR2_X1 U10220 ( .A(n8793), .B(n4609), .ZN(n8794) );
  OAI222_X1 U10221 ( .A1(n8864), .A2(n8796), .B1(n8866), .B2(n8795), .C1(n8862), .C2(n8794), .ZN(n8922) );
  NAND2_X1 U10222 ( .A1(n8922), .A2(n9837), .ZN(n8802) );
  INV_X1 U10223 ( .A(n8797), .ZN(n8799) );
  OAI22_X1 U10224 ( .A1(n8799), .A2(n9821), .B1(n8894), .B2(n8798), .ZN(n8800)
         );
  AOI21_X1 U10225 ( .B1(n8923), .B2(n8899), .A(n8800), .ZN(n8801) );
  OAI211_X1 U10226 ( .C1(n8988), .C2(n8903), .A(n8802), .B(n8801), .ZN(
        P2_U3211) );
  XNOR2_X1 U10227 ( .A(n8803), .B(n8804), .ZN(n8994) );
  XNOR2_X1 U10228 ( .A(n8805), .B(n8804), .ZN(n8808) );
  AOI222_X1 U10229 ( .A1(n9829), .A2(n8808), .B1(n8807), .B2(n9824), .C1(n8806), .C2(n9826), .ZN(n8989) );
  MUX2_X1 U10230 ( .A(n8809), .B(n8989), .S(n8894), .Z(n8812) );
  AOI22_X1 U10231 ( .A1(n8991), .A2(n8899), .B1(n8898), .B2(n8810), .ZN(n8811)
         );
  OAI211_X1 U10232 ( .C1(n8994), .C2(n8903), .A(n8812), .B(n8811), .ZN(
        P2_U3212) );
  XNOR2_X1 U10233 ( .A(n8813), .B(n8819), .ZN(n8997) );
  NAND2_X1 U10234 ( .A1(n8814), .A2(n8815), .ZN(n8859) );
  OR2_X1 U10235 ( .A1(n8859), .A2(n8816), .ZN(n8818) );
  AND2_X1 U10236 ( .A1(n8818), .A2(n8817), .ZN(n8820) );
  NAND2_X1 U10237 ( .A1(n8820), .A2(n8819), .ZN(n8821) );
  NAND2_X1 U10238 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U10239 ( .A1(n8823), .A2(n9829), .ZN(n8827) );
  AOI22_X1 U10240 ( .A1(n8825), .A2(n9824), .B1(n9826), .B2(n8824), .ZN(n8826)
         );
  NAND2_X1 U10241 ( .A1(n8827), .A2(n8826), .ZN(n8995) );
  MUX2_X1 U10242 ( .A(n8995), .B(P2_REG2_REG_20__SCAN_IN), .S(n9839), .Z(n8828) );
  INV_X1 U10243 ( .A(n8828), .ZN(n8832) );
  AOI22_X1 U10244 ( .A1(n8830), .A2(n8899), .B1(n8898), .B2(n8829), .ZN(n8831)
         );
  OAI211_X1 U10245 ( .C1(n8997), .C2(n8903), .A(n8832), .B(n8831), .ZN(
        P2_U3213) );
  OR2_X1 U10246 ( .A1(n8833), .A2(n8837), .ZN(n8834) );
  NAND2_X1 U10247 ( .A1(n8835), .A2(n8834), .ZN(n9003) );
  NAND2_X1 U10248 ( .A1(n8857), .A2(n8836), .ZN(n8838) );
  NAND2_X1 U10249 ( .A1(n8838), .A2(n8837), .ZN(n8841) );
  NAND2_X1 U10250 ( .A1(n8857), .A2(n8839), .ZN(n8840) );
  NAND3_X1 U10251 ( .A1(n8841), .A2(n9829), .A3(n8840), .ZN(n8846) );
  OAI22_X1 U10252 ( .A1(n8843), .A2(n8866), .B1(n8842), .B2(n8864), .ZN(n8844)
         );
  INV_X1 U10253 ( .A(n8844), .ZN(n8845) );
  MUX2_X1 U10254 ( .A(n9000), .B(n8847), .S(n9839), .Z(n8850) );
  AOI22_X1 U10255 ( .A1(n5985), .A2(n8899), .B1(n8898), .B2(n8848), .ZN(n8849)
         );
  OAI211_X1 U10256 ( .C1(n9003), .C2(n8903), .A(n8850), .B(n8849), .ZN(
        P2_U3214) );
  NAND2_X1 U10257 ( .A1(n8851), .A2(n8852), .ZN(n8854) );
  NAND2_X1 U10258 ( .A1(n8854), .A2(n8853), .ZN(n8856) );
  NAND2_X1 U10259 ( .A1(n8856), .A2(n8855), .ZN(n9007) );
  INV_X1 U10260 ( .A(n8857), .ZN(n8858) );
  AOI21_X1 U10261 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n8861) );
  OAI222_X1 U10262 ( .A1(n8866), .A2(n8865), .B1(n8864), .B2(n8863), .C1(n8862), .C2(n8861), .ZN(n8934) );
  NAND2_X1 U10263 ( .A1(n8934), .A2(n9837), .ZN(n8872) );
  INV_X1 U10264 ( .A(n8867), .ZN(n8868) );
  OAI22_X1 U10265 ( .A1(n8894), .A2(n8869), .B1(n8868), .B2(n9821), .ZN(n8870)
         );
  AOI21_X1 U10266 ( .B1(n8935), .B2(n8899), .A(n8870), .ZN(n8871) );
  OAI211_X1 U10267 ( .C1(n9007), .C2(n8903), .A(n8872), .B(n8871), .ZN(
        P2_U3215) );
  INV_X1 U10268 ( .A(n8851), .ZN(n8874) );
  AOI21_X1 U10269 ( .B1(n8875), .B2(n8873), .A(n8874), .ZN(n9014) );
  NAND3_X1 U10270 ( .A1(n8887), .A2(n6142), .A3(n8876), .ZN(n8877) );
  NAND3_X1 U10271 ( .A1(n8814), .A2(n9829), .A3(n8877), .ZN(n8881) );
  AOI22_X1 U10272 ( .A1(n8879), .A2(n9826), .B1(n8878), .B2(n9824), .ZN(n8880)
         );
  MUX2_X1 U10273 ( .A(n9009), .B(n8882), .S(n9839), .Z(n8885) );
  AOI22_X1 U10274 ( .A1(n9011), .A2(n8899), .B1(n8898), .B2(n8883), .ZN(n8884)
         );
  OAI211_X1 U10275 ( .C1(n9014), .C2(n8903), .A(n8885), .B(n8884), .ZN(
        P2_U3216) );
  XOR2_X1 U10276 ( .A(n8886), .B(n8889), .Z(n9019) );
  OAI211_X1 U10277 ( .C1(n8889), .C2(n8888), .A(n8887), .B(n9829), .ZN(n8893)
         );
  AOI22_X1 U10278 ( .A1(n9826), .A2(n8891), .B1(n8890), .B2(n9824), .ZN(n8892)
         );
  NAND2_X1 U10279 ( .A1(n8893), .A2(n8892), .ZN(n9015) );
  MUX2_X1 U10280 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9015), .S(n8894), .Z(n8895) );
  INV_X1 U10281 ( .A(n8895), .ZN(n8902) );
  INV_X1 U10282 ( .A(n8896), .ZN(n8897) );
  AOI22_X1 U10283 ( .A1(n8900), .A2(n8899), .B1(n8898), .B2(n8897), .ZN(n8901)
         );
  OAI211_X1 U10284 ( .C1(n9019), .C2(n8903), .A(n8902), .B(n8901), .ZN(
        P2_U3217) );
  NOR2_X1 U10285 ( .A1(n8951), .A2(n9913), .ZN(n8906) );
  AOI21_X1 U10286 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9913), .A(n8906), .ZN(
        n8904) );
  OAI21_X1 U10287 ( .B1(n8905), .B2(n8942), .A(n8904), .ZN(P2_U3490) );
  AOI21_X1 U10288 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9913), .A(n8906), .ZN(
        n8907) );
  OAI21_X1 U10289 ( .B1(n8908), .B2(n8942), .A(n8907), .ZN(P2_U3489) );
  INV_X1 U10290 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8909) );
  MUX2_X1 U10291 ( .A(n8909), .B(n8956), .S(n9915), .Z(n8911) );
  NAND2_X1 U10292 ( .A1(n8958), .A2(n8939), .ZN(n8910) );
  OAI211_X1 U10293 ( .C1(n8961), .C2(n8943), .A(n8911), .B(n8910), .ZN(
        P2_U3486) );
  MUX2_X1 U10294 ( .A(n10077), .B(n8962), .S(n9915), .Z(n8913) );
  NAND2_X1 U10295 ( .A1(n8964), .A2(n8939), .ZN(n8912) );
  OAI211_X1 U10296 ( .C1(n8943), .C2(n8967), .A(n8913), .B(n8912), .ZN(
        P2_U3485) );
  MUX2_X1 U10297 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8968), .S(n9915), .Z(n8915) );
  OAI22_X1 U10298 ( .A1(n8970), .A2(n8943), .B1(n8969), .B2(n8942), .ZN(n8914)
         );
  OR2_X1 U10299 ( .A1(n8915), .A2(n8914), .ZN(P2_U3484) );
  MUX2_X1 U10300 ( .A(n8916), .B(n8973), .S(n9915), .Z(n8918) );
  NAND2_X1 U10301 ( .A1(n8975), .A2(n8939), .ZN(n8917) );
  OAI211_X1 U10302 ( .C1(n8943), .C2(n8978), .A(n8918), .B(n8917), .ZN(
        P2_U3483) );
  INV_X1 U10303 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8919) );
  MUX2_X1 U10304 ( .A(n8919), .B(n8979), .S(n9915), .Z(n8921) );
  NAND2_X1 U10305 ( .A1(n8981), .A2(n8939), .ZN(n8920) );
  OAI211_X1 U10306 ( .C1(n8984), .C2(n8943), .A(n8921), .B(n8920), .ZN(
        P2_U3482) );
  INV_X1 U10307 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8924) );
  AOI21_X1 U10308 ( .B1(n9892), .B2(n8923), .A(n8922), .ZN(n8985) );
  MUX2_X1 U10309 ( .A(n8924), .B(n8985), .S(n9915), .Z(n8925) );
  OAI21_X1 U10310 ( .B1(n8988), .B2(n8943), .A(n8925), .ZN(P2_U3481) );
  INV_X1 U10311 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8926) );
  MUX2_X1 U10312 ( .A(n8926), .B(n8989), .S(n9915), .Z(n8928) );
  NAND2_X1 U10313 ( .A1(n8991), .A2(n8939), .ZN(n8927) );
  OAI211_X1 U10314 ( .C1(n8943), .C2(n8994), .A(n8928), .B(n8927), .ZN(
        P2_U3480) );
  MUX2_X1 U10315 ( .A(n8995), .B(P2_REG1_REG_20__SCAN_IN), .S(n9913), .Z(n8930) );
  OAI22_X1 U10316 ( .A1(n8997), .A2(n8943), .B1(n8996), .B2(n8942), .ZN(n8929)
         );
  OR2_X1 U10317 ( .A1(n8930), .A2(n8929), .ZN(P2_U3479) );
  MUX2_X1 U10318 ( .A(n9000), .B(n8931), .S(n9913), .Z(n8933) );
  NAND2_X1 U10319 ( .A1(n5985), .A2(n8939), .ZN(n8932) );
  OAI211_X1 U10320 ( .C1(n8943), .C2(n9003), .A(n8933), .B(n8932), .ZN(
        P2_U3478) );
  AOI21_X1 U10321 ( .B1(n9892), .B2(n8935), .A(n8934), .ZN(n9004) );
  MUX2_X1 U10322 ( .A(n8936), .B(n9004), .S(n9915), .Z(n8937) );
  OAI21_X1 U10323 ( .B1(n8943), .B2(n9007), .A(n8937), .ZN(P2_U3477) );
  MUX2_X1 U10324 ( .A(n9009), .B(n8938), .S(n9913), .Z(n8941) );
  NAND2_X1 U10325 ( .A1(n9011), .A2(n8939), .ZN(n8940) );
  OAI211_X1 U10326 ( .C1(n9014), .C2(n8943), .A(n8941), .B(n8940), .ZN(
        P2_U3476) );
  MUX2_X1 U10327 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9015), .S(n9915), .Z(n8945) );
  OAI22_X1 U10328 ( .A1(n9019), .A2(n8943), .B1(n9017), .B2(n8942), .ZN(n8944)
         );
  OR2_X1 U10329 ( .A1(n8945), .A2(n8944), .ZN(P2_U3475) );
  AOI22_X1 U10330 ( .A1(n8947), .A2(n9895), .B1(n9892), .B2(n8946), .ZN(n8949)
         );
  AND2_X1 U10331 ( .A1(n8949), .A2(n8948), .ZN(n9840) );
  INV_X1 U10332 ( .A(n9840), .ZN(n8950) );
  MUX2_X1 U10333 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8950), .S(n9915), .Z(
        P2_U3460) );
  NAND2_X1 U10334 ( .A1(n8319), .A2(n9010), .ZN(n8953) );
  INV_X1 U10335 ( .A(n8951), .ZN(n8952) );
  NAND2_X1 U10336 ( .A1(n8952), .A2(n9899), .ZN(n8954) );
  OAI211_X1 U10337 ( .C1(n8306), .C2(n9899), .A(n8953), .B(n8954), .ZN(
        P2_U3458) );
  NAND2_X1 U10338 ( .A1(n8318), .A2(n9010), .ZN(n8955) );
  OAI211_X1 U10339 ( .C1(n6545), .C2(n9899), .A(n8955), .B(n8954), .ZN(
        P2_U3457) );
  INV_X1 U10340 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8957) );
  MUX2_X1 U10341 ( .A(n8957), .B(n8956), .S(n9899), .Z(n8960) );
  NAND2_X1 U10342 ( .A1(n8958), .A2(n9010), .ZN(n8959) );
  OAI211_X1 U10343 ( .C1(n8961), .C2(n9018), .A(n8960), .B(n8959), .ZN(
        P2_U3454) );
  INV_X1 U10344 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8963) );
  MUX2_X1 U10345 ( .A(n8963), .B(n8962), .S(n9899), .Z(n8966) );
  NAND2_X1 U10346 ( .A1(n8964), .A2(n9010), .ZN(n8965) );
  OAI211_X1 U10347 ( .C1(n8967), .C2(n9018), .A(n8966), .B(n8965), .ZN(
        P2_U3453) );
  MUX2_X1 U10348 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8968), .S(n9899), .Z(n8972) );
  OAI22_X1 U10349 ( .A1(n8970), .A2(n9018), .B1(n8969), .B2(n9016), .ZN(n8971)
         );
  OR2_X1 U10350 ( .A1(n8972), .A2(n8971), .ZN(P2_U3452) );
  INV_X1 U10351 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8974) );
  MUX2_X1 U10352 ( .A(n8974), .B(n8973), .S(n9899), .Z(n8977) );
  NAND2_X1 U10353 ( .A1(n8975), .A2(n9010), .ZN(n8976) );
  OAI211_X1 U10354 ( .C1(n8978), .C2(n9018), .A(n8977), .B(n8976), .ZN(
        P2_U3451) );
  INV_X1 U10355 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8980) );
  MUX2_X1 U10356 ( .A(n8980), .B(n8979), .S(n9899), .Z(n8983) );
  NAND2_X1 U10357 ( .A1(n8981), .A2(n9010), .ZN(n8982) );
  OAI211_X1 U10358 ( .C1(n8984), .C2(n9018), .A(n8983), .B(n8982), .ZN(
        P2_U3450) );
  INV_X1 U10359 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U10360 ( .A(n8986), .B(n8985), .S(n9899), .Z(n8987) );
  OAI21_X1 U10361 ( .B1(n8988), .B2(n9018), .A(n8987), .ZN(P2_U3449) );
  INV_X1 U10362 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8990) );
  MUX2_X1 U10363 ( .A(n8990), .B(n8989), .S(n9899), .Z(n8993) );
  NAND2_X1 U10364 ( .A1(n8991), .A2(n9010), .ZN(n8992) );
  OAI211_X1 U10365 ( .C1(n8994), .C2(n9018), .A(n8993), .B(n8992), .ZN(
        P2_U3448) );
  MUX2_X1 U10366 ( .A(n8995), .B(P2_REG0_REG_20__SCAN_IN), .S(n9901), .Z(n8999) );
  OAI22_X1 U10367 ( .A1(n8997), .A2(n9018), .B1(n8996), .B2(n9016), .ZN(n8998)
         );
  OR2_X1 U10368 ( .A1(n8999), .A2(n8998), .ZN(P2_U3447) );
  MUX2_X1 U10369 ( .A(n9000), .B(n9982), .S(n9901), .Z(n9002) );
  NAND2_X1 U10370 ( .A1(n5985), .A2(n9010), .ZN(n9001) );
  OAI211_X1 U10371 ( .C1(n9003), .C2(n9018), .A(n9002), .B(n9001), .ZN(
        P2_U3446) );
  MUX2_X1 U10372 ( .A(n9005), .B(n9004), .S(n9899), .Z(n9006) );
  OAI21_X1 U10373 ( .B1(n9007), .B2(n9018), .A(n9006), .ZN(P2_U3444) );
  MUX2_X1 U10374 ( .A(n9009), .B(n9008), .S(n9901), .Z(n9013) );
  NAND2_X1 U10375 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  OAI211_X1 U10376 ( .C1(n9014), .C2(n9018), .A(n9013), .B(n9012), .ZN(
        P2_U3441) );
  MUX2_X1 U10377 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9015), .S(n9899), .Z(n9021) );
  OAI22_X1 U10378 ( .A1(n9019), .A2(n9018), .B1(n9017), .B2(n9016), .ZN(n9020)
         );
  OR2_X1 U10379 ( .A1(n9021), .A2(n9020), .ZN(P2_U3438) );
  INV_X1 U10380 ( .A(n9022), .ZN(n9725) );
  NAND3_X1 U10381 ( .A1(n9024), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9027) );
  OAI22_X1 U10382 ( .A1(n9023), .A2(n9027), .B1(n9026), .B2(n9025), .ZN(n9028)
         );
  INV_X1 U10383 ( .A(n9028), .ZN(n9029) );
  OAI21_X1 U10384 ( .B1(n9725), .B2(n9034), .A(n9029), .ZN(P2_U3264) );
  INV_X1 U10385 ( .A(n9030), .ZN(n9727) );
  OAI222_X1 U10386 ( .A1(n9034), .A2(n9727), .B1(n9033), .B2(P2_U3151), .C1(
        n9032), .C2(n9031), .ZN(P2_U3266) );
  INV_X1 U10387 ( .A(n9035), .ZN(n9036) );
  MUX2_X1 U10388 ( .A(n9036), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10389 ( .A(n9039), .B(n9038), .ZN(n9040) );
  XNOR2_X1 U10390 ( .A(n9037), .B(n9040), .ZN(n9047) );
  AOI22_X1 U10391 ( .A1(n9041), .A2(n9224), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n9042) );
  OAI21_X1 U10392 ( .B1(n9226), .B2(n9043), .A(n9042), .ZN(n9044) );
  AOI21_X1 U10393 ( .B1(n9045), .B2(n9228), .A(n9044), .ZN(n9046) );
  OAI21_X1 U10394 ( .B1(n9047), .B2(n10103), .A(n9046), .ZN(P1_U3215) );
  NAND2_X1 U10395 ( .A1(n9049), .A2(n9050), .ZN(n9053) );
  NAND2_X1 U10396 ( .A1(n9051), .A2(n9154), .ZN(n9052) );
  XNOR2_X1 U10397 ( .A(n9053), .B(n9052), .ZN(n9059) );
  NAND2_X1 U10398 ( .A1(n9250), .A2(n9196), .ZN(n9055) );
  OR2_X1 U10399 ( .A1(n9109), .A2(n9220), .ZN(n9054) );
  NAND2_X1 U10400 ( .A1(n9055), .A2(n9054), .ZN(n9450) );
  AOI22_X1 U10401 ( .A1(n9450), .A2(n9224), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9056) );
  OAI21_X1 U10402 ( .B1(n9226), .B2(n9453), .A(n9056), .ZN(n9057) );
  AOI21_X1 U10403 ( .B1(n9609), .B2(n9228), .A(n9057), .ZN(n9058) );
  OAI21_X1 U10404 ( .B1(n9059), .B2(n10103), .A(n9058), .ZN(P1_U3216) );
  XNOR2_X1 U10405 ( .A(n9060), .B(n9205), .ZN(n9062) );
  NOR2_X1 U10406 ( .A1(n9062), .A2(n9061), .ZN(n9204) );
  AOI21_X1 U10407 ( .B1(n9062), .B2(n9061), .A(n9204), .ZN(n9069) );
  AOI22_X1 U10408 ( .A1(n9063), .A2(n9224), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n9064) );
  OAI21_X1 U10409 ( .B1(n9226), .B2(n9065), .A(n9064), .ZN(n9066) );
  AOI21_X1 U10410 ( .B1(n9067), .B2(n9228), .A(n9066), .ZN(n9068) );
  OAI21_X1 U10411 ( .B1(n9069), .B2(n10103), .A(n9068), .ZN(P1_U3217) );
  NAND2_X1 U10412 ( .A1(n9071), .A2(n9072), .ZN(n9074) );
  NAND2_X1 U10413 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  NAND2_X1 U10414 ( .A1(n9070), .A2(n9075), .ZN(n9218) );
  OR2_X1 U10415 ( .A1(n9218), .A2(n9219), .ZN(n9216) );
  NAND2_X1 U10416 ( .A1(n9216), .A2(n9070), .ZN(n9078) );
  NAND2_X1 U10417 ( .A1(n9172), .A2(n9076), .ZN(n9077) );
  XNOR2_X1 U10418 ( .A(n9078), .B(n9077), .ZN(n9084) );
  NAND2_X1 U10419 ( .A1(n9256), .A2(n9237), .ZN(n9080) );
  NAND2_X1 U10420 ( .A1(n9254), .A2(n9196), .ZN(n9079) );
  NAND2_X1 U10421 ( .A1(n9080), .A2(n9079), .ZN(n9513) );
  AOI22_X1 U10422 ( .A1(n9513), .A2(n9224), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9081) );
  OAI21_X1 U10423 ( .B1(n9226), .B2(n9506), .A(n9081), .ZN(n9082) );
  AOI21_X1 U10424 ( .B1(n9630), .B2(n9228), .A(n9082), .ZN(n9083) );
  OAI21_X1 U10425 ( .B1(n9084), .B2(n10103), .A(n9083), .ZN(P1_U3219) );
  NAND2_X1 U10426 ( .A1(n9380), .A2(n6205), .ZN(n9087) );
  OR2_X1 U10427 ( .A1(n9090), .A2(n9085), .ZN(n9086) );
  NAND2_X1 U10428 ( .A1(n9087), .A2(n9086), .ZN(n9089) );
  XNOR2_X1 U10429 ( .A(n9089), .B(n9088), .ZN(n9094) );
  NOR2_X1 U10430 ( .A1(n9090), .A2(n6264), .ZN(n9091) );
  AOI21_X1 U10431 ( .B1(n9380), .B2(n9092), .A(n9091), .ZN(n9093) );
  XNOR2_X1 U10432 ( .A(n9094), .B(n9093), .ZN(n9100) );
  INV_X1 U10433 ( .A(n9100), .ZN(n9095) );
  NAND2_X1 U10434 ( .A1(n9095), .A2(n6436), .ZN(n9106) );
  NAND4_X1 U10435 ( .A1(n9105), .A2(n6436), .A3(n9099), .A4(n9100), .ZN(n9104)
         );
  INV_X1 U10436 ( .A(n9379), .ZN(n9098) );
  AOI22_X1 U10437 ( .A1(n9096), .A2(n9224), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9097) );
  OAI21_X1 U10438 ( .B1(n9226), .B2(n9098), .A(n9097), .ZN(n9102) );
  NOR3_X1 U10439 ( .A1(n9100), .A2(n9099), .A3(n10103), .ZN(n9101) );
  AOI211_X1 U10440 ( .C1(n9228), .C2(n9380), .A(n9102), .B(n9101), .ZN(n9103)
         );
  OAI211_X1 U10441 ( .C1(n9106), .C2(n9105), .A(n9104), .B(n9103), .ZN(
        P1_U3220) );
  XOR2_X1 U10442 ( .A(n9107), .B(n9108), .Z(n9115) );
  OR2_X1 U10443 ( .A1(n9109), .A2(n9235), .ZN(n9111) );
  NAND2_X1 U10444 ( .A1(n9254), .A2(n9237), .ZN(n9110) );
  NAND2_X1 U10445 ( .A1(n9111), .A2(n9110), .ZN(n9477) );
  AOI22_X1 U10446 ( .A1(n9477), .A2(n9224), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9112) );
  OAI21_X1 U10447 ( .B1(n9226), .B2(n9482), .A(n9112), .ZN(n9113) );
  AOI21_X1 U10448 ( .B1(n9618), .B2(n9228), .A(n9113), .ZN(n9114) );
  OAI21_X1 U10449 ( .B1(n9115), .B2(n10103), .A(n9114), .ZN(P1_U3223) );
  XOR2_X1 U10450 ( .A(n9116), .B(n9117), .Z(n9126) );
  INV_X1 U10451 ( .A(n9118), .ZN(n9119) );
  NAND2_X1 U10452 ( .A1(n9242), .A2(n9119), .ZN(n9121) );
  OAI211_X1 U10453 ( .C1(n9122), .C2(n10098), .A(n9121), .B(n9120), .ZN(n9123)
         );
  AOI21_X1 U10454 ( .B1(n9124), .B2(n9228), .A(n9123), .ZN(n9125) );
  OAI21_X1 U10455 ( .B1(n9126), .B2(n10103), .A(n9125), .ZN(P1_U3224) );
  OAI21_X1 U10456 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9130) );
  NAND2_X1 U10457 ( .A1(n9130), .A2(n6436), .ZN(n9134) );
  AOI22_X1 U10458 ( .A1(n9249), .A2(n9196), .B1(n9237), .B2(n9250), .ZN(n9420)
         );
  OAI22_X1 U10459 ( .A1(n9420), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9131), .ZN(n9132) );
  AOI21_X1 U10460 ( .B1(n9424), .B2(n9242), .A(n9132), .ZN(n9133) );
  OAI211_X1 U10461 ( .C1(n9427), .C2(n10096), .A(n9134), .B(n9133), .ZN(
        P1_U3225) );
  XOR2_X1 U10462 ( .A(n9135), .B(n9136), .Z(n9144) );
  OR2_X1 U10463 ( .A1(n9137), .A2(n9220), .ZN(n9139) );
  OR2_X1 U10464 ( .A1(n9221), .A2(n9235), .ZN(n9138) );
  NAND2_X1 U10465 ( .A1(n9139), .A2(n9138), .ZN(n9565) );
  NAND2_X1 U10466 ( .A1(n9565), .A2(n9224), .ZN(n9141) );
  OAI211_X1 U10467 ( .C1(n9226), .C2(n9558), .A(n9141), .B(n9140), .ZN(n9142)
         );
  AOI21_X1 U10468 ( .B1(n9644), .B2(n9228), .A(n9142), .ZN(n9143) );
  OAI21_X1 U10469 ( .B1(n9144), .B2(n10103), .A(n9143), .ZN(P1_U3226) );
  AOI21_X1 U10470 ( .B1(n9146), .B2(n9145), .A(n10103), .ZN(n9147) );
  NAND2_X1 U10471 ( .A1(n9147), .A2(n9071), .ZN(n9153) );
  OR2_X1 U10472 ( .A1(n9236), .A2(n9220), .ZN(n9149) );
  NAND2_X1 U10473 ( .A1(n9256), .A2(n9196), .ZN(n9148) );
  NAND2_X1 U10474 ( .A1(n9149), .A2(n9148), .ZN(n9546) );
  NOR2_X1 U10475 ( .A1(n9226), .A2(n9538), .ZN(n9150) );
  AOI211_X1 U10476 ( .C1(n9224), .C2(n9546), .A(n9151), .B(n9150), .ZN(n9152)
         );
  OAI211_X1 U10477 ( .C1(n9537), .C2(n10096), .A(n9153), .B(n9152), .ZN(
        P1_U3228) );
  AND2_X1 U10478 ( .A1(n9155), .A2(n9154), .ZN(n9157) );
  OAI21_X1 U10479 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9165) );
  NAND2_X1 U10480 ( .A1(n9678), .A2(n9228), .ZN(n9163) );
  OR2_X1 U10481 ( .A1(n9159), .A2(n9235), .ZN(n9161) );
  NAND2_X1 U10482 ( .A1(n9251), .A2(n9237), .ZN(n9160) );
  NAND2_X1 U10483 ( .A1(n9161), .A2(n9160), .ZN(n9432) );
  AOI22_X1 U10484 ( .A1(n9432), .A2(n9224), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9162) );
  OAI211_X1 U10485 ( .C1(n9226), .C2(n9438), .A(n9163), .B(n9162), .ZN(n9164)
         );
  AOI21_X1 U10486 ( .B1(n9165), .B2(n6436), .A(n9164), .ZN(n9166) );
  INV_X1 U10487 ( .A(n9166), .ZN(P1_U3229) );
  NAND2_X1 U10488 ( .A1(n9071), .A2(n9168), .ZN(n9170) );
  NAND2_X1 U10489 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  NAND2_X1 U10490 ( .A1(n9167), .A2(n9171), .ZN(n9173) );
  AND2_X1 U10491 ( .A1(n9173), .A2(n9172), .ZN(n9176) );
  AOI21_X1 U10492 ( .B1(n9177), .B2(n9176), .A(n4378), .ZN(n9182) );
  NOR2_X1 U10493 ( .A1(n9226), .A2(n9499), .ZN(n9180) );
  INV_X1 U10494 ( .A(n9223), .ZN(n9255) );
  AOI22_X1 U10495 ( .A1(n9196), .A2(n9253), .B1(n9255), .B2(n9237), .ZN(n9496)
         );
  OAI22_X1 U10496 ( .A1(n9496), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9178), .ZN(n9179) );
  AOI211_X1 U10497 ( .C1(n9625), .C2(n9228), .A(n9180), .B(n9179), .ZN(n9181)
         );
  OAI21_X1 U10498 ( .B1(n9182), .B2(n10103), .A(n9181), .ZN(P1_U3233) );
  XOR2_X1 U10499 ( .A(n9184), .B(n9183), .Z(n9192) );
  NOR2_X1 U10500 ( .A1(n9226), .A2(n9185), .ZN(n9189) );
  OAI22_X1 U10501 ( .A1(n9187), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9186), .ZN(n9188) );
  AOI211_X1 U10502 ( .C1(n9190), .C2(n9228), .A(n9189), .B(n9188), .ZN(n9191)
         );
  OAI21_X1 U10503 ( .B1(n9192), .B2(n10103), .A(n9191), .ZN(P1_U3234) );
  OAI21_X1 U10504 ( .B1(n9194), .B2(n9193), .A(n9049), .ZN(n9202) );
  NAND2_X1 U10505 ( .A1(n9614), .A2(n9228), .ZN(n9200) );
  OR2_X1 U10506 ( .A1(n9195), .A2(n9220), .ZN(n9198) );
  NAND2_X1 U10507 ( .A1(n9251), .A2(n9196), .ZN(n9197) );
  NAND2_X1 U10508 ( .A1(n9198), .A2(n9197), .ZN(n9468) );
  AOI22_X1 U10509 ( .A1(n9468), .A2(n9224), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9199) );
  OAI211_X1 U10510 ( .C1(n9226), .C2(n9471), .A(n9200), .B(n9199), .ZN(n9201)
         );
  AOI21_X1 U10511 ( .B1(n9202), .B2(n6436), .A(n9201), .ZN(n9203) );
  INV_X1 U10512 ( .A(n9203), .ZN(P1_U3235) );
  AOI21_X1 U10513 ( .B1(n9205), .B2(n9060), .A(n9204), .ZN(n9209) );
  XNOR2_X1 U10514 ( .A(n9207), .B(n9206), .ZN(n9208) );
  XNOR2_X1 U10515 ( .A(n9209), .B(n9208), .ZN(n9215) );
  AOI22_X1 U10516 ( .A1(n9210), .A2(n9224), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9211) );
  OAI21_X1 U10517 ( .B1(n9226), .B2(n9212), .A(n9211), .ZN(n9213) );
  AOI21_X1 U10518 ( .B1(n9662), .B2(n9228), .A(n9213), .ZN(n9214) );
  OAI21_X1 U10519 ( .B1(n9215), .B2(n10103), .A(n9214), .ZN(P1_U3236) );
  INV_X1 U10520 ( .A(n9216), .ZN(n9217) );
  AOI21_X1 U10521 ( .B1(n9219), .B2(n9218), .A(n9217), .ZN(n9230) );
  OR2_X1 U10522 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  OAI21_X1 U10523 ( .B1(n9223), .B2(n9235), .A(n9222), .ZN(n9521) );
  NAND2_X1 U10524 ( .A1(n9521), .A2(n9224), .ZN(n9225) );
  NAND2_X1 U10525 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9334) );
  OAI211_X1 U10526 ( .C1(n9226), .C2(n9526), .A(n9225), .B(n9334), .ZN(n9227)
         );
  AOI21_X1 U10527 ( .B1(n9697), .B2(n9228), .A(n9227), .ZN(n9229) );
  OAI21_X1 U10528 ( .B1(n9230), .B2(n10103), .A(n9229), .ZN(P1_U3238) );
  OAI21_X1 U10529 ( .B1(n9233), .B2(n9232), .A(n9231), .ZN(n9234) );
  NAND2_X1 U10530 ( .A1(n9234), .A2(n6436), .ZN(n9245) );
  INV_X1 U10531 ( .A(n9582), .ZN(n9243) );
  OR2_X1 U10532 ( .A1(n9236), .A2(n9235), .ZN(n9239) );
  NAND2_X1 U10533 ( .A1(n9259), .A2(n9237), .ZN(n9238) );
  AND2_X1 U10534 ( .A1(n9239), .A2(n9238), .ZN(n9577) );
  OAI22_X1 U10535 ( .A1(n9577), .A2(n10098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9240), .ZN(n9241) );
  AOI21_X1 U10536 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9244) );
  OAI211_X1 U10537 ( .C1(n9648), .C2(n10096), .A(n9245), .B(n9244), .ZN(
        P1_U3241) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9246), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9247), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10540 ( .A(n9248), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9272), .Z(
        P1_U3581) );
  MUX2_X1 U10541 ( .A(n9249), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9272), .Z(
        P1_U3580) );
  MUX2_X1 U10542 ( .A(n9250), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9272), .Z(
        P1_U3578) );
  MUX2_X1 U10543 ( .A(n9251), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9272), .Z(
        P1_U3577) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9252), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9253), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10546 ( .A(n9254), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9272), .Z(
        P1_U3574) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9255), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10548 ( .A(n9256), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9272), .Z(
        P1_U3572) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9257), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10550 ( .A(n9258), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9272), .Z(
        P1_U3569) );
  MUX2_X1 U10551 ( .A(n9259), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9272), .Z(
        P1_U3568) );
  MUX2_X1 U10552 ( .A(n9260), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9272), .Z(
        P1_U3567) );
  MUX2_X1 U10553 ( .A(n9261), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9272), .Z(
        P1_U3566) );
  MUX2_X1 U10554 ( .A(n9262), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9272), .Z(
        P1_U3565) );
  MUX2_X1 U10555 ( .A(n9263), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9272), .Z(
        P1_U3564) );
  MUX2_X1 U10556 ( .A(n9264), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9272), .Z(
        P1_U3563) );
  MUX2_X1 U10557 ( .A(n9265), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9272), .Z(
        P1_U3562) );
  MUX2_X1 U10558 ( .A(n9266), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9272), .Z(
        P1_U3561) );
  MUX2_X1 U10559 ( .A(n9267), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9272), .Z(
        P1_U3560) );
  MUX2_X1 U10560 ( .A(n9268), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9272), .Z(
        P1_U3559) );
  MUX2_X1 U10561 ( .A(n9269), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9272), .Z(
        P1_U3558) );
  MUX2_X1 U10562 ( .A(n9270), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9272), .Z(
        P1_U3557) );
  MUX2_X1 U10563 ( .A(n9271), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9272), .Z(
        P1_U3556) );
  MUX2_X1 U10564 ( .A(n6942), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9272), .Z(
        P1_U3555) );
  OAI211_X1 U10565 ( .C1(n9275), .C2(n9274), .A(n9354), .B(n9273), .ZN(n9282)
         );
  AOI22_X1 U10566 ( .A1(n9739), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9281) );
  NAND2_X1 U10567 ( .A1(n9359), .A2(n9276), .ZN(n9280) );
  OAI211_X1 U10568 ( .C1(n9278), .C2(n9284), .A(n9360), .B(n9277), .ZN(n9279)
         );
  NAND4_X1 U10569 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(
        P1_U3244) );
  AOI21_X1 U10570 ( .B1(n9735), .B2(n4892), .A(n5672), .ZN(n9734) );
  MUX2_X1 U10571 ( .A(n9284), .B(n9283), .S(n5673), .Z(n9286) );
  NAND2_X1 U10572 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  OAI211_X1 U10573 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9734), .A(n9287), .B(
        P1_U3973), .ZN(n9328) );
  INV_X1 U10574 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9289) );
  OAI22_X1 U10575 ( .A1(n9366), .A2(n9289), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9288), .ZN(n9290) );
  AOI21_X1 U10576 ( .B1(n9359), .B2(n9291), .A(n9290), .ZN(n9300) );
  OAI211_X1 U10577 ( .C1(n9294), .C2(n9293), .A(n9360), .B(n9292), .ZN(n9299)
         );
  OAI211_X1 U10578 ( .C1(n9297), .C2(n9296), .A(n9354), .B(n9295), .ZN(n9298)
         );
  NAND4_X1 U10579 ( .A1(n9328), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(
        P1_U3245) );
  INV_X1 U10580 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U10581 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9301) );
  OAI21_X1 U10582 ( .B1(n9366), .B2(n9302), .A(n9301), .ZN(n9303) );
  AOI21_X1 U10583 ( .B1(n9359), .B2(n9304), .A(n9303), .ZN(n9313) );
  OAI211_X1 U10584 ( .C1(n9307), .C2(n9306), .A(n9360), .B(n9305), .ZN(n9312)
         );
  OAI211_X1 U10585 ( .C1(n9310), .C2(n9309), .A(n9354), .B(n9308), .ZN(n9311)
         );
  NAND3_X1 U10586 ( .A1(n9313), .A2(n9312), .A3(n9311), .ZN(P1_U3246) );
  INV_X1 U10587 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9316) );
  INV_X1 U10588 ( .A(n9314), .ZN(n9315) );
  OAI21_X1 U10589 ( .B1(n9366), .B2(n9316), .A(n9315), .ZN(n9317) );
  AOI21_X1 U10590 ( .B1(n9359), .B2(n9318), .A(n9317), .ZN(n9327) );
  OAI211_X1 U10591 ( .C1(n9321), .C2(n9320), .A(n9354), .B(n9319), .ZN(n9326)
         );
  OAI211_X1 U10592 ( .C1(n9324), .C2(n9323), .A(n9360), .B(n9322), .ZN(n9325)
         );
  NAND4_X1 U10593 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(
        P1_U3247) );
  AND2_X1 U10594 ( .A1(n9330), .A2(n9329), .ZN(n9333) );
  OR2_X1 U10595 ( .A1(n9341), .A2(n9527), .ZN(n9347) );
  NAND2_X1 U10596 ( .A1(n9341), .A2(n9527), .ZN(n9331) );
  AND2_X1 U10597 ( .A1(n9347), .A2(n9331), .ZN(n9332) );
  NAND2_X1 U10598 ( .A1(n9333), .A2(n9332), .ZN(n9348) );
  OAI211_X1 U10599 ( .C1(n9333), .C2(n9332), .A(n9348), .B(n9360), .ZN(n9346)
         );
  INV_X1 U10600 ( .A(n9341), .ZN(n9336) );
  OAI21_X1 U10601 ( .B1(n9366), .B2(n9922), .A(n9334), .ZN(n9335) );
  AOI21_X1 U10602 ( .B1(n9359), .B2(n9336), .A(n9335), .ZN(n9345) );
  INV_X1 U10603 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9340) );
  NOR2_X1 U10604 ( .A1(n9341), .A2(n9340), .ZN(n9350) );
  AOI21_X1 U10605 ( .B1(n9341), .B2(n9340), .A(n9350), .ZN(n9342) );
  NAND2_X1 U10606 ( .A1(n9343), .A2(n9342), .ZN(n9352) );
  OAI211_X1 U10607 ( .C1(n9343), .C2(n9342), .A(n9352), .B(n9354), .ZN(n9344)
         );
  NAND3_X1 U10608 ( .A1(n9346), .A2(n9345), .A3(n9344), .ZN(P1_U3261) );
  NAND2_X1 U10609 ( .A1(n9348), .A2(n9347), .ZN(n9349) );
  XNOR2_X1 U10610 ( .A(n9349), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9361) );
  INV_X1 U10611 ( .A(n9361), .ZN(n9355) );
  INV_X1 U10612 ( .A(n9350), .ZN(n9351) );
  NAND2_X1 U10613 ( .A1(n9352), .A2(n9351), .ZN(n9353) );
  XNOR2_X1 U10614 ( .A(n9353), .B(n9631), .ZN(n9357) );
  AOI22_X1 U10615 ( .A1(n9355), .A2(n9360), .B1(n9354), .B2(n9357), .ZN(n9363)
         );
  NOR2_X1 U10616 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  AOI211_X1 U10617 ( .C1(n9361), .C2(n9360), .A(n9359), .B(n9358), .ZN(n9362)
         );
  MUX2_X1 U10618 ( .A(n9363), .B(n9362), .S(n5619), .Z(n9365) );
  NAND2_X1 U10619 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9364) );
  OAI211_X1 U10620 ( .C1(n4880), .C2(n9366), .A(n9365), .B(n9364), .ZN(
        P1_U3262) );
  NOR2_X1 U10621 ( .A1(n9367), .A2(n9778), .ZN(n9375) );
  NOR2_X1 U10622 ( .A1(n9745), .A2(n9368), .ZN(n9369) );
  AOI211_X1 U10623 ( .C1(n9370), .C2(n9769), .A(n9375), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10624 ( .B1(n9372), .B2(n9760), .A(n9371), .ZN(P1_U3263) );
  NOR2_X1 U10625 ( .A1(n9373), .A2(n9556), .ZN(n9374) );
  AOI211_X1 U10626 ( .C1(n9778), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9375), .B(
        n9374), .ZN(n9376) );
  OAI21_X1 U10627 ( .B1(n9760), .B2(n9377), .A(n9376), .ZN(P1_U3264) );
  INV_X1 U10628 ( .A(n9378), .ZN(n9385) );
  AOI22_X1 U10629 ( .A1(n9379), .A2(n9767), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9778), .ZN(n9382) );
  NAND2_X1 U10630 ( .A1(n9380), .A2(n9769), .ZN(n9381) );
  OAI211_X1 U10631 ( .C1(n9383), .C2(n9760), .A(n9382), .B(n9381), .ZN(n9384)
         );
  AOI21_X1 U10632 ( .B1(n9385), .B2(n9568), .A(n9384), .ZN(n9386) );
  OAI21_X1 U10633 ( .B1(n9387), .B2(n9589), .A(n9386), .ZN(P1_U3265) );
  INV_X1 U10634 ( .A(n9388), .ZN(n9397) );
  NAND2_X1 U10635 ( .A1(n9389), .A2(n9772), .ZN(n9392) );
  AOI22_X1 U10636 ( .A1(n9390), .A2(n9767), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9778), .ZN(n9391) );
  OAI211_X1 U10637 ( .C1(n9393), .C2(n9556), .A(n9392), .B(n9391), .ZN(n9394)
         );
  AOI21_X1 U10638 ( .B1(n9395), .B2(n9568), .A(n9394), .ZN(n9396) );
  OAI21_X1 U10639 ( .B1(n9397), .B2(n9589), .A(n9396), .ZN(P1_U3266) );
  OR2_X1 U10640 ( .A1(n9398), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U10641 ( .A1(n9401), .A2(n9400), .ZN(n9402) );
  XOR2_X1 U10642 ( .A(n9403), .B(n9402), .Z(n9671) );
  XNOR2_X1 U10643 ( .A(n9404), .B(n9403), .ZN(n9407) );
  INV_X1 U10644 ( .A(n9405), .ZN(n9406) );
  AOI21_X1 U10645 ( .B1(n9407), .B2(n9575), .A(n9406), .ZN(n9595) );
  INV_X1 U10646 ( .A(n9595), .ZN(n9415) );
  INV_X1 U10647 ( .A(n9408), .ZN(n9423) );
  OAI211_X1 U10648 ( .C1(n9423), .C2(n9410), .A(n6447), .B(n9409), .ZN(n9594)
         );
  AOI22_X1 U10649 ( .A1(n9411), .A2(n9767), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9778), .ZN(n9413) );
  NAND2_X1 U10650 ( .A1(n9669), .A2(n9769), .ZN(n9412) );
  OAI211_X1 U10651 ( .C1(n9594), .C2(n9760), .A(n9413), .B(n9412), .ZN(n9414)
         );
  AOI21_X1 U10652 ( .B1(n9415), .B2(n9568), .A(n9414), .ZN(n9416) );
  OAI21_X1 U10653 ( .B1(n9671), .B2(n9589), .A(n9416), .ZN(P1_U3267) );
  XOR2_X1 U10654 ( .A(n9398), .B(n9418), .Z(n9675) );
  OAI211_X1 U10655 ( .C1(n9419), .C2(n9418), .A(n9417), .B(n9575), .ZN(n9421)
         );
  NAND2_X1 U10656 ( .A1(n9421), .A2(n9420), .ZN(n9599) );
  INV_X1 U10657 ( .A(n9422), .ZN(n9440) );
  AOI211_X1 U10658 ( .C1(n9600), .C2(n9440), .A(n9579), .B(n9423), .ZN(n9598)
         );
  NAND2_X1 U10659 ( .A1(n9598), .A2(n9772), .ZN(n9426) );
  AOI22_X1 U10660 ( .A1(n9424), .A2(n9767), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9778), .ZN(n9425) );
  OAI211_X1 U10661 ( .C1(n9427), .C2(n9556), .A(n9426), .B(n9425), .ZN(n9428)
         );
  AOI21_X1 U10662 ( .B1(n9568), .B2(n9599), .A(n9428), .ZN(n9429) );
  OAI21_X1 U10663 ( .B1(n9675), .B2(n9589), .A(n9429), .ZN(P1_U3268) );
  AOI21_X1 U10664 ( .B1(n9431), .B2(n9430), .A(n9497), .ZN(n9434) );
  AOI21_X1 U10665 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9604) );
  XNOR2_X1 U10666 ( .A(n9435), .B(n9436), .ZN(n9680) );
  INV_X1 U10667 ( .A(n9680), .ZN(n9437) );
  NAND2_X1 U10668 ( .A1(n9437), .A2(n9763), .ZN(n9445) );
  OAI22_X1 U10669 ( .A1(n9568), .A2(n9439), .B1(n9438), .B2(n9754), .ZN(n9443)
         );
  OAI211_X1 U10670 ( .C1(n9441), .C2(n4395), .A(n9440), .B(n6447), .ZN(n9603)
         );
  NOR2_X1 U10671 ( .A1(n9603), .A2(n9760), .ZN(n9442) );
  AOI211_X1 U10672 ( .C1(n9769), .C2(n9678), .A(n9443), .B(n9442), .ZN(n9444)
         );
  OAI211_X1 U10673 ( .C1(n9778), .C2(n9604), .A(n9445), .B(n9444), .ZN(
        P1_U3269) );
  XOR2_X1 U10674 ( .A(n9446), .B(n9447), .Z(n9684) );
  XNOR2_X1 U10675 ( .A(n9448), .B(n9447), .ZN(n9449) );
  NAND2_X1 U10676 ( .A1(n9449), .A2(n9575), .ZN(n9452) );
  INV_X1 U10677 ( .A(n9450), .ZN(n9451) );
  NAND2_X1 U10678 ( .A1(n9452), .A2(n9451), .ZN(n9608) );
  AOI211_X1 U10679 ( .C1(n9609), .C2(n9460), .A(n9579), .B(n4395), .ZN(n9607)
         );
  NAND2_X1 U10680 ( .A1(n9607), .A2(n9772), .ZN(n9456) );
  INV_X1 U10681 ( .A(n9453), .ZN(n9454) );
  AOI22_X1 U10682 ( .A1(n9778), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9454), .B2(
        n9767), .ZN(n9455) );
  OAI211_X1 U10683 ( .C1(n4514), .C2(n9556), .A(n9456), .B(n9455), .ZN(n9457)
         );
  AOI21_X1 U10684 ( .B1(n9568), .B2(n9608), .A(n9457), .ZN(n9458) );
  OAI21_X1 U10685 ( .B1(n9684), .B2(n9589), .A(n9458), .ZN(P1_U3270) );
  XOR2_X1 U10686 ( .A(n9459), .B(n9466), .Z(n9616) );
  INV_X1 U10687 ( .A(n9460), .ZN(n9461) );
  AOI211_X1 U10688 ( .C1(n9614), .C2(n9485), .A(n9579), .B(n9461), .ZN(n9612)
         );
  OAI22_X1 U10689 ( .A1(n9463), .A2(n9556), .B1(n9462), .B2(n9568), .ZN(n9464)
         );
  AOI21_X1 U10690 ( .B1(n9612), .B2(n9772), .A(n9464), .ZN(n9474) );
  OAI211_X1 U10691 ( .C1(n9467), .C2(n9466), .A(n9465), .B(n9575), .ZN(n9470)
         );
  INV_X1 U10692 ( .A(n9468), .ZN(n9469) );
  NAND2_X1 U10693 ( .A1(n9470), .A2(n9469), .ZN(n9613) );
  NOR2_X1 U10694 ( .A1(n9471), .A2(n9754), .ZN(n9472) );
  OAI21_X1 U10695 ( .B1(n9613), .B2(n9472), .A(n9745), .ZN(n9473) );
  OAI211_X1 U10696 ( .C1(n9616), .C2(n9589), .A(n9474), .B(n9473), .ZN(
        P1_U3271) );
  OAI21_X1 U10697 ( .B1(n6509), .B2(n9495), .A(n9475), .ZN(n9476) );
  XNOR2_X1 U10698 ( .A(n9476), .B(n9479), .ZN(n9478) );
  AOI21_X1 U10699 ( .B1(n9478), .B2(n9575), .A(n9477), .ZN(n9621) );
  OR2_X1 U10700 ( .A1(n9480), .A2(n9479), .ZN(n9617) );
  NAND3_X1 U10701 ( .A1(n9617), .A2(n9481), .A3(n9763), .ZN(n9490) );
  OAI22_X1 U10702 ( .A1(n9568), .A2(n9483), .B1(n9482), .B2(n9754), .ZN(n9488)
         );
  OAI211_X1 U10703 ( .C1(n9484), .C2(n9486), .A(n6447), .B(n9485), .ZN(n9620)
         );
  NOR2_X1 U10704 ( .A1(n9620), .A2(n9760), .ZN(n9487) );
  AOI211_X1 U10705 ( .C1(n9769), .C2(n9618), .A(n9488), .B(n9487), .ZN(n9489)
         );
  OAI211_X1 U10706 ( .C1(n9778), .C2(n9621), .A(n9490), .B(n9489), .ZN(
        P1_U3272) );
  XOR2_X1 U10707 ( .A(n9495), .B(n9491), .Z(n9690) );
  INV_X1 U10708 ( .A(n9504), .ZN(n9492) );
  AOI211_X1 U10709 ( .C1(n9625), .C2(n9492), .A(n9579), .B(n9484), .ZN(n9624)
         );
  OAI22_X1 U10710 ( .A1(n9493), .A2(n9556), .B1(n10060), .B2(n9568), .ZN(n9494) );
  AOI21_X1 U10711 ( .B1(n9624), .B2(n9772), .A(n9494), .ZN(n9502) );
  XNOR2_X1 U10712 ( .A(n6509), .B(n9495), .ZN(n9498) );
  OAI21_X1 U10713 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9623) );
  NOR2_X1 U10714 ( .A1(n9754), .A2(n9499), .ZN(n9500) );
  OAI21_X1 U10715 ( .B1(n9623), .B2(n9500), .A(n9745), .ZN(n9501) );
  OAI211_X1 U10716 ( .C1(n9690), .C2(n9589), .A(n9502), .B(n9501), .ZN(
        P1_U3273) );
  XOR2_X1 U10717 ( .A(n9503), .B(n9510), .Z(n9694) );
  AOI211_X1 U10718 ( .C1(n9630), .C2(n9528), .A(n9579), .B(n9504), .ZN(n9628)
         );
  NOR2_X1 U10719 ( .A1(n9505), .A2(n9556), .ZN(n9509) );
  OAI22_X1 U10720 ( .A1(n9568), .A2(n9507), .B1(n9506), .B2(n9754), .ZN(n9508)
         );
  AOI211_X1 U10721 ( .C1(n9628), .C2(n9772), .A(n9509), .B(n9508), .ZN(n9517)
         );
  XNOR2_X1 U10722 ( .A(n9511), .B(n9510), .ZN(n9512) );
  NAND2_X1 U10723 ( .A1(n9512), .A2(n9575), .ZN(n9515) );
  INV_X1 U10724 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U10725 ( .A1(n9515), .A2(n9514), .ZN(n9629) );
  NAND2_X1 U10726 ( .A1(n9629), .A2(n9568), .ZN(n9516) );
  OAI211_X1 U10727 ( .C1(n9694), .C2(n9589), .A(n9517), .B(n9516), .ZN(
        P1_U3274) );
  NAND2_X1 U10728 ( .A1(n9542), .A2(n9518), .ZN(n9520) );
  XNOR2_X1 U10729 ( .A(n9520), .B(n9519), .ZN(n9522) );
  AOI21_X1 U10730 ( .B1(n9522), .B2(n9575), .A(n9521), .ZN(n9634) );
  XNOR2_X1 U10731 ( .A(n9524), .B(n9523), .ZN(n9699) );
  INV_X1 U10732 ( .A(n9699), .ZN(n9525) );
  NAND2_X1 U10733 ( .A1(n9525), .A2(n9763), .ZN(n9533) );
  OAI22_X1 U10734 ( .A1(n9568), .A2(n9527), .B1(n9526), .B2(n9754), .ZN(n9531)
         );
  OAI211_X1 U10735 ( .C1(n4394), .C2(n9529), .A(n6447), .B(n9528), .ZN(n9633)
         );
  NOR2_X1 U10736 ( .A1(n9633), .A2(n9760), .ZN(n9530) );
  AOI211_X1 U10737 ( .C1(n9769), .C2(n9697), .A(n9531), .B(n9530), .ZN(n9532)
         );
  OAI211_X1 U10738 ( .C1(n9778), .C2(n9634), .A(n9533), .B(n9532), .ZN(
        P1_U3275) );
  XNOR2_X1 U10739 ( .A(n9535), .B(n9534), .ZN(n9703) );
  INV_X1 U10740 ( .A(n9555), .ZN(n9536) );
  AOI211_X1 U10741 ( .C1(n9639), .C2(n9536), .A(n9579), .B(n4394), .ZN(n9637)
         );
  NOR2_X1 U10742 ( .A1(n9537), .A2(n9556), .ZN(n9541) );
  OAI22_X1 U10743 ( .A1(n9568), .A2(n9539), .B1(n9538), .B2(n9754), .ZN(n9540)
         );
  AOI211_X1 U10744 ( .C1(n9637), .C2(n9772), .A(n9541), .B(n9540), .ZN(n9551)
         );
  NAND2_X1 U10745 ( .A1(n9542), .A2(n9575), .ZN(n9549) );
  AOI21_X1 U10746 ( .B1(n9543), .B2(n9545), .A(n9544), .ZN(n9548) );
  INV_X1 U10747 ( .A(n9546), .ZN(n9547) );
  OAI21_X1 U10748 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(n9638) );
  NAND2_X1 U10749 ( .A1(n9638), .A2(n9568), .ZN(n9550) );
  OAI211_X1 U10750 ( .C1(n9703), .C2(n9589), .A(n9551), .B(n9550), .ZN(
        P1_U3276) );
  OAI21_X1 U10751 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9707) );
  AOI211_X1 U10752 ( .C1(n9644), .C2(n9580), .A(n9579), .B(n9555), .ZN(n9643)
         );
  NOR2_X1 U10753 ( .A1(n9557), .A2(n9556), .ZN(n9561) );
  OAI22_X1 U10754 ( .A1(n9568), .A2(n9559), .B1(n9558), .B2(n9754), .ZN(n9560)
         );
  AOI211_X1 U10755 ( .C1(n9643), .C2(n9772), .A(n9561), .B(n9560), .ZN(n9570)
         );
  OAI21_X1 U10756 ( .B1(n9563), .B2(n9562), .A(n9543), .ZN(n9564) );
  NAND2_X1 U10757 ( .A1(n9564), .A2(n9575), .ZN(n9567) );
  INV_X1 U10758 ( .A(n9565), .ZN(n9566) );
  NAND2_X1 U10759 ( .A1(n9567), .A2(n9566), .ZN(n9642) );
  NAND2_X1 U10760 ( .A1(n9642), .A2(n9568), .ZN(n9569) );
  OAI211_X1 U10761 ( .C1(n9707), .C2(n9589), .A(n9570), .B(n9569), .ZN(
        P1_U3277) );
  XNOR2_X1 U10762 ( .A(n9571), .B(n9573), .ZN(n9712) );
  NAND2_X1 U10763 ( .A1(n8059), .A2(n9572), .ZN(n9574) );
  XNOR2_X1 U10764 ( .A(n9574), .B(n9573), .ZN(n9576) );
  NAND2_X1 U10765 ( .A1(n9576), .A2(n9575), .ZN(n9578) );
  NAND2_X1 U10766 ( .A1(n9578), .A2(n9577), .ZN(n9650) );
  AOI21_X1 U10767 ( .B1(n8070), .B2(n9585), .A(n9579), .ZN(n9581) );
  NAND2_X1 U10768 ( .A1(n9581), .A2(n9580), .ZN(n9647) );
  OAI22_X1 U10769 ( .A1(n9745), .A2(n9583), .B1(n9582), .B2(n9754), .ZN(n9584)
         );
  AOI21_X1 U10770 ( .B1(n9585), .B2(n9769), .A(n9584), .ZN(n9586) );
  OAI21_X1 U10771 ( .B1(n9647), .B2(n9760), .A(n9586), .ZN(n9587) );
  AOI21_X1 U10772 ( .B1(n9650), .B2(n9745), .A(n9587), .ZN(n9588) );
  OAI21_X1 U10773 ( .B1(n9712), .B2(n9589), .A(n9588), .ZN(P1_U3278) );
  INV_X1 U10774 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9590) );
  OAI21_X1 U10775 ( .B1(n9593), .B2(n9659), .A(n9592), .ZN(P1_U3553) );
  NAND2_X1 U10776 ( .A1(n9595), .A2(n9594), .ZN(n9667) );
  MUX2_X1 U10777 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9667), .S(n9818), .Z(n9596) );
  AOI21_X1 U10778 ( .B1(n6535), .B2(n9669), .A(n9596), .ZN(n9597) );
  OAI21_X1 U10779 ( .B1(n9671), .B2(n9653), .A(n9597), .ZN(P1_U3548) );
  AOI211_X1 U10780 ( .C1(n9788), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9672)
         );
  MUX2_X1 U10781 ( .A(n9601), .B(n9672), .S(n9818), .Z(n9602) );
  OAI21_X1 U10782 ( .B1(n9675), .B2(n9653), .A(n9602), .ZN(P1_U3547) );
  NAND2_X1 U10783 ( .A1(n9604), .A2(n9603), .ZN(n9676) );
  MUX2_X1 U10784 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9676), .S(n9818), .Z(n9605) );
  AOI21_X1 U10785 ( .B1(n6535), .B2(n9678), .A(n9605), .ZN(n9606) );
  OAI21_X1 U10786 ( .B1(n9680), .B2(n9653), .A(n9606), .ZN(P1_U3546) );
  AOI211_X1 U10787 ( .C1(n9788), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9681)
         );
  MUX2_X1 U10788 ( .A(n9610), .B(n9681), .S(n9818), .Z(n9611) );
  OAI21_X1 U10789 ( .B1(n9684), .B2(n9653), .A(n9611), .ZN(P1_U3545) );
  AOI211_X1 U10790 ( .C1(n9788), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9615)
         );
  OAI21_X1 U10791 ( .B1(n9616), .B2(n9792), .A(n9615), .ZN(n9685) );
  MUX2_X1 U10792 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9685), .S(n9818), .Z(
        P1_U3544) );
  NAND3_X1 U10793 ( .A1(n9617), .A2(n9481), .A3(n9801), .ZN(n9622) );
  NAND2_X1 U10794 ( .A1(n9618), .A2(n9788), .ZN(n9619) );
  NAND4_X1 U10795 ( .A1(n9622), .A2(n9621), .A3(n9620), .A4(n9619), .ZN(n9686)
         );
  MUX2_X1 U10796 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9686), .S(n9818), .Z(
        P1_U3543) );
  INV_X1 U10797 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9626) );
  AOI211_X1 U10798 ( .C1(n9788), .C2(n9625), .A(n9624), .B(n9623), .ZN(n9687)
         );
  MUX2_X1 U10799 ( .A(n9626), .B(n9687), .S(n9818), .Z(n9627) );
  OAI21_X1 U10800 ( .B1(n9690), .B2(n9653), .A(n9627), .ZN(P1_U3542) );
  AOI211_X1 U10801 ( .C1(n9788), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9691)
         );
  MUX2_X1 U10802 ( .A(n9631), .B(n9691), .S(n9818), .Z(n9632) );
  OAI21_X1 U10803 ( .B1(n9694), .B2(n9653), .A(n9632), .ZN(P1_U3541) );
  NAND2_X1 U10804 ( .A1(n9634), .A2(n9633), .ZN(n9695) );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9695), .S(n9818), .Z(n9635) );
  AOI21_X1 U10806 ( .B1(n6535), .B2(n9697), .A(n9635), .ZN(n9636) );
  OAI21_X1 U10807 ( .B1(n9699), .B2(n9653), .A(n9636), .ZN(P1_U3540) );
  AOI211_X1 U10808 ( .C1(n9788), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9700)
         );
  MUX2_X1 U10809 ( .A(n9640), .B(n9700), .S(n9818), .Z(n9641) );
  OAI21_X1 U10810 ( .B1(n9703), .B2(n9653), .A(n9641), .ZN(P1_U3539) );
  AOI211_X1 U10811 ( .C1(n9788), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9704)
         );
  MUX2_X1 U10812 ( .A(n9645), .B(n9704), .S(n9818), .Z(n9646) );
  OAI21_X1 U10813 ( .B1(n9707), .B2(n9653), .A(n9646), .ZN(P1_U3538) );
  OAI21_X1 U10814 ( .B1(n9648), .B2(n9804), .A(n9647), .ZN(n9649) );
  NOR2_X1 U10815 ( .A1(n9650), .A2(n9649), .ZN(n9708) );
  MUX2_X1 U10816 ( .A(n9651), .B(n9708), .S(n9818), .Z(n9652) );
  OAI21_X1 U10817 ( .B1(n9712), .B2(n9653), .A(n9652), .ZN(P1_U3537) );
  OAI211_X1 U10818 ( .C1(n9656), .C2(n9792), .A(n9655), .B(n9654), .ZN(n9657)
         );
  INV_X1 U10819 ( .A(n9657), .ZN(n9714) );
  MUX2_X1 U10820 ( .A(n10041), .B(n9714), .S(n9818), .Z(n9658) );
  OAI21_X1 U10821 ( .B1(n9718), .B2(n9659), .A(n9658), .ZN(P1_U3536) );
  INV_X1 U10822 ( .A(n9660), .ZN(n9665) );
  AOI21_X1 U10823 ( .B1(n9788), .B2(n9662), .A(n9661), .ZN(n9663) );
  OAI211_X1 U10824 ( .C1(n9665), .C2(n9781), .A(n9664), .B(n9663), .ZN(n9719)
         );
  MUX2_X1 U10825 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9719), .S(n9818), .Z(
        P1_U3533) );
  MUX2_X1 U10826 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9666), .S(n9818), .Z(
        P1_U3522) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9667), .S(n9794), .Z(n9668) );
  AOI21_X1 U10828 ( .B1(n6528), .B2(n9669), .A(n9668), .ZN(n9670) );
  OAI21_X1 U10829 ( .B1(n9671), .B2(n9711), .A(n9670), .ZN(P1_U3516) );
  INV_X1 U10830 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9673) );
  MUX2_X1 U10831 ( .A(n9673), .B(n9672), .S(n9794), .Z(n9674) );
  OAI21_X1 U10832 ( .B1(n9675), .B2(n9711), .A(n9674), .ZN(P1_U3515) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9676), .S(n9794), .Z(n9677) );
  AOI21_X1 U10834 ( .B1(n6528), .B2(n9678), .A(n9677), .ZN(n9679) );
  OAI21_X1 U10835 ( .B1(n9680), .B2(n9711), .A(n9679), .ZN(P1_U3514) );
  INV_X1 U10836 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U10837 ( .A(n9682), .B(n9681), .S(n9794), .Z(n9683) );
  OAI21_X1 U10838 ( .B1(n9684), .B2(n9711), .A(n9683), .ZN(P1_U3513) );
  MUX2_X1 U10839 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9685), .S(n9713), .Z(
        P1_U3512) );
  MUX2_X1 U10840 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9686), .S(n9713), .Z(
        P1_U3511) );
  MUX2_X1 U10841 ( .A(n9688), .B(n9687), .S(n9794), .Z(n9689) );
  OAI21_X1 U10842 ( .B1(n9690), .B2(n9711), .A(n9689), .ZN(P1_U3510) );
  INV_X1 U10843 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9692) );
  MUX2_X1 U10844 ( .A(n9692), .B(n9691), .S(n9794), .Z(n9693) );
  OAI21_X1 U10845 ( .B1(n9694), .B2(n9711), .A(n9693), .ZN(P1_U3509) );
  MUX2_X1 U10846 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9695), .S(n9794), .Z(n9696) );
  AOI21_X1 U10847 ( .B1(n6528), .B2(n9697), .A(n9696), .ZN(n9698) );
  OAI21_X1 U10848 ( .B1(n9699), .B2(n9711), .A(n9698), .ZN(P1_U3507) );
  INV_X1 U10849 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9701) );
  MUX2_X1 U10850 ( .A(n9701), .B(n9700), .S(n9713), .Z(n9702) );
  OAI21_X1 U10851 ( .B1(n9703), .B2(n9711), .A(n9702), .ZN(P1_U3504) );
  INV_X1 U10852 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9705) );
  MUX2_X1 U10853 ( .A(n9705), .B(n9704), .S(n9713), .Z(n9706) );
  OAI21_X1 U10854 ( .B1(n9707), .B2(n9711), .A(n9706), .ZN(P1_U3501) );
  INV_X1 U10855 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9709) );
  MUX2_X1 U10856 ( .A(n9709), .B(n9708), .S(n9794), .Z(n9710) );
  OAI21_X1 U10857 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(P1_U3498) );
  MUX2_X1 U10858 ( .A(n9715), .B(n9714), .S(n9713), .Z(n9716) );
  OAI21_X1 U10859 ( .B1(n9718), .B2(n9717), .A(n9716), .ZN(P1_U3495) );
  MUX2_X1 U10860 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9719), .S(n9794), .Z(
        P1_U3486) );
  MUX2_X1 U10861 ( .A(n9720), .B(P1_D_REG_1__SCAN_IN), .S(n9780), .Z(P1_U3440)
         );
  MUX2_X1 U10862 ( .A(n9721), .B(P1_D_REG_0__SCAN_IN), .S(n9780), .Z(P1_U3439)
         );
  NOR4_X1 U10863 ( .A1(n4433), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4862), .A4(
        P1_U3086), .ZN(n9722) );
  AOI21_X1 U10864 ( .B1(n9723), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9722), .ZN(
        n9724) );
  OAI21_X1 U10865 ( .B1(n9725), .B2(n9732), .A(n9724), .ZN(P1_U3324) );
  OAI222_X1 U10866 ( .A1(n9728), .A2(n9727), .B1(P1_U3086), .B2(n9726), .C1(
        n10021), .C2(n9729), .ZN(P1_U3326) );
  OAI222_X1 U10867 ( .A1(n5672), .A2(P1_U3086), .B1(n9732), .B2(n9731), .C1(
        n9730), .C2(n9729), .ZN(P1_U3327) );
  MUX2_X1 U10868 ( .A(n9733), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10869 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10870 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10871 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9735), .A(n9734), .ZN(
        n9736) );
  XOR2_X1 U10872 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9736), .Z(n9742) );
  INV_X1 U10873 ( .A(n9737), .ZN(n9738) );
  AOI21_X1 U10874 ( .B1(n9739), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n9738), .ZN(
        n9740) );
  OAI21_X1 U10875 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(P1_U3243) );
  OAI22_X1 U10876 ( .A1(n9745), .A2(n9744), .B1(n9743), .B2(n9754), .ZN(n9746)
         );
  AOI21_X1 U10877 ( .B1(n9769), .B2(n9747), .A(n9746), .ZN(n9748) );
  OAI21_X1 U10878 ( .B1(n9749), .B2(n9760), .A(n9748), .ZN(n9750) );
  AOI21_X1 U10879 ( .B1(n9751), .B2(n9773), .A(n9750), .ZN(n9752) );
  OAI21_X1 U10880 ( .B1(n9778), .B2(n9753), .A(n9752), .ZN(P1_U3286) );
  OAI22_X1 U10881 ( .A1(n9745), .A2(n9756), .B1(n9755), .B2(n9754), .ZN(n9757)
         );
  AOI21_X1 U10882 ( .B1(n9769), .B2(n9758), .A(n9757), .ZN(n9759) );
  OAI21_X1 U10883 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(n9762) );
  AOI21_X1 U10884 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  OAI21_X1 U10885 ( .B1(n9778), .B2(n9766), .A(n9765), .ZN(P1_U3288) );
  AOI22_X1 U10886 ( .A1(n9767), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n9778), .ZN(n9776) );
  INV_X1 U10887 ( .A(n9768), .ZN(n9771) );
  AOI222_X1 U10888 ( .A1(n9774), .A2(n9773), .B1(n9772), .B2(n9771), .C1(n9770), .C2(n9769), .ZN(n9775) );
  OAI211_X1 U10889 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(
        P1_U3292) );
  AND2_X1 U10890 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9780), .ZN(P1_U3294) );
  AND2_X1 U10891 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9780), .ZN(P1_U3295) );
  AND2_X1 U10892 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9780), .ZN(P1_U3296) );
  AND2_X1 U10893 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9780), .ZN(P1_U3297) );
  INV_X1 U10894 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U10895 ( .A1(n9779), .A2(n10038), .ZN(P1_U3298) );
  AND2_X1 U10896 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9780), .ZN(P1_U3299) );
  AND2_X1 U10897 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9780), .ZN(P1_U3300) );
  AND2_X1 U10898 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9780), .ZN(P1_U3301) );
  AND2_X1 U10899 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9780), .ZN(P1_U3302) );
  AND2_X1 U10900 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9780), .ZN(P1_U3303) );
  AND2_X1 U10901 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9780), .ZN(P1_U3304) );
  INV_X1 U10902 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9994) );
  NOR2_X1 U10903 ( .A1(n9779), .A2(n9994), .ZN(P1_U3305) );
  INV_X1 U10904 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U10905 ( .A1(n9779), .A2(n10017), .ZN(P1_U3306) );
  AND2_X1 U10906 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9780), .ZN(P1_U3307) );
  AND2_X1 U10907 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9780), .ZN(P1_U3308) );
  INV_X1 U10908 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10084) );
  NOR2_X1 U10909 ( .A1(n9779), .A2(n10084), .ZN(P1_U3309) );
  AND2_X1 U10910 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9780), .ZN(P1_U3310) );
  AND2_X1 U10911 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9780), .ZN(P1_U3311) );
  AND2_X1 U10912 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9780), .ZN(P1_U3312) );
  INV_X1 U10913 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10914 ( .A1(n9779), .A2(n10049), .ZN(P1_U3313) );
  AND2_X1 U10915 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9780), .ZN(P1_U3314) );
  AND2_X1 U10916 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9780), .ZN(P1_U3315) );
  AND2_X1 U10917 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9780), .ZN(P1_U3316) );
  AND2_X1 U10918 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9780), .ZN(P1_U3317) );
  AND2_X1 U10919 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9780), .ZN(P1_U3318) );
  AND2_X1 U10920 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9780), .ZN(P1_U3319) );
  AND2_X1 U10921 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9780), .ZN(P1_U3320) );
  INV_X1 U10922 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U10923 ( .A1(n9779), .A2(n10039), .ZN(P1_U3321) );
  AND2_X1 U10924 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9780), .ZN(P1_U3322) );
  AND2_X1 U10925 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9780), .ZN(P1_U3323) );
  INV_X1 U10926 ( .A(n9781), .ZN(n9800) );
  OAI21_X1 U10927 ( .B1(n10097), .B2(n9804), .A(n9782), .ZN(n9784) );
  AOI211_X1 U10928 ( .C1(n9800), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9812)
         );
  AOI22_X1 U10929 ( .A1(n9794), .A2(n9812), .B1(n4902), .B2(n9809), .ZN(
        P1_U3459) );
  AOI21_X1 U10930 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  OAI211_X1 U10931 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9793)
         );
  INV_X1 U10932 ( .A(n9793), .ZN(n9813) );
  AOI22_X1 U10933 ( .A1(n9794), .A2(n9813), .B1(n4943), .B2(n9809), .ZN(
        P1_U3465) );
  OAI21_X1 U10934 ( .B1(n9796), .B2(n9804), .A(n9795), .ZN(n9798) );
  AOI211_X1 U10935 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9815)
         );
  AOI22_X1 U10936 ( .A1(n9713), .A2(n9815), .B1(n5033), .B2(n9809), .ZN(
        P1_U3477) );
  AND2_X1 U10937 ( .A1(n9802), .A2(n9801), .ZN(n9808) );
  OAI21_X1 U10938 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9806) );
  NOR3_X1 U10939 ( .A1(n9808), .A2(n9807), .A3(n9806), .ZN(n9817) );
  INV_X1 U10940 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9810) );
  AOI22_X1 U10941 ( .A1(n9713), .A2(n9817), .B1(n9810), .B2(n9809), .ZN(
        P1_U3480) );
  AOI22_X1 U10942 ( .A1(n9818), .A2(n9812), .B1(n9811), .B2(n9816), .ZN(
        P1_U3524) );
  AOI22_X1 U10943 ( .A1(n9818), .A2(n9813), .B1(n9990), .B2(n9816), .ZN(
        P1_U3526) );
  INV_X1 U10944 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10945 ( .A1(n9818), .A2(n9815), .B1(n9814), .B2(n9816), .ZN(
        P1_U3530) );
  AOI22_X1 U10946 ( .A1(n9818), .A2(n9817), .B1(n4541), .B2(n9816), .ZN(
        P1_U3531) );
  INV_X1 U10947 ( .A(n7182), .ZN(n9819) );
  AOI21_X1 U10948 ( .B1(n9827), .B2(n9820), .A(n9819), .ZN(n9842) );
  INV_X1 U10949 ( .A(n9842), .ZN(n9835) );
  OAI22_X1 U10950 ( .A1(n9841), .A2(n9823), .B1(n9822), .B2(n9821), .ZN(n9834)
         );
  AOI22_X1 U10951 ( .A1(n9826), .A2(n5704), .B1(n9825), .B2(n9824), .ZN(n9832)
         );
  XNOR2_X1 U10952 ( .A(n9828), .B(n9827), .ZN(n9830) );
  NAND2_X1 U10953 ( .A1(n9830), .A2(n9829), .ZN(n9831) );
  OAI211_X1 U10954 ( .C1(n9842), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9844)
         );
  AOI211_X1 U10955 ( .C1(n9836), .C2(n9835), .A(n9834), .B(n9844), .ZN(n9838)
         );
  AOI22_X1 U10956 ( .A1(n9839), .A2(n6715), .B1(n9838), .B2(n9837), .ZN(
        P2_U3231) );
  AOI22_X1 U10957 ( .A1(n9901), .A2(n5685), .B1(n9840), .B2(n9899), .ZN(
        P2_U3393) );
  OAI22_X1 U10958 ( .A1(n9842), .A2(n9874), .B1(n9841), .B2(n9886), .ZN(n9843)
         );
  NOR2_X1 U10959 ( .A1(n9844), .A2(n9843), .ZN(n9902) );
  AOI22_X1 U10960 ( .A1(n9901), .A2(n5715), .B1(n9902), .B2(n9899), .ZN(
        P2_U3396) );
  INV_X1 U10961 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9848) );
  OAI21_X1 U10962 ( .B1(n6839), .B2(n9886), .A(n9845), .ZN(n9846) );
  AOI21_X1 U10963 ( .B1(n9895), .B2(n9847), .A(n9846), .ZN(n9903) );
  AOI22_X1 U10964 ( .A1(n9901), .A2(n9848), .B1(n9903), .B2(n9899), .ZN(
        P2_U3399) );
  INV_X1 U10965 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9853) );
  NOR2_X1 U10966 ( .A1(n9849), .A2(n9886), .ZN(n9851) );
  AOI211_X1 U10967 ( .C1(n9895), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9905)
         );
  AOI22_X1 U10968 ( .A1(n9901), .A2(n9853), .B1(n9905), .B2(n9899), .ZN(
        P2_U3402) );
  INV_X1 U10969 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9858) );
  OAI21_X1 U10970 ( .B1(n9855), .B2(n9886), .A(n9854), .ZN(n9856) );
  AOI21_X1 U10971 ( .B1(n9857), .B2(n9895), .A(n9856), .ZN(n9906) );
  AOI22_X1 U10972 ( .A1(n9901), .A2(n9858), .B1(n9906), .B2(n9899), .ZN(
        P2_U3405) );
  INV_X1 U10973 ( .A(n9859), .ZN(n9863) );
  OAI21_X1 U10974 ( .B1(n9861), .B2(n9886), .A(n9860), .ZN(n9862) );
  AOI21_X1 U10975 ( .B1(n9863), .B2(n9895), .A(n9862), .ZN(n9907) );
  AOI22_X1 U10976 ( .A1(n9901), .A2(n5769), .B1(n9907), .B2(n9899), .ZN(
        P2_U3408) );
  INV_X1 U10977 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9868) );
  OAI22_X1 U10978 ( .A1(n9865), .A2(n9874), .B1(n9864), .B2(n9886), .ZN(n9866)
         );
  NOR2_X1 U10979 ( .A1(n9867), .A2(n9866), .ZN(n9908) );
  AOI22_X1 U10980 ( .A1(n9901), .A2(n9868), .B1(n9908), .B2(n9899), .ZN(
        P2_U3411) );
  INV_X1 U10981 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9873) );
  OAI21_X1 U10982 ( .B1(n9870), .B2(n9886), .A(n9869), .ZN(n9871) );
  AOI21_X1 U10983 ( .B1(n9895), .B2(n9872), .A(n9871), .ZN(n9909) );
  AOI22_X1 U10984 ( .A1(n9901), .A2(n9873), .B1(n9909), .B2(n9899), .ZN(
        P2_U3414) );
  INV_X1 U10985 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9879) );
  NOR2_X1 U10986 ( .A1(n9875), .A2(n9874), .ZN(n9877) );
  AOI211_X1 U10987 ( .C1(n9892), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9910)
         );
  AOI22_X1 U10988 ( .A1(n9901), .A2(n9879), .B1(n9910), .B2(n9899), .ZN(
        P2_U3417) );
  INV_X1 U10989 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9885) );
  INV_X1 U10990 ( .A(n9895), .ZN(n9880) );
  NOR2_X1 U10991 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  AOI211_X1 U10992 ( .C1(n9892), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9911)
         );
  AOI22_X1 U10993 ( .A1(n9901), .A2(n9885), .B1(n9911), .B2(n9899), .ZN(
        P2_U3420) );
  INV_X1 U10994 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U10995 ( .A1(n9887), .A2(n9886), .ZN(n9889) );
  AOI211_X1 U10996 ( .C1(n9895), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9912)
         );
  AOI22_X1 U10997 ( .A1(n9901), .A2(n9891), .B1(n9912), .B2(n9899), .ZN(
        P2_U3423) );
  INV_X1 U10998 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9900) );
  AND2_X1 U10999 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  AOI21_X1 U11000 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9897) );
  AND2_X1 U11001 ( .A1(n9898), .A2(n9897), .ZN(n9914) );
  AOI22_X1 U11002 ( .A1(n9901), .A2(n9900), .B1(n9914), .B2(n9899), .ZN(
        P2_U3426) );
  AOI22_X1 U11003 ( .A1(n9915), .A2(n9902), .B1(n6724), .B2(n9913), .ZN(
        P2_U3461) );
  AOI22_X1 U11004 ( .A1(n9915), .A2(n9903), .B1(n10082), .B2(n9913), .ZN(
        P2_U3462) );
  AOI22_X1 U11005 ( .A1(n9915), .A2(n9905), .B1(n9904), .B2(n9913), .ZN(
        P2_U3463) );
  AOI22_X1 U11006 ( .A1(n9915), .A2(n9906), .B1(n6849), .B2(n9913), .ZN(
        P2_U3464) );
  AOI22_X1 U11007 ( .A1(n9915), .A2(n9907), .B1(n6968), .B2(n9913), .ZN(
        P2_U3465) );
  AOI22_X1 U11008 ( .A1(n9915), .A2(n9908), .B1(n5783), .B2(n9913), .ZN(
        P2_U3466) );
  AOI22_X1 U11009 ( .A1(n9915), .A2(n9909), .B1(n5799), .B2(n9913), .ZN(
        P2_U3467) );
  AOI22_X1 U11010 ( .A1(n9915), .A2(n9910), .B1(n5828), .B2(n9913), .ZN(
        P2_U3468) );
  AOI22_X1 U11011 ( .A1(n9915), .A2(n9911), .B1(n5840), .B2(n9913), .ZN(
        P2_U3469) );
  AOI22_X1 U11012 ( .A1(n9915), .A2(n9912), .B1(n5855), .B2(n9913), .ZN(
        P2_U3470) );
  AOI22_X1 U11013 ( .A1(n9915), .A2(n9914), .B1(n7827), .B2(n9913), .ZN(
        P2_U3471) );
  OAI222_X1 U11014 ( .A1(n9920), .A2(n9919), .B1(n9920), .B2(n9918), .C1(n9917), .C2(n9916), .ZN(ADD_1068_U5) );
  XOR2_X1 U11015 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11016 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9924) );
  XNOR2_X1 U11017 ( .A(n9924), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11018 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(ADD_1068_U56) );
  OAI21_X1 U11019 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(ADD_1068_U57) );
  OAI21_X1 U11020 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(ADD_1068_U58) );
  OAI21_X1 U11021 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1068_U59) );
  OAI21_X1 U11022 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(ADD_1068_U60) );
  OAI21_X1 U11023 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(ADD_1068_U61) );
  OAI21_X1 U11024 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(ADD_1068_U62) );
  OAI21_X1 U11025 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(ADD_1068_U63) );
  NAND4_X1 U11026 ( .A1(keyinput54), .A2(keyinput34), .A3(keyinput63), .A4(
        keyinput4), .ZN(n9953) );
  NAND3_X1 U11027 ( .A1(keyinput22), .A2(keyinput37), .A3(keyinput32), .ZN(
        n9952) );
  NOR2_X1 U11028 ( .A1(keyinput9), .A2(keyinput62), .ZN(n9950) );
  NOR4_X1 U11029 ( .A1(keyinput30), .A2(keyinput5), .A3(keyinput29), .A4(
        keyinput41), .ZN(n9949) );
  NAND4_X1 U11030 ( .A1(keyinput43), .A2(keyinput51), .A3(n9950), .A4(n9949), 
        .ZN(n9951) );
  NOR4_X1 U11031 ( .A1(keyinput25), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(
        n10095) );
  NOR2_X1 U11032 ( .A1(keyinput56), .A2(keyinput48), .ZN(n9956) );
  INV_X1 U11033 ( .A(keyinput28), .ZN(n9954) );
  NOR4_X1 U11034 ( .A1(keyinput26), .A2(keyinput10), .A3(keyinput58), .A4(
        n9954), .ZN(n9955) );
  NAND4_X1 U11035 ( .A1(keyinput1), .A2(keyinput11), .A3(n9956), .A4(n9955), 
        .ZN(n9975) );
  NOR2_X1 U11036 ( .A1(keyinput45), .A2(keyinput50), .ZN(n9958) );
  NOR4_X1 U11037 ( .A1(keyinput59), .A2(keyinput18), .A3(keyinput44), .A4(
        keyinput16), .ZN(n9957) );
  NAND4_X1 U11038 ( .A1(keyinput13), .A2(keyinput61), .A3(n9958), .A4(n9957), 
        .ZN(n9974) );
  NOR3_X1 U11039 ( .A1(keyinput35), .A2(keyinput2), .A3(keyinput27), .ZN(n9964) );
  NAND2_X1 U11040 ( .A1(keyinput33), .A2(keyinput57), .ZN(n9959) );
  NOR3_X1 U11041 ( .A1(keyinput42), .A2(keyinput36), .A3(n9959), .ZN(n9963) );
  NAND3_X1 U11042 ( .A1(keyinput47), .A2(keyinput19), .A3(keyinput23), .ZN(
        n9961) );
  NAND3_X1 U11043 ( .A1(keyinput52), .A2(keyinput6), .A3(keyinput49), .ZN(
        n9960) );
  NOR4_X1 U11044 ( .A1(keyinput24), .A2(keyinput55), .A3(n9961), .A4(n9960), 
        .ZN(n9962) );
  NAND4_X1 U11045 ( .A1(keyinput60), .A2(n9964), .A3(n9963), .A4(n9962), .ZN(
        n9973) );
  NOR4_X1 U11046 ( .A1(keyinput8), .A2(keyinput46), .A3(keyinput17), .A4(
        keyinput21), .ZN(n9971) );
  INV_X1 U11047 ( .A(keyinput20), .ZN(n9965) );
  NOR3_X1 U11048 ( .A1(keyinput12), .A2(keyinput53), .A3(n9965), .ZN(n9970) );
  NAND3_X1 U11049 ( .A1(keyinput14), .A2(keyinput39), .A3(keyinput40), .ZN(
        n9968) );
  INV_X1 U11050 ( .A(keyinput38), .ZN(n9966) );
  NAND3_X1 U11051 ( .A1(keyinput3), .A2(keyinput0), .A3(n9966), .ZN(n9967) );
  NOR4_X1 U11052 ( .A1(keyinput31), .A2(keyinput7), .A3(n9968), .A4(n9967), 
        .ZN(n9969) );
  NAND4_X1 U11053 ( .A1(n9971), .A2(keyinput15), .A3(n9970), .A4(n9969), .ZN(
        n9972) );
  NOR4_X1 U11054 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n10094)
         );
  AOI22_X1 U11055 ( .A1(n9978), .A2(keyinput13), .B1(n9977), .B2(keyinput61), 
        .ZN(n9976) );
  OAI221_X1 U11056 ( .B1(n9978), .B2(keyinput13), .C1(n9977), .C2(keyinput61), 
        .A(n9976), .ZN(n9988) );
  INV_X1 U11057 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11058 ( .A1(n6810), .A2(keyinput45), .B1(keyinput50), .B2(n9980), 
        .ZN(n9979) );
  OAI221_X1 U11059 ( .B1(n6810), .B2(keyinput45), .C1(n9980), .C2(keyinput50), 
        .A(n9979), .ZN(n9987) );
  AOI22_X1 U11060 ( .A1(n9983), .A2(keyinput56), .B1(keyinput1), .B2(n9982), 
        .ZN(n9981) );
  OAI221_X1 U11061 ( .B1(n9983), .B2(keyinput56), .C1(n9982), .C2(keyinput1), 
        .A(n9981), .ZN(n9986) );
  AOI22_X1 U11062 ( .A1(n8597), .A2(keyinput11), .B1(n8798), .B2(keyinput48), 
        .ZN(n9984) );
  OAI221_X1 U11063 ( .B1(n8597), .B2(keyinput11), .C1(n8798), .C2(keyinput48), 
        .A(n9984), .ZN(n9985) );
  NOR4_X1 U11064 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n10031)
         );
  AOI22_X1 U11065 ( .A1(n9991), .A2(keyinput26), .B1(keyinput58), .B2(n9990), 
        .ZN(n9989) );
  OAI221_X1 U11066 ( .B1(n9991), .B2(keyinput26), .C1(n9990), .C2(keyinput58), 
        .A(n9989), .ZN(n10001) );
  AOI22_X1 U11067 ( .A1(n5740), .A2(keyinput28), .B1(n9993), .B2(keyinput10), 
        .ZN(n9992) );
  OAI221_X1 U11068 ( .B1(n5740), .B2(keyinput28), .C1(n9993), .C2(keyinput10), 
        .A(n9992), .ZN(n10000) );
  XNOR2_X1 U11069 ( .A(n9994), .B(keyinput44), .ZN(n9999) );
  XNOR2_X1 U11070 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput16), .ZN(n9997) );
  XNOR2_X1 U11071 ( .A(P1_REG1_REG_20__SCAN_IN), .B(keyinput18), .ZN(n9996) );
  XNOR2_X1 U11072 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput59), .ZN(n9995) );
  NAND3_X1 U11073 ( .A1(n9997), .A2(n9996), .A3(n9995), .ZN(n9998) );
  NOR4_X1 U11074 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10030) );
  INV_X1 U11075 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11076 ( .A1(n10004), .A2(keyinput32), .B1(n10003), .B2(keyinput25), 
        .ZN(n10002) );
  OAI221_X1 U11077 ( .B1(n10004), .B2(keyinput32), .C1(n10003), .C2(keyinput25), .A(n10002), .ZN(n10015) );
  AOI22_X1 U11078 ( .A1(n5410), .A2(keyinput63), .B1(keyinput4), .B2(n10006), 
        .ZN(n10005) );
  OAI221_X1 U11079 ( .B1(n5410), .B2(keyinput63), .C1(n10006), .C2(keyinput4), 
        .A(n10005), .ZN(n10014) );
  AOI22_X1 U11080 ( .A1(n10009), .A2(keyinput54), .B1(n10008), .B2(keyinput34), 
        .ZN(n10007) );
  OAI221_X1 U11081 ( .B1(n10009), .B2(keyinput54), .C1(n10008), .C2(keyinput34), .A(n10007), .ZN(n10013) );
  XNOR2_X1 U11082 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput22), .ZN(n10011)
         );
  XNOR2_X1 U11083 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput37), .ZN(n10010) );
  NAND2_X1 U11084 ( .A1(n10011), .A2(n10010), .ZN(n10012) );
  NOR4_X1 U11085 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(n10012), .ZN(
        n10029) );
  AOI22_X1 U11086 ( .A1(n10017), .A2(keyinput29), .B1(n5007), .B2(keyinput41), 
        .ZN(n10016) );
  OAI221_X1 U11087 ( .B1(n10017), .B2(keyinput29), .C1(n5007), .C2(keyinput41), 
        .A(n10016), .ZN(n10027) );
  AOI22_X1 U11088 ( .A1(n10019), .A2(keyinput9), .B1(n5685), .B2(keyinput62), 
        .ZN(n10018) );
  OAI221_X1 U11089 ( .B1(n10019), .B2(keyinput9), .C1(n5685), .C2(keyinput62), 
        .A(n10018), .ZN(n10026) );
  AOI22_X1 U11090 ( .A1(n9583), .A2(keyinput43), .B1(keyinput51), .B2(n10021), 
        .ZN(n10020) );
  OAI221_X1 U11091 ( .B1(n9583), .B2(keyinput43), .C1(n10021), .C2(keyinput51), 
        .A(n10020), .ZN(n10025) );
  XNOR2_X1 U11092 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput30), .ZN(n10023)
         );
  XNOR2_X1 U11093 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput5), .ZN(n10022) );
  NAND2_X1 U11094 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  NOR4_X1 U11095 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        n10028) );
  NAND4_X1 U11096 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10093) );
  AOI22_X1 U11097 ( .A1(n10034), .A2(keyinput49), .B1(keyinput55), .B2(n10033), 
        .ZN(n10032) );
  OAI221_X1 U11098 ( .B1(n10034), .B2(keyinput49), .C1(n10033), .C2(keyinput55), .A(n10032), .ZN(n10046) );
  AOI22_X1 U11099 ( .A1(n10036), .A2(keyinput52), .B1(keyinput6), .B2(n7624), 
        .ZN(n10035) );
  OAI221_X1 U11100 ( .B1(n10036), .B2(keyinput52), .C1(n7624), .C2(keyinput6), 
        .A(n10035), .ZN(n10045) );
  AOI22_X1 U11101 ( .A1(n10039), .A2(keyinput36), .B1(keyinput33), .B2(n10038), 
        .ZN(n10037) );
  OAI221_X1 U11102 ( .B1(n10039), .B2(keyinput36), .C1(n10038), .C2(keyinput33), .A(n10037), .ZN(n10044) );
  AOI22_X1 U11103 ( .A1(n10042), .A2(keyinput42), .B1(n10041), .B2(keyinput57), 
        .ZN(n10040) );
  OAI221_X1 U11104 ( .B1(n10042), .B2(keyinput42), .C1(n10041), .C2(keyinput57), .A(n10040), .ZN(n10043) );
  NOR4_X1 U11105 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10091) );
  AOI22_X1 U11106 ( .A1(n10049), .A2(keyinput19), .B1(keyinput23), .B2(n10048), 
        .ZN(n10047) );
  OAI221_X1 U11107 ( .B1(n10049), .B2(keyinput19), .C1(n10048), .C2(keyinput23), .A(n10047), .ZN(n10058) );
  AOI22_X1 U11108 ( .A1(n8809), .A2(keyinput24), .B1(n10051), .B2(keyinput47), 
        .ZN(n10050) );
  OAI221_X1 U11109 ( .B1(n8809), .B2(keyinput24), .C1(n10051), .C2(keyinput47), 
        .A(n10050), .ZN(n10057) );
  XNOR2_X1 U11110 ( .A(SI_19_), .B(keyinput27), .ZN(n10055) );
  XNOR2_X1 U11111 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput2), .ZN(n10054) );
  XNOR2_X1 U11112 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput60), .ZN(n10053)
         );
  XNOR2_X1 U11113 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput35), .ZN(n10052) );
  NAND4_X1 U11114 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10056) );
  NOR3_X1 U11115 ( .A1(n10058), .A2(n10057), .A3(n10056), .ZN(n10090) );
  AOI22_X1 U11116 ( .A1(n9507), .A2(keyinput12), .B1(n10060), .B2(keyinput53), 
        .ZN(n10059) );
  OAI221_X1 U11117 ( .B1(n9507), .B2(keyinput12), .C1(n10060), .C2(keyinput53), 
        .A(n10059), .ZN(n10065) );
  XNOR2_X1 U11118 ( .A(n10061), .B(keyinput38), .ZN(n10064) );
  XNOR2_X1 U11119 ( .A(n10062), .B(keyinput7), .ZN(n10063) );
  OR3_X1 U11120 ( .A1(n10065), .A2(n10064), .A3(n10063), .ZN(n10072) );
  AOI22_X1 U11121 ( .A1(n4854), .A2(keyinput0), .B1(keyinput3), .B2(n6545), 
        .ZN(n10066) );
  OAI221_X1 U11122 ( .B1(n4854), .B2(keyinput0), .C1(n6545), .C2(keyinput3), 
        .A(n10066), .ZN(n10071) );
  AOI22_X1 U11123 ( .A1(n10069), .A2(keyinput15), .B1(n10068), .B2(keyinput20), 
        .ZN(n10067) );
  OAI221_X1 U11124 ( .B1(n10069), .B2(keyinput15), .C1(n10068), .C2(keyinput20), .A(n10067), .ZN(n10070) );
  NOR3_X1 U11125 ( .A1(n10072), .A2(n10071), .A3(n10070), .ZN(n10089) );
  AOI22_X1 U11126 ( .A1(n10074), .A2(keyinput17), .B1(keyinput21), .B2(n6894), 
        .ZN(n10073) );
  OAI221_X1 U11127 ( .B1(n10074), .B2(keyinput17), .C1(n6894), .C2(keyinput21), 
        .A(n10073), .ZN(n10080) );
  INV_X1 U11128 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11129 ( .A1(n10077), .A2(keyinput39), .B1(n10076), .B2(keyinput40), 
        .ZN(n10075) );
  OAI221_X1 U11130 ( .B1(n10077), .B2(keyinput39), .C1(n10076), .C2(keyinput40), .A(n10075), .ZN(n10079) );
  XOR2_X1 U11131 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput14), .Z(n10078) );
  OR3_X1 U11132 ( .A1(n10080), .A2(n10079), .A3(n10078), .ZN(n10087) );
  AOI22_X1 U11133 ( .A1(n10083), .A2(keyinput8), .B1(keyinput46), .B2(n10082), 
        .ZN(n10081) );
  OAI221_X1 U11134 ( .B1(n10083), .B2(keyinput8), .C1(n10082), .C2(keyinput46), 
        .A(n10081), .ZN(n10086) );
  XNOR2_X1 U11135 ( .A(n10084), .B(keyinput31), .ZN(n10085) );
  NOR3_X1 U11136 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10088) );
  NAND4_X1 U11137 ( .A1(n10091), .A2(n10090), .A3(n10089), .A4(n10088), .ZN(
        n10092) );
  AOI211_X1 U11138 ( .C1(n10095), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        n10109) );
  OAI22_X1 U11139 ( .A1(n10099), .A2(n10098), .B1(n10097), .B2(n10096), .ZN(
        n10106) );
  AOI21_X1 U11140 ( .B1(n10102), .B2(n10101), .A(n10100), .ZN(n10104) );
  NOR2_X1 U11141 ( .A1(n10104), .A2(n10103), .ZN(n10105) );
  AOI211_X1 U11142 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n10107), .A(n10106), .B(
        n10105), .ZN(n10108) );
  XNOR2_X1 U11143 ( .A(n10109), .B(n10108), .ZN(P1_U3237) );
  OAI21_X1 U11144 ( .B1(n10112), .B2(n10111), .A(n10110), .ZN(ADD_1068_U50) );
  OAI21_X1 U11145 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(ADD_1068_U51) );
  OAI21_X1 U11146 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(ADD_1068_U47) );
  OAI21_X1 U11147 ( .B1(n10121), .B2(n10120), .A(n10119), .ZN(ADD_1068_U49) );
  OAI21_X1 U11148 ( .B1(n10124), .B2(n10123), .A(n10122), .ZN(ADD_1068_U48) );
  AOI21_X1 U11149 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(ADD_1068_U54) );
  AOI21_X1 U11150 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(ADD_1068_U53) );
  OAI21_X1 U11151 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(ADD_1068_U52) );
  INV_X1 U4811 ( .A(n5688), .ZN(n5686) );
  INV_X1 U4847 ( .A(n5827), .ZN(n8303) );
  INV_X1 U4867 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U4878 ( .A(n5684), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5687) );
  NAND2_X2 U5036 ( .A1(n4469), .A2(n4468), .ZN(n4907) );
  CLKBUF_X1 U7388 ( .A(n6127), .Z(n4316) );
endmodule

