

module b14_C_AntiSAT_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704;

  AND2_X1 U2293 ( .A1(n4115), .A2(n4125), .ZN(n4117) );
  CLKBUF_X1 U2294 ( .A(n2053), .Z(n2051) );
  CLKBUF_X1 U2295 ( .A(n2356), .Z(n2432) );
  CLKBUF_X2 U2296 ( .A(n2355), .Z(n2525) );
  INV_X2 U2297 ( .A(n2917), .ZN(n2897) );
  INV_X2 U2298 ( .A(n2909), .ZN(n2914) );
  NAND3_X1 U2299 ( .A1(n2178), .A2(n2353), .A3(n2170), .ZN(n2697) );
  NAND4_X1 U2300 ( .A1(n2363), .A2(n2362), .A3(n2361), .A4(n2360), .ZN(n2364)
         );
  XNOR2_X1 U2301 ( .A(n2221), .B(IR_REG_1__SCAN_IN), .ZN(n4425) );
  INV_X1 U2302 ( .A(n2354), .ZN(n2053) );
  XNOR2_X1 U2303 ( .A(n2333), .B(IR_REG_29__SCAN_IN), .ZN(n2357) );
  XNOR2_X1 U2304 ( .A(n2331), .B(IR_REG_30__SCAN_IN), .ZN(n2338) );
  NAND2_X1 U2305 ( .A1(n2169), .A2(IR_REG_31__SCAN_IN), .ZN(n2331) );
  NOR2_X2 U2306 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2184)
         );
  INV_X1 U2307 ( .A(n2913), .ZN(n2906) );
  NAND2_X1 U2308 ( .A1(n3348), .A2(n3801), .ZN(n3249) );
  INV_X1 U2309 ( .A(IR_REG_7__SCAN_IN), .ZN(n2212) );
  NAND2_X1 U2310 ( .A1(n3796), .A2(n3798), .ZN(n3330) );
  INV_X1 U2311 ( .A(n4188), .ZN(n4304) );
  INV_X2 U2312 ( .A(n2911), .ZN(n2942) );
  INV_X1 U2313 ( .A(n4203), .ZN(n4158) );
  CLKBUF_X2 U2314 ( .A(n2366), .Z(n3857) );
  NAND2_X1 U2315 ( .A1(n2219), .A2(n2180), .ZN(n2224) );
  NAND2_X1 U2317 ( .A1(n2274), .A2(IR_REG_31__SCAN_IN), .ZN(n2275) );
  NAND2_X2 U2318 ( .A1(n3126), .A2(n3132), .ZN(n2913) );
  NAND2_X2 U2319 ( .A1(n3131), .A2(n4225), .ZN(n4227) );
  INV_X1 U2320 ( .A(n2338), .ZN(n2359) );
  INV_X1 U2321 ( .A(n2913), .ZN(n2052) );
  NAND2_X1 U2322 ( .A1(n2372), .A2(n3332), .ZN(n3796) );
  AND2_X1 U2323 ( .A1(n2351), .A2(n2350), .ZN(n2178) );
  BUF_X4 U2324 ( .A(n2720), .Z(n2911) );
  INV_X1 U2325 ( .A(n4223), .ZN(n4200) );
  NOR2_X1 U2326 ( .A1(n3629), .A2(n2783), .ZN(n2152) );
  CLKBUF_X3 U2327 ( .A(n2393), .Z(n2586) );
  INV_X1 U2328 ( .A(n3671), .ZN(n2707) );
  NAND2_X1 U2329 ( .A1(n2334), .A2(n3153), .ZN(n2393) );
  NAND2_X1 U2330 ( .A1(n2089), .A2(n2088), .ZN(n2366) );
  NAND2_X1 U2331 ( .A1(n2063), .A2(IR_REG_31__SCAN_IN), .ZN(n2278) );
  OAI21_X1 U2332 ( .B1(n2279), .B2(n2100), .A(n2093), .ZN(n2092) );
  NAND2_X1 U2333 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2334 ( .A1(n2163), .A2(n2162), .ZN(n2161) );
  INV_X1 U2335 ( .A(n2094), .ZN(n2093) );
  OAI21_X1 U2336 ( .B1(n2100), .B2(IR_REG_31__SCAN_IN), .A(n2069), .ZN(n2094)
         );
  AND2_X1 U2337 ( .A1(n2080), .A2(n2183), .ZN(n2188) );
  AND4_X1 U2338 ( .A1(n2187), .A2(n2186), .A3(n2185), .A4(n2184), .ZN(n2194)
         );
  AND2_X1 U2339 ( .A1(n2227), .A2(n2181), .ZN(n2175) );
  INV_X1 U2340 ( .A(IR_REG_14__SCAN_IN), .ZN(n2198) );
  INV_X1 U2341 ( .A(IR_REG_15__SCAN_IN), .ZN(n2259) );
  INV_X1 U2342 ( .A(IR_REG_23__SCAN_IN), .ZN(n2277) );
  NOR2_X1 U2343 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2266)
         );
  INV_X1 U2344 ( .A(IR_REG_21__SCAN_IN), .ZN(n2166) );
  INV_X1 U2345 ( .A(IR_REG_3__SCAN_IN), .ZN(n2227) );
  NOR2_X1 U2346 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2187)
         );
  NOR2_X1 U2347 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2185)
         );
  NOR2_X1 U2348 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2186)
         );
  CLKBUF_X1 U2349 ( .A(n3448), .Z(n2054) );
  NAND2_X1 U2350 ( .A1(n2446), .A2(n2070), .ZN(n3534) );
  OAI21_X1 U2351 ( .B1(n2686), .B2(n3850), .A(n2640), .ZN(n2641) );
  OAI21_X2 U2352 ( .B1(n3362), .B2(n3361), .A(n3809), .ZN(n3389) );
  OAI21_X2 U2353 ( .B1(n3606), .B2(n3608), .A(n3607), .ZN(n3659) );
  NOR2_X2 U2354 ( .A1(n4056), .A2(n3792), .ZN(n2637) );
  OAI21_X2 U2355 ( .B1(n4070), .B2(n2635), .A(n3871), .ZN(n4056) );
  AOI21_X2 U2356 ( .B1(n4217), .B2(n2540), .A(n2173), .ZN(n4135) );
  NOR2_X2 U2357 ( .A1(n2559), .A2(n2558), .ZN(n4069) );
  OAI22_X1 U2359 ( .A1(n2684), .A2(n3901), .B1(n4014), .B2(n2916), .ZN(n2592)
         );
  NOR2_X2 U2360 ( .A1(n2637), .A2(n3852), .ZN(n4039) );
  INV_X1 U2361 ( .A(n2266), .ZN(n2162) );
  NAND2_X1 U2362 ( .A1(n2164), .A2(n2067), .ZN(n2163) );
  INV_X1 U2363 ( .A(IR_REG_17__SCAN_IN), .ZN(n2183) );
  INV_X1 U2364 ( .A(IR_REG_5__SCAN_IN), .ZN(n2137) );
  AND2_X1 U2365 ( .A1(n2566), .A2(REG3_REG_26__SCAN_IN), .ZN(n2570) );
  AND2_X1 U2366 ( .A1(n2570), .A2(REG3_REG_27__SCAN_IN), .ZN(n2578) );
  AND2_X1 U2367 ( .A1(n3280), .A2(n3277), .ZN(n3281) );
  NAND2_X1 U2369 ( .A1(n2123), .A2(n2122), .ZN(n2121) );
  INV_X1 U2370 ( .A(n4441), .ZN(n2122) );
  NAND2_X1 U2371 ( .A1(n4506), .A2(n4507), .ZN(n4505) );
  NOR2_X1 U2372 ( .A1(n3931), .A2(n3850), .ZN(n3901) );
  NOR3_X1 U2373 ( .A1(n4091), .A2(n4029), .A3(n2104), .ZN(n2692) );
  NAND2_X1 U2374 ( .A1(n4280), .A2(n2105), .ZN(n2104) );
  NOR2_X1 U2375 ( .A1(n4049), .A2(n4061), .ZN(n2105) );
  AND2_X1 U2376 ( .A1(n2083), .A2(n2271), .ZN(n2082) );
  INV_X1 U2377 ( .A(IR_REG_25__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2378 ( .A1(n3985), .A2(n2108), .ZN(n2290) );
  NAND2_X1 U2379 ( .A1(n2507), .A2(n2109), .ZN(n2108) );
  NOR2_X1 U2380 ( .A1(n2290), .A2(n2291), .ZN(n3994) );
  INV_X1 U2381 ( .A(n4234), .ZN(n4429) );
  OR2_X1 U2382 ( .A1(n2522), .A2(n2521), .ZN(n2533) );
  INV_X1 U2383 ( .A(n4172), .ZN(n2669) );
  AND2_X1 U2384 ( .A1(n3650), .A2(n3651), .ZN(n2871) );
  INV_X1 U2385 ( .A(n2157), .ZN(n2155) );
  INV_X1 U2386 ( .A(n2881), .ZN(n2154) );
  INV_X1 U2387 ( .A(n2871), .ZN(n2156) );
  NAND2_X1 U2388 ( .A1(IR_REG_28__SCAN_IN), .A2(n2101), .ZN(n2100) );
  NAND2_X1 U2389 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2101) );
  NOR2_X1 U2390 ( .A1(n2560), .A2(n3691), .ZN(n2566) );
  NAND2_X1 U2391 ( .A1(n3717), .A2(n3254), .ZN(n3805) );
  NAND2_X1 U2392 ( .A1(n4418), .A2(n2670), .ZN(n3132) );
  NAND2_X1 U2393 ( .A1(n3573), .A2(n3479), .ZN(n2103) );
  INV_X1 U2394 ( .A(IR_REG_18__SCAN_IN), .ZN(n2083) );
  INV_X1 U2395 ( .A(IR_REG_19__SCAN_IN), .ZN(n2593) );
  NOR2_X1 U2396 ( .A1(n3753), .A2(n2158), .ZN(n2157) );
  INV_X1 U2397 ( .A(n2860), .ZN(n2158) );
  OAI211_X1 U2398 ( .C1(n2140), .C2(n2911), .A(n2138), .B(n2726), .ZN(n2727)
         );
  NAND2_X1 U2399 ( .A1(n2141), .A2(n2942), .ZN(n2138) );
  AOI21_X1 U2400 ( .B1(n2697), .B2(n2942), .A(n2062), .ZN(n2703) );
  NAND2_X1 U2401 ( .A1(n2735), .A2(n2725), .ZN(n2736) );
  XNOR2_X1 U2402 ( .A(n2723), .B(n2914), .ZN(n2742) );
  INV_X1 U2403 ( .A(n2732), .ZN(n2733) );
  NAND2_X1 U2404 ( .A1(n3260), .A2(n2753), .ZN(n2144) );
  AND2_X1 U2405 ( .A1(n4417), .A2(n4418), .ZN(n2925) );
  AND2_X1 U2406 ( .A1(n2096), .A2(IR_REG_31__SCAN_IN), .ZN(n2095) );
  INV_X1 U2407 ( .A(IR_REG_27__SCAN_IN), .ZN(n2096) );
  INV_X1 U2408 ( .A(n2092), .ZN(n2089) );
  OR2_X1 U2409 ( .A1(n2600), .A2(n2917), .ZN(n2702) );
  OR2_X1 U2410 ( .A1(n3945), .A2(n4420), .ZN(n2939) );
  NAND2_X1 U2411 ( .A1(n2053), .A2(REG1_REG_1__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U2412 ( .A1(n2359), .A2(n2357), .ZN(n2354) );
  NAND2_X1 U2413 ( .A1(n4445), .A2(n2235), .ZN(n2236) );
  NAND2_X1 U2414 ( .A1(n4623), .A2(REG1_REG_5__SCAN_IN), .ZN(n2120) );
  NAND2_X1 U2415 ( .A1(n4468), .A2(n2238), .ZN(n2239) );
  XNOR2_X1 U2416 ( .A(n2117), .B(n4473), .ZN(n4475) );
  INV_X1 U2417 ( .A(n2301), .ZN(n2117) );
  NAND2_X1 U2418 ( .A1(n4486), .A2(n2241), .ZN(n2242) );
  NAND2_X1 U2419 ( .A1(n4505), .A2(n2306), .ZN(n2307) );
  NAND2_X1 U2420 ( .A1(n4518), .A2(n2246), .ZN(n3380) );
  NAND2_X1 U2421 ( .A1(n2126), .A2(n2076), .ZN(n2309) );
  NAND2_X1 U2422 ( .A1(n3373), .A2(n2127), .ZN(n2126) );
  INV_X1 U2423 ( .A(n3372), .ZN(n2127) );
  AOI21_X1 U2424 ( .B1(n4037), .B2(n2577), .A(n2576), .ZN(n2684) );
  AND2_X1 U2425 ( .A1(n3954), .A2(n4049), .ZN(n2576) );
  AND2_X1 U2426 ( .A1(n2579), .A2(n4019), .ZN(n4028) );
  OR2_X1 U2427 ( .A1(n2465), .A2(n3374), .ZN(n2482) );
  OR2_X1 U2428 ( .A1(n2440), .A2(n3442), .ZN(n2448) );
  INV_X1 U2429 ( .A(n3962), .ZN(n3533) );
  NOR2_X1 U2430 ( .A1(n3863), .A2(n2644), .ZN(n2645) );
  INV_X1 U2431 ( .A(n3901), .ZN(n2685) );
  NOR2_X1 U2432 ( .A1(n4120), .A2(n4110), .ZN(n4103) );
  OR2_X1 U2433 ( .A1(n2061), .A2(n4253), .ZN(n4344) );
  AND2_X1 U2434 ( .A1(n4426), .A2(n2925), .ZN(n4644) );
  NAND2_X1 U2435 ( .A1(n2086), .A2(n2098), .ZN(n2097) );
  INV_X1 U2436 ( .A(IR_REG_26__SCAN_IN), .ZN(n2098) );
  INV_X1 U2437 ( .A(n2279), .ZN(n2086) );
  NOR2_X1 U2438 ( .A1(n2946), .A2(n4426), .ZN(n3690) );
  NAND4_X1 U2439 ( .A1(n2436), .A2(n2435), .A3(n2434), .A4(n2433), .ZN(n3483)
         );
  AND2_X1 U2440 ( .A1(n2321), .A2(n2320), .ZN(n4436) );
  XNOR2_X1 U2441 ( .A(n2236), .B(n4622), .ZN(n4457) );
  NAND2_X1 U2442 ( .A1(n4457), .A2(REG2_REG_6__SCAN_IN), .ZN(n4456) );
  XNOR2_X1 U2443 ( .A(n2242), .B(n2115), .ZN(n4499) );
  NAND2_X1 U2444 ( .A1(n4499), .A2(REG2_REG_10__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U2445 ( .A1(n4509), .A2(n4510), .ZN(n4508) );
  XNOR2_X1 U2446 ( .A(n2307), .B(n2119), .ZN(n4525) );
  XNOR2_X1 U2447 ( .A(n2309), .B(n2125), .ZN(n4535) );
  NAND2_X1 U2448 ( .A1(n2132), .A2(n2133), .ZN(n3997) );
  NOR2_X1 U2449 ( .A1(n3981), .A2(n2316), .ZN(n2318) );
  OR2_X1 U2450 ( .A1(n3994), .A2(n2078), .ZN(n2107) );
  OAI21_X1 U2451 ( .B1(n2130), .B2(n2129), .A(n2128), .ZN(n4000) );
  INV_X1 U2452 ( .A(n2133), .ZN(n2129) );
  INV_X1 U2453 ( .A(n4519), .ZN(n4548) );
  AND4_X1 U2454 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n3621)
         );
  NAND2_X1 U2455 ( .A1(n4227), .A2(n3141), .ZN(n4234) );
  OR2_X1 U2456 ( .A1(n2692), .A2(n2691), .ZN(n4027) );
  INV_X1 U2457 ( .A(IR_REG_29__SCAN_IN), .ZN(n2167) );
  XNOR2_X1 U2458 ( .A(n2594), .B(IR_REG_19__SCAN_IN), .ZN(n4420) );
  CLKBUF_X1 U2459 ( .A(n2601), .Z(n3795) );
  INV_X1 U2460 ( .A(IR_REG_24__SCAN_IN), .ZN(n2268) );
  INV_X1 U2461 ( .A(n2165), .ZN(n2164) );
  INV_X1 U2462 ( .A(IR_REG_6__SCAN_IN), .ZN(n2210) );
  INV_X1 U2463 ( .A(IR_REG_8__SCAN_IN), .ZN(n3040) );
  INV_X1 U2464 ( .A(n3546), .ZN(n2159) );
  NOR2_X1 U2465 ( .A1(n3547), .A2(n3546), .ZN(n2160) );
  NAND2_X1 U2466 ( .A1(n2356), .A2(REG0_REG_1__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U2467 ( .A1(n4508), .A2(n2176), .ZN(n2245) );
  AND2_X1 U2468 ( .A1(n4041), .A2(n2916), .ZN(n3850) );
  AND2_X1 U2469 ( .A1(n4014), .A2(n4029), .ZN(n3931) );
  OR2_X1 U2470 ( .A1(n2536), .A2(n2534), .ZN(n2535) );
  NOR2_X1 U2471 ( .A1(n2528), .A2(n2336), .ZN(n2541) );
  OR2_X1 U2472 ( .A1(n4211), .A2(n4212), .ZN(n4209) );
  AND2_X1 U2473 ( .A1(n3827), .A2(n3835), .ZN(n3134) );
  INV_X1 U2474 ( .A(n3450), .ZN(n3457) );
  AND2_X1 U2475 ( .A1(n3421), .A2(n3254), .ZN(n2081) );
  NAND2_X1 U2476 ( .A1(n2267), .A2(n2166), .ZN(n2165) );
  INV_X1 U2477 ( .A(IR_REG_16__SCAN_IN), .ZN(n2182) );
  CLKBUF_X1 U2478 ( .A(n2192), .Z(n2193) );
  AND2_X1 U2479 ( .A1(n2057), .A2(n2901), .ZN(n2147) );
  NAND2_X1 U2480 ( .A1(n2149), .A2(n2057), .ZN(n2146) );
  OAI21_X1 U2481 ( .B1(n2861), .B2(n2156), .A(n2153), .ZN(n2884) );
  AOI21_X1 U2482 ( .B1(n2871), .B2(n2155), .A(n2154), .ZN(n2153) );
  OR2_X1 U2483 ( .A1(n2552), .A2(n3735), .ZN(n2560) );
  OR2_X1 U2484 ( .A1(n2943), .A2(n3949), .ZN(n2946) );
  OR2_X1 U2485 ( .A1(n2578), .A2(n2571), .ZN(n3642) );
  NAND2_X1 U2486 ( .A1(n2355), .A2(REG2_REG_3__SCAN_IN), .ZN(n2376) );
  OAI21_X1 U2487 ( .B1(n2586), .B2(REG3_REG_3__SCAN_IN), .A(n2375), .ZN(n2142)
         );
  NAND2_X1 U2488 ( .A1(n3238), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2489 ( .A1(n4475), .A2(REG1_REG_8__SCAN_IN), .ZN(n4474) );
  NAND2_X1 U2490 ( .A1(n4476), .A2(n2240), .ZN(n4488) );
  NAND2_X1 U2491 ( .A1(n4496), .A2(n2305), .ZN(n4506) );
  XNOR2_X1 U2492 ( .A(n2245), .B(n2119), .ZN(n4520) );
  NAND2_X1 U2493 ( .A1(n4520), .A2(REG2_REG_12__SCAN_IN), .ZN(n4518) );
  OR2_X1 U2494 ( .A1(n2206), .A2(IR_REG_9__SCAN_IN), .ZN(n2251) );
  XNOR2_X1 U2495 ( .A(n2110), .B(n2479), .ZN(n4529) );
  NOR2_X1 U2496 ( .A1(n4529), .A2(n4530), .ZN(n4528) );
  NAND2_X1 U2497 ( .A1(n4542), .A2(n2311), .ZN(n2312) );
  NAND2_X1 U2498 ( .A1(n2130), .A2(n2131), .ZN(n2132) );
  NOR2_X1 U2499 ( .A1(n2134), .A2(n2316), .ZN(n2133) );
  INV_X1 U2500 ( .A(n2319), .ZN(n2134) );
  AOI21_X1 U2501 ( .B1(n3982), .B2(n2133), .A(n2079), .ZN(n2128) );
  NAND2_X1 U2502 ( .A1(n2692), .A2(n3849), .ZN(n4263) );
  XOR2_X1 U2503 ( .A(n3849), .B(n3953), .Z(n3902) );
  AND2_X1 U2504 ( .A1(n2638), .A2(n2639), .ZN(n4038) );
  OAI22_X2 U2505 ( .A1(n4098), .A2(n2557), .B1(n3736), .B2(n4291), .ZN(n4083)
         );
  AND2_X1 U2506 ( .A1(n2541), .A2(REG3_REG_21__SCAN_IN), .ZN(n2543) );
  INV_X1 U2507 ( .A(n3918), .ZN(n2629) );
  NOR2_X1 U2508 ( .A1(n3836), .A2(n4154), .ZN(n2630) );
  AND2_X1 U2509 ( .A1(n4181), .A2(n4182), .ZN(n4212) );
  NAND2_X1 U2510 ( .A1(n2500), .A2(REG3_REG_17__SCAN_IN), .ZN(n2526) );
  OR2_X1 U2511 ( .A1(n2526), .A2(n3027), .ZN(n2528) );
  INV_X1 U2512 ( .A(n3701), .ZN(n3140) );
  NOR2_X1 U2513 ( .A1(n2482), .A2(n2335), .ZN(n2493) );
  AND4_X1 U2514 ( .A1(n2505), .A2(n2504), .A3(n2503), .A4(n2502), .ZN(n4205)
         );
  CLKBUF_X1 U2515 ( .A(n3584), .Z(n3585) );
  NAND2_X1 U2516 ( .A1(n2618), .A2(n3829), .ZN(n4240) );
  AND4_X1 U2517 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n4244)
         );
  NOR2_X1 U2518 ( .A1(n2448), .A2(n3634), .ZN(n2458) );
  INV_X1 U2519 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3634) );
  CLKBUF_X1 U2520 ( .A(n3516), .Z(n3517) );
  OR2_X1 U2521 ( .A1(n3963), .A2(n3450), .ZN(n2427) );
  AND4_X1 U2522 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n3452)
         );
  INV_X1 U2523 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2410) );
  NOR2_X1 U2524 ( .A1(n2411), .A2(n2410), .ZN(n2421) );
  INV_X1 U2525 ( .A(n4567), .ZN(n4241) );
  NAND2_X1 U2526 ( .A1(n3812), .A2(n3814), .ZN(n3908) );
  OR2_X1 U2527 ( .A1(n3365), .A2(n3390), .ZN(n3405) );
  NOR2_X1 U2528 ( .A1(n3405), .A2(n3409), .ZN(n3458) );
  AND3_X1 U2529 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2399) );
  CLKBUF_X1 U2530 ( .A(n3247), .Z(n3248) );
  NOR2_X1 U2531 ( .A1(n3339), .A2(n4643), .ZN(n3351) );
  AND4_X1 U2532 ( .A1(n2367), .A2(n2370), .A3(n2368), .A4(n2369), .ZN(n2372)
         );
  CLKBUF_X1 U2533 ( .A(n3328), .Z(n3329) );
  INV_X1 U2534 ( .A(n3330), .ZN(n3874) );
  NOR2_X1 U2535 ( .A1(n4263), .A2(n4266), .ZN(n4262) );
  INV_X1 U2536 ( .A(n3935), .ZN(n4266) );
  NOR2_X1 U2537 ( .A1(n2106), .A2(n4049), .ZN(n4044) );
  INV_X1 U2538 ( .A(n4062), .ZN(n2106) );
  NOR3_X1 U2539 ( .A1(n4091), .A2(n4078), .A3(n4061), .ZN(n4062) );
  NAND2_X1 U2540 ( .A1(n3856), .A2(DATAI_24_), .ZN(n4092) );
  NAND2_X1 U2541 ( .A1(n4197), .A2(n2077), .ZN(n4120) );
  NAND2_X1 U2542 ( .A1(n4197), .A2(n2059), .ZN(n4142) );
  NAND2_X1 U2543 ( .A1(n4197), .A2(n2058), .ZN(n4310) );
  OR2_X1 U2544 ( .A1(n4328), .A2(n4231), .ZN(n4223) );
  AND4_X1 U2545 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n4323)
         );
  NOR2_X1 U2546 ( .A1(n4344), .A2(n3782), .ZN(n3593) );
  NAND2_X1 U2547 ( .A1(n2786), .A2(n2800), .ZN(n2102) );
  NOR3_X1 U2548 ( .A1(n3491), .A2(n3633), .A3(n3490), .ZN(n3540) );
  INV_X1 U2549 ( .A(n3620), .ZN(n3573) );
  NOR2_X1 U2550 ( .A1(n3491), .A2(n3490), .ZN(n4677) );
  OR2_X1 U2551 ( .A1(n3459), .A2(n3473), .ZN(n3491) );
  NAND2_X1 U2552 ( .A1(n3351), .A2(n3254), .ZN(n3366) );
  INV_X1 U2553 ( .A(n3714), .ZN(n3421) );
  OR2_X1 U2554 ( .A1(n2393), .A2(n3290), .ZN(n2379) );
  INV_X1 U2555 ( .A(n4644), .ZN(n4336) );
  NAND2_X1 U2556 ( .A1(n4248), .A2(n4347), .ZN(n4664) );
  INV_X1 U2557 ( .A(n4334), .ZN(n4642) );
  INV_X1 U2558 ( .A(n4674), .ZN(n4667) );
  NAND2_X1 U2559 ( .A1(n4562), .A2(n2707), .ZN(n3298) );
  AND2_X1 U2560 ( .A1(n2665), .A2(n3129), .ZN(n2677) );
  INV_X1 U2561 ( .A(n2161), .ZN(n2084) );
  AND2_X1 U2562 ( .A1(n2284), .A2(n2329), .ZN(n2168) );
  XNOR2_X1 U2563 ( .A(n2282), .B(n2166), .ZN(n2653) );
  XNOR2_X1 U2564 ( .A(n2597), .B(n2596), .ZN(n2670) );
  INV_X1 U2565 ( .A(IR_REG_20__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U2566 ( .A1(n2085), .A2(IR_REG_31__SCAN_IN), .ZN(n2594) );
  INV_X1 U2567 ( .A(n4291), .ZN(n4110) );
  CLKBUF_X1 U2568 ( .A(n3659), .Z(n3660) );
  MUX2_X1 U2569 ( .A(n4473), .B(DATAI_8_), .S(n3857), .Z(n3450) );
  NAND2_X1 U2570 ( .A1(n2737), .A2(n2736), .ZN(n2738) );
  INV_X1 U2571 ( .A(n4322), .ZN(n4231) );
  AND2_X1 U2572 ( .A1(n2758), .A2(n2764), .ZN(n2143) );
  AND2_X1 U2573 ( .A1(n2931), .A2(n2930), .ZN(n3710) );
  NAND2_X1 U2574 ( .A1(n2090), .A2(n2087), .ZN(n3296) );
  AOI22_X1 U2575 ( .A1(n2092), .A2(DATAI_0_), .B1(n2097), .B2(n2091), .ZN(
        n2090) );
  AND2_X1 U2576 ( .A1(n2095), .A2(DATAI_0_), .ZN(n2091) );
  NAND2_X1 U2577 ( .A1(n2861), .A2(n2860), .ZN(n3752) );
  OAI21_X1 U2578 ( .B1(n2945), .B2(n4334), .A(n4225), .ZN(n3733) );
  INV_X1 U2579 ( .A(n3784), .ZN(n3772) );
  INV_X1 U2580 ( .A(n2636), .ZN(n4061) );
  MUX2_X1 U2581 ( .A(n4611), .B(DATAI_15_), .S(n3856), .Z(n3782) );
  CLKBUF_X1 U2582 ( .A(n3733), .Z(n3781) );
  BUF_X1 U2583 ( .A(n3690), .Z(n3780) );
  XNOR2_X1 U2584 ( .A(n2280), .B(n2267), .ZN(n3945) );
  INV_X1 U2585 ( .A(n4292), .ZN(n4139) );
  NAND4_X1 U2586 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2544), .ZN(n4156)
         );
  INV_X1 U2587 ( .A(n4323), .ZN(n3779) );
  NAND4_X1 U2588 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n4242)
         );
  INV_X1 U2589 ( .A(n4337), .ZN(n3786) );
  INV_X1 U2590 ( .A(n4244), .ZN(n3959) );
  NAND4_X1 U2591 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n3632)
         );
  OR2_X1 U2592 ( .A1(n2586), .A2(n3523), .ZN(n2462) );
  NAND4_X1 U2593 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n3962)
         );
  INV_X1 U2594 ( .A(n3452), .ZN(n3964) );
  NAND2_X1 U2595 ( .A1(n2396), .A2(n2395), .ZN(n3965) );
  CLKBUF_X1 U2596 ( .A(n2364), .Z(n3172) );
  OR2_X1 U2597 ( .A1(n2354), .A2(n4686), .ZN(n2170) );
  NAND2_X1 U2598 ( .A1(n2352), .A2(REG3_REG_0__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U2599 ( .A1(n4456), .A2(n2237), .ZN(n4469) );
  XNOR2_X1 U2600 ( .A(n2239), .B(n2114), .ZN(n4477) );
  NAND2_X1 U2601 ( .A1(n4477), .A2(REG2_REG_8__SCAN_IN), .ZN(n4476) );
  INV_X1 U2602 ( .A(n2302), .ZN(n2118) );
  AOI21_X1 U2603 ( .B1(n2302), .B2(n2420), .A(n2293), .ZN(n2116) );
  NAND2_X1 U2604 ( .A1(n4474), .A2(n2302), .ZN(n4485) );
  NAND2_X1 U2605 ( .A1(n4498), .A2(n2243), .ZN(n4509) );
  AND2_X1 U2606 ( .A1(n4436), .A2(n2289), .ZN(n4519) );
  NAND2_X1 U2607 ( .A1(n4524), .A2(n2308), .ZN(n3373) );
  NAND2_X1 U2608 ( .A1(n4534), .A2(n2310), .ZN(n4543) );
  NAND2_X1 U2609 ( .A1(n4543), .A2(n4544), .ZN(n4542) );
  OAI21_X1 U2610 ( .B1(n4529), .B2(n2112), .A(n2111), .ZN(n4538) );
  NAND2_X1 U2611 ( .A1(n2113), .A2(REG2_REG_14__SCAN_IN), .ZN(n2112) );
  NAND2_X1 U2612 ( .A1(n2257), .A2(n2113), .ZN(n2111) );
  INV_X1 U2613 ( .A(n4539), .ZN(n2113) );
  XNOR2_X1 U2614 ( .A(n2312), .B(n2499), .ZN(n4556) );
  INV_X1 U2615 ( .A(n2132), .ZN(n3981) );
  CLKBUF_X1 U2616 ( .A(n4017), .Z(n4018) );
  NAND2_X1 U2617 ( .A1(n3593), .A2(n3140), .ZN(n4328) );
  AND2_X1 U2618 ( .A1(n3489), .A2(n3488), .ZN(n4682) );
  OR2_X1 U2619 ( .A1(n3158), .A2(n2944), .ZN(n4225) );
  NAND2_X1 U2620 ( .A1(n4685), .A2(n4674), .ZN(n4633) );
  XNOR2_X1 U2621 ( .A(n2287), .B(IR_REG_28__SCAN_IN), .ZN(n4426) );
  AND2_X1 U2622 ( .A1(n2285), .A2(n2284), .ZN(n2330) );
  NAND2_X1 U2623 ( .A1(n2097), .A2(IR_REG_31__SCAN_IN), .ZN(n2288) );
  XNOR2_X1 U2624 ( .A(n2276), .B(IR_REG_26__SCAN_IN), .ZN(n4415) );
  AND2_X1 U2625 ( .A1(n2937), .A2(STATE_REG_SCAN_IN), .ZN(n4605) );
  INV_X1 U2626 ( .A(n2653), .ZN(n4418) );
  INV_X1 U2627 ( .A(n2224), .ZN(n2135) );
  OR2_X1 U2628 ( .A1(n2328), .A2(n2327), .ZN(U3258) );
  NAND2_X1 U2629 ( .A1(n2326), .A2(n2325), .ZN(n2327) );
  XNOR2_X1 U2630 ( .A(n2107), .B(n3996), .ZN(n4007) );
  AOI211_X1 U2631 ( .C1(n4429), .C2(n4035), .A(n4034), .B(n4033), .ZN(n4036)
         );
  AND2_X1 U2632 ( .A1(n2674), .A2(n2673), .ZN(n2675) );
  NAND2_X1 U2633 ( .A1(n3965), .A2(n3714), .ZN(n2055) );
  AND2_X1 U2634 ( .A1(n2168), .A2(n2167), .ZN(n2056) );
  AOI21_X1 U2635 ( .B1(n2798), .B2(n2072), .A(n2177), .ZN(n3507) );
  AND2_X1 U2636 ( .A1(n2933), .A2(n2932), .ZN(n2057) );
  INV_X1 U2637 ( .A(n2800), .ZN(n3566) );
  AND2_X1 U2638 ( .A1(n4191), .A2(n2669), .ZN(n2058) );
  AND2_X1 U2639 ( .A1(n2058), .A2(n4303), .ZN(n2059) );
  INV_X1 U2640 ( .A(n2479), .ZN(n2125) );
  INV_X1 U2641 ( .A(n3982), .ZN(n2131) );
  AND2_X1 U2642 ( .A1(n2121), .A2(n2120), .ZN(n2060) );
  OR3_X1 U2643 ( .A1(n3491), .A2(n2103), .A3(n2102), .ZN(n2061) );
  AND2_X1 U2644 ( .A1(n3296), .A2(n2052), .ZN(n2062) );
  NAND2_X1 U2645 ( .A1(n2151), .A2(n3763), .ZN(n3640) );
  OR2_X1 U2646 ( .A1(n2281), .A2(n2165), .ZN(n2063) );
  NOR2_X1 U2647 ( .A1(n2085), .A2(n2084), .ZN(n2272) );
  OR2_X1 U2648 ( .A1(n2281), .A2(IR_REG_21__SCAN_IN), .ZN(n2064) );
  NOR2_X1 U2649 ( .A1(n4528), .A2(n2257), .ZN(n2065) );
  NAND2_X1 U2650 ( .A1(n2135), .A2(n2175), .ZN(n2217) );
  NAND2_X1 U2651 ( .A1(n3688), .A2(n3687), .ZN(n3761) );
  NOR2_X1 U2652 ( .A1(n2393), .A2(n3715), .ZN(n2066) );
  AND2_X1 U2653 ( .A1(n2277), .A2(n2268), .ZN(n2067) );
  NOR2_X1 U2654 ( .A1(n2782), .A2(n2781), .ZN(n2783) );
  AND2_X1 U2655 ( .A1(n2151), .A2(n2148), .ZN(n2068) );
  NAND2_X1 U2656 ( .A1(n2329), .A2(IR_REG_27__SCAN_IN), .ZN(n2069) );
  INV_X1 U2657 ( .A(n2141), .ZN(n2139) );
  OAI21_X1 U2658 ( .B1(n2398), .B2(n2374), .A(n2376), .ZN(n2141) );
  INV_X1 U2659 ( .A(IR_REG_28__SCAN_IN), .ZN(n2329) );
  NAND2_X1 U2660 ( .A1(n3962), .A2(n3490), .ZN(n2070) );
  NAND2_X1 U2661 ( .A1(n4197), .A2(n4191), .ZN(n2071) );
  MUX2_X1 U2662 ( .A(n4495), .B(DATAI_10_), .S(n3856), .Z(n3490) );
  NAND2_X1 U2663 ( .A1(n3617), .A2(n3616), .ZN(n2072) );
  OR2_X1 U2664 ( .A1(n2951), .A2(n2950), .ZN(n2073) );
  OR2_X1 U2665 ( .A1(n4091), .A2(n4078), .ZN(n2074) );
  INV_X1 U2666 ( .A(n3633), .ZN(n2786) );
  INV_X1 U2667 ( .A(n2149), .ZN(n2148) );
  OR2_X1 U2668 ( .A1(n3641), .A2(n2150), .ZN(n2149) );
  INV_X1 U2669 ( .A(n3763), .ZN(n2150) );
  NAND2_X1 U2670 ( .A1(n2189), .A2(n2192), .ZN(n2265) );
  NAND2_X1 U2671 ( .A1(n2144), .A2(n2758), .ZN(n3267) );
  NAND2_X1 U2672 ( .A1(n3439), .A2(n2784), .ZN(n3627) );
  NAND2_X1 U2673 ( .A1(n3856), .A2(DATAI_21_), .ZN(n4303) );
  INV_X1 U2674 ( .A(n3163), .ZN(n2652) );
  OR3_X1 U2675 ( .A1(n3491), .A2(n2103), .A3(n3633), .ZN(n2075) );
  OR2_X1 U2676 ( .A1(n3377), .A2(n4352), .ZN(n2076) );
  AND2_X1 U2677 ( .A1(n3856), .A2(DATAI_22_), .ZN(n4118) );
  AND2_X1 U2678 ( .A1(n2059), .A2(n4130), .ZN(n2077) );
  AND2_X1 U2679 ( .A1(n3856), .A2(DATAI_28_), .ZN(n4029) );
  INV_X1 U2680 ( .A(n4280), .ZN(n4078) );
  INV_X1 U2681 ( .A(n3332), .ZN(n3340) );
  INV_X1 U2682 ( .A(n4473), .ZN(n2114) );
  INV_X1 U2683 ( .A(n4517), .ZN(n2119) );
  INV_X1 U2684 ( .A(n4495), .ZN(n2115) );
  INV_X1 U2685 ( .A(IR_REG_2__SCAN_IN), .ZN(n2180) );
  AND2_X1 U2686 ( .A1(n3995), .A2(REG2_REG_18__SCAN_IN), .ZN(n2078) );
  NOR2_X1 U2687 ( .A1(n4608), .A2(n3998), .ZN(n2079) );
  INV_X1 U2688 ( .A(IR_REG_0__SCAN_IN), .ZN(n2099) );
  INV_X1 U2689 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2109) );
  OAI22_X1 U2690 ( .A1(n3721), .A2(n2828), .B1(n3723), .B2(n3722), .ZN(n3606)
         );
  NAND2_X4 U2691 ( .A1(n2052), .A2(n4667), .ZN(n2917) );
  NAND2_X1 U2692 ( .A1(n3649), .A2(n2871), .ZN(n3648) );
  NAND2_X1 U2693 ( .A1(n3281), .A2(n2735), .ZN(n2737) );
  XNOR2_X1 U2694 ( .A(n2742), .B(n2740), .ZN(n2735) );
  AND3_X2 U2695 ( .A1(n2182), .A2(n2259), .A3(n2198), .ZN(n2080) );
  NAND2_X1 U2696 ( .A1(n2253), .A2(n2080), .ZN(n2195) );
  NAND3_X1 U2697 ( .A1(n4562), .A2(n2707), .A3(n3340), .ZN(n3339) );
  AND2_X1 U2698 ( .A1(n3298), .A2(n3332), .ZN(n4637) );
  NAND2_X1 U2699 ( .A1(n3351), .A2(n2081), .ZN(n3365) );
  AND4_X2 U2700 ( .A1(n2161), .A2(n2189), .A3(n2082), .A4(n2192), .ZN(n2285)
         );
  NAND3_X1 U2701 ( .A1(n2189), .A2(n2192), .A3(n2083), .ZN(n2085) );
  INV_X1 U2702 ( .A(n2085), .ZN(n2520) );
  NAND2_X1 U2703 ( .A1(n2097), .A2(n2095), .ZN(n2088) );
  NAND3_X1 U2704 ( .A1(n2089), .A2(n2088), .A3(IR_REG_0__SCAN_IN), .ZN(n2087)
         );
  INV_X1 U2705 ( .A(n2256), .ZN(n2110) );
  OAI21_X1 U2706 ( .B1(n2118), .B2(n4475), .A(n2116), .ZN(n4483) );
  INV_X1 U2707 ( .A(n2123), .ZN(n4442) );
  INV_X1 U2708 ( .A(n2121), .ZN(n4440) );
  NAND2_X1 U2709 ( .A1(n2298), .A2(n2383), .ZN(n2124) );
  INV_X1 U2710 ( .A(n3983), .ZN(n2130) );
  NAND2_X1 U2711 ( .A1(n2175), .A2(n2137), .ZN(n2136) );
  NOR2_X2 U2712 ( .A1(n2136), .A2(n2224), .ZN(n2192) );
  NAND2_X2 U2713 ( .A1(n2140), .A2(n2139), .ZN(n3966) );
  INV_X1 U2714 ( .A(n2142), .ZN(n2140) );
  NAND2_X1 U2715 ( .A1(n2144), .A2(n2143), .ZN(n2769) );
  NAND2_X1 U2716 ( .A1(n2145), .A2(n2146), .ZN(n2952) );
  NAND2_X1 U2717 ( .A1(n3761), .A2(n2147), .ZN(n2145) );
  NAND2_X1 U2718 ( .A1(n3761), .A2(n2901), .ZN(n2151) );
  NAND2_X1 U2719 ( .A1(n3439), .A2(n2152), .ZN(n2791) );
  NAND2_X2 U2720 ( .A1(n3431), .A2(n2779), .ZN(n3439) );
  NAND2_X1 U2721 ( .A1(n2861), .A2(n2157), .ZN(n3649) );
  OAI22_X2 U2722 ( .A1(n3545), .A2(n2160), .B1(n2808), .B2(n2159), .ZN(n2818)
         );
  INV_X1 U2723 ( .A(n2818), .ZN(n2813) );
  NAND2_X1 U2724 ( .A1(n2520), .A2(n2266), .ZN(n2281) );
  NAND2_X1 U2725 ( .A1(n2285), .A2(n2168), .ZN(n2332) );
  NAND2_X1 U2726 ( .A1(n2285), .A2(n2056), .ZN(n2169) );
  NAND2_X1 U2727 ( .A1(n4103), .A2(n4092), .ZN(n4091) );
  INV_X1 U2728 ( .A(n2339), .ZN(n3153) );
  INV_X1 U2729 ( .A(n2357), .ZN(n2339) );
  AND2_X1 U2730 ( .A1(n2697), .A2(n3296), .ZN(n3293) );
  CLKBUF_X1 U2731 ( .A(n3260), .Z(n3313) );
  OR2_X1 U2732 ( .A1(n4020), .A2(n4690), .ZN(n2681) );
  OR2_X1 U2733 ( .A1(n4020), .A2(n4633), .ZN(n2674) );
  NOR2_X2 U2734 ( .A1(n2630), .A2(n2629), .ZN(n4137) );
  NAND2_X1 U2735 ( .A1(n3648), .A2(n2878), .ZN(n3730) );
  AND2_X1 U2736 ( .A1(n2188), .A2(n2194), .ZN(n2189) );
  XNOR2_X1 U2737 ( .A(n3966), .B(n4643), .ZN(n3912) );
  OAI21_X2 U2738 ( .B1(n4084), .B2(n3880), .A(n3879), .ZN(n4070) );
  AOI21_X2 U2739 ( .B1(n4054), .B2(n3867), .A(n3869), .ZN(n4037) );
  AOI21_X2 U2740 ( .B1(n4069), .B2(n2565), .A(n2564), .ZN(n4054) );
  OAI22_X2 U2741 ( .A1(n3127), .A2(n3134), .B1(n4323), .B2(n3140), .ZN(n4217)
         );
  OR2_X1 U2742 ( .A1(n4027), .A2(n4690), .ZN(n2171) );
  AND2_X2 U2743 ( .A1(n2677), .A2(n2924), .ZN(n4704) );
  OR2_X1 U2744 ( .A1(n4027), .A2(n4633), .ZN(n2172) );
  AND2_X2 U2745 ( .A1(n2677), .A2(n3130), .ZN(n4685) );
  NOR2_X1 U2746 ( .A1(n2539), .A2(n2538), .ZN(n2173) );
  NOR2_X1 U2747 ( .A1(n2455), .A2(n3909), .ZN(n2174) );
  NAND2_X1 U2748 ( .A1(n3295), .A2(n2365), .ZN(n3326) );
  INV_X1 U2749 ( .A(IR_REG_22__SCAN_IN), .ZN(n2267) );
  INV_X1 U2750 ( .A(IR_REG_31__SCAN_IN), .ZN(n2286) );
  OR2_X1 U2751 ( .A1(n4513), .A2(n3015), .ZN(n2176) );
  AND2_X1 U2752 ( .A1(n3590), .A2(n3834), .ZN(n4247) );
  INV_X1 U2753 ( .A(n4247), .ZN(n2480) );
  AND2_X1 U2754 ( .A1(n2797), .A2(n2796), .ZN(n2177) );
  OR2_X1 U2755 ( .A1(n3126), .A2(n3125), .ZN(n3967) );
  INV_X1 U2756 ( .A(n2953), .ZN(n2933) );
  OR2_X1 U2757 ( .A1(n3849), .A2(n4334), .ZN(n2179) );
  NAND2_X1 U2758 ( .A1(n2634), .A2(n3891), .ZN(n4084) );
  NAND2_X1 U2759 ( .A1(n2371), .A2(n3330), .ZN(n3325) );
  INV_X1 U2760 ( .A(IR_REG_4__SCAN_IN), .ZN(n2181) );
  NAND2_X1 U2761 ( .A1(n2397), .A2(n2055), .ZN(n3386) );
  OAI21_X1 U2762 ( .B1(n3311), .B2(n3312), .A(n2757), .ZN(n2752) );
  NAND2_X1 U2763 ( .A1(n3965), .A2(n2942), .ZN(n2721) );
  INV_X1 U2764 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2429) );
  INV_X1 U2765 ( .A(n2817), .ZN(n2812) );
  OR2_X1 U2766 ( .A1(n2359), .A2(n2358), .ZN(n2360) );
  AND2_X1 U2767 ( .A1(n2736), .A2(n3278), .ZN(n2728) );
  OR2_X1 U2768 ( .A1(n2430), .A2(n2429), .ZN(n2440) );
  INV_X1 U2769 ( .A(n2783), .ZN(n2784) );
  OR2_X1 U2770 ( .A1(n2550), .A2(n3652), .ZN(n2552) );
  OR2_X1 U2771 ( .A1(n2393), .A2(n3205), .ZN(n2369) );
  AND2_X1 U2772 ( .A1(n3953), .A2(n4241), .ZN(n2687) );
  AND2_X1 U2773 ( .A1(n4281), .A2(n4092), .ZN(n2558) );
  NAND2_X1 U2774 ( .A1(n2543), .A2(REG3_REG_22__SCAN_IN), .ZN(n2550) );
  OR2_X1 U2775 ( .A1(n2586), .A2(n3703), .ZN(n2495) );
  AND2_X1 U2776 ( .A1(n2647), .A2(n2179), .ZN(n2648) );
  NAND2_X1 U2777 ( .A1(n2481), .A2(n2480), .ZN(n3584) );
  INV_X1 U2778 ( .A(n3286), .ZN(n3254) );
  OR2_X1 U2779 ( .A1(n2251), .A2(IR_REG_10__SCAN_IN), .ZN(n2202) );
  NAND2_X1 U2780 ( .A1(n3856), .A2(DATAI_25_), .ZN(n4280) );
  INV_X1 U2781 ( .A(n3787), .ZN(n3770) );
  OR2_X1 U2782 ( .A1(n2586), .A2(n3681), .ZN(n2546) );
  AND4_X1 U2783 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(n4337)
         );
  NAND4_X1 U2784 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .ZN(n3169)
         );
  AOI21_X1 U2785 ( .B1(n4424), .B2(REG2_REG_2__SCAN_IN), .A(n3209), .ZN(n2225)
         );
  NOR2_X1 U2786 ( .A1(n2300), .A2(n4452), .ZN(n4465) );
  INV_X1 U2787 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U2788 ( .A1(n4551), .A2(n4549), .ZN(n4550) );
  XNOR2_X1 U2789 ( .A(n2263), .B(n2499), .ZN(n4551) );
  AND2_X1 U2790 ( .A1(n2493), .A2(REG3_REG_16__SCAN_IN), .ZN(n2500) );
  AND2_X1 U2791 ( .A1(n3164), .A2(n3160), .ZN(n2666) );
  INV_X1 U2792 ( .A(n4202), .ZN(n4199) );
  OR2_X1 U2793 ( .A1(n4561), .A2(n2670), .ZN(n4334) );
  NAND2_X1 U2794 ( .A1(n3202), .A2(n2925), .ZN(n4567) );
  AND2_X1 U2795 ( .A1(n2208), .A2(n2251), .ZN(n3148) );
  INV_X1 U2796 ( .A(n4303), .ZN(n4147) );
  NAND2_X1 U2797 ( .A1(n2938), .A2(STATE_REG_SCAN_IN), .ZN(n3784) );
  AND2_X1 U2798 ( .A1(n3856), .A2(DATAI_20_), .ZN(n4172) );
  AND2_X1 U2799 ( .A1(n2585), .A2(n2584), .ZN(n4014) );
  AND4_X1 U2800 ( .A1(n2349), .A2(n2348), .A3(n2347), .A4(n2346), .ZN(n4292)
         );
  AND4_X1 U2801 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n4220)
         );
  NAND2_X1 U2802 ( .A1(n2234), .A2(n2233), .ZN(n4446) );
  INV_X1 U2803 ( .A(n4426), .ZN(n3202) );
  AND2_X1 U2804 ( .A1(n4436), .A2(n2317), .ZN(n4555) );
  INV_X1 U2805 ( .A(n4420), .ZN(n4003) );
  INV_X1 U2806 ( .A(n4256), .ZN(n4570) );
  AOI21_X1 U2807 ( .B1(n2668), .B2(n2667), .A(n2666), .ZN(n2924) );
  INV_X1 U2808 ( .A(n4187), .ZN(n4191) );
  AND2_X1 U2809 ( .A1(n4563), .A2(n3945), .ZN(n4679) );
  AND2_X1 U2810 ( .A1(n2322), .A2(n2321), .ZN(n4554) );
  INV_X1 U2811 ( .A(n3122), .ZN(n3123) );
  INV_X1 U2812 ( .A(n3710), .ZN(n3740) );
  INV_X1 U2813 ( .A(n4014), .ZN(n4041) );
  OAI211_X1 U2814 ( .C1(n4074), .C2(n2586), .A(n2563), .B(n2562), .ZN(n4087)
         );
  INV_X1 U2815 ( .A(n4205), .ZN(n3958) );
  NAND2_X1 U2816 ( .A1(n4436), .A2(n3202), .ZN(n4560) );
  INV_X1 U2817 ( .A(n4227), .ZN(n4259) );
  NAND2_X1 U2818 ( .A1(n4227), .A2(n3133), .ZN(n4237) );
  AND2_X1 U2819 ( .A1(n2681), .A2(n2680), .ZN(n2682) );
  NAND2_X1 U2820 ( .A1(n4704), .A2(n4674), .ZN(n4690) );
  INV_X1 U2821 ( .A(n4704), .ZN(n4702) );
  AND2_X1 U2822 ( .A1(n4682), .A2(n4681), .ZN(n4703) );
  INV_X1 U2823 ( .A(n4685), .ZN(n4683) );
  INV_X2 U2824 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X2 U2825 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2219)
         );
  NAND2_X1 U2826 ( .A1(n2265), .A2(IR_REG_31__SCAN_IN), .ZN(n2190) );
  XNOR2_X1 U2827 ( .A(n2190), .B(IR_REG_18__SCAN_IN), .ZN(n3995) );
  INV_X1 U2828 ( .A(n3995), .ZN(n4608) );
  INV_X1 U2829 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2191) );
  AOI22_X1 U2830 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4608), .B1(n3995), .B2(
        n2191), .ZN(n2291) );
  AND2_X1 U2831 ( .A1(n2193), .A2(n2194), .ZN(n2253) );
  NAND2_X1 U2832 ( .A1(n2195), .A2(IR_REG_31__SCAN_IN), .ZN(n2196) );
  MUX2_X1 U2833 ( .A(IR_REG_31__SCAN_IN), .B(n2196), .S(IR_REG_17__SCAN_IN), 
        .Z(n2197) );
  NAND2_X1 U2834 ( .A1(n2197), .A2(n2265), .ZN(n2507) );
  INV_X1 U2835 ( .A(n2507), .ZN(n4421) );
  NAND2_X1 U2836 ( .A1(n2253), .A2(n2198), .ZN(n2199) );
  NAND2_X1 U2837 ( .A1(n2199), .A2(IR_REG_31__SCAN_IN), .ZN(n2260) );
  XNOR2_X1 U2838 ( .A(n2260), .B(IR_REG_15__SCAN_IN), .ZN(n4611) );
  INV_X1 U2839 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4530) );
  OR2_X1 U2840 ( .A1(n2253), .A2(n2286), .ZN(n2200) );
  XNOR2_X1 U2841 ( .A(n2200), .B(IR_REG_14__SCAN_IN), .ZN(n2479) );
  AND3_X1 U2842 ( .A1(n3040), .A2(n2210), .A3(n2212), .ZN(n2201) );
  NAND2_X1 U2843 ( .A1(n2193), .A2(n2201), .ZN(n2206) );
  NAND2_X1 U2844 ( .A1(n2202), .A2(IR_REG_31__SCAN_IN), .ZN(n2244) );
  INV_X1 U2845 ( .A(IR_REG_11__SCAN_IN), .ZN(n2249) );
  NAND2_X1 U2846 ( .A1(n2244), .A2(n2249), .ZN(n2203) );
  NAND2_X1 U2847 ( .A1(n2203), .A2(IR_REG_31__SCAN_IN), .ZN(n2204) );
  XNOR2_X1 U2848 ( .A(n2204), .B(IR_REG_12__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U2849 ( .A1(n2251), .A2(IR_REG_31__SCAN_IN), .ZN(n2205) );
  XNOR2_X1 U2850 ( .A(n2205), .B(IR_REG_10__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U2851 ( .A1(n2206), .A2(IR_REG_31__SCAN_IN), .ZN(n2207) );
  MUX2_X1 U2852 ( .A(IR_REG_31__SCAN_IN), .B(n2207), .S(IR_REG_9__SCAN_IN), 
        .Z(n2208) );
  NAND2_X1 U2853 ( .A1(n3148), .A2(REG2_REG_9__SCAN_IN), .ZN(n2241) );
  INV_X1 U2854 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2209) );
  MUX2_X1 U2855 ( .A(REG2_REG_9__SCAN_IN), .B(n2209), .S(n3148), .Z(n4487) );
  NAND2_X1 U2856 ( .A1(n2193), .A2(n2210), .ZN(n2211) );
  NAND2_X1 U2857 ( .A1(n2211), .A2(IR_REG_31__SCAN_IN), .ZN(n2215) );
  NAND2_X1 U2858 ( .A1(n2215), .A2(n2212), .ZN(n2213) );
  NAND2_X1 U2859 ( .A1(n2213), .A2(IR_REG_31__SCAN_IN), .ZN(n2214) );
  XNOR2_X1 U2860 ( .A(n2214), .B(IR_REG_8__SCAN_IN), .ZN(n4473) );
  XNOR2_X1 U2861 ( .A(n2215), .B(IR_REG_7__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U2862 ( .A1(REG2_REG_7__SCAN_IN), .A2(n2417), .ZN(n2238) );
  INV_X1 U2863 ( .A(n2417), .ZN(n4620) );
  INV_X1 U2864 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U2865 ( .A1(REG2_REG_7__SCAN_IN), .A2(n2417), .B1(n4620), .B2(n3415), .ZN(n4470) );
  OR2_X1 U2866 ( .A1(n2193), .A2(n2286), .ZN(n2216) );
  XNOR2_X1 U2867 ( .A(n2216), .B(IR_REG_6__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U2868 ( .A1(n2217), .A2(IR_REG_31__SCAN_IN), .ZN(n2218) );
  XNOR2_X1 U2869 ( .A(n2218), .B(IR_REG_5__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U2870 ( .A1(n4623), .A2(REG2_REG_5__SCAN_IN), .ZN(n2235) );
  INV_X1 U2871 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3423) );
  INV_X1 U2872 ( .A(n4623), .ZN(n4450) );
  AOI22_X1 U2873 ( .A1(n4623), .A2(REG2_REG_5__SCAN_IN), .B1(n3423), .B2(n4450), .ZN(n4447) );
  OR2_X1 U2874 ( .A1(n2219), .A2(n2286), .ZN(n2220) );
  XNOR2_X2 U2875 ( .A(n2220), .B(IR_REG_2__SCAN_IN), .ZN(n4424) );
  INV_X1 U2876 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2222) );
  NAND2_X1 U2877 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2221)
         );
  MUX2_X1 U2878 ( .A(REG2_REG_1__SCAN_IN), .B(n2222), .S(n4425), .Z(n3973) );
  NAND3_X1 U2879 ( .A1(n3973), .A2(REG2_REG_0__SCAN_IN), .A3(IR_REG_0__SCAN_IN), .ZN(n3972) );
  NAND2_X1 U2880 ( .A1(n4425), .A2(REG2_REG_1__SCAN_IN), .ZN(n3210) );
  INV_X1 U2881 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2223) );
  MUX2_X1 U2882 ( .A(n2223), .B(REG2_REG_2__SCAN_IN), .S(n4424), .Z(n3211) );
  AOI21_X1 U2883 ( .B1(n3972), .B2(n3210), .A(n3211), .ZN(n3209) );
  NAND2_X1 U2884 ( .A1(n2224), .A2(IR_REG_31__SCAN_IN), .ZN(n2228) );
  XNOR2_X1 U2885 ( .A(n2228), .B(IR_REG_3__SCAN_IN), .ZN(n4423) );
  XNOR2_X1 U2886 ( .A(n2225), .B(n4423), .ZN(n3183) );
  INV_X1 U2887 ( .A(n2225), .ZN(n2226) );
  AOI22_X1 U2888 ( .A1(n3183), .A2(REG2_REG_3__SCAN_IN), .B1(n4423), .B2(n2226), .ZN(n2231) );
  NAND2_X1 U2889 ( .A1(n2228), .A2(n2227), .ZN(n2229) );
  NAND2_X1 U2890 ( .A1(n2229), .A2(IR_REG_31__SCAN_IN), .ZN(n2230) );
  XNOR2_X1 U2891 ( .A(n2230), .B(IR_REG_4__SCAN_IN), .ZN(n2383) );
  XNOR2_X1 U2892 ( .A(n2231), .B(n2383), .ZN(n3237) );
  NAND2_X1 U2893 ( .A1(n3237), .A2(REG2_REG_4__SCAN_IN), .ZN(n2234) );
  INV_X1 U2894 ( .A(n2231), .ZN(n2232) );
  INV_X1 U2895 ( .A(n2383), .ZN(n3242) );
  NAND2_X1 U2896 ( .A1(n2232), .A2(n2383), .ZN(n2233) );
  NAND2_X1 U2897 ( .A1(n4447), .A2(n4446), .ZN(n4445) );
  NAND2_X1 U2898 ( .A1(n2404), .A2(n2236), .ZN(n2237) );
  NAND2_X1 U2899 ( .A1(n4470), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U2900 ( .A1(n4473), .A2(n2239), .ZN(n2240) );
  NAND2_X1 U2901 ( .A1(n4487), .A2(n4488), .ZN(n4486) );
  NAND2_X1 U2902 ( .A1(n4495), .A2(n2242), .ZN(n2243) );
  XNOR2_X1 U2903 ( .A(n2244), .B(IR_REG_11__SCAN_IN), .ZN(n4615) );
  INV_X1 U2904 ( .A(n4615), .ZN(n4513) );
  INV_X1 U2905 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3015) );
  AOI22_X1 U2906 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4615), .B1(n4513), .B2(
        n3015), .ZN(n4510) );
  NAND2_X1 U2907 ( .A1(n4517), .A2(n2245), .ZN(n2246) );
  INV_X1 U2908 ( .A(IR_REG_10__SCAN_IN), .ZN(n2248) );
  INV_X1 U2909 ( .A(IR_REG_12__SCAN_IN), .ZN(n2247) );
  NAND3_X1 U2910 ( .A1(n2249), .A2(n2248), .A3(n2247), .ZN(n2250) );
  OAI21_X1 U2911 ( .B1(n2251), .B2(n2250), .A(IR_REG_31__SCAN_IN), .ZN(n2252)
         );
  MUX2_X1 U2912 ( .A(IR_REG_31__SCAN_IN), .B(n2252), .S(IR_REG_13__SCAN_IN), 
        .Z(n2255) );
  INV_X1 U2913 ( .A(n2253), .ZN(n2254) );
  NAND2_X1 U2914 ( .A1(n2255), .A2(n2254), .ZN(n3377) );
  INV_X1 U2915 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3378) );
  NOR2_X1 U2916 ( .A1(n3377), .A2(n3378), .ZN(n3376) );
  INV_X1 U2917 ( .A(n3377), .ZN(n4422) );
  OAI22_X1 U2918 ( .A1(n3380), .A2(n3376), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4422), .ZN(n2256) );
  NOR2_X1 U2919 ( .A1(n2125), .A2(n2256), .ZN(n2257) );
  NAND2_X1 U2920 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4611), .ZN(n2258) );
  OAI21_X1 U2921 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4611), .A(n2258), .ZN(n4539) );
  AOI21_X1 U2922 ( .B1(n4611), .B2(REG2_REG_15__SCAN_IN), .A(n4538), .ZN(n2263) );
  NAND2_X1 U2923 ( .A1(n2260), .A2(n2259), .ZN(n2261) );
  NAND2_X1 U2924 ( .A1(n2261), .A2(IR_REG_31__SCAN_IN), .ZN(n2262) );
  XNOR2_X1 U2925 ( .A(n2262), .B(IR_REG_16__SCAN_IN), .ZN(n2499) );
  INV_X1 U2926 ( .A(n2499), .ZN(n4610) );
  NAND2_X1 U2927 ( .A1(n2263), .A2(n4610), .ZN(n2264) );
  INV_X1 U2928 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U2929 ( .A1(n2264), .A2(n4550), .ZN(n3984) );
  XNOR2_X1 U2930 ( .A(n2507), .B(REG2_REG_17__SCAN_IN), .ZN(n3986) );
  NAND2_X1 U2931 ( .A1(n3984), .A2(n3986), .ZN(n3985) );
  NOR2_X1 U2932 ( .A1(n2272), .A2(n2286), .ZN(n2269) );
  MUX2_X1 U2933 ( .A(n2286), .B(n2269), .S(IR_REG_25__SCAN_IN), .Z(n2270) );
  INV_X1 U2934 ( .A(n2270), .ZN(n2273) );
  INV_X1 U2935 ( .A(n2285), .ZN(n2279) );
  NAND2_X1 U2936 ( .A1(n2273), .A2(n2279), .ZN(n3163) );
  NAND2_X1 U2937 ( .A1(n2278), .A2(n2277), .ZN(n2274) );
  XNOR2_X2 U2938 ( .A(n2275), .B(IR_REG_24__SCAN_IN), .ZN(n4416) );
  OR2_X1 U2939 ( .A1(n2086), .A2(n2286), .ZN(n2276) );
  NAND3_X2 U2940 ( .A1(n2652), .A2(n4416), .A3(n4415), .ZN(n3126) );
  XNOR2_X1 U2941 ( .A(n2278), .B(n2277), .ZN(n2937) );
  NAND2_X1 U2942 ( .A1(n3126), .A2(n4605), .ZN(n3158) );
  NOR2_X1 U2943 ( .A1(n2937), .A2(U3149), .ZN(n3946) );
  INV_X1 U2944 ( .A(n3946), .ZN(n3951) );
  NAND2_X1 U2945 ( .A1(n3158), .A2(n3951), .ZN(n2321) );
  NAND2_X1 U2946 ( .A1(n2064), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  INV_X1 U2947 ( .A(n3945), .ZN(n4417) );
  NAND2_X1 U2948 ( .A1(n2281), .A2(IR_REG_31__SCAN_IN), .ZN(n2282) );
  NAND2_X1 U2949 ( .A1(n2925), .A2(n2937), .ZN(n2283) );
  AND2_X1 U2950 ( .A1(n3856), .A2(n2283), .ZN(n2320) );
  NOR2_X1 U2951 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2284)
         );
  OR2_X1 U2952 ( .A1(n2330), .A2(n2286), .ZN(n2287) );
  XNOR2_X1 U2953 ( .A(n2288), .B(IR_REG_27__SCAN_IN), .ZN(n4434) );
  NAND2_X1 U2954 ( .A1(n4426), .A2(n4434), .ZN(n3948) );
  INV_X1 U2955 ( .A(n3948), .ZN(n2289) );
  AOI211_X1 U2956 ( .C1(n2291), .C2(n2290), .A(n3994), .B(n4548), .ZN(n2328)
         );
  INV_X1 U2957 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U2958 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3995), .B1(n4608), .B2(
        n3998), .ZN(n2319) );
  NOR2_X1 U2959 ( .A1(n4421), .A2(REG1_REG_17__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2960 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4611), .ZN(n2311) );
  INV_X1 U2961 ( .A(n4611), .ZN(n4547) );
  AOI22_X1 U2962 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4611), .B1(n4547), .B2(
        n4341), .ZN(n4544) );
  NAND2_X1 U2963 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4615), .ZN(n2306) );
  INV_X1 U2964 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2447) );
  AOI22_X1 U2965 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4615), .B1(n4513), .B2(
        n2447), .ZN(n4507) );
  NAND2_X1 U2966 ( .A1(n3148), .A2(REG1_REG_9__SCAN_IN), .ZN(n2303) );
  INV_X1 U2967 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2292) );
  MUX2_X1 U2968 ( .A(n2292), .B(REG1_REG_9__SCAN_IN), .S(n3148), .Z(n2293) );
  INV_X1 U2969 ( .A(n2293), .ZN(n4484) );
  INV_X1 U2970 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4694) );
  MUX2_X1 U2971 ( .A(REG1_REG_2__SCAN_IN), .B(n4694), .S(n4424), .Z(n3208) );
  INV_X1 U2972 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4688) );
  XNOR2_X1 U2973 ( .A(n4425), .B(n4688), .ZN(n3970) );
  AND2_X1 U2974 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3969)
         );
  NAND2_X1 U2975 ( .A1(n3970), .A2(n3969), .ZN(n3968) );
  NAND2_X1 U2976 ( .A1(n4425), .A2(REG1_REG_1__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2977 ( .A1(n3968), .A2(n2294), .ZN(n3207) );
  NAND2_X1 U2978 ( .A1(n3208), .A2(n3207), .ZN(n3206) );
  NAND2_X1 U2979 ( .A1(n4424), .A2(REG1_REG_2__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2980 ( .A1(n3206), .A2(n2295), .ZN(n2296) );
  INV_X1 U2981 ( .A(n4423), .ZN(n3184) );
  XNOR2_X1 U2982 ( .A(n2296), .B(n3184), .ZN(n3187) );
  NAND2_X1 U2983 ( .A1(n3187), .A2(REG1_REG_3__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U2984 ( .A1(n2296), .A2(n4423), .ZN(n2297) );
  NAND2_X1 U2985 ( .A1(n3186), .A2(n2297), .ZN(n2298) );
  XNOR2_X1 U2986 ( .A(n2298), .B(n3242), .ZN(n3239) );
  NAND2_X1 U2987 ( .A1(n3239), .A2(REG1_REG_4__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U2988 ( .A1(n4623), .A2(REG1_REG_5__SCAN_IN), .ZN(n2299) );
  OAI21_X1 U2989 ( .B1(n4623), .B2(REG1_REG_5__SCAN_IN), .A(n2299), .ZN(n4441)
         );
  INV_X1 U2990 ( .A(n2404), .ZN(n4622) );
  NOR2_X1 U2991 ( .A1(n2060), .A2(n4622), .ZN(n2300) );
  INV_X1 U2992 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4698) );
  XNOR2_X1 U2993 ( .A(n2060), .B(n4622), .ZN(n4453) );
  NOR2_X1 U2994 ( .A1(n4698), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U2995 ( .A1(REG1_REG_7__SCAN_IN), .A2(n2417), .ZN(n4461) );
  NOR2_X1 U2996 ( .A1(REG1_REG_7__SCAN_IN), .A2(n2417), .ZN(n4460) );
  AOI21_X1 U2997 ( .B1(n4465), .B2(n4461), .A(n4460), .ZN(n2301) );
  NAND2_X1 U2998 ( .A1(n4473), .A2(n2301), .ZN(n2302) );
  NAND2_X1 U2999 ( .A1(n2303), .A2(n4483), .ZN(n2304) );
  NAND2_X1 U3000 ( .A1(n4495), .A2(n2304), .ZN(n2305) );
  XOR2_X1 U3001 ( .A(n2304), .B(n4495), .Z(n4497) );
  NAND2_X1 U3002 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4497), .ZN(n4496) );
  NAND2_X1 U3003 ( .A1(n4517), .A2(n2307), .ZN(n2308) );
  NAND2_X1 U3004 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4525), .ZN(n4524) );
  INV_X1 U3005 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4352) );
  XNOR2_X1 U3006 ( .A(n3377), .B(n4352), .ZN(n3372) );
  NAND2_X1 U3007 ( .A1(n2479), .A2(n2309), .ZN(n2310) );
  NAND2_X1 U3008 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4535), .ZN(n4534) );
  NOR2_X1 U3009 ( .A1(n2499), .A2(n2312), .ZN(n2313) );
  NOR2_X1 U3010 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4556), .ZN(n4557) );
  NOR2_X1 U3011 ( .A1(n2313), .A2(n4557), .ZN(n3983) );
  INV_X1 U3012 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2315) );
  INV_X1 U3013 ( .A(n2316), .ZN(n2314) );
  OAI21_X1 U3014 ( .B1(n2315), .B2(n2507), .A(n2314), .ZN(n3982) );
  INV_X1 U3015 ( .A(n4434), .ZN(n2317) );
  OAI211_X1 U3016 ( .C1(n2319), .C2(n2318), .A(n4555), .B(n3997), .ZN(n2326)
         );
  INV_X1 U3017 ( .A(n2320), .ZN(n2322) );
  INV_X1 U3018 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3027) );
  NOR2_X1 U3019 ( .A1(n3027), .A2(STATE_REG_SCAN_IN), .ZN(n3612) );
  AOI21_X1 U3020 ( .B1(n4554), .B2(ADDR_REG_18__SCAN_IN), .A(n3612), .ZN(n2323) );
  OAI21_X1 U3021 ( .B1(n4560), .B2(n4608), .A(n2323), .ZN(n2324) );
  INV_X1 U3022 ( .A(n2324), .ZN(n2325) );
  INV_X1 U3023 ( .A(n4092), .ZN(n3734) );
  INV_X1 U3024 ( .A(n2359), .ZN(n2334) );
  NAND2_X1 U3025 ( .A1(n2399), .A2(REG3_REG_6__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3026 ( .A1(n2421), .A2(REG3_REG_8__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3027 ( .A1(n2458), .A2(REG3_REG_12__SCAN_IN), .ZN(n2465) );
  INV_X1 U3028 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U3029 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2335) );
  NAND2_X1 U3030 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2336) );
  INV_X1 U3031 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3652) );
  INV_X1 U3032 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U3033 ( .A1(n2552), .A2(n3735), .ZN(n2337) );
  AND2_X1 U3034 ( .A1(n2560), .A2(n2337), .ZN(n4093) );
  NAND2_X1 U3035 ( .A1(n2352), .A2(n4093), .ZN(n2343) );
  INV_X4 U3036 ( .A(n2053), .ZN(n2398) );
  INV_X1 U3037 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4289) );
  OR2_X1 U3038 ( .A1(n2398), .A2(n4289), .ZN(n2342) );
  AND2_X2 U3039 ( .A1(n2359), .A2(n2339), .ZN(n2356) );
  NAND2_X1 U3040 ( .A1(n2432), .A2(REG0_REG_24__SCAN_IN), .ZN(n2341) );
  AND2_X2 U3041 ( .A1(n2338), .A2(n2339), .ZN(n2355) );
  NAND2_X1 U3042 ( .A1(n2525), .A2(REG2_REG_24__SCAN_IN), .ZN(n2340) );
  NAND4_X1 U3043 ( .A1(n2343), .A2(n2342), .A3(n2341), .A4(n2340), .ZN(n3956)
         );
  NAND2_X1 U3044 ( .A1(n2525), .A2(REG2_REG_22__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3045 ( .A1(n2432), .A2(REG0_REG_22__SCAN_IN), .ZN(n2348) );
  INV_X1 U3046 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2344) );
  OR2_X1 U3047 ( .A1(n2398), .A2(n2344), .ZN(n2347) );
  OR2_X1 U3048 ( .A1(n2543), .A2(REG3_REG_22__SCAN_IN), .ZN(n2345) );
  NAND2_X1 U3049 ( .A1(n2550), .A2(n2345), .ZN(n4121) );
  OR2_X1 U3050 ( .A1(n2586), .A2(n4121), .ZN(n2346) );
  NAND2_X1 U3051 ( .A1(n2356), .A2(REG0_REG_0__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3052 ( .A1(n2355), .A2(REG2_REG_0__SCAN_IN), .ZN(n2350) );
  INV_X1 U3053 ( .A(n2393), .ZN(n2352) );
  INV_X1 U3054 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U3055 ( .A1(n2355), .A2(REG2_REG_1__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3056 ( .A1(n2357), .A2(REG3_REG_1__SCAN_IN), .ZN(n2358) );
  INV_X2 U3057 ( .A(n2364), .ZN(n2705) );
  MUX2_X1 U3058 ( .A(n4425), .B(DATAI_1_), .S(n2366), .Z(n3671) );
  NAND2_X1 U3059 ( .A1(n2705), .A2(n3671), .ZN(n2601) );
  NAND2_X1 U3060 ( .A1(n2707), .A2(n2364), .ZN(n3793) );
  NAND2_X2 U3061 ( .A1(n2601), .A2(n3793), .ZN(n2599) );
  NAND2_X1 U3062 ( .A1(n3293), .A2(n2599), .ZN(n3295) );
  NAND2_X1 U3063 ( .A1(n3172), .A2(n3671), .ZN(n2365) );
  INV_X1 U3064 ( .A(n3326), .ZN(n2371) );
  NAND2_X1 U3065 ( .A1(n2356), .A2(REG0_REG_2__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3066 ( .A1(n2355), .A2(REG2_REG_2__SCAN_IN), .ZN(n2370) );
  OR2_X1 U3067 ( .A1(n2354), .A2(n4694), .ZN(n2368) );
  INV_X1 U3068 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3205) );
  MUX2_X1 U3069 ( .A(n4424), .B(DATAI_2_), .S(n2366), .Z(n3332) );
  NAND2_X1 U3070 ( .A1(n3169), .A2(n3340), .ZN(n3798) );
  NAND2_X1 U3071 ( .A1(n2372), .A2(n3340), .ZN(n2373) );
  NAND2_X1 U3072 ( .A1(n3325), .A2(n2373), .ZN(n3345) );
  INV_X1 U3073 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U3074 ( .A1(n2356), .A2(REG0_REG_3__SCAN_IN), .ZN(n2375) );
  MUX2_X1 U3075 ( .A(n4423), .B(DATAI_3_), .S(n3857), .Z(n4643) );
  NOR2_X1 U3076 ( .A1(n3966), .A2(n4643), .ZN(n2377) );
  INV_X1 U3077 ( .A(n3966), .ZN(n3800) );
  INV_X1 U3078 ( .A(n4643), .ZN(n3355) );
  OAI22_X1 U3079 ( .A1(n3345), .A2(n2377), .B1(n3800), .B2(n3355), .ZN(n3247)
         );
  NAND2_X1 U3080 ( .A1(n2355), .A2(REG2_REG_4__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3081 ( .A1(n2356), .A2(REG0_REG_4__SCAN_IN), .ZN(n2381) );
  INV_X1 U3082 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2378) );
  OR2_X1 U3083 ( .A1(n2398), .A2(n2378), .ZN(n2380) );
  XNOR2_X1 U3084 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3290) );
  AND4_X2 U3085 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .ZN(n3420)
         );
  MUX2_X1 U3086 ( .A(n2383), .B(DATAI_4_), .S(n3857), .Z(n3286) );
  NAND2_X1 U3087 ( .A1(n3420), .A2(n3286), .ZN(n3802) );
  INV_X1 U3088 ( .A(n3420), .ZN(n3717) );
  NAND2_X1 U3089 ( .A1(n3802), .A2(n3805), .ZN(n3907) );
  NAND2_X1 U3090 ( .A1(n3247), .A2(n3907), .ZN(n2385) );
  NAND2_X1 U3091 ( .A1(n3717), .A2(n3286), .ZN(n2384) );
  NAND2_X1 U3092 ( .A1(n2385), .A2(n2384), .ZN(n3360) );
  INV_X1 U3093 ( .A(n3360), .ZN(n2397) );
  INV_X1 U3094 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2386) );
  OR2_X1 U3095 ( .A1(n2398), .A2(n2386), .ZN(n2396) );
  NAND2_X1 U3096 ( .A1(n2355), .A2(REG2_REG_5__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U3097 ( .A1(n2356), .A2(REG0_REG_5__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U3098 ( .A1(n2388), .A2(n2387), .ZN(n2394) );
  INV_X1 U3099 ( .A(n2399), .ZN(n2392) );
  INV_X1 U3100 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3101 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2389) );
  NAND2_X1 U3102 ( .A1(n2390), .A2(n2389), .ZN(n2391) );
  NAND2_X1 U3103 ( .A1(n2392), .A2(n2391), .ZN(n3715) );
  NOR2_X1 U3104 ( .A1(n2394), .A2(n2066), .ZN(n2395) );
  MUX2_X1 U3105 ( .A(n4623), .B(DATAI_5_), .S(n3857), .Z(n3714) );
  OR2_X1 U3106 ( .A1(n2398), .A2(n4698), .ZN(n2403) );
  OAI21_X1 U3107 ( .B1(n2399), .B2(REG3_REG_6__SCAN_IN), .A(n2411), .ZN(n3399)
         );
  OR2_X1 U3108 ( .A1(n2586), .A2(n3399), .ZN(n2402) );
  NAND2_X1 U3109 ( .A1(n2525), .A2(REG2_REG_6__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3110 ( .A1(n2356), .A2(REG0_REG_6__SCAN_IN), .ZN(n2400) );
  NAND4_X1 U3111 ( .A1(n2403), .A2(n2402), .A3(n2401), .A4(n2400), .ZN(n3713)
         );
  MUX2_X1 U3112 ( .A(n2404), .B(DATAI_6_), .S(n3857), .Z(n3390) );
  OR2_X1 U3113 ( .A1(n3713), .A2(n3390), .ZN(n2405) );
  INV_X1 U3114 ( .A(n3965), .ZN(n3392) );
  NAND2_X1 U3115 ( .A1(n3392), .A2(n3421), .ZN(n3387) );
  AND2_X1 U3116 ( .A1(n2405), .A2(n3387), .ZN(n2406) );
  NAND2_X1 U3117 ( .A1(n3386), .A2(n2406), .ZN(n2408) );
  NAND2_X1 U3118 ( .A1(n3713), .A2(n3390), .ZN(n2407) );
  NAND2_X1 U3119 ( .A1(n2408), .A2(n2407), .ZN(n3413) );
  NAND2_X1 U3120 ( .A1(n2525), .A2(REG2_REG_7__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U3121 ( .A1(n2356), .A2(REG0_REG_7__SCAN_IN), .ZN(n2415) );
  INV_X1 U3122 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2409) );
  OR2_X1 U3123 ( .A1(n2398), .A2(n2409), .ZN(n2414) );
  AND2_X1 U3124 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  OR2_X1 U3125 ( .A1(n2412), .A2(n2421), .ZN(n3414) );
  OR2_X1 U3126 ( .A1(n2586), .A2(n3414), .ZN(n2413) );
  MUX2_X1 U3127 ( .A(n2417), .B(DATAI_7_), .S(n3857), .Z(n3409) );
  NAND2_X1 U3128 ( .A1(n3452), .A2(n3409), .ZN(n3812) );
  INV_X1 U3129 ( .A(n3409), .ZN(n2749) );
  NAND2_X1 U3130 ( .A1(n3964), .A2(n2749), .ZN(n3814) );
  NAND2_X1 U3131 ( .A1(n3413), .A2(n3908), .ZN(n2419) );
  NAND2_X1 U3132 ( .A1(n3964), .A2(n3409), .ZN(n2418) );
  NAND2_X1 U3133 ( .A1(n2419), .A2(n2418), .ZN(n3448) );
  INV_X1 U3134 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2420) );
  OR2_X1 U3135 ( .A1(n2398), .A2(n2420), .ZN(n2426) );
  OR2_X1 U3136 ( .A1(n2421), .A2(REG3_REG_8__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3137 ( .A1(n2430), .A2(n2422), .ZN(n3460) );
  OR2_X1 U3138 ( .A1(n2586), .A2(n3460), .ZN(n2425) );
  NAND2_X1 U3139 ( .A1(n2432), .A2(REG0_REG_8__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3140 ( .A1(n2525), .A2(REG2_REG_8__SCAN_IN), .ZN(n2423) );
  NAND4_X1 U3141 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(n3963)
         );
  AND2_X1 U3142 ( .A1(n3963), .A2(n3450), .ZN(n2428) );
  OAI21_X2 U3143 ( .B1(n3448), .B2(n2428), .A(n2427), .ZN(n3469) );
  NAND2_X1 U3144 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  NAND2_X1 U3145 ( .A1(n2440), .A2(n2431), .ZN(n3470) );
  OR2_X1 U3146 ( .A1(n2586), .A2(n3470), .ZN(n2436) );
  OR2_X1 U3147 ( .A1(n2398), .A2(n2292), .ZN(n2435) );
  NAND2_X1 U31480 ( .A1(n2525), .A2(REG2_REG_9__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U31490 ( .A1(n2432), .A2(REG0_REG_9__SCAN_IN), .ZN(n2433) );
  MUX2_X1 U3150 ( .A(n3148), .B(DATAI_9_), .S(n3856), .Z(n3473) );
  NOR2_X1 U3151 ( .A1(n3483), .A2(n3473), .ZN(n2438) );
  NAND2_X1 U3152 ( .A1(n3483), .A2(n3473), .ZN(n2437) );
  OAI21_X2 U3153 ( .B1(n3469), .B2(n2438), .A(n2437), .ZN(n3480) );
  INV_X1 U3154 ( .A(n3480), .ZN(n2446) );
  INV_X1 U3155 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2439) );
  OR2_X1 U3156 ( .A1(n2398), .A2(n2439), .ZN(n2445) );
  NAND2_X1 U3157 ( .A1(n2440), .A2(n3442), .ZN(n2441) );
  NAND2_X1 U3158 ( .A1(n2448), .A2(n2441), .ZN(n3492) );
  OR2_X1 U3159 ( .A1(n2586), .A2(n3492), .ZN(n2444) );
  NAND2_X1 U3160 ( .A1(n2432), .A2(REG0_REG_10__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3161 ( .A1(n2525), .A2(REG2_REG_10__SCAN_IN), .ZN(n2442) );
  INV_X1 U3162 ( .A(n3490), .ZN(n3479) );
  NAND2_X1 U3163 ( .A1(n3533), .A2(n3479), .ZN(n3535) );
  NAND2_X1 U3164 ( .A1(n2432), .A2(REG0_REG_11__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3165 ( .A1(n2525), .A2(REG2_REG_11__SCAN_IN), .ZN(n2452) );
  OR2_X1 U3166 ( .A1(n2398), .A2(n2447), .ZN(n2451) );
  AND2_X1 U3167 ( .A1(n2448), .A2(n3634), .ZN(n2449) );
  OR2_X1 U3168 ( .A1(n2449), .A2(n2458), .ZN(n3635) );
  OR2_X1 U3169 ( .A1(n2586), .A2(n3635), .ZN(n2450) );
  MUX2_X1 U3170 ( .A(n4615), .B(DATAI_11_), .S(n3856), .Z(n3633) );
  NAND2_X1 U3171 ( .A1(n3621), .A2(n2786), .ZN(n2454) );
  AND2_X1 U3172 ( .A1(n3535), .A2(n2454), .ZN(n2456) );
  INV_X1 U3173 ( .A(n2454), .ZN(n2455) );
  NAND2_X1 U3174 ( .A1(n3621), .A2(n3633), .ZN(n3518) );
  INV_X1 U3175 ( .A(n3621), .ZN(n3961) );
  NAND2_X1 U3176 ( .A1(n3961), .A2(n2786), .ZN(n3520) );
  NAND2_X1 U3177 ( .A1(n3518), .A2(n3520), .ZN(n3909) );
  AOI21_X2 U3178 ( .B1(n3534), .B2(n2456), .A(n2174), .ZN(n3526) );
  INV_X1 U3179 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3180 ( .A1(n2398), .A2(n2457), .ZN(n2463) );
  OR2_X1 U3181 ( .A1(n2458), .A2(REG3_REG_12__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3182 ( .A1(n2465), .A2(n2459), .ZN(n3523) );
  NAND2_X1 U3183 ( .A1(n2525), .A2(REG2_REG_12__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3184 ( .A1(n2432), .A2(REG0_REG_12__SCAN_IN), .ZN(n2460) );
  MUX2_X1 U3185 ( .A(n4517), .B(DATAI_12_), .S(n3856), .Z(n3620) );
  NOR2_X1 U3186 ( .A1(n3632), .A2(n3620), .ZN(n2464) );
  INV_X1 U3187 ( .A(n3632), .ZN(n2613) );
  OAI22_X1 U3188 ( .A1(n3526), .A2(n2464), .B1(n2613), .B2(n3573), .ZN(n3556)
         );
  NAND2_X1 U3189 ( .A1(n2525), .A2(REG2_REG_13__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3190 ( .A1(n2432), .A2(REG0_REG_13__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3191 ( .A1(n2398), .A2(n4352), .ZN(n2468) );
  NAND2_X1 U3192 ( .A1(n2465), .A2(n3374), .ZN(n2466) );
  NAND2_X1 U3193 ( .A1(n2482), .A2(n2466), .ZN(n3568) );
  OR2_X1 U3194 ( .A1(n2586), .A2(n3568), .ZN(n2467) );
  INV_X1 U3195 ( .A(DATAI_13_), .ZN(n2471) );
  MUX2_X1 U3196 ( .A(n3377), .B(n2471), .S(n3856), .Z(n2800) );
  NAND2_X1 U3197 ( .A1(n4244), .A2(n2800), .ZN(n3555) );
  NAND2_X1 U3198 ( .A1(n3556), .A2(n3555), .ZN(n2472) );
  NAND2_X1 U3199 ( .A1(n3959), .A2(n3566), .ZN(n3554) );
  NAND2_X1 U3200 ( .A1(n2472), .A2(n3554), .ZN(n4245) );
  INV_X1 U3201 ( .A(n4245), .ZN(n2481) );
  NAND2_X1 U3202 ( .A1(n2525), .A2(REG2_REG_14__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U3203 ( .A1(n2432), .A2(REG0_REG_14__SCAN_IN), .ZN(n2477) );
  INV_X1 U3204 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3205 ( .A1(n2398), .A2(n2473), .ZN(n2476) );
  INV_X1 U3206 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2474) );
  XNOR2_X1 U3207 ( .A(n2482), .B(n2474), .ZN(n3549) );
  OR2_X1 U3208 ( .A1(n2586), .A2(n3549), .ZN(n2475) );
  MUX2_X1 U3209 ( .A(n2479), .B(DATAI_14_), .S(n3856), .Z(n4253) );
  NAND2_X1 U32100 ( .A1(n4337), .A2(n4253), .ZN(n3590) );
  INV_X1 U32110 ( .A(n4253), .ZN(n2807) );
  NAND2_X1 U32120 ( .A1(n3786), .A2(n2807), .ZN(n3834) );
  INV_X1 U32130 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4341) );
  OR2_X1 U32140 ( .A1(n2398), .A2(n4341), .ZN(n2488) );
  INV_X1 U32150 ( .A(n2482), .ZN(n2483) );
  AOI21_X1 U32160 ( .B1(n2483), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2484) );
  OR2_X1 U32170 ( .A1(n2484), .A2(n2493), .ZN(n3783) );
  OR2_X1 U32180 ( .A1(n2586), .A2(n3783), .ZN(n2487) );
  NAND2_X1 U32190 ( .A1(n2432), .A2(REG0_REG_15__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U32200 ( .A1(n2525), .A2(REG2_REG_15__SCAN_IN), .ZN(n2485) );
  AND2_X1 U32210 ( .A1(n4242), .A2(n3782), .ZN(n2491) );
  NOR2_X1 U32220 ( .A1(n3786), .A2(n4253), .ZN(n3586) );
  INV_X1 U32230 ( .A(n2491), .ZN(n2489) );
  INV_X1 U32240 ( .A(n4242), .ZN(n2619) );
  INV_X1 U32250 ( .A(n3782), .ZN(n4335) );
  AOI22_X1 U32260 ( .A1(n3586), .A2(n2489), .B1(n2619), .B2(n4335), .ZN(n2490)
         );
  OAI21_X2 U32270 ( .B1(n3584), .B2(n2491), .A(n2490), .ZN(n3127) );
  NAND2_X1 U32280 ( .A1(n2432), .A2(REG0_REG_16__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U32290 ( .A1(n2525), .A2(REG2_REG_16__SCAN_IN), .ZN(n2497) );
  INV_X1 U32300 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2492) );
  OR2_X1 U32310 ( .A1(n2398), .A2(n2492), .ZN(n2496) );
  NOR2_X1 U32320 ( .A1(n2493), .A2(REG3_REG_16__SCAN_IN), .ZN(n2494) );
  OR2_X1 U32330 ( .A1(n2500), .A2(n2494), .ZN(n3703) );
  MUX2_X1 U32340 ( .A(n2499), .B(DATAI_16_), .S(n3856), .Z(n3701) );
  NAND2_X1 U32350 ( .A1(n4323), .A2(n3701), .ZN(n3827) );
  NAND2_X1 U32360 ( .A1(n3779), .A2(n3140), .ZN(n3835) );
  NAND2_X1 U32370 ( .A1(n2525), .A2(REG2_REG_17__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32380 ( .A1(n2432), .A2(REG0_REG_17__SCAN_IN), .ZN(n2504) );
  OR2_X1 U32390 ( .A1(n2398), .A2(n2315), .ZN(n2503) );
  OR2_X1 U32400 ( .A1(n2500), .A2(REG3_REG_17__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U32410 ( .A1(n2526), .A2(n2501), .ZN(n4226) );
  OR2_X1 U32420 ( .A1(n2586), .A2(n4226), .ZN(n2502) );
  INV_X1 U32430 ( .A(DATAI_17_), .ZN(n2506) );
  MUX2_X1 U32440 ( .A(n2507), .B(n2506), .S(n3856), .Z(n4322) );
  NAND2_X1 U32450 ( .A1(n4205), .A2(n4322), .ZN(n4159) );
  INV_X1 U32460 ( .A(REG1_REG_20__SCAN_IN), .ZN(n2508) );
  OR2_X1 U32470 ( .A1(n2398), .A2(n2508), .ZN(n2514) );
  INV_X1 U32480 ( .A(n2528), .ZN(n2509) );
  AOI21_X1 U32490 ( .B1(n2509), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2510) );
  OR2_X1 U32500 ( .A1(n2510), .A2(n2541), .ZN(n3745) );
  OR2_X1 U32510 ( .A1(n2586), .A2(n3745), .ZN(n2513) );
  NAND2_X1 U32520 ( .A1(n2432), .A2(REG0_REG_20__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32530 ( .A1(n2525), .A2(REG2_REG_20__SCAN_IN), .ZN(n2511) );
  NAND4_X1 U32540 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n4188)
         );
  NAND2_X1 U32550 ( .A1(n4188), .A2(n4172), .ZN(n3888) );
  INV_X1 U32560 ( .A(n3888), .ZN(n2522) );
  INV_X1 U32570 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4317) );
  OR2_X1 U32580 ( .A1(n2398), .A2(n4317), .ZN(n2519) );
  INV_X1 U32590 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2515) );
  XNOR2_X1 U32600 ( .A(n2528), .B(n2515), .ZN(n4192) );
  OR2_X1 U32610 ( .A1(n2586), .A2(n4192), .ZN(n2518) );
  NAND2_X1 U32620 ( .A1(n2432), .A2(REG0_REG_19__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32630 ( .A1(n2525), .A2(REG2_REG_19__SCAN_IN), .ZN(n2516) );
  NAND4_X1 U32640 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n4203)
         );
  MUX2_X1 U32650 ( .A(n4420), .B(DATAI_19_), .S(n3856), .Z(n4187) );
  NAND2_X1 U32660 ( .A1(n4158), .A2(n4191), .ZN(n4164) );
  NAND2_X1 U32670 ( .A1(n4304), .A2(n2669), .ZN(n3889) );
  AND2_X1 U32680 ( .A1(n4164), .A2(n3889), .ZN(n2521) );
  INV_X1 U32690 ( .A(n2533), .ZN(n2524) );
  NAND2_X1 U32700 ( .A1(n4203), .A2(n4187), .ZN(n4163) );
  AND2_X1 U32710 ( .A1(n4163), .A2(n3888), .ZN(n2523) );
  NOR2_X1 U32720 ( .A1(n2524), .A2(n2523), .ZN(n2536) );
  NAND2_X1 U32730 ( .A1(n2525), .A2(REG2_REG_18__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32740 ( .A1(n2432), .A2(REG0_REG_18__SCAN_IN), .ZN(n2531) );
  OR2_X1 U32750 ( .A1(n2398), .A2(n3998), .ZN(n2530) );
  NAND2_X1 U32760 ( .A1(n2526), .A2(n3027), .ZN(n2527) );
  NAND2_X1 U32770 ( .A1(n2528), .A2(n2527), .ZN(n4208) );
  OR2_X1 U32780 ( .A1(n2586), .A2(n4208), .ZN(n2529) );
  MUX2_X1 U32790 ( .A(n3995), .B(DATAI_18_), .S(n3857), .Z(n4202) );
  NAND2_X1 U32800 ( .A1(n4220), .A2(n4199), .ZN(n4162) );
  AND2_X1 U32810 ( .A1(n4162), .A2(n2533), .ZN(n2534) );
  AND2_X1 U32820 ( .A1(n4159), .A2(n2535), .ZN(n2540) );
  INV_X1 U32830 ( .A(n2535), .ZN(n2539) );
  NAND2_X1 U32840 ( .A1(n3958), .A2(n4231), .ZN(n4160) );
  NAND2_X1 U32850 ( .A1(n4220), .A2(n4202), .ZN(n4181) );
  INV_X1 U32860 ( .A(n4220), .ZN(n3957) );
  NAND2_X1 U32870 ( .A1(n3957), .A2(n4199), .ZN(n4182) );
  NOR2_X1 U32880 ( .A1(n4212), .A2(n2536), .ZN(n2537) );
  AND2_X1 U32890 ( .A1(n4160), .A2(n2537), .ZN(n2538) );
  INV_X1 U32900 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4308) );
  OR2_X1 U32910 ( .A1(n2398), .A2(n4308), .ZN(n2547) );
  NOR2_X1 U32920 ( .A1(n2541), .A2(REG3_REG_21__SCAN_IN), .ZN(n2542) );
  OR2_X1 U32930 ( .A1(n2543), .A2(n2542), .ZN(n3681) );
  NAND2_X1 U32940 ( .A1(n2355), .A2(REG2_REG_21__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U32950 ( .A1(n2432), .A2(REG0_REG_21__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32960 ( .A1(n4156), .A2(n4147), .ZN(n2549) );
  NOR2_X1 U32970 ( .A1(n4156), .A2(n4147), .ZN(n2548) );
  AOI21_X1 U32980 ( .B1(n4135), .B2(n2549), .A(n2548), .ZN(n4115) );
  INV_X1 U32990 ( .A(n4118), .ZN(n4130) );
  NAND2_X1 U33000 ( .A1(n4139), .A2(n4130), .ZN(n2632) );
  NAND2_X1 U33010 ( .A1(n4292), .A2(n4118), .ZN(n4099) );
  NAND2_X1 U33020 ( .A1(n2632), .A2(n4099), .ZN(n4125) );
  AOI21_X1 U33030 ( .B1(n4118), .B2(n4139), .A(n4117), .ZN(n4098) );
  INV_X1 U33040 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4296) );
  OR2_X1 U33050 ( .A1(n2398), .A2(n4296), .ZN(n2556) );
  NAND2_X1 U33060 ( .A1(n2550), .A2(n3652), .ZN(n2551) );
  NAND2_X1 U33070 ( .A1(n2552), .A2(n2551), .ZN(n4106) );
  OR2_X1 U33080 ( .A1(n2586), .A2(n4106), .ZN(n2555) );
  NAND2_X1 U33090 ( .A1(n2432), .A2(REG0_REG_23__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U33100 ( .A1(n2525), .A2(REG2_REG_23__SCAN_IN), .ZN(n2553) );
  NAND4_X1 U33110 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n4127)
         );
  NAND2_X1 U33120 ( .A1(n3857), .A2(DATAI_23_), .ZN(n4291) );
  NOR2_X1 U33130 ( .A1(n4127), .A2(n4110), .ZN(n2557) );
  INV_X1 U33140 ( .A(n4127), .ZN(n3736) );
  INV_X1 U33150 ( .A(n3956), .ZN(n4281) );
  INV_X1 U33160 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3691) );
  AND2_X1 U33170 ( .A1(n2560), .A2(n3691), .ZN(n2561) );
  OR2_X1 U33180 ( .A1(n2561), .A2(n2566), .ZN(n4074) );
  AOI22_X1 U33190 ( .A1(n2051), .A2(REG1_REG_25__SCAN_IN), .B1(n2432), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U33200 ( .A1(n2525), .A2(REG2_REG_25__SCAN_IN), .ZN(n2562) );
  INV_X1 U33210 ( .A(n4087), .ZN(n3769) );
  NAND2_X1 U33220 ( .A1(n3769), .A2(n4280), .ZN(n2565) );
  NOR2_X1 U33230 ( .A1(n3769), .A2(n4280), .ZN(n2564) );
  NOR2_X1 U33240 ( .A1(n2566), .A2(REG3_REG_26__SCAN_IN), .ZN(n2567) );
  OR2_X1 U33250 ( .A1(n2570), .A2(n2567), .ZN(n3767) );
  AOI22_X1 U33260 ( .A1(n2051), .A2(REG1_REG_26__SCAN_IN), .B1(n2432), .B2(
        REG0_REG_26__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U33270 ( .A1(n2525), .A2(REG2_REG_26__SCAN_IN), .ZN(n2568) );
  OAI211_X1 U33280 ( .C1(n3767), .C2(n2586), .A(n2569), .B(n2568), .ZN(n3955)
         );
  NAND2_X1 U33290 ( .A1(n3857), .A2(DATAI_26_), .ZN(n2636) );
  NAND2_X1 U33300 ( .A1(n3955), .A2(n4061), .ZN(n3867) );
  NOR2_X1 U33310 ( .A1(n3955), .A2(n4061), .ZN(n3869) );
  NOR2_X1 U33320 ( .A1(n2570), .A2(REG3_REG_27__SCAN_IN), .ZN(n2571) );
  INV_X1 U33330 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U33340 ( .A1(n2525), .A2(REG2_REG_27__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U33350 ( .A1(n2432), .A2(REG0_REG_27__SCAN_IN), .ZN(n2572) );
  OAI211_X1 U33360 ( .C1(n2398), .C2(n4274), .A(n2573), .B(n2572), .ZN(n2574)
         );
  INV_X1 U33370 ( .A(n2574), .ZN(n2575) );
  OAI21_X1 U33380 ( .B1(n3642), .B2(n2586), .A(n2575), .ZN(n3954) );
  INV_X1 U33390 ( .A(n3954), .ZN(n4060) );
  NAND2_X1 U33400 ( .A1(n3857), .A2(DATAI_27_), .ZN(n4269) );
  NAND2_X1 U33410 ( .A1(n4060), .A2(n4269), .ZN(n2577) );
  INV_X1 U33420 ( .A(n4269), .ZN(n4049) );
  OR2_X1 U33430 ( .A1(n2578), .A2(REG3_REG_28__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33440 ( .A1(n2578), .A2(REG3_REG_28__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U33450 ( .A1(n4028), .A2(n2352), .ZN(n2585) );
  INV_X1 U33460 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33470 ( .A1(n2525), .A2(REG2_REG_28__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33480 ( .A1(n2432), .A2(REG0_REG_28__SCAN_IN), .ZN(n2580) );
  OAI211_X1 U33490 ( .C1(n2398), .C2(n2582), .A(n2581), .B(n2580), .ZN(n2583)
         );
  INV_X1 U33500 ( .A(n2583), .ZN(n2584) );
  INV_X1 U33510 ( .A(n4029), .ZN(n2916) );
  NAND2_X1 U33520 ( .A1(n3857), .A2(DATAI_29_), .ZN(n3849) );
  OR2_X1 U3353 ( .A1(n4019), .A2(n2586), .ZN(n2591) );
  INV_X1 U33540 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2679) );
  NAND2_X1 U3355 ( .A1(n2432), .A2(REG0_REG_29__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U3356 ( .A1(n2525), .A2(REG2_REG_29__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U3357 ( .C1(n2679), .C2(n2398), .A(n2588), .B(n2587), .ZN(n2589)
         );
  INV_X1 U3358 ( .A(n2589), .ZN(n2590) );
  NAND2_X1 U3359 ( .A1(n2591), .A2(n2590), .ZN(n3953) );
  XNOR2_X1 U3360 ( .A(n2592), .B(n3902), .ZN(n4013) );
  NAND2_X1 U3361 ( .A1(n2594), .A2(n2593), .ZN(n2595) );
  NAND2_X1 U3362 ( .A1(n2595), .A2(IR_REG_31__SCAN_IN), .ZN(n2597) );
  XNOR2_X1 U3363 ( .A(n4417), .B(n3132), .ZN(n2598) );
  NAND2_X1 U3364 ( .A1(n2598), .A2(n4003), .ZN(n4248) );
  AND2_X1 U3365 ( .A1(n2670), .A2(n4420), .ZN(n4563) );
  INV_X1 U3366 ( .A(n4679), .ZN(n4347) );
  AND2_X1 U3367 ( .A1(n4188), .A2(n2669), .ZN(n3836) );
  INV_X1 U3368 ( .A(n2599), .ZN(n3873) );
  INV_X1 U3369 ( .A(n2697), .ZN(n2600) );
  NAND2_X1 U3370 ( .A1(n2600), .A2(n3296), .ZN(n3300) );
  INV_X1 U3371 ( .A(n3300), .ZN(n3794) );
  NAND2_X1 U3372 ( .A1(n3873), .A2(n3794), .ZN(n3299) );
  NAND2_X1 U3373 ( .A1(n3299), .A2(n3795), .ZN(n2602) );
  NAND2_X1 U3374 ( .A1(n2602), .A2(n3874), .ZN(n3328) );
  NAND2_X1 U3375 ( .A1(n3328), .A2(n3796), .ZN(n2603) );
  NAND2_X1 U3376 ( .A1(n2603), .A2(n3912), .ZN(n3348) );
  NAND2_X1 U3377 ( .A1(n3800), .A2(n4643), .ZN(n3801) );
  INV_X1 U3378 ( .A(n3249), .ZN(n2604) );
  NAND2_X1 U3379 ( .A1(n2604), .A2(n3802), .ZN(n2605) );
  NAND2_X1 U3380 ( .A1(n2605), .A2(n3805), .ZN(n3362) );
  AND2_X1 U3381 ( .A1(n3965), .A2(n3421), .ZN(n3361) );
  NAND2_X1 U3382 ( .A1(n3392), .A2(n3714), .ZN(n3809) );
  INV_X1 U3383 ( .A(n3390), .ZN(n3397) );
  NAND2_X1 U3384 ( .A1(n3713), .A2(n3397), .ZN(n3807) );
  NAND2_X1 U3385 ( .A1(n3389), .A2(n3807), .ZN(n2606) );
  INV_X1 U3386 ( .A(n3713), .ZN(n3412) );
  NAND2_X1 U3387 ( .A1(n3412), .A2(n3390), .ZN(n3811) );
  NAND2_X1 U3388 ( .A1(n2606), .A2(n3811), .ZN(n3407) );
  INV_X1 U3389 ( .A(n3812), .ZN(n2607) );
  OAI21_X1 U3390 ( .B1(n3407), .B2(n2607), .A(n3814), .ZN(n3449) );
  INV_X1 U3391 ( .A(n3963), .ZN(n3498) );
  NAND2_X1 U3392 ( .A1(n3498), .A2(n3450), .ZN(n3817) );
  NAND2_X1 U3393 ( .A1(n3449), .A2(n3817), .ZN(n2608) );
  NAND2_X1 U3394 ( .A1(n3963), .A2(n3457), .ZN(n3813) );
  NAND2_X1 U3395 ( .A1(n2608), .A2(n3813), .ZN(n3467) );
  INV_X1 U3396 ( .A(n3473), .ZN(n3497) );
  AND2_X1 U3397 ( .A1(n3483), .A2(n3497), .ZN(n3821) );
  INV_X1 U3398 ( .A(n3483), .ZN(n2609) );
  NAND2_X1 U3399 ( .A1(n2609), .A2(n3473), .ZN(n3818) );
  OAI21_X2 U3400 ( .B1(n3467), .B2(n3821), .A(n3818), .ZN(n3482) );
  NAND2_X1 U3401 ( .A1(n3962), .A2(n3479), .ZN(n3823) );
  NAND2_X1 U3402 ( .A1(n3482), .A2(n3823), .ZN(n2610) );
  NAND2_X1 U3403 ( .A1(n3533), .A2(n3490), .ZN(n3820) );
  NAND2_X1 U3404 ( .A1(n2610), .A2(n3820), .ZN(n3516) );
  NAND2_X1 U3405 ( .A1(n3632), .A2(n3573), .ZN(n3557) );
  NAND2_X1 U3406 ( .A1(n3959), .A2(n2800), .ZN(n2611) );
  NAND2_X1 U3407 ( .A1(n3557), .A2(n2611), .ZN(n2614) );
  INV_X1 U3408 ( .A(n3520), .ZN(n2612) );
  NOR2_X1 U3409 ( .A1(n2614), .A2(n2612), .ZN(n3824) );
  NAND2_X1 U3410 ( .A1(n3516), .A2(n3824), .ZN(n2618) );
  NAND2_X1 U3411 ( .A1(n2613), .A2(n3620), .ZN(n3559) );
  NAND2_X1 U3412 ( .A1(n3518), .A2(n3559), .ZN(n2617) );
  INV_X1 U3413 ( .A(n2614), .ZN(n2616) );
  NOR2_X1 U3414 ( .A1(n3959), .A2(n2800), .ZN(n2615) );
  AOI21_X1 U3415 ( .B1(n2617), .B2(n2616), .A(n2615), .ZN(n3829) );
  NAND2_X2 U3416 ( .A1(n4240), .A2(n4247), .ZN(n4239) );
  NAND2_X1 U3417 ( .A1(n2619), .A2(n3782), .ZN(n3826) );
  NAND2_X1 U3418 ( .A1(n4242), .A2(n4335), .ZN(n3833) );
  NAND2_X1 U3419 ( .A1(n3826), .A2(n3833), .ZN(n3589) );
  INV_X1 U3420 ( .A(n3590), .ZN(n3828) );
  NOR2_X1 U3421 ( .A1(n3589), .A2(n3828), .ZN(n2620) );
  NAND2_X1 U3422 ( .A1(n4239), .A2(n2620), .ZN(n3588) );
  NAND2_X1 U3423 ( .A1(n3588), .A2(n3833), .ZN(n3135) );
  NAND2_X1 U3424 ( .A1(n3135), .A2(n3134), .ZN(n2621) );
  NAND2_X1 U3425 ( .A1(n2621), .A2(n3835), .ZN(n4218) );
  NAND2_X1 U3426 ( .A1(n4203), .A2(n4191), .ZN(n2622) );
  AND2_X1 U3427 ( .A1(n4182), .A2(n2622), .ZN(n2623) );
  NAND2_X1 U3428 ( .A1(n3958), .A2(n4322), .ZN(n4178) );
  NAND2_X1 U3429 ( .A1(n2623), .A2(n4178), .ZN(n3838) );
  OR2_X2 U3430 ( .A1(n4218), .A2(n3838), .ZN(n4154) );
  NAND2_X1 U3431 ( .A1(n4205), .A2(n4231), .ZN(n4179) );
  NAND2_X1 U3432 ( .A1(n4181), .A2(n4179), .ZN(n2624) );
  NAND2_X1 U3433 ( .A1(n2624), .A2(n2623), .ZN(n2626) );
  NAND2_X1 U3434 ( .A1(n4158), .A2(n4187), .ZN(n2625) );
  NAND2_X1 U3435 ( .A1(n2626), .A2(n2625), .ZN(n4152) );
  NOR2_X1 U3436 ( .A1(n4188), .A2(n2669), .ZN(n2628) );
  INV_X1 U3437 ( .A(n3836), .ZN(n2627) );
  OAI21_X1 U3438 ( .B1(n4152), .B2(n2628), .A(n2627), .ZN(n3918) );
  INV_X1 U3439 ( .A(n4156), .ZN(n3755) );
  NAND2_X1 U3440 ( .A1(n3755), .A2(n4147), .ZN(n3919) );
  NAND2_X1 U3441 ( .A1(n4137), .A2(n3919), .ZN(n2631) );
  NAND2_X1 U3442 ( .A1(n4156), .A2(n4303), .ZN(n3924) );
  NAND2_X1 U3443 ( .A1(n2631), .A2(n3924), .ZN(n4126) );
  NAND2_X1 U3444 ( .A1(n4126), .A2(n4099), .ZN(n2633) );
  NAND2_X1 U3445 ( .A1(n4127), .A2(n4291), .ZN(n3890) );
  AND2_X1 U3446 ( .A1(n2632), .A2(n3890), .ZN(n3845) );
  NAND2_X1 U3447 ( .A1(n2633), .A2(n3845), .ZN(n2634) );
  NAND2_X1 U3448 ( .A1(n3736), .A2(n4110), .ZN(n3891) );
  NOR2_X1 U3449 ( .A1(n3956), .A2(n4092), .ZN(n3880) );
  NAND2_X1 U3450 ( .A1(n3956), .A2(n4092), .ZN(n3879) );
  NAND2_X1 U3451 ( .A1(n4087), .A2(n4280), .ZN(n3870) );
  INV_X1 U3452 ( .A(n3870), .ZN(n2635) );
  OR2_X1 U3453 ( .A1(n4087), .A2(n4280), .ZN(n3871) );
  NOR2_X1 U3454 ( .A1(n3955), .A2(n2636), .ZN(n3792) );
  AND2_X1 U3455 ( .A1(n3955), .A2(n2636), .ZN(n3852) );
  AND2_X1 U3456 ( .A1(n3954), .A2(n4269), .ZN(n3854) );
  INV_X1 U3457 ( .A(n3854), .ZN(n2638) );
  OR2_X1 U34580 ( .A1(n3954), .A2(n4269), .ZN(n2639) );
  INV_X1 U34590 ( .A(n2639), .ZN(n3930) );
  AOI21_X1 U3460 ( .B1(n4039), .B2(n4038), .A(n3930), .ZN(n2686) );
  INV_X1 U3461 ( .A(n3931), .ZN(n2640) );
  XNOR2_X1 U3462 ( .A(n2641), .B(n3902), .ZN(n2646) );
  NAND2_X1 U3463 ( .A1(n4417), .A2(n4420), .ZN(n2643) );
  INV_X1 U3464 ( .A(n2670), .ZN(n4419) );
  NAND2_X1 U3465 ( .A1(n4418), .A2(n4419), .ZN(n2642) );
  NAND2_X2 U3466 ( .A1(n2643), .A2(n2642), .ZN(n4564) );
  AOI222_X1 U34670 ( .A1(n2525), .A2(REG2_REG_30__SCAN_IN), .B1(n2051), .B2(
        REG1_REG_30__SCAN_IN), .C1(n2432), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n3863) );
  INV_X1 U3468 ( .A(n3863), .ZN(n3858) );
  AOI21_X1 U34690 ( .B1(B_REG_SCAN_IN), .B2(n4434), .A(n4567), .ZN(n4008) );
  INV_X1 U3470 ( .A(n4008), .ZN(n2644) );
  AOI21_X2 U34710 ( .B1(n2646), .B2(n4564), .A(n2645), .ZN(n4017) );
  NAND2_X1 U3472 ( .A1(n4041), .A2(n4644), .ZN(n2647) );
  NAND2_X1 U34730 ( .A1(n3945), .A2(n2653), .ZN(n4561) );
  NAND2_X1 U3474 ( .A1(n4017), .A2(n2648), .ZN(n2649) );
  AOI21_X1 U34750 ( .B1(n4013), .B2(n4664), .A(n2649), .ZN(n2678) );
  NAND2_X1 U3476 ( .A1(n3163), .A2(B_REG_SCAN_IN), .ZN(n2650) );
  MUX2_X1 U34770 ( .A(n2650), .B(B_REG_SCAN_IN), .S(n4416), .Z(n2651) );
  NAND2_X1 U3478 ( .A1(n2651), .A2(n4415), .ZN(n3159) );
  OAI22_X1 U34790 ( .A1(n3159), .A2(D_REG_1__SCAN_IN), .B1(n2652), .B2(n4415), 
        .ZN(n2922) );
  NAND2_X1 U3480 ( .A1(n4679), .A2(n2653), .ZN(n2944) );
  AND2_X1 U34810 ( .A1(n2922), .A2(n2944), .ZN(n2665) );
  NOR4_X1 U3482 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2657) );
  NOR4_X1 U34830 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2656) );
  NOR4_X1 U3484 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2655) );
  NOR4_X1 U34850 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2654) );
  NAND4_X1 U3486 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n2663)
         );
  NOR2_X1 U34870 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_8__SCAN_IN), .ZN(n2661)
         );
  NOR4_X1 U3488 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2660) );
  NOR4_X1 U34890 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2659) );
  NOR4_X1 U3490 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2658) );
  NAND4_X1 U34910 ( .A1(n2661), .A2(n2660), .A3(n2659), .A4(n2658), .ZN(n2662)
         );
  INV_X1 U3492 ( .A(n3159), .ZN(n2668) );
  OAI21_X1 U34930 ( .B1(n2663), .B2(n2662), .A(n2668), .ZN(n2923) );
  NAND2_X1 U3494 ( .A1(n2670), .A2(n4003), .ZN(n2926) );
  AND2_X1 U34950 ( .A1(n2925), .A2(n2926), .ZN(n2936) );
  NOR2_X1 U3496 ( .A1(n3158), .A2(n2936), .ZN(n2664) );
  AND2_X1 U34970 ( .A1(n2923), .A2(n2664), .ZN(n3129) );
  INV_X1 U3498 ( .A(D_REG_0__SCAN_IN), .ZN(n2667) );
  INV_X1 U34990 ( .A(n4415), .ZN(n3164) );
  INV_X1 U3500 ( .A(n4416), .ZN(n3160) );
  INV_X1 U35010 ( .A(n2924), .ZN(n3130) );
  OR2_X1 U3502 ( .A1(n2678), .A2(n4683), .ZN(n2676) );
  INV_X1 U35030 ( .A(n3296), .ZN(n4562) );
  NAND2_X1 U3504 ( .A1(n3458), .A2(n3457), .ZN(n3459) );
  OAI21_X1 U35050 ( .B1(n2692), .B2(n3849), .A(n4263), .ZN(n4020) );
  INV_X1 U35060 ( .A(n4561), .ZN(n2671) );
  INV_X1 U35080 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2672) );
  OR2_X1 U35090 ( .A1(n4685), .A2(n2672), .ZN(n2673) );
  NAND2_X1 U35100 ( .A1(n2676), .A2(n2675), .ZN(U3515) );
  OR2_X1 U35110 ( .A1(n2678), .A2(n4702), .ZN(n2683) );
  OR2_X1 U35120 ( .A1(n4704), .A2(n2679), .ZN(n2680) );
  NAND2_X1 U35130 ( .A1(n2683), .A2(n2682), .ZN(U3547) );
  XNOR2_X1 U35140 ( .A(n2684), .B(n3901), .ZN(n4026) );
  INV_X1 U35150 ( .A(n4664), .ZN(n4332) );
  XNOR2_X1 U35160 ( .A(n2686), .B(n2685), .ZN(n2688) );
  AOI21_X2 U35170 ( .B1(n2688), .B2(n4564), .A(n2687), .ZN(n4032) );
  AOI22_X1 U35180 ( .A1(n3954), .A2(n4644), .B1(n4029), .B2(n4642), .ZN(n2689)
         );
  OAI211_X1 U35190 ( .C1(n4026), .C2(n4332), .A(n4032), .B(n2689), .ZN(n2694)
         );
  MUX2_X1 U35200 ( .A(REG1_REG_28__SCAN_IN), .B(n2694), .S(n4704), .Z(n2690)
         );
  INV_X1 U35210 ( .A(n2690), .ZN(n2693) );
  NOR2_X1 U35220 ( .A1(n4044), .A2(n2916), .ZN(n2691) );
  NAND2_X1 U35230 ( .A1(n2693), .A2(n2171), .ZN(U3546) );
  MUX2_X1 U35240 ( .A(REG0_REG_28__SCAN_IN), .B(n2694), .S(n4685), .Z(n2695)
         );
  INV_X1 U35250 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U35260 ( .A1(n2696), .A2(n2172), .ZN(U3514) );
  INV_X1 U35270 ( .A(n3132), .ZN(n2698) );
  NAND2_X1 U35280 ( .A1(n3126), .A2(n2698), .ZN(n2720) );
  INV_X1 U35290 ( .A(n3126), .ZN(n2700) );
  NAND2_X1 U35300 ( .A1(n2700), .A2(REG1_REG_0__SCAN_IN), .ZN(n2699) );
  NAND2_X1 U35310 ( .A1(n2703), .A2(n2699), .ZN(n3200) );
  AOI22_X1 U35320 ( .A1(n3296), .A2(n2942), .B1(IR_REG_0__SCAN_IN), .B2(n2700), 
        .ZN(n2701) );
  NAND2_X1 U35330 ( .A1(n2702), .A2(n2701), .ZN(n3199) );
  NAND2_X1 U35340 ( .A1(n3200), .A2(n3199), .ZN(n3198) );
  NAND2_X1 U35360 ( .A1(n2703), .A2(n2909), .ZN(n2704) );
  NAND2_X1 U35370 ( .A1(n3198), .A2(n2704), .ZN(n3669) );
  OAI22_X1 U35380 ( .A1(n2705), .A2(n2911), .B1(n2707), .B2(n2913), .ZN(n2706)
         );
  XNOR2_X1 U35390 ( .A(n2706), .B(n2909), .ZN(n2708) );
  OAI22_X1 U35400 ( .A1(n2705), .A2(n2917), .B1(n2707), .B2(n2911), .ZN(n2709)
         );
  XNOR2_X1 U35410 ( .A(n2708), .B(n2709), .ZN(n3667) );
  NAND2_X1 U35420 ( .A1(n3669), .A2(n3667), .ZN(n3668) );
  INV_X1 U35430 ( .A(n2708), .ZN(n2710) );
  NAND2_X1 U35440 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND2_X1 U35450 ( .A1(n3668), .A2(n2711), .ZN(n3222) );
  INV_X1 U35460 ( .A(n3222), .ZN(n2714) );
  OAI22_X1 U35480 ( .A1(n2372), .A2(n2825), .B1(n3340), .B2(n2913), .ZN(n2712)
         );
  XNOR2_X1 U35490 ( .A(n2712), .B(n2914), .ZN(n2715) );
  OAI22_X1 U35500 ( .A1(n2372), .A2(n2917), .B1(n3340), .B2(n2911), .ZN(n2716)
         );
  XNOR2_X1 U35510 ( .A(n2715), .B(n2716), .ZN(n3223) );
  INV_X1 U35520 ( .A(n3223), .ZN(n2713) );
  NAND2_X1 U35530 ( .A1(n2714), .A2(n2713), .ZN(n3220) );
  INV_X1 U35540 ( .A(n2715), .ZN(n2718) );
  INV_X1 U35550 ( .A(n2716), .ZN(n2717) );
  NAND2_X1 U35560 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  NAND2_X2 U35570 ( .A1(n3220), .A2(n2719), .ZN(n3279) );
  NAND2_X1 U35580 ( .A1(n3714), .A2(n2906), .ZN(n2722) );
  NAND2_X1 U35590 ( .A1(n2722), .A2(n2721), .ZN(n2723) );
  AOI22_X1 U35600 ( .A1(n3965), .A2(n2897), .B1(n3714), .B2(n2942), .ZN(n2740)
         );
  OAI22_X1 U35610 ( .A1(n3420), .A2(n2825), .B1(n2913), .B2(n3254), .ZN(n2724)
         );
  XNOR2_X1 U35620 ( .A(n2724), .B(n2914), .ZN(n2734) );
  OAI22_X1 U35630 ( .A1(n3420), .A2(n2917), .B1(n2825), .B2(n3254), .ZN(n2732)
         );
  NAND2_X1 U35640 ( .A1(n2734), .A2(n2732), .ZN(n3708) );
  INV_X1 U35650 ( .A(n3708), .ZN(n2725) );
  NAND2_X1 U35660 ( .A1(n4643), .A2(n2906), .ZN(n2726) );
  XNOR2_X1 U35670 ( .A(n2727), .B(n2914), .ZN(n2729) );
  AOI22_X1 U35680 ( .A1(n3966), .A2(n2897), .B1(n4643), .B2(n2942), .ZN(n2730)
         );
  XNOR2_X1 U35690 ( .A(n2729), .B(n2730), .ZN(n3278) );
  NAND2_X1 U35700 ( .A1(n3279), .A2(n2728), .ZN(n2739) );
  INV_X1 U35710 ( .A(n2729), .ZN(n2731) );
  NAND2_X1 U35720 ( .A1(n2731), .A2(n2730), .ZN(n3280) );
  XNOR2_X1 U35730 ( .A(n2734), .B(n2733), .ZN(n3277) );
  NAND2_X1 U35740 ( .A1(n2739), .A2(n2738), .ZN(n3711) );
  INV_X1 U35750 ( .A(n2740), .ZN(n2741) );
  NAND2_X1 U35760 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  NAND2_X1 U35770 ( .A1(n3711), .A2(n2743), .ZN(n3260) );
  NAND2_X1 U35780 ( .A1(n3713), .A2(n2942), .ZN(n2745) );
  NAND2_X1 U35790 ( .A1(n3390), .A2(n2906), .ZN(n2744) );
  NAND2_X1 U35800 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  XNOR2_X1 U35810 ( .A(n2746), .B(n2914), .ZN(n3311) );
  NAND2_X1 U3582 ( .A1(n3713), .A2(n2897), .ZN(n2748) );
  NAND2_X1 U3583 ( .A1(n3390), .A2(n2942), .ZN(n2747) );
  NAND2_X1 U3584 ( .A1(n2748), .A2(n2747), .ZN(n3312) );
  OAI22_X1 U3585 ( .A1(n3452), .A2(n2911), .B1(n2749), .B2(n2913), .ZN(n2750)
         );
  XNOR2_X1 U3586 ( .A(n2750), .B(n2909), .ZN(n3318) );
  AND2_X1 U3587 ( .A1(n3409), .A2(n2942), .ZN(n2751) );
  AOI21_X1 U3588 ( .B1(n3964), .B2(n2897), .A(n2751), .ZN(n2754) );
  NAND2_X1 U3589 ( .A1(n3318), .A2(n2754), .ZN(n2757) );
  INV_X1 U3590 ( .A(n2752), .ZN(n2753) );
  AND2_X1 U3591 ( .A1(n3311), .A2(n3312), .ZN(n2756) );
  INV_X1 U3592 ( .A(n3318), .ZN(n2755) );
  INV_X1 U3593 ( .A(n2754), .ZN(n3317) );
  AOI22_X1 U3594 ( .A1(n2757), .A2(n2756), .B1(n2755), .B2(n3317), .ZN(n2758)
         );
  NAND2_X1 U3595 ( .A1(n3963), .A2(n2942), .ZN(n2760) );
  NAND2_X1 U3596 ( .A1(n3450), .A2(n2906), .ZN(n2759) );
  NAND2_X1 U3597 ( .A1(n2760), .A2(n2759), .ZN(n2761) );
  XNOR2_X1 U3598 ( .A(n2761), .B(n2914), .ZN(n2765) );
  NAND2_X1 U3599 ( .A1(n3963), .A2(n2897), .ZN(n2763) );
  NAND2_X1 U3600 ( .A1(n3450), .A2(n2942), .ZN(n2762) );
  NAND2_X1 U3601 ( .A1(n2763), .A2(n2762), .ZN(n2766) );
  AND2_X1 U3602 ( .A1(n2765), .A2(n2766), .ZN(n3269) );
  INV_X1 U3603 ( .A(n3269), .ZN(n2764) );
  INV_X1 U3604 ( .A(n2765), .ZN(n2768) );
  INV_X1 U3605 ( .A(n2766), .ZN(n2767) );
  NAND2_X1 U3606 ( .A1(n2768), .A2(n2767), .ZN(n3268) );
  NAND2_X1 U3607 ( .A1(n2769), .A2(n3268), .ZN(n3432) );
  NAND2_X1 U3608 ( .A1(n3483), .A2(n2942), .ZN(n2771) );
  NAND2_X1 U3609 ( .A1(n3473), .A2(n2906), .ZN(n2770) );
  NAND2_X1 U3610 ( .A1(n2771), .A2(n2770), .ZN(n2772) );
  XNOR2_X1 U3611 ( .A(n2772), .B(n2914), .ZN(n2776) );
  AOI22_X1 U3612 ( .A1(n3483), .A2(n2897), .B1(n3473), .B2(n2942), .ZN(n2777)
         );
  XNOR2_X1 U3613 ( .A(n2776), .B(n2777), .ZN(n3433) );
  NAND2_X1 U3614 ( .A1(n3432), .A2(n3433), .ZN(n3431) );
  NAND2_X1 U3615 ( .A1(n3962), .A2(n2942), .ZN(n2774) );
  NAND2_X1 U3616 ( .A1(n3490), .A2(n2906), .ZN(n2773) );
  NAND2_X1 U3617 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  XNOR2_X1 U3618 ( .A(n2775), .B(n2914), .ZN(n2780) );
  AOI22_X1 U3619 ( .A1(n3962), .A2(n2897), .B1(n2942), .B2(n3490), .ZN(n2781)
         );
  XNOR2_X1 U3620 ( .A(n2780), .B(n2781), .ZN(n3440) );
  INV_X1 U3621 ( .A(n2776), .ZN(n2778) );
  NAND2_X1 U3622 ( .A1(n2778), .A2(n2777), .ZN(n3441) );
  AND2_X1 U3623 ( .A1(n3440), .A2(n3441), .ZN(n2779) );
  INV_X1 U3624 ( .A(n2780), .ZN(n2782) );
  OAI22_X1 U3625 ( .A1(n3621), .A2(n2825), .B1(n2786), .B2(n2913), .ZN(n2785)
         );
  XNOR2_X1 U3626 ( .A(n2785), .B(n2914), .ZN(n2787) );
  OAI22_X1 U3627 ( .A1(n3621), .A2(n2917), .B1(n2786), .B2(n2911), .ZN(n2788)
         );
  AND2_X1 U3628 ( .A1(n2787), .A2(n2788), .ZN(n3629) );
  INV_X1 U3629 ( .A(n2787), .ZN(n2790) );
  INV_X1 U3630 ( .A(n2788), .ZN(n2789) );
  NAND2_X1 U3631 ( .A1(n2790), .A2(n2789), .ZN(n3628) );
  NAND2_X1 U3632 ( .A1(n2791), .A2(n3628), .ZN(n3619) );
  INV_X1 U3633 ( .A(n3619), .ZN(n2798) );
  NAND2_X1 U3634 ( .A1(n3632), .A2(n2942), .ZN(n2793) );
  NAND2_X1 U3635 ( .A1(n3620), .A2(n2906), .ZN(n2792) );
  NAND2_X1 U3636 ( .A1(n2793), .A2(n2792), .ZN(n2794) );
  XNOR2_X1 U3637 ( .A(n2794), .B(n2909), .ZN(n3617) );
  AND2_X1 U3638 ( .A1(n3620), .A2(n2942), .ZN(n2795) );
  AOI21_X1 U3639 ( .B1(n3632), .B2(n2897), .A(n2795), .ZN(n3616) );
  INV_X1 U3640 ( .A(n3617), .ZN(n2797) );
  INV_X1 U3641 ( .A(n3616), .ZN(n2796) );
  OAI22_X1 U3642 ( .A1(n4244), .A2(n2825), .B1(n2913), .B2(n2800), .ZN(n2799)
         );
  XNOR2_X1 U3643 ( .A(n2799), .B(n2914), .ZN(n2801) );
  OAI22_X1 U3644 ( .A1(n4244), .A2(n2917), .B1(n2825), .B2(n2800), .ZN(n2802)
         );
  NAND2_X1 U3645 ( .A1(n2801), .A2(n2802), .ZN(n3509) );
  NAND2_X1 U3646 ( .A1(n3507), .A2(n3509), .ZN(n2805) );
  INV_X1 U3647 ( .A(n2801), .ZN(n2804) );
  INV_X1 U3648 ( .A(n2802), .ZN(n2803) );
  NAND2_X1 U3649 ( .A1(n2804), .A2(n2803), .ZN(n3508) );
  NAND2_X1 U3650 ( .A1(n2805), .A2(n3508), .ZN(n3545) );
  OAI22_X1 U3651 ( .A1(n4337), .A2(n2825), .B1(n2913), .B2(n2807), .ZN(n2806)
         );
  XNOR2_X1 U3652 ( .A(n2806), .B(n2909), .ZN(n2808) );
  OAI22_X1 U3653 ( .A1(n4337), .A2(n2917), .B1(n2825), .B2(n2807), .ZN(n3546)
         );
  INV_X1 U3654 ( .A(n2808), .ZN(n3547) );
  NAND2_X1 U3655 ( .A1(n4242), .A2(n2942), .ZN(n2810) );
  NAND2_X1 U3656 ( .A1(n3782), .A2(n2906), .ZN(n2809) );
  NAND2_X1 U3657 ( .A1(n2810), .A2(n2809), .ZN(n2811) );
  XNOR2_X1 U3658 ( .A(n2811), .B(n2914), .ZN(n2817) );
  NAND2_X1 U3659 ( .A1(n2813), .A2(n2812), .ZN(n3697) );
  NAND2_X1 U3660 ( .A1(n4242), .A2(n2897), .ZN(n2815) );
  NAND2_X1 U3661 ( .A1(n3782), .A2(n2942), .ZN(n2814) );
  NAND2_X1 U3662 ( .A1(n2815), .A2(n2814), .ZN(n3777) );
  NAND2_X1 U3663 ( .A1(n3697), .A2(n3777), .ZN(n2819) );
  OAI22_X1 U3664 ( .A1(n4323), .A2(n2825), .B1(n2913), .B2(n3140), .ZN(n2816)
         );
  XNOR2_X1 U3665 ( .A(n2816), .B(n2909), .ZN(n2822) );
  OAI22_X1 U3666 ( .A1(n4323), .A2(n2917), .B1(n2825), .B2(n3140), .ZN(n2820)
         );
  XNOR2_X1 U3667 ( .A(n2822), .B(n2820), .ZN(n3700) );
  NAND2_X1 U3668 ( .A1(n2818), .A2(n2817), .ZN(n3776) );
  NAND3_X1 U3669 ( .A1(n2819), .A2(n3700), .A3(n3776), .ZN(n2824) );
  INV_X1 U3670 ( .A(n2820), .ZN(n2821) );
  NAND2_X1 U3671 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  NAND2_X1 U3672 ( .A1(n2824), .A2(n2823), .ZN(n3721) );
  OAI22_X1 U3673 ( .A1(n4205), .A2(n2825), .B1(n4322), .B2(n2913), .ZN(n2826)
         );
  XNOR2_X1 U3674 ( .A(n2826), .B(n2909), .ZN(n3723) );
  NOR2_X1 U3675 ( .A1(n4322), .A2(n2911), .ZN(n2827) );
  AOI21_X1 U3676 ( .B1(n3958), .B2(n2897), .A(n2827), .ZN(n3722) );
  AND2_X1 U3677 ( .A1(n3723), .A2(n3722), .ZN(n2828) );
  OAI22_X1 U3678 ( .A1(n4220), .A2(n2825), .B1(n2913), .B2(n4199), .ZN(n2829)
         );
  XNOR2_X1 U3679 ( .A(n2829), .B(n2914), .ZN(n2830) );
  OAI22_X1 U3680 ( .A1(n4220), .A2(n2917), .B1(n2825), .B2(n4199), .ZN(n2831)
         );
  AND2_X1 U3681 ( .A1(n2830), .A2(n2831), .ZN(n3608) );
  INV_X1 U3682 ( .A(n2830), .ZN(n2833) );
  INV_X1 U3683 ( .A(n2831), .ZN(n2832) );
  NAND2_X1 U3684 ( .A1(n2833), .A2(n2832), .ZN(n3607) );
  NAND2_X1 U3685 ( .A1(n4203), .A2(n2942), .ZN(n2835) );
  NAND2_X1 U3686 ( .A1(n4187), .A2(n2906), .ZN(n2834) );
  NAND2_X1 U3687 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  XNOR2_X1 U3688 ( .A(n2836), .B(n2914), .ZN(n2837) );
  AOI22_X1 U3689 ( .A1(n4203), .A2(n2897), .B1(n2942), .B2(n4187), .ZN(n2838)
         );
  XNOR2_X1 U3690 ( .A(n2837), .B(n2838), .ZN(n3661) );
  NAND2_X1 U3691 ( .A1(n3659), .A2(n3661), .ZN(n2841) );
  INV_X1 U3692 ( .A(n2837), .ZN(n2839) );
  NAND2_X1 U3693 ( .A1(n2839), .A2(n2838), .ZN(n2840) );
  NAND2_X1 U3694 ( .A1(n2841), .A2(n2840), .ZN(n3675) );
  NAND2_X1 U3695 ( .A1(n4188), .A2(n2942), .ZN(n2843) );
  NAND2_X1 U3696 ( .A1(n4172), .A2(n2906), .ZN(n2842) );
  NAND2_X1 U3697 ( .A1(n2843), .A2(n2842), .ZN(n2844) );
  XNOR2_X1 U3698 ( .A(n2844), .B(n2914), .ZN(n2847) );
  NAND2_X1 U3699 ( .A1(n4188), .A2(n2897), .ZN(n2846) );
  NAND2_X1 U3700 ( .A1(n4172), .A2(n2942), .ZN(n2845) );
  NAND2_X1 U3701 ( .A1(n2846), .A2(n2845), .ZN(n2848) );
  NAND2_X1 U3702 ( .A1(n2847), .A2(n2848), .ZN(n3743) );
  NAND2_X1 U3703 ( .A1(n3675), .A2(n3743), .ZN(n2857) );
  INV_X1 U3704 ( .A(n2847), .ZN(n2850) );
  INV_X1 U3705 ( .A(n2848), .ZN(n2849) );
  NAND2_X1 U3706 ( .A1(n2850), .A2(n2849), .ZN(n3742) );
  NAND2_X1 U3707 ( .A1(n4156), .A2(n2942), .ZN(n2852) );
  NAND2_X1 U3708 ( .A1(n4147), .A2(n2906), .ZN(n2851) );
  NAND2_X1 U3709 ( .A1(n2852), .A2(n2851), .ZN(n2853) );
  XNOR2_X1 U3710 ( .A(n2853), .B(n2909), .ZN(n3678) );
  NOR2_X1 U3711 ( .A1(n4303), .A2(n2911), .ZN(n2854) );
  AOI21_X1 U3712 ( .B1(n4156), .B2(n2897), .A(n2854), .ZN(n2858) );
  NAND2_X1 U3713 ( .A1(n3678), .A2(n2858), .ZN(n2855) );
  AND2_X1 U3714 ( .A1(n3742), .A2(n2855), .ZN(n2856) );
  NAND2_X1 U3715 ( .A1(n2857), .A2(n2856), .ZN(n2861) );
  INV_X1 U3716 ( .A(n3678), .ZN(n2859) );
  INV_X1 U3717 ( .A(n2858), .ZN(n3677) );
  NAND2_X1 U3718 ( .A1(n2859), .A2(n3677), .ZN(n2860) );
  OAI22_X1 U3719 ( .A1(n4292), .A2(n2911), .B1(n2913), .B2(n4130), .ZN(n2862)
         );
  XNOR2_X1 U3720 ( .A(n2862), .B(n2914), .ZN(n2867) );
  OAI22_X1 U3721 ( .A1(n4292), .A2(n2917), .B1(n2825), .B2(n4130), .ZN(n2868)
         );
  XNOR2_X1 U3722 ( .A(n2867), .B(n2868), .ZN(n3753) );
  NAND2_X1 U3723 ( .A1(n4127), .A2(n2942), .ZN(n2864) );
  NAND2_X1 U3724 ( .A1(n4110), .A2(n2906), .ZN(n2863) );
  NAND2_X1 U3725 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
  XNOR2_X1 U3726 ( .A(n2865), .B(n2914), .ZN(n2874) );
  NOR2_X1 U3727 ( .A1(n4291), .A2(n2825), .ZN(n2866) );
  AOI21_X1 U3728 ( .B1(n4127), .B2(n2897), .A(n2866), .ZN(n2872) );
  XNOR2_X1 U3729 ( .A(n2874), .B(n2872), .ZN(n3650) );
  INV_X1 U3730 ( .A(n2867), .ZN(n2870) );
  INV_X1 U3731 ( .A(n2868), .ZN(n2869) );
  NAND2_X1 U3732 ( .A1(n2870), .A2(n2869), .ZN(n3651) );
  INV_X1 U3733 ( .A(n2872), .ZN(n2873) );
  NAND2_X1 U3734 ( .A1(n2874), .A2(n2873), .ZN(n2881) );
  NAND2_X1 U3735 ( .A1(n3956), .A2(n2942), .ZN(n2876) );
  NAND2_X1 U3736 ( .A1(n3734), .A2(n2906), .ZN(n2875) );
  NAND2_X1 U3737 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  XNOR2_X1 U3738 ( .A(n2877), .B(n2909), .ZN(n2882) );
  AND2_X1 U3739 ( .A1(n2881), .A2(n2882), .ZN(n2878) );
  NAND2_X1 U3740 ( .A1(n3956), .A2(n2897), .ZN(n2880) );
  NAND2_X1 U3741 ( .A1(n3734), .A2(n2942), .ZN(n2879) );
  NAND2_X1 U3742 ( .A1(n2880), .A2(n2879), .ZN(n3732) );
  NAND2_X1 U3743 ( .A1(n3730), .A2(n3732), .ZN(n2885) );
  INV_X1 U3744 ( .A(n2882), .ZN(n2883) );
  NAND2_X1 U3745 ( .A1(n2884), .A2(n2883), .ZN(n3729) );
  NAND2_X1 U3746 ( .A1(n2885), .A2(n3729), .ZN(n3688) );
  NAND2_X1 U3747 ( .A1(n4087), .A2(n2942), .ZN(n2887) );
  NAND2_X1 U3748 ( .A1(n4078), .A2(n2906), .ZN(n2886) );
  NAND2_X1 U3749 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  XNOR2_X1 U3750 ( .A(n2888), .B(n2909), .ZN(n2890) );
  NOR2_X1 U3751 ( .A1(n4280), .A2(n2911), .ZN(n2889) );
  AOI21_X1 U3752 ( .B1(n4087), .B2(n2897), .A(n2889), .ZN(n2891) );
  NAND2_X1 U3753 ( .A1(n2890), .A2(n2891), .ZN(n3687) );
  INV_X1 U3754 ( .A(n2890), .ZN(n2893) );
  INV_X1 U3755 ( .A(n2891), .ZN(n2892) );
  NAND2_X1 U3756 ( .A1(n2893), .A2(n2892), .ZN(n3762) );
  NAND2_X1 U3757 ( .A1(n3955), .A2(n2942), .ZN(n2895) );
  NAND2_X1 U3758 ( .A1(n4061), .A2(n2906), .ZN(n2894) );
  NAND2_X1 U3759 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  XNOR2_X1 U3760 ( .A(n2896), .B(n2914), .ZN(n2902) );
  NAND2_X1 U3761 ( .A1(n3955), .A2(n2897), .ZN(n2899) );
  NAND2_X1 U3762 ( .A1(n4061), .A2(n2942), .ZN(n2898) );
  NAND2_X1 U3763 ( .A1(n2899), .A2(n2898), .ZN(n2903) );
  AND2_X1 U3764 ( .A1(n2902), .A2(n2903), .ZN(n3764) );
  INV_X1 U3765 ( .A(n3764), .ZN(n2900) );
  AND2_X1 U3766 ( .A1(n3762), .A2(n2900), .ZN(n2901) );
  INV_X1 U3767 ( .A(n2902), .ZN(n2905) );
  INV_X1 U3768 ( .A(n2903), .ZN(n2904) );
  NAND2_X1 U3769 ( .A1(n2905), .A2(n2904), .ZN(n3763) );
  NAND2_X1 U3770 ( .A1(n3954), .A2(n2942), .ZN(n2908) );
  NAND2_X1 U3771 ( .A1(n4049), .A2(n2906), .ZN(n2907) );
  NAND2_X1 U3772 ( .A1(n2908), .A2(n2907), .ZN(n2910) );
  XNOR2_X1 U3773 ( .A(n2910), .B(n2909), .ZN(n2921) );
  NOR2_X1 U3774 ( .A1(n4269), .A2(n2911), .ZN(n2912) );
  AOI21_X1 U3775 ( .B1(n3954), .B2(n2897), .A(n2912), .ZN(n2920) );
  XNOR2_X1 U3776 ( .A(n2921), .B(n2920), .ZN(n3641) );
  OAI22_X1 U3777 ( .A1(n4014), .A2(n2911), .B1(n2913), .B2(n2916), .ZN(n2915)
         );
  XNOR2_X1 U3778 ( .A(n2915), .B(n2914), .ZN(n2919) );
  OAI22_X1 U3779 ( .A1(n4014), .A2(n2917), .B1(n2825), .B2(n2916), .ZN(n2918)
         );
  XNOR2_X1 U3780 ( .A(n2919), .B(n2918), .ZN(n2953) );
  NOR2_X1 U3781 ( .A1(n2921), .A2(n2920), .ZN(n2934) );
  INV_X1 U3782 ( .A(n2922), .ZN(n3128) );
  NAND3_X1 U3783 ( .A1(n3128), .A2(n2924), .A3(n2923), .ZN(n2943) );
  OR2_X1 U3784 ( .A1(n2943), .A2(n3158), .ZN(n2945) );
  INV_X1 U3785 ( .A(n2945), .ZN(n2931) );
  INV_X1 U3786 ( .A(n2925), .ZN(n2929) );
  INV_X1 U3787 ( .A(n2926), .ZN(n2927) );
  OR2_X1 U3788 ( .A1(n4561), .A2(n2927), .ZN(n2928) );
  AND2_X1 U3789 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  NOR2_X1 U3790 ( .A1(n2934), .A2(n3740), .ZN(n2932) );
  INV_X1 U3791 ( .A(n2934), .ZN(n2935) );
  NOR3_X1 U3792 ( .A1(n2933), .A2(n3740), .A3(n2935), .ZN(n2951) );
  INV_X1 U3793 ( .A(n4028), .ZN(n2949) );
  AOI21_X1 U3794 ( .B1(n2943), .B2(n2944), .A(n2936), .ZN(n3225) );
  NAND3_X1 U3795 ( .A1(n3225), .A2(n3126), .A3(n2937), .ZN(n2938) );
  INV_X1 U3796 ( .A(n2939), .ZN(n2940) );
  AND2_X1 U3797 ( .A1(n4605), .A2(n2940), .ZN(n2941) );
  NAND2_X1 U3798 ( .A1(n2942), .A2(n2941), .ZN(n3949) );
  NOR2_X2 U3799 ( .A1(n2946), .A2(n3202), .ZN(n3787) );
  AOI22_X1 U3800 ( .A1(n3954), .A2(n3787), .B1(n3781), .B2(n4029), .ZN(n2948)
         );
  AOI22_X1 U3801 ( .A1(n3953), .A2(n3780), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2947) );
  OAI211_X1 U3802 ( .C1(n2949), .C2(n3784), .A(n2948), .B(n2947), .ZN(n2950)
         );
  NOR2_X1 U3803 ( .A1(n2952), .A2(n2073), .ZN(n2955) );
  NAND3_X1 U3804 ( .A1(n2068), .A2(n3710), .A3(n2953), .ZN(n2954) );
  NAND2_X1 U3805 ( .A1(n2955), .A2(n2954), .ZN(n3124) );
  OAI22_X1 U3806 ( .A1(DATAI_16_), .A2(keyinput102), .B1(DATAI_18_), .B2(
        keyinput110), .ZN(n2956) );
  AOI221_X1 U3807 ( .B1(DATAI_16_), .B2(keyinput102), .C1(keyinput110), .C2(
        DATAI_18_), .A(n2956), .ZN(n2963) );
  OAI22_X1 U3808 ( .A1(DATAI_3_), .A2(keyinput85), .B1(keyinput100), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n2957) );
  AOI221_X1 U3809 ( .B1(DATAI_3_), .B2(keyinput85), .C1(DATAO_REG_9__SCAN_IN), 
        .C2(keyinput100), .A(n2957), .ZN(n2962) );
  OAI22_X1 U3810 ( .A1(DATAI_29_), .A2(keyinput115), .B1(keyinput87), .B2(
        DATAI_30_), .ZN(n2958) );
  AOI221_X1 U3811 ( .B1(DATAI_29_), .B2(keyinput115), .C1(DATAI_30_), .C2(
        keyinput87), .A(n2958), .ZN(n2961) );
  OAI22_X1 U3812 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput123), .B1(DATAI_26_), 
        .B2(keyinput74), .ZN(n2959) );
  AOI221_X1 U3813 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput123), .C1(keyinput74), 
        .C2(DATAI_26_), .A(n2959), .ZN(n2960) );
  NAND4_X1 U3814 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), .ZN(n2972)
         );
  INV_X1 U3815 ( .A(DATAI_20_), .ZN(n3107) );
  INV_X1 U3816 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U3817 ( .A1(n3107), .A2(keyinput69), .B1(keyinput64), .B2(n4650), 
        .ZN(n2964) );
  OAI221_X1 U3818 ( .B1(n3107), .B2(keyinput69), .C1(n4650), .C2(keyinput64), 
        .A(n2964), .ZN(n2971) );
  INV_X1 U3819 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U3820 ( .A1(n3180), .A2(keyinput122), .B1(n3652), .B2(keyinput75), 
        .ZN(n2965) );
  OAI221_X1 U3821 ( .B1(n3180), .B2(keyinput122), .C1(n3652), .C2(keyinput75), 
        .A(n2965), .ZN(n2970) );
  XNOR2_X1 U3822 ( .A(IR_REG_6__SCAN_IN), .B(keyinput88), .ZN(n2968) );
  XNOR2_X1 U3823 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput68), .ZN(n2967) );
  XNOR2_X1 U3824 ( .A(IR_REG_25__SCAN_IN), .B(keyinput78), .ZN(n2966) );
  NAND3_X1 U3825 ( .A1(n2968), .A2(n2967), .A3(n2966), .ZN(n2969) );
  OR4_X1 U3826 ( .A1(n2972), .A2(n2971), .A3(n2970), .A4(n2969), .ZN(n2986) );
  OAI22_X1 U3827 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput107), .B1(keyinput105), .B2(DATAI_24_), .ZN(n2973) );
  AOI221_X1 U3828 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput107), .C1(DATAI_24_), 
        .C2(keyinput105), .A(n2973), .ZN(n2980) );
  OAI22_X1 U3829 ( .A1(DATAI_25_), .A2(keyinput106), .B1(keyinput96), .B2(
        DATAI_23_), .ZN(n2974) );
  AOI221_X1 U3830 ( .B1(DATAI_25_), .B2(keyinput106), .C1(DATAI_23_), .C2(
        keyinput96), .A(n2974), .ZN(n2979) );
  OAI22_X1 U3831 ( .A1(REG0_REG_20__SCAN_IN), .A2(keyinput108), .B1(
        REG0_REG_17__SCAN_IN), .B2(keyinput109), .ZN(n2975) );
  AOI221_X1 U3832 ( .B1(REG0_REG_20__SCAN_IN), .B2(keyinput108), .C1(
        keyinput109), .C2(REG0_REG_17__SCAN_IN), .A(n2975), .ZN(n2978) );
  OAI22_X1 U3833 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput118), .B1(
        REG0_REG_24__SCAN_IN), .B2(keyinput113), .ZN(n2976) );
  AOI221_X1 U3834 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput118), .C1(keyinput113), 
        .C2(REG0_REG_24__SCAN_IN), .A(n2976), .ZN(n2977) );
  NAND4_X1 U3835 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n2985)
         );
  INV_X1 U3836 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3174) );
  INV_X1 U3837 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U3838 ( .A1(n3174), .A2(keyinput84), .B1(keyinput82), .B2(n3194), 
        .ZN(n2981) );
  OAI221_X1 U3839 ( .B1(n3174), .B2(keyinput84), .C1(n3194), .C2(keyinput82), 
        .A(n2981), .ZN(n2984) );
  AOI22_X1 U3840 ( .A1(n2593), .A2(keyinput104), .B1(n3040), .B2(keyinput91), 
        .ZN(n2982) );
  OAI221_X1 U3841 ( .B1(n2593), .B2(keyinput104), .C1(n3040), .C2(keyinput91), 
        .A(n2982), .ZN(n2983) );
  NOR4_X1 U3842 ( .A1(n2986), .A2(n2985), .A3(n2984), .A4(n2983), .ZN(n3024)
         );
  INV_X1 U3843 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n2988) );
  AOI22_X1 U3844 ( .A1(n2988), .A2(keyinput71), .B1(n3998), .B2(keyinput77), 
        .ZN(n2987) );
  OAI221_X1 U3845 ( .B1(n2988), .B2(keyinput71), .C1(n3998), .C2(keyinput77), 
        .A(n2987), .ZN(n2996) );
  INV_X1 U3846 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n3097) );
  INV_X1 U3847 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2990) );
  AOI22_X1 U3848 ( .A1(n3097), .A2(keyinput79), .B1(n2990), .B2(keyinput125), 
        .ZN(n2989) );
  OAI221_X1 U3849 ( .B1(n3097), .B2(keyinput79), .C1(n2990), .C2(keyinput125), 
        .A(n2989), .ZN(n2995) );
  AOI22_X1 U3850 ( .A1(n3493), .A2(keyinput117), .B1(n2679), .B2(keyinput103), 
        .ZN(n2991) );
  OAI221_X1 U3851 ( .B1(n3493), .B2(keyinput117), .C1(n2679), .C2(keyinput103), 
        .A(n2991), .ZN(n2994) );
  INV_X1 U3852 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U3853 ( .A1(n4308), .A2(keyinput83), .B1(n4371), .B2(keyinput95), 
        .ZN(n2992) );
  OAI221_X1 U3854 ( .B1(n4308), .B2(keyinput83), .C1(n4371), .C2(keyinput95), 
        .A(n2992), .ZN(n2993) );
  NOR4_X1 U3855 ( .A1(n2996), .A2(n2995), .A3(n2994), .A4(n2993), .ZN(n3023)
         );
  OAI22_X1 U3856 ( .A1(REG2_REG_9__SCAN_IN), .A2(keyinput80), .B1(
        REG2_REG_0__SCAN_IN), .B2(keyinput67), .ZN(n2997) );
  AOI221_X1 U3857 ( .B1(REG2_REG_9__SCAN_IN), .B2(keyinput80), .C1(keyinput67), 
        .C2(REG2_REG_0__SCAN_IN), .A(n2997), .ZN(n3004) );
  OAI22_X1 U3858 ( .A1(REG1_REG_4__SCAN_IN), .A2(keyinput97), .B1(keyinput101), 
        .B2(ADDR_REG_5__SCAN_IN), .ZN(n2998) );
  AOI221_X1 U3859 ( .B1(REG1_REG_4__SCAN_IN), .B2(keyinput97), .C1(
        ADDR_REG_5__SCAN_IN), .C2(keyinput101), .A(n2998), .ZN(n3003) );
  OAI22_X1 U3860 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput89), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput73), .ZN(n2999) );
  AOI221_X1 U3861 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput89), .C1(keyinput73), .C2(DATAO_REG_16__SCAN_IN), .A(n2999), .ZN(n3002) );
  OAI22_X1 U3862 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput114), .B1(keyinput126), 
        .B2(REG3_REG_11__SCAN_IN), .ZN(n3000) );
  AOI221_X1 U3863 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput114), .C1(
        REG3_REG_11__SCAN_IN), .C2(keyinput126), .A(n3000), .ZN(n3001) );
  NAND4_X1 U3864 ( .A1(n3004), .A2(n3003), .A3(n3002), .A4(n3001), .ZN(n3010)
         );
  INV_X1 U3865 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3975) );
  INV_X1 U3866 ( .A(DATAI_27_), .ZN(n3157) );
  AOI22_X1 U3867 ( .A1(n3975), .A2(keyinput92), .B1(n3157), .B2(keyinput116), 
        .ZN(n3005) );
  OAI221_X1 U3868 ( .B1(n3975), .B2(keyinput92), .C1(n3157), .C2(keyinput116), 
        .A(n3005), .ZN(n3009) );
  INV_X1 U3869 ( .A(D_REG_31__SCAN_IN), .ZN(n4574) );
  INV_X1 U3870 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U3871 ( .A1(n4574), .A2(keyinput124), .B1(keyinput90), .B2(n4411), 
        .ZN(n3006) );
  OAI221_X1 U3872 ( .B1(n4574), .B2(keyinput124), .C1(n4411), .C2(keyinput90), 
        .A(n3006), .ZN(n3008) );
  INV_X1 U3873 ( .A(D_REG_10__SCAN_IN), .ZN(n4595) );
  XNOR2_X1 U3874 ( .A(n4595), .B(keyinput93), .ZN(n3007) );
  NOR4_X1 U3875 ( .A1(n3010), .A2(n3009), .A3(n3008), .A4(n3007), .ZN(n3022)
         );
  OAI22_X1 U3876 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput112), .B1(keyinput111), 
        .B2(D_REG_16__SCAN_IN), .ZN(n3011) );
  AOI221_X1 U3877 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput112), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput111), .A(n3011), .ZN(n3020) );
  OAI22_X1 U3878 ( .A1(IR_REG_21__SCAN_IN), .A2(keyinput121), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput127), .ZN(n3012) );
  AOI221_X1 U3879 ( .B1(IR_REG_21__SCAN_IN), .B2(keyinput121), .C1(keyinput127), .C2(IR_REG_16__SCAN_IN), .A(n3012), .ZN(n3019) );
  INV_X1 U3880 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3035) );
  OAI22_X1 U3881 ( .A1(n3035), .A2(keyinput94), .B1(n4549), .B2(keyinput81), 
        .ZN(n3013) );
  AOI221_X1 U3882 ( .B1(n3035), .B2(keyinput94), .C1(keyinput81), .C2(n4549), 
        .A(n3013), .ZN(n3018) );
  INV_X1 U3883 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3016) );
  OAI22_X1 U3884 ( .A1(n3016), .A2(keyinput76), .B1(n3015), .B2(keyinput120), 
        .ZN(n3014) );
  AOI221_X1 U3885 ( .B1(n3016), .B2(keyinput76), .C1(keyinput120), .C2(n3015), 
        .A(n3014), .ZN(n3017) );
  AND4_X1 U3886 ( .A1(n3020), .A2(n3019), .A3(n3018), .A4(n3017), .ZN(n3021)
         );
  AND4_X1 U3887 ( .A1(n3024), .A2(n3023), .A3(n3022), .A4(n3021), .ZN(n3121)
         );
  INV_X1 U3888 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3176) );
  INV_X1 U3889 ( .A(IR_REG_30__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U3890 ( .A1(n3176), .A2(keyinput98), .B1(n3603), .B2(keyinput72), 
        .ZN(n3025) );
  OAI221_X1 U3891 ( .B1(n3176), .B2(keyinput98), .C1(n3603), .C2(keyinput72), 
        .A(n3025), .ZN(n3033) );
  INV_X1 U3892 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U3893 ( .A1(n3027), .A2(keyinput119), .B1(keyinput99), .B2(n3192), 
        .ZN(n3026) );
  OAI221_X1 U3894 ( .B1(n3027), .B2(keyinput119), .C1(n3192), .C2(keyinput99), 
        .A(n3026), .ZN(n3032) );
  INV_X1 U3895 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3168) );
  INV_X1 U3896 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U3897 ( .A1(n3168), .A2(keyinput86), .B1(keyinput65), .B2(n3178), 
        .ZN(n3028) );
  OAI221_X1 U3898 ( .B1(n3168), .B2(keyinput86), .C1(n3178), .C2(keyinput65), 
        .A(n3028), .ZN(n3031) );
  INV_X1 U3899 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n3082) );
  INV_X1 U3900 ( .A(D_REG_8__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U3901 ( .A1(n3082), .A2(keyinput70), .B1(n4597), .B2(keyinput66), 
        .ZN(n3029) );
  OAI221_X1 U3902 ( .B1(n3082), .B2(keyinput70), .C1(n4597), .C2(keyinput66), 
        .A(n3029), .ZN(n3030) );
  NOR4_X1 U3903 ( .A1(n3033), .A2(n3032), .A3(n3031), .A4(n3030), .ZN(n3120)
         );
  INV_X1 U3904 ( .A(DATAI_16_), .ZN(n4609) );
  AOI22_X1 U3905 ( .A1(n4609), .A2(keyinput38), .B1(n3035), .B2(keyinput30), 
        .ZN(n3034) );
  OAI221_X1 U3906 ( .B1(n4609), .B2(keyinput38), .C1(n3035), .C2(keyinput30), 
        .A(n3034), .ZN(n3044) );
  INV_X1 U3907 ( .A(DATAI_18_), .ZN(n4607) );
  INV_X1 U3908 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U3909 ( .A1(n4607), .A2(keyinput46), .B1(n4661), .B2(keyinput43), 
        .ZN(n3036) );
  OAI221_X1 U3910 ( .B1(n4607), .B2(keyinput46), .C1(n4661), .C2(keyinput43), 
        .A(n3036), .ZN(n3043) );
  AOI22_X1 U3911 ( .A1(n3194), .A2(keyinput18), .B1(n4308), .B2(keyinput19), 
        .ZN(n3037) );
  OAI221_X1 U3912 ( .B1(n3194), .B2(keyinput18), .C1(n4308), .C2(keyinput19), 
        .A(n3037), .ZN(n3042) );
  INV_X1 U3913 ( .A(DATAI_30_), .ZN(n3039) );
  AOI22_X1 U3914 ( .A1(n3040), .A2(keyinput27), .B1(keyinput23), .B2(n3039), 
        .ZN(n3038) );
  OAI221_X1 U3915 ( .B1(n3040), .B2(keyinput27), .C1(n3039), .C2(keyinput23), 
        .A(n3038), .ZN(n3041) );
  NOR4_X1 U3916 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3063)
         );
  AOI22_X1 U3917 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput25), .B1(
        REG2_REG_29__SCAN_IN), .B2(keyinput61), .ZN(n3045) );
  OAI221_X1 U3918 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput25), .C1(
        REG2_REG_29__SCAN_IN), .C2(keyinput61), .A(n3045), .ZN(n3052) );
  AOI22_X1 U3919 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput13), .B1(DATAI_3_), 
        .B2(keyinput21), .ZN(n3046) );
  OAI221_X1 U3920 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput13), .C1(DATAI_3_), 
        .C2(keyinput21), .A(n3046), .ZN(n3051) );
  AOI22_X1 U3921 ( .A1(REG0_REG_24__SCAN_IN), .A2(keyinput49), .B1(
        REG0_REG_17__SCAN_IN), .B2(keyinput45), .ZN(n3047) );
  OAI221_X1 U3922 ( .B1(REG0_REG_24__SCAN_IN), .B2(keyinput49), .C1(
        REG0_REG_17__SCAN_IN), .C2(keyinput45), .A(n3047), .ZN(n3050) );
  AOI22_X1 U3923 ( .A1(DATAO_REG_16__SCAN_IN), .A2(keyinput9), .B1(
        D_REG_10__SCAN_IN), .B2(keyinput29), .ZN(n3048) );
  OAI221_X1 U3924 ( .B1(DATAO_REG_16__SCAN_IN), .B2(keyinput9), .C1(
        D_REG_10__SCAN_IN), .C2(keyinput29), .A(n3048), .ZN(n3049) );
  NOR4_X1 U3925 ( .A1(n3052), .A2(n3051), .A3(n3050), .A4(n3049), .ZN(n3062)
         );
  AOI22_X1 U3926 ( .A1(ADDR_REG_16__SCAN_IN), .A2(keyinput7), .B1(
        REG2_REG_0__SCAN_IN), .B2(keyinput3), .ZN(n3053) );
  OAI221_X1 U3927 ( .B1(ADDR_REG_16__SCAN_IN), .B2(keyinput7), .C1(
        REG2_REG_0__SCAN_IN), .C2(keyinput3), .A(n3053), .ZN(n3060) );
  AOI22_X1 U3928 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput56), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput47), .ZN(n3054) );
  OAI221_X1 U3929 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput56), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput47), .A(n3054), .ZN(n3059) );
  AOI22_X1 U3930 ( .A1(DATAO_REG_30__SCAN_IN), .A2(keyinput35), .B1(
        REG3_REG_18__SCAN_IN), .B2(keyinput55), .ZN(n3055) );
  OAI221_X1 U3931 ( .B1(DATAO_REG_30__SCAN_IN), .B2(keyinput35), .C1(
        REG3_REG_18__SCAN_IN), .C2(keyinput55), .A(n3055), .ZN(n3058) );
  AOI22_X1 U3932 ( .A1(DATAI_27_), .A2(keyinput52), .B1(REG1_REG_29__SCAN_IN), 
        .B2(keyinput39), .ZN(n3056) );
  OAI221_X1 U3933 ( .B1(DATAI_27_), .B2(keyinput52), .C1(REG1_REG_29__SCAN_IN), 
        .C2(keyinput39), .A(n3056), .ZN(n3057) );
  NOR4_X1 U3934 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), .ZN(n3061)
         );
  AND3_X1 U3935 ( .A1(n3063), .A2(n3062), .A3(n3061), .ZN(n3118) );
  AOI22_X1 U3936 ( .A1(DATAO_REG_12__SCAN_IN), .A2(keyinput58), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput54), .ZN(n3064) );
  OAI221_X1 U3937 ( .B1(DATAO_REG_12__SCAN_IN), .B2(keyinput58), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput54), .A(n3064), .ZN(n3071) );
  AOI22_X1 U3938 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput34), .B1(DATAI_25_), 
        .B2(keyinput42), .ZN(n3065) );
  OAI221_X1 U3939 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput34), .C1(DATAI_25_), .C2(keyinput42), .A(n3065), .ZN(n3070) );
  AOI22_X1 U3940 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput22), .B1(
        REG0_REG_13__SCAN_IN), .B2(keyinput26), .ZN(n3066) );
  OAI221_X1 U3941 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput22), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput26), .A(n3066), .ZN(n3069) );
  AOI22_X1 U3942 ( .A1(DATAI_26_), .A2(keyinput10), .B1(REG3_REG_23__SCAN_IN), 
        .B2(keyinput11), .ZN(n3067) );
  OAI221_X1 U3943 ( .B1(DATAI_26_), .B2(keyinput10), .C1(REG3_REG_23__SCAN_IN), 
        .C2(keyinput11), .A(n3067), .ZN(n3068) );
  NOR4_X1 U3944 ( .A1(n3071), .A2(n3070), .A3(n3069), .A4(n3068), .ZN(n3117)
         );
  AOI22_X1 U3945 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput36), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput4), .ZN(n3072) );
  OAI221_X1 U3946 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput36), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput4), .A(n3072), .ZN(n3079) );
  AOI22_X1 U3947 ( .A1(REG0_REG_20__SCAN_IN), .A2(keyinput44), .B1(
        REG2_REG_21__SCAN_IN), .B2(keyinput12), .ZN(n3073) );
  OAI221_X1 U3948 ( .B1(REG0_REG_20__SCAN_IN), .B2(keyinput44), .C1(
        REG2_REG_21__SCAN_IN), .C2(keyinput12), .A(n3073), .ZN(n3078) );
  AOI22_X1 U3949 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput20), .B1(
        REG2_REG_9__SCAN_IN), .B2(keyinput16), .ZN(n3074) );
  OAI221_X1 U3950 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput20), .C1(
        REG2_REG_9__SCAN_IN), .C2(keyinput16), .A(n3074), .ZN(n3077) );
  AOI22_X1 U3951 ( .A1(REG2_REG_16__SCAN_IN), .A2(keyinput17), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput40), .ZN(n3075) );
  OAI221_X1 U3952 ( .B1(REG2_REG_16__SCAN_IN), .B2(keyinput17), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput40), .A(n3075), .ZN(n3076) );
  NOR4_X1 U3953 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3116)
         );
  INV_X1 U3954 ( .A(DATAI_23_), .ZN(n4606) );
  AOI22_X1 U3955 ( .A1(n4574), .A2(keyinput60), .B1(keyinput32), .B2(n4606), 
        .ZN(n3080) );
  OAI221_X1 U3956 ( .B1(n4574), .B2(keyinput60), .C1(n4606), .C2(keyinput32), 
        .A(n3080), .ZN(n3084) );
  AOI22_X1 U3957 ( .A1(n3082), .A2(keyinput6), .B1(n4597), .B2(keyinput2), 
        .ZN(n3081) );
  OAI221_X1 U3958 ( .B1(n3082), .B2(keyinput6), .C1(n4597), .C2(keyinput2), 
        .A(n3081), .ZN(n3083) );
  NOR2_X1 U3959 ( .A1(n3084), .A2(n3083), .ZN(n3091) );
  AOI22_X1 U3960 ( .A1(REG0_REG_26__SCAN_IN), .A2(keyinput31), .B1(n3493), 
        .B2(keyinput53), .ZN(n3085) );
  OAI221_X1 U3961 ( .B1(REG0_REG_26__SCAN_IN), .B2(keyinput31), .C1(n3493), 
        .C2(keyinput53), .A(n3085), .ZN(n3089) );
  INV_X1 U3962 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U3963 ( .A1(n2378), .A2(keyinput33), .B1(keyinput37), .B2(n3087), 
        .ZN(n3086) );
  OAI221_X1 U3964 ( .B1(n2378), .B2(keyinput33), .C1(n3087), .C2(keyinput37), 
        .A(n3086), .ZN(n3088) );
  NOR2_X1 U3965 ( .A1(n3089), .A2(n3088), .ZN(n3090) );
  AND2_X1 U3966 ( .A1(n3091), .A2(n3090), .ZN(n3114) );
  AOI22_X1 U3967 ( .A1(n3603), .A2(keyinput8), .B1(keyinput28), .B2(n3975), 
        .ZN(n3092) );
  OAI221_X1 U3968 ( .B1(n3603), .B2(keyinput8), .C1(n3975), .C2(keyinput28), 
        .A(n3092), .ZN(n3095) );
  INV_X1 U3969 ( .A(DATAI_29_), .ZN(n3155) );
  AOI22_X1 U3970 ( .A1(n2180), .A2(keyinput50), .B1(keyinput51), .B2(n3155), 
        .ZN(n3093) );
  OAI221_X1 U3971 ( .B1(n2180), .B2(keyinput50), .C1(n3155), .C2(keyinput51), 
        .A(n3093), .ZN(n3094) );
  NOR2_X1 U3972 ( .A1(n3095), .A2(n3094), .ZN(n3113) );
  AOI22_X1 U3973 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput63), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput59), .ZN(n3096) );
  OAI221_X1 U3974 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput63), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput59), .A(n3096), .ZN(n3104) );
  XNOR2_X1 U3975 ( .A(n3097), .B(keyinput15), .ZN(n3103) );
  XNOR2_X1 U3976 ( .A(DATAI_24_), .B(keyinput41), .ZN(n3101) );
  XNOR2_X1 U3977 ( .A(IR_REG_21__SCAN_IN), .B(keyinput57), .ZN(n3100) );
  XNOR2_X1 U3978 ( .A(IR_REG_6__SCAN_IN), .B(keyinput24), .ZN(n3099) );
  XNOR2_X1 U3979 ( .A(IR_REG_25__SCAN_IN), .B(keyinput14), .ZN(n3098) );
  NAND4_X1 U3980 ( .A1(n3101), .A2(n3100), .A3(n3099), .A4(n3098), .ZN(n3102)
         );
  NOR3_X1 U3981 ( .A1(n3104), .A2(n3103), .A3(n3102), .ZN(n3112) );
  AOI22_X1 U3982 ( .A1(n4650), .A2(keyinput0), .B1(n3634), .B2(keyinput62), 
        .ZN(n3105) );
  OAI221_X1 U3983 ( .B1(n4650), .B2(keyinput0), .C1(n3634), .C2(keyinput62), 
        .A(n3105), .ZN(n3110) );
  AOI22_X1 U3984 ( .A1(n3178), .A2(keyinput1), .B1(n3107), .B2(keyinput5), 
        .ZN(n3106) );
  OAI221_X1 U3985 ( .B1(n3178), .B2(keyinput1), .C1(n3107), .C2(keyinput5), 
        .A(n3106), .ZN(n3109) );
  INV_X1 U3986 ( .A(D_REG_21__SCAN_IN), .ZN(n4584) );
  XNOR2_X1 U3987 ( .A(n4584), .B(keyinput48), .ZN(n3108) );
  NOR3_X1 U3988 ( .A1(n3110), .A2(n3109), .A3(n3108), .ZN(n3111) );
  AND4_X1 U3989 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3115)
         );
  NAND4_X1 U3990 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3119)
         );
  AOI21_X1 U3991 ( .B1(n3121), .B2(n3120), .A(n3119), .ZN(n3122) );
  XNOR2_X1 U3992 ( .A(n3124), .B(n3123), .ZN(U3217) );
  INV_X1 U3993 ( .A(n4605), .ZN(n3125) );
  XNOR2_X1 U3994 ( .A(n3127), .B(n3134), .ZN(n4333) );
  NAND3_X1 U3995 ( .A1(n3130), .A2(n3129), .A3(n3128), .ZN(n3131) );
  OR2_X1 U3996 ( .A1(n3132), .A2(n4003), .ZN(n3257) );
  NAND2_X1 U3997 ( .A1(n4248), .A2(n3257), .ZN(n3133) );
  NOR2_X1 U3998 ( .A1(n4333), .A2(n4237), .ZN(n3145) );
  INV_X1 U3999 ( .A(n3134), .ZN(n3883) );
  XNOR2_X1 U4000 ( .A(n3135), .B(n3883), .ZN(n3139) );
  NAND2_X1 U4001 ( .A1(n3701), .A2(n4642), .ZN(n3137) );
  NAND2_X1 U4002 ( .A1(n4242), .A2(n4644), .ZN(n3136) );
  OAI211_X1 U4003 ( .C1(n4205), .C2(n4567), .A(n3137), .B(n3136), .ZN(n3138)
         );
  AOI21_X1 U4004 ( .B1(n3139), .B2(n4564), .A(n3138), .ZN(n4331) );
  NOR2_X1 U4005 ( .A1(n4331), .A2(n4259), .ZN(n3144) );
  OR2_X1 U4006 ( .A1(n3593), .A2(n3140), .ZN(n4329) );
  AND2_X1 U4007 ( .A1(n4674), .A2(n4003), .ZN(n3141) );
  AND3_X1 U4008 ( .A1(n4328), .A2(n4329), .A3(n4429), .ZN(n3143) );
  OAI22_X1 U4009 ( .A1(n4227), .A2(n4549), .B1(n3703), .B2(n4225), .ZN(n3142)
         );
  OR4_X1 U4010 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(U3274) );
  INV_X1 U4011 ( .A(DATAI_4_), .ZN(n3146) );
  MUX2_X1 U4012 ( .A(n3146), .B(n3242), .S(STATE_REG_SCAN_IN), .Z(n3147) );
  INV_X1 U4013 ( .A(n3147), .ZN(U3348) );
  INV_X1 U4014 ( .A(n3148), .ZN(n4491) );
  INV_X1 U4015 ( .A(DATAI_9_), .ZN(n3149) );
  MUX2_X1 U4016 ( .A(n4491), .B(n3149), .S(U3149), .Z(n3150) );
  INV_X1 U4017 ( .A(n3150), .ZN(U3343) );
  INV_X1 U4018 ( .A(DATAI_25_), .ZN(n3152) );
  NAND2_X1 U4019 ( .A1(n2652), .A2(STATE_REG_SCAN_IN), .ZN(n3151) );
  OAI21_X1 U4020 ( .B1(STATE_REG_SCAN_IN), .B2(n3152), .A(n3151), .ZN(U3327)
         );
  NAND2_X1 U4021 ( .A1(n3153), .A2(STATE_REG_SCAN_IN), .ZN(n3154) );
  OAI21_X1 U4022 ( .B1(STATE_REG_SCAN_IN), .B2(n3155), .A(n3154), .ZN(U3323)
         );
  NAND2_X1 U4023 ( .A1(n4434), .A2(STATE_REG_SCAN_IN), .ZN(n3156) );
  OAI21_X1 U4024 ( .B1(STATE_REG_SCAN_IN), .B2(n3157), .A(n3156), .ZN(U3325)
         );
  INV_X1 U4025 ( .A(n3158), .ZN(n3224) );
  AND2_X2 U4026 ( .A1(n3224), .A2(n3159), .ZN(n4604) );
  NAND3_X1 U4027 ( .A1(n3164), .A2(n4605), .A3(n3160), .ZN(n3161) );
  OAI21_X1 U4028 ( .B1(n4604), .B2(D_REG_0__SCAN_IN), .A(n3161), .ZN(n3162) );
  INV_X1 U4029 ( .A(n3162), .ZN(U3458) );
  NAND3_X1 U4030 ( .A1(n3164), .A2(n4605), .A3(n3163), .ZN(n3165) );
  OAI21_X1 U4031 ( .B1(n4604), .B2(D_REG_1__SCAN_IN), .A(n3165), .ZN(n3166) );
  INV_X1 U4032 ( .A(n3166), .ZN(U3459) );
  NOR2_X1 U4033 ( .A1(n4554), .A2(U4043), .ZN(U3148) );
  INV_X2 U4034 ( .A(n3967), .ZN(U4043) );
  NAND2_X1 U4035 ( .A1(n3717), .A2(U4043), .ZN(n3167) );
  OAI21_X1 U4036 ( .B1(U4043), .B2(n3168), .A(n3167), .ZN(U3554) );
  INV_X1 U4037 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4038 ( .A1(n3169), .A2(U4043), .ZN(n3170) );
  OAI21_X1 U4039 ( .B1(U4043), .B2(n3171), .A(n3170), .ZN(U3552) );
  NAND2_X1 U4040 ( .A1(n3172), .A2(U4043), .ZN(n3173) );
  OAI21_X1 U4041 ( .B1(U4043), .B2(n3174), .A(n3173), .ZN(U3551) );
  NAND2_X1 U4042 ( .A1(n4156), .A2(U4043), .ZN(n3175) );
  OAI21_X1 U40430 ( .B1(U4043), .B2(n3176), .A(n3175), .ZN(U3571) );
  NAND2_X1 U4044 ( .A1(n3713), .A2(U4043), .ZN(n3177) );
  OAI21_X1 U4045 ( .B1(U4043), .B2(n3178), .A(n3177), .ZN(U3556) );
  NAND2_X1 U4046 ( .A1(n3632), .A2(U4043), .ZN(n3179) );
  OAI21_X1 U4047 ( .B1(U4043), .B2(n3180), .A(n3179), .ZN(U3562) );
  INV_X1 U4048 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4049 ( .A1(n3483), .A2(U4043), .ZN(n3181) );
  OAI21_X1 U4050 ( .B1(U4043), .B2(n3182), .A(n3181), .ZN(U3559) );
  XNOR2_X1 U4051 ( .A(n3183), .B(REG2_REG_3__SCAN_IN), .ZN(n3190) );
  INV_X1 U4052 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3353) );
  NOR2_X1 U4053 ( .A1(STATE_REG_SCAN_IN), .A2(n3353), .ZN(n3230) );
  NOR2_X1 U4054 ( .A1(n4560), .A2(n3184), .ZN(n3185) );
  AOI211_X1 U4055 ( .C1(n4554), .C2(ADDR_REG_3__SCAN_IN), .A(n3230), .B(n3185), 
        .ZN(n3189) );
  OAI211_X1 U4056 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3187), .A(n4555), .B(n3186), 
        .ZN(n3188) );
  OAI211_X1 U4057 ( .C1(n3190), .C2(n4548), .A(n3189), .B(n3188), .ZN(U3243)
         );
  NAND2_X1 U4058 ( .A1(n3858), .A2(U4043), .ZN(n3191) );
  OAI21_X1 U4059 ( .B1(U4043), .B2(n3192), .A(n3191), .ZN(U3580) );
  NAND2_X1 U4060 ( .A1(n3786), .A2(U4043), .ZN(n3193) );
  OAI21_X1 U4061 ( .B1(U4043), .B2(n3194), .A(n3193), .ZN(U3564) );
  INV_X1 U4062 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4063 ( .A1(n3779), .A2(U4043), .ZN(n3195) );
  OAI21_X1 U4064 ( .B1(U4043), .B2(n3196), .A(n3195), .ZN(U3566) );
  INV_X1 U4065 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U4066 ( .A1(n4434), .A2(n4572), .ZN(n3197) );
  NAND2_X1 U4067 ( .A1(n4426), .A2(n3197), .ZN(n4435) );
  NAND2_X1 U4068 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3971) );
  OAI21_X1 U4069 ( .B1(n3200), .B2(n3199), .A(n3198), .ZN(n3236) );
  NOR2_X1 U4070 ( .A1(n3236), .A2(n4434), .ZN(n3201) );
  AOI211_X1 U4071 ( .C1(n4434), .C2(n3971), .A(n3202), .B(n3201), .ZN(n3203)
         );
  AOI211_X1 U4072 ( .C1(n2099), .C2(n4435), .A(n3967), .B(n3203), .ZN(n3243)
         );
  INV_X1 U4073 ( .A(n3243), .ZN(n3219) );
  INV_X1 U4074 ( .A(n4560), .ZN(n3989) );
  NAND2_X1 U4075 ( .A1(n4554), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3204) );
  OAI21_X1 U4076 ( .B1(STATE_REG_SCAN_IN), .B2(n3205), .A(n3204), .ZN(n3217)
         );
  OAI211_X1 U4077 ( .C1(n3208), .C2(n3207), .A(n4555), .B(n3206), .ZN(n3215)
         );
  INV_X1 U4078 ( .A(n3209), .ZN(n3213) );
  NAND3_X1 U4079 ( .A1(n3211), .A2(n3972), .A3(n3210), .ZN(n3212) );
  NAND3_X1 U4080 ( .A1(n4519), .A2(n3213), .A3(n3212), .ZN(n3214) );
  NAND2_X1 U4081 ( .A1(n3215), .A2(n3214), .ZN(n3216) );
  AOI211_X1 U4082 ( .C1(n4424), .C2(n3989), .A(n3217), .B(n3216), .ZN(n3218)
         );
  NAND2_X1 U4083 ( .A1(n3219), .A2(n3218), .ZN(U3242) );
  INV_X1 U4084 ( .A(n3220), .ZN(n3221) );
  AOI21_X1 U4085 ( .B1(n3223), .B2(n3222), .A(n3221), .ZN(n3228) );
  AOI22_X1 U4086 ( .A1(n3787), .A2(n3172), .B1(n3780), .B2(n3966), .ZN(n3227)
         );
  NAND2_X1 U4087 ( .A1(n3225), .A2(n3224), .ZN(n3670) );
  AOI22_X1 U4088 ( .A1(n3332), .A2(n3733), .B1(n3670), .B2(REG3_REG_2__SCAN_IN), .ZN(n3226) );
  OAI211_X1 U4089 ( .C1(n3228), .C2(n3740), .A(n3227), .B(n3226), .ZN(U3234)
         );
  XOR2_X1 U4090 ( .A(n3278), .B(n3279), .Z(n3233) );
  AOI22_X1 U4091 ( .A1(n4643), .A2(n3733), .B1(n3780), .B2(n3717), .ZN(n3232)
         );
  NOR2_X1 U4092 ( .A1(n3784), .A2(REG3_REG_3__SCAN_IN), .ZN(n3229) );
  AOI211_X1 U4093 ( .C1(n3787), .C2(n3169), .A(n3230), .B(n3229), .ZN(n3231)
         );
  OAI211_X1 U4094 ( .C1(n3233), .C2(n3740), .A(n3232), .B(n3231), .ZN(U3215)
         );
  AOI22_X1 U4095 ( .A1(n3780), .A2(n3172), .B1(n3670), .B2(REG3_REG_0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4096 ( .A1(n3781), .A2(n3296), .ZN(n3234) );
  OAI211_X1 U4097 ( .C1(n3236), .C2(n3740), .A(n3235), .B(n3234), .ZN(U3229)
         );
  XOR2_X1 U4098 ( .A(REG2_REG_4__SCAN_IN), .B(n3237), .Z(n3245) );
  OAI211_X1 U4099 ( .C1(n3239), .C2(REG1_REG_4__SCAN_IN), .A(n4555), .B(n3238), 
        .ZN(n3241) );
  AND2_X1 U4100 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3287) );
  AOI21_X1 U4101 ( .B1(n4554), .B2(ADDR_REG_4__SCAN_IN), .A(n3287), .ZN(n3240)
         );
  OAI211_X1 U4102 ( .C1(n4560), .C2(n3242), .A(n3241), .B(n3240), .ZN(n3244)
         );
  AOI211_X1 U4103 ( .C1(n4519), .C2(n3245), .A(n3244), .B(n3243), .ZN(n3246)
         );
  INV_X1 U4104 ( .A(n3246), .ZN(U3244) );
  XNOR2_X1 U4105 ( .A(n3907), .B(n3248), .ZN(n3256) );
  XOR2_X1 U4106 ( .A(n3249), .B(n3907), .Z(n3252) );
  AOI22_X1 U4107 ( .A1(n3965), .A2(n4241), .B1(n4642), .B2(n3286), .ZN(n3250)
         );
  OAI21_X1 U4108 ( .B1(n3800), .B2(n4336), .A(n3250), .ZN(n3251) );
  AOI21_X1 U4109 ( .B1(n3252), .B2(n4564), .A(n3251), .ZN(n3253) );
  OAI21_X1 U4110 ( .B1(n3256), .B2(n4248), .A(n3253), .ZN(n4652) );
  OAI211_X1 U4111 ( .C1(n3351), .C2(n3254), .A(n3366), .B(n4674), .ZN(n4651)
         );
  OAI22_X1 U4112 ( .A1(n4651), .A2(n4420), .B1(n4225), .B2(n3290), .ZN(n3255)
         );
  OAI21_X1 U4113 ( .B1(n4652), .B2(n3255), .A(n4227), .ZN(n3259) );
  INV_X1 U4114 ( .A(n3256), .ZN(n4654) );
  OR2_X1 U4115 ( .A1(n4259), .A2(n3257), .ZN(n4256) );
  INV_X1 U4116 ( .A(n4227), .ZN(n4428) );
  AOI22_X1 U4117 ( .A1(n4654), .A2(n4570), .B1(REG2_REG_4__SCAN_IN), .B2(n4428), .ZN(n3258) );
  NAND2_X1 U4118 ( .A1(n3259), .A2(n3258), .ZN(U3286) );
  INV_X1 U4119 ( .A(n3312), .ZN(n3315) );
  XNOR2_X1 U4120 ( .A(n3311), .B(n3315), .ZN(n3261) );
  XNOR2_X1 U4121 ( .A(n3313), .B(n3261), .ZN(n3266) );
  AOI22_X1 U4122 ( .A1(n3390), .A2(n3733), .B1(n3780), .B2(n3964), .ZN(n3265)
         );
  INV_X1 U4123 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3262) );
  NOR2_X1 U4124 ( .A1(STATE_REG_SCAN_IN), .A2(n3262), .ZN(n4454) );
  NOR2_X1 U4125 ( .A1(n3784), .A2(n3399), .ZN(n3263) );
  AOI211_X1 U4126 ( .C1(n3787), .C2(n3965), .A(n4454), .B(n3263), .ZN(n3264)
         );
  OAI211_X1 U4127 ( .C1(n3266), .C2(n3740), .A(n3265), .B(n3264), .ZN(U3236)
         );
  INV_X1 U4128 ( .A(n3268), .ZN(n3270) );
  NOR2_X1 U4129 ( .A1(n3270), .A2(n3269), .ZN(n3271) );
  XNOR2_X1 U4130 ( .A(n3267), .B(n3271), .ZN(n3276) );
  AOI22_X1 U4131 ( .A1(n3450), .A2(n3733), .B1(n3690), .B2(n3483), .ZN(n3275)
         );
  INV_X1 U4132 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3272) );
  NOR2_X1 U4133 ( .A1(STATE_REG_SCAN_IN), .A2(n3272), .ZN(n4481) );
  NOR2_X1 U4134 ( .A1(n3784), .A2(n3460), .ZN(n3273) );
  AOI211_X1 U4135 ( .C1(n3787), .C2(n3964), .A(n4481), .B(n3273), .ZN(n3274)
         );
  OAI211_X1 U4136 ( .C1(n3276), .C2(n3740), .A(n3275), .B(n3274), .ZN(U3218)
         );
  INV_X1 U4137 ( .A(n3277), .ZN(n3285) );
  NAND2_X1 U4138 ( .A1(n3279), .A2(n3278), .ZN(n3282) );
  NAND2_X1 U4139 ( .A1(n3282), .A2(n3280), .ZN(n3284) );
  NAND2_X1 U4140 ( .A1(n3282), .A2(n3281), .ZN(n3709) );
  INV_X1 U4141 ( .A(n3709), .ZN(n3283) );
  AOI211_X1 U4142 ( .C1(n3285), .C2(n3284), .A(n3740), .B(n3283), .ZN(n3292)
         );
  AOI22_X1 U4143 ( .A1(n3286), .A2(n3733), .B1(n3690), .B2(n3965), .ZN(n3289)
         );
  AOI21_X1 U4144 ( .B1(n3787), .B2(n3966), .A(n3287), .ZN(n3288) );
  OAI211_X1 U4145 ( .C1(n3290), .C2(n3784), .A(n3289), .B(n3288), .ZN(n3291)
         );
  OR2_X1 U4146 ( .A1(n3292), .A2(n3291), .ZN(U3227) );
  OR2_X1 U4147 ( .A1(n3293), .A2(n2599), .ZN(n3294) );
  AND2_X1 U4148 ( .A1(n3295), .A2(n3294), .ZN(n4631) );
  NAND2_X1 U4149 ( .A1(n3671), .A2(n3296), .ZN(n3297) );
  NAND2_X1 U4150 ( .A1(n3298), .A2(n3297), .ZN(n4689) );
  OAI22_X1 U4151 ( .A1(n4234), .A2(n4689), .B1(n3975), .B2(n4225), .ZN(n3309)
         );
  NAND2_X1 U4152 ( .A1(n2599), .A2(n3300), .ZN(n3301) );
  NAND2_X1 U4153 ( .A1(n3299), .A2(n3301), .ZN(n3305) );
  NAND2_X1 U4154 ( .A1(n3671), .A2(n4642), .ZN(n3303) );
  NAND2_X1 U4155 ( .A1(n2697), .A2(n4644), .ZN(n3302) );
  OAI211_X1 U4156 ( .C1(n2372), .C2(n4567), .A(n3303), .B(n3302), .ZN(n3304)
         );
  AOI21_X1 U4157 ( .B1(n3305), .B2(n4564), .A(n3304), .ZN(n3307) );
  INV_X1 U4158 ( .A(n4248), .ZN(n4565) );
  NAND2_X1 U4159 ( .A1(n4631), .A2(n4565), .ZN(n3306) );
  NAND2_X1 U4160 ( .A1(n3307), .A2(n3306), .ZN(n4630) );
  MUX2_X1 U4161 ( .A(n4630), .B(REG2_REG_1__SCAN_IN), .S(n4259), .Z(n3308) );
  AOI211_X1 U4162 ( .C1(n4631), .C2(n4570), .A(n3309), .B(n3308), .ZN(n3310)
         );
  INV_X1 U4163 ( .A(n3310), .ZN(U3289) );
  INV_X1 U4164 ( .A(n3313), .ZN(n3316) );
  OAI21_X1 U4165 ( .B1(n3313), .B2(n3312), .A(n3311), .ZN(n3314) );
  OAI21_X1 U4166 ( .B1(n3316), .B2(n3315), .A(n3314), .ZN(n3320) );
  XNOR2_X1 U4167 ( .A(n3318), .B(n3317), .ZN(n3319) );
  XNOR2_X1 U4168 ( .A(n3320), .B(n3319), .ZN(n3324) );
  AOI22_X1 U4169 ( .A1(n3409), .A2(n3733), .B1(n3780), .B2(n3963), .ZN(n3323)
         );
  AND2_X1 U4170 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4466) );
  NOR2_X1 U4171 ( .A1(n3784), .A2(n3414), .ZN(n3321) );
  AOI211_X1 U4172 ( .C1(n3787), .C2(n3713), .A(n4466), .B(n3321), .ZN(n3322)
         );
  OAI211_X1 U4173 ( .C1(n3324), .C2(n3740), .A(n3323), .B(n3322), .ZN(U3210)
         );
  NAND2_X1 U4174 ( .A1(n3326), .A2(n3874), .ZN(n3327) );
  NAND2_X1 U4175 ( .A1(n3325), .A2(n3327), .ZN(n4640) );
  INV_X1 U4176 ( .A(n4640), .ZN(n3344) );
  NAND3_X1 U4177 ( .A1(n3330), .A2(n3795), .A3(n3299), .ZN(n3331) );
  NAND2_X1 U4178 ( .A1(n3329), .A2(n3331), .ZN(n3335) );
  AOI22_X1 U4179 ( .A1(n3966), .A2(n4241), .B1(n4642), .B2(n3332), .ZN(n3333)
         );
  OAI21_X1 U4180 ( .B1(n2705), .B2(n4336), .A(n3333), .ZN(n3334) );
  AOI21_X1 U4181 ( .B1(n3335), .B2(n4564), .A(n3334), .ZN(n3337) );
  NAND2_X1 U4182 ( .A1(n4640), .A2(n4565), .ZN(n3336) );
  NAND2_X1 U4183 ( .A1(n3337), .A2(n3336), .ZN(n4638) );
  MUX2_X1 U4184 ( .A(n4638), .B(REG2_REG_2__SCAN_IN), .S(n4259), .Z(n3338) );
  INV_X1 U4185 ( .A(n3338), .ZN(n3343) );
  INV_X1 U4186 ( .A(n4225), .ZN(n4569) );
  INV_X1 U4187 ( .A(n3339), .ZN(n4636) );
  NOR3_X1 U4188 ( .A1(n4234), .A2(n4636), .A3(n4637), .ZN(n3341) );
  AOI21_X1 U4189 ( .B1(n4569), .B2(REG3_REG_2__SCAN_IN), .A(n3341), .ZN(n3342)
         );
  OAI211_X1 U4190 ( .C1(n3344), .C2(n4256), .A(n3343), .B(n3342), .ZN(U3288)
         );
  XNOR2_X1 U4191 ( .A(n3912), .B(n3345), .ZN(n3350) );
  INV_X1 U4192 ( .A(n4564), .ZN(n4221) );
  INV_X1 U4193 ( .A(n3912), .ZN(n3346) );
  NAND3_X1 U4194 ( .A1(n3329), .A2(n3796), .A3(n3346), .ZN(n3347) );
  AND2_X1 U4195 ( .A1(n3348), .A2(n3347), .ZN(n3349) );
  OAI222_X1 U4196 ( .A1(n4567), .A2(n3420), .B1(n4248), .B2(n3350), .C1(n4221), 
        .C2(n3349), .ZN(n4647) );
  INV_X1 U4197 ( .A(n4647), .ZN(n3359) );
  INV_X1 U4198 ( .A(n3350), .ZN(n4649) );
  INV_X1 U4199 ( .A(n3351), .ZN(n3352) );
  OAI21_X1 U4200 ( .B1(n4636), .B2(n3355), .A(n3352), .ZN(n4646) );
  AOI22_X1 U4201 ( .A1(n4259), .A2(REG2_REG_3__SCAN_IN), .B1(n4569), .B2(n3353), .ZN(n3354) );
  OAI21_X1 U4202 ( .B1(n4646), .B2(n4234), .A(n3354), .ZN(n3357) );
  AND2_X1 U4203 ( .A1(n4227), .A2(n4642), .ZN(n4232) );
  INV_X1 U4204 ( .A(n4232), .ZN(n3422) );
  NAND2_X1 U4205 ( .A1(n4227), .A2(n4644), .ZN(n4228) );
  OAI22_X1 U4206 ( .A1(n3422), .A2(n3355), .B1(n2372), .B2(n4228), .ZN(n3356)
         );
  AOI211_X1 U4207 ( .C1(n4649), .C2(n4570), .A(n3357), .B(n3356), .ZN(n3358)
         );
  OAI21_X1 U4208 ( .B1(n3359), .B2(n4428), .A(n3358), .ZN(U3287) );
  INV_X1 U4209 ( .A(n3361), .ZN(n3804) );
  NAND2_X1 U4210 ( .A1(n3804), .A2(n3809), .ZN(n3877) );
  XOR2_X1 U4211 ( .A(n3360), .B(n3877), .Z(n3419) );
  OAI22_X1 U4212 ( .A1(n3420), .A2(n4336), .B1(n3421), .B2(n4334), .ZN(n3364)
         );
  XOR2_X1 U4213 ( .A(n3362), .B(n3877), .Z(n3363) );
  OAI22_X1 U4214 ( .A1(n3363), .A2(n4221), .B1(n3412), .B2(n4567), .ZN(n3427)
         );
  AOI211_X1 U4215 ( .C1(n3419), .C2(n4664), .A(n3364), .B(n3427), .ZN(n3371)
         );
  INV_X1 U4216 ( .A(n3365), .ZN(n3398) );
  AOI21_X1 U4217 ( .B1(n3714), .B2(n3366), .A(n3398), .ZN(n3426) );
  INV_X1 U4218 ( .A(n4690), .ZN(n3367) );
  AOI22_X1 U4219 ( .A1(n3426), .A2(n3367), .B1(REG1_REG_5__SCAN_IN), .B2(n4702), .ZN(n3368) );
  OAI21_X1 U4220 ( .B1(n3371), .B2(n4702), .A(n3368), .ZN(U3523) );
  INV_X1 U4221 ( .A(n4633), .ZN(n3369) );
  AOI22_X1 U4222 ( .A1(n3426), .A2(n3369), .B1(REG0_REG_5__SCAN_IN), .B2(n4683), .ZN(n3370) );
  OAI21_X1 U4223 ( .B1(n3371), .B2(n4683), .A(n3370), .ZN(U3477) );
  XNOR2_X1 U4224 ( .A(n3373), .B(n3372), .ZN(n3384) );
  NOR2_X1 U4225 ( .A1(STATE_REG_SCAN_IN), .A2(n3374), .ZN(n3512) );
  AOI21_X1 U4226 ( .B1(n4554), .B2(ADDR_REG_13__SCAN_IN), .A(n3512), .ZN(n3375) );
  OAI21_X1 U4227 ( .B1(n4560), .B2(n3377), .A(n3375), .ZN(n3383) );
  AOI21_X1 U4228 ( .B1(n3378), .B2(n3377), .A(n3376), .ZN(n3381) );
  OAI21_X1 U4229 ( .B1(n3381), .B2(n3380), .A(n4519), .ZN(n3379) );
  AOI21_X1 U4230 ( .B1(n3381), .B2(n3380), .A(n3379), .ZN(n3382) );
  AOI211_X1 U4231 ( .C1(n3384), .C2(n4555), .A(n3383), .B(n3382), .ZN(n3385)
         );
  INV_X1 U4232 ( .A(n3385), .ZN(U3253) );
  NAND2_X1 U4233 ( .A1(n3811), .A2(n3807), .ZN(n3878) );
  NAND2_X1 U4234 ( .A1(n3386), .A2(n3387), .ZN(n3388) );
  XOR2_X1 U4235 ( .A(n3878), .B(n3388), .Z(n3396) );
  XOR2_X1 U4236 ( .A(n3389), .B(n3878), .Z(n3394) );
  AOI22_X1 U4237 ( .A1(n3964), .A2(n4241), .B1(n4642), .B2(n3390), .ZN(n3391)
         );
  OAI21_X1 U4238 ( .B1(n3392), .B2(n4336), .A(n3391), .ZN(n3393) );
  AOI21_X1 U4239 ( .B1(n3394), .B2(n4564), .A(n3393), .ZN(n3395) );
  OAI21_X1 U4240 ( .B1(n3396), .B2(n4248), .A(n3395), .ZN(n4658) );
  INV_X1 U4241 ( .A(n4658), .ZN(n3404) );
  INV_X1 U4242 ( .A(n3396), .ZN(n4660) );
  NOR2_X1 U4243 ( .A1(n3398), .A2(n3397), .ZN(n4657) );
  INV_X1 U4244 ( .A(n3405), .ZN(n4656) );
  NOR3_X1 U4245 ( .A1(n4657), .A2(n4656), .A3(n4234), .ZN(n3402) );
  INV_X1 U4246 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3400) );
  OAI22_X1 U4247 ( .A1(n4227), .A2(n3400), .B1(n3399), .B2(n4225), .ZN(n3401)
         );
  AOI211_X1 U4248 ( .C1(n4660), .C2(n4570), .A(n3402), .B(n3401), .ZN(n3403)
         );
  OAI21_X1 U4249 ( .B1(n3404), .B2(n4428), .A(n3403), .ZN(U3284) );
  AOI211_X1 U4250 ( .C1(n3409), .C2(n3405), .A(n4667), .B(n3458), .ZN(n4663)
         );
  INV_X1 U4251 ( .A(n3908), .ZN(n3406) );
  XNOR2_X1 U4252 ( .A(n3407), .B(n3406), .ZN(n3408) );
  NAND2_X1 U4253 ( .A1(n3408), .A2(n4564), .ZN(n3411) );
  AOI22_X1 U4254 ( .A1(n3963), .A2(n4241), .B1(n4642), .B2(n3409), .ZN(n3410)
         );
  OAI211_X1 U4255 ( .C1(n3412), .C2(n4336), .A(n3411), .B(n3410), .ZN(n4662)
         );
  AOI21_X1 U4256 ( .B1(n4663), .B2(n4003), .A(n4662), .ZN(n3418) );
  XOR2_X1 U4257 ( .A(n3413), .B(n3908), .Z(n4665) );
  INV_X1 U4258 ( .A(n4237), .ZN(n3476) );
  OAI22_X1 U4259 ( .A1(n4227), .A2(n3415), .B1(n3414), .B2(n4225), .ZN(n3416)
         );
  AOI21_X1 U4260 ( .B1(n4665), .B2(n3476), .A(n3416), .ZN(n3417) );
  OAI21_X1 U4261 ( .B1(n3418), .B2(n4428), .A(n3417), .ZN(U3283) );
  INV_X1 U4262 ( .A(n3419), .ZN(n3430) );
  OAI22_X1 U4263 ( .A1(n3422), .A2(n3421), .B1(n3420), .B2(n4228), .ZN(n3425)
         );
  OAI22_X1 U4264 ( .A1(n3715), .A2(n4225), .B1(n3423), .B2(n4227), .ZN(n3424)
         );
  AOI211_X1 U4265 ( .C1(n3426), .C2(n4429), .A(n3425), .B(n3424), .ZN(n3429)
         );
  NAND2_X1 U4266 ( .A1(n3427), .A2(n4227), .ZN(n3428) );
  OAI211_X1 U4267 ( .C1(n3430), .C2(n4237), .A(n3429), .B(n3428), .ZN(U3285)
         );
  OAI21_X1 U4268 ( .B1(n3433), .B2(n3432), .A(n3431), .ZN(n3437) );
  AOI22_X1 U4269 ( .A1(n3473), .A2(n3781), .B1(n3780), .B2(n3962), .ZN(n3435)
         );
  AND2_X1 U4270 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4493) );
  AOI21_X1 U4271 ( .B1(n3787), .B2(n3963), .A(n4493), .ZN(n3434) );
  OAI211_X1 U4272 ( .C1(n3470), .C2(n3784), .A(n3435), .B(n3434), .ZN(n3436)
         );
  AOI21_X1 U4273 ( .B1(n3437), .B2(n3710), .A(n3436), .ZN(n3438) );
  INV_X1 U4274 ( .A(n3438), .ZN(U3228) );
  NAND2_X1 U4275 ( .A1(n3439), .A2(n3710), .ZN(n3447) );
  AOI21_X1 U4276 ( .B1(n3431), .B2(n3441), .A(n3440), .ZN(n3446) );
  AOI22_X1 U4277 ( .A1(n3490), .A2(n3781), .B1(n3690), .B2(n3961), .ZN(n3445)
         );
  NOR2_X1 U4278 ( .A1(STATE_REG_SCAN_IN), .A2(n3442), .ZN(n4503) );
  NOR2_X1 U4279 ( .A1(n3784), .A2(n3492), .ZN(n3443) );
  AOI211_X1 U4280 ( .C1(n3787), .C2(n3483), .A(n4503), .B(n3443), .ZN(n3444)
         );
  OAI211_X1 U4281 ( .C1(n3447), .C2(n3446), .A(n3445), .B(n3444), .ZN(U3214)
         );
  NAND2_X1 U4282 ( .A1(n3817), .A2(n3813), .ZN(n3892) );
  XNOR2_X1 U4283 ( .A(n2054), .B(n3892), .ZN(n3456) );
  XNOR2_X1 U4284 ( .A(n3449), .B(n3892), .ZN(n3454) );
  AOI22_X1 U4285 ( .A1(n3483), .A2(n4241), .B1(n4642), .B2(n3450), .ZN(n3451)
         );
  OAI21_X1 U4286 ( .B1(n3452), .B2(n4336), .A(n3451), .ZN(n3453) );
  AOI21_X1 U4287 ( .B1(n3454), .B2(n4564), .A(n3453), .ZN(n3455) );
  OAI21_X1 U4288 ( .B1(n3456), .B2(n4248), .A(n3455), .ZN(n4670) );
  INV_X1 U4289 ( .A(n4670), .ZN(n3465) );
  INV_X1 U4290 ( .A(n3456), .ZN(n4672) );
  NOR2_X1 U4291 ( .A1(n3458), .A2(n3457), .ZN(n4669) );
  INV_X1 U4292 ( .A(n3459), .ZN(n4668) );
  NOR3_X1 U4293 ( .A1(n4669), .A2(n4668), .A3(n4234), .ZN(n3463) );
  INV_X1 U4294 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3461) );
  OAI22_X1 U4295 ( .A1(n4227), .A2(n3461), .B1(n3460), .B2(n4225), .ZN(n3462)
         );
  AOI211_X1 U4296 ( .C1(n4672), .C2(n4570), .A(n3463), .B(n3462), .ZN(n3464)
         );
  OAI21_X1 U4297 ( .B1(n3465), .B2(n4428), .A(n3464), .ZN(U3282) );
  INV_X1 U4298 ( .A(n3821), .ZN(n3466) );
  NAND2_X1 U4299 ( .A1(n3466), .A2(n3818), .ZN(n3905) );
  XOR2_X1 U4300 ( .A(n3467), .B(n3905), .Z(n3468) );
  OAI22_X1 U4301 ( .A1(n3468), .A2(n4221), .B1(n3533), .B2(n4567), .ZN(n3499)
         );
  INV_X1 U4302 ( .A(n3499), .ZN(n3478) );
  XNOR2_X1 U4303 ( .A(n3469), .B(n3905), .ZN(n3501) );
  OAI21_X1 U4304 ( .B1(n4668), .B2(n3497), .A(n3491), .ZN(n3506) );
  OAI22_X1 U4305 ( .A1(n3470), .A2(n4225), .B1(n2209), .B2(n4227), .ZN(n3472)
         );
  NOR2_X1 U4306 ( .A1(n4228), .A2(n3498), .ZN(n3471) );
  AOI211_X1 U4307 ( .C1(n4232), .C2(n3473), .A(n3472), .B(n3471), .ZN(n3474)
         );
  OAI21_X1 U4308 ( .B1(n3506), .B2(n4234), .A(n3474), .ZN(n3475) );
  AOI21_X1 U4309 ( .B1(n3501), .B2(n3476), .A(n3475), .ZN(n3477) );
  OAI21_X1 U4310 ( .B1(n3478), .B2(n4428), .A(n3477), .ZN(U3281) );
  XNOR2_X1 U4311 ( .A(n3962), .B(n3479), .ZN(n3875) );
  INV_X1 U4312 ( .A(n3875), .ZN(n3481) );
  XNOR2_X1 U4313 ( .A(n3480), .B(n3481), .ZN(n4680) );
  NAND2_X1 U4314 ( .A1(n4680), .A2(n4565), .ZN(n3489) );
  XNOR2_X1 U4315 ( .A(n3482), .B(n3481), .ZN(n3487) );
  NAND2_X1 U4316 ( .A1(n3490), .A2(n4642), .ZN(n3485) );
  NAND2_X1 U4317 ( .A1(n3483), .A2(n4644), .ZN(n3484) );
  OAI211_X1 U4318 ( .C1(n3621), .C2(n4567), .A(n3485), .B(n3484), .ZN(n3486)
         );
  AOI21_X1 U4319 ( .B1(n3487), .B2(n4564), .A(n3486), .ZN(n3488) );
  INV_X1 U4320 ( .A(n4677), .ZN(n3541) );
  NAND2_X1 U4321 ( .A1(n3491), .A2(n3490), .ZN(n4675) );
  AND3_X1 U4322 ( .A1(n3541), .A2(n4429), .A3(n4675), .ZN(n3495) );
  INV_X1 U4323 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3493) );
  OAI22_X1 U4324 ( .A1(n4227), .A2(n3493), .B1(n3492), .B2(n4225), .ZN(n3494)
         );
  AOI211_X1 U4325 ( .C1(n4680), .C2(n4570), .A(n3495), .B(n3494), .ZN(n3496)
         );
  OAI21_X1 U4326 ( .B1(n4682), .B2(n4259), .A(n3496), .ZN(U3280) );
  INV_X1 U4327 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3502) );
  OAI22_X1 U4328 ( .A1(n3498), .A2(n4336), .B1(n3497), .B2(n4334), .ZN(n3500)
         );
  AOI211_X1 U4329 ( .C1(n4664), .C2(n3501), .A(n3500), .B(n3499), .ZN(n3504)
         );
  MUX2_X1 U4330 ( .A(n3502), .B(n3504), .S(n4685), .Z(n3503) );
  OAI21_X1 U4331 ( .B1(n3506), .B2(n4633), .A(n3503), .ZN(U3485) );
  MUX2_X1 U4332 ( .A(n2292), .B(n3504), .S(n4704), .Z(n3505) );
  OAI21_X1 U4333 ( .B1(n4690), .B2(n3506), .A(n3505), .ZN(U3527) );
  NAND2_X1 U4334 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  XNOR2_X1 U4335 ( .A(n3507), .B(n3510), .ZN(n3515) );
  AOI22_X1 U4336 ( .A1(n3566), .A2(n3733), .B1(n3690), .B2(n3786), .ZN(n3514)
         );
  NOR2_X1 U4337 ( .A1(n3784), .A2(n3568), .ZN(n3511) );
  AOI211_X1 U4338 ( .C1(n3787), .C2(n3632), .A(n3512), .B(n3511), .ZN(n3513)
         );
  OAI211_X1 U4339 ( .C1(n3515), .C2(n3740), .A(n3514), .B(n3513), .ZN(U3231)
         );
  INV_X1 U4340 ( .A(n3518), .ZN(n3519) );
  AOI21_X1 U4341 ( .B1(n3517), .B2(n3520), .A(n3519), .ZN(n3560) );
  NAND2_X1 U4342 ( .A1(n3559), .A2(n3557), .ZN(n3904) );
  XNOR2_X1 U4343 ( .A(n3560), .B(n3904), .ZN(n3522) );
  NOR2_X1 U4344 ( .A1(n4244), .A2(n4567), .ZN(n3521) );
  AOI21_X1 U4345 ( .B1(n3522), .B2(n4564), .A(n3521), .ZN(n3576) );
  OAI21_X1 U4346 ( .B1(n3540), .B2(n3573), .A(n2075), .ZN(n3583) );
  INV_X1 U4347 ( .A(n3583), .ZN(n3530) );
  INV_X1 U4348 ( .A(n3523), .ZN(n3623) );
  AOI22_X1 U4349 ( .A1(n4259), .A2(REG2_REG_12__SCAN_IN), .B1(n3623), .B2(
        n4569), .ZN(n3525) );
  NAND2_X1 U4350 ( .A1(n4232), .A2(n3620), .ZN(n3524) );
  OAI211_X1 U4351 ( .C1(n3621), .C2(n4228), .A(n3525), .B(n3524), .ZN(n3529)
         );
  INV_X1 U4352 ( .A(n3904), .ZN(n3527) );
  XNOR2_X1 U4353 ( .A(n3526), .B(n3527), .ZN(n3577) );
  NOR2_X1 U4354 ( .A1(n3577), .A2(n4237), .ZN(n3528) );
  AOI211_X1 U4355 ( .C1(n3530), .C2(n4429), .A(n3529), .B(n3528), .ZN(n3531)
         );
  OAI21_X1 U4356 ( .B1(n4259), .B2(n3576), .A(n3531), .ZN(U3278) );
  XOR2_X1 U4357 ( .A(n3517), .B(n3909), .Z(n3539) );
  AOI22_X1 U4358 ( .A1(n3632), .A2(n4241), .B1(n4642), .B2(n3633), .ZN(n3532)
         );
  OAI21_X1 U4359 ( .B1(n3533), .B2(n4336), .A(n3532), .ZN(n3538) );
  NAND2_X1 U4360 ( .A1(n3534), .A2(n3535), .ZN(n3536) );
  XOR2_X1 U4361 ( .A(n3909), .B(n3536), .Z(n4354) );
  NOR2_X1 U4362 ( .A1(n4354), .A2(n4248), .ZN(n3537) );
  AOI211_X1 U4363 ( .C1(n3539), .C2(n4564), .A(n3538), .B(n3537), .ZN(n4358)
         );
  AOI21_X1 U4364 ( .B1(n3633), .B2(n3541), .A(n3540), .ZN(n4355) );
  OAI22_X1 U4365 ( .A1(n4227), .A2(n3015), .B1(n3635), .B2(n4225), .ZN(n3543)
         );
  NOR2_X1 U4366 ( .A1(n4354), .A2(n4256), .ZN(n3542) );
  AOI211_X1 U4367 ( .C1(n4355), .C2(n4429), .A(n3543), .B(n3542), .ZN(n3544)
         );
  OAI21_X1 U4368 ( .B1(n4358), .B2(n4259), .A(n3544), .ZN(U3279) );
  XNOR2_X1 U4369 ( .A(n3547), .B(n3546), .ZN(n3548) );
  XNOR2_X1 U4370 ( .A(n3545), .B(n3548), .ZN(n3553) );
  AOI22_X1 U4371 ( .A1(n4253), .A2(n3733), .B1(n3690), .B2(n4242), .ZN(n3552)
         );
  INV_X1 U4372 ( .A(n3549), .ZN(n4252) );
  NAND2_X1 U4373 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4531) );
  OAI21_X1 U4374 ( .B1(n3770), .B2(n4244), .A(n4531), .ZN(n3550) );
  AOI21_X1 U4375 ( .B1(n4252), .B2(n3772), .A(n3550), .ZN(n3551) );
  OAI211_X1 U4376 ( .C1(n3553), .C2(n3740), .A(n3552), .B(n3551), .ZN(U3212)
         );
  AND2_X1 U4377 ( .A1(n3555), .A2(n3554), .ZN(n3906) );
  XNOR2_X1 U4378 ( .A(n3556), .B(n3906), .ZN(n4349) );
  INV_X1 U4379 ( .A(n3557), .ZN(n3558) );
  AOI21_X1 U4380 ( .B1(n3560), .B2(n3559), .A(n3558), .ZN(n3561) );
  XOR2_X1 U4381 ( .A(n3906), .B(n3561), .Z(n3564) );
  AOI22_X1 U4382 ( .A1(n3632), .A2(n4644), .B1(n3566), .B2(n4642), .ZN(n3562)
         );
  OAI21_X1 U4383 ( .B1(n4337), .B2(n4567), .A(n3562), .ZN(n3563) );
  AOI21_X1 U4384 ( .B1(n3564), .B2(n4564), .A(n3563), .ZN(n3565) );
  OAI21_X1 U4385 ( .B1(n4349), .B2(n4248), .A(n3565), .ZN(n4350) );
  NAND2_X1 U4386 ( .A1(n4350), .A2(n4227), .ZN(n3572) );
  NAND2_X1 U4387 ( .A1(n2075), .A2(n3566), .ZN(n3567) );
  NAND2_X1 U4388 ( .A1(n2061), .A2(n3567), .ZN(n4413) );
  INV_X1 U4389 ( .A(n4413), .ZN(n3570) );
  OAI22_X1 U4390 ( .A1(n4227), .A2(n3378), .B1(n3568), .B2(n4225), .ZN(n3569)
         );
  AOI21_X1 U4391 ( .B1(n3570), .B2(n4429), .A(n3569), .ZN(n3571) );
  OAI211_X1 U4392 ( .C1(n4349), .C2(n4256), .A(n3572), .B(n3571), .ZN(U3277)
         );
  OAI22_X1 U4393 ( .A1(n3621), .A2(n4336), .B1(n3573), .B2(n4334), .ZN(n3574)
         );
  INV_X1 U4394 ( .A(n3574), .ZN(n3575) );
  OAI211_X1 U4395 ( .C1(n4332), .C2(n3577), .A(n3576), .B(n3575), .ZN(n3580)
         );
  MUX2_X1 U4396 ( .A(REG1_REG_12__SCAN_IN), .B(n3580), .S(n4704), .Z(n3578) );
  INV_X1 U4397 ( .A(n3578), .ZN(n3579) );
  OAI21_X1 U4398 ( .B1(n4690), .B2(n3583), .A(n3579), .ZN(U3530) );
  MUX2_X1 U4399 ( .A(REG0_REG_12__SCAN_IN), .B(n3580), .S(n4685), .Z(n3581) );
  INV_X1 U4400 ( .A(n3581), .ZN(n3582) );
  OAI21_X1 U4401 ( .B1(n3583), .B2(n4633), .A(n3582), .ZN(U3491) );
  INV_X1 U4402 ( .A(n3585), .ZN(n4246) );
  NOR2_X1 U4403 ( .A1(n4246), .A2(n3586), .ZN(n3587) );
  XOR2_X1 U4404 ( .A(n3589), .B(n3587), .Z(n4340) );
  INV_X1 U4405 ( .A(n4340), .ZN(n3602) );
  NAND2_X1 U4406 ( .A1(n3588), .A2(n4564), .ZN(n3592) );
  INV_X1 U4407 ( .A(n3589), .ZN(n3886) );
  AOI21_X1 U4408 ( .B1(n4239), .B2(n3590), .A(n3886), .ZN(n3591) );
  OAI22_X1 U4409 ( .A1(n3592), .A2(n3591), .B1(n4323), .B2(n4567), .ZN(n4339)
         );
  INV_X1 U4410 ( .A(n4344), .ZN(n3595) );
  INV_X1 U4411 ( .A(n3593), .ZN(n3594) );
  OAI21_X1 U4412 ( .B1(n3595), .B2(n4335), .A(n3594), .ZN(n4408) );
  INV_X1 U4413 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3596) );
  OAI22_X1 U4414 ( .A1(n4227), .A2(n3596), .B1(n3783), .B2(n4225), .ZN(n3598)
         );
  NOR2_X1 U4415 ( .A1(n4228), .A2(n4337), .ZN(n3597) );
  AOI211_X1 U4416 ( .C1(n4232), .C2(n3782), .A(n3598), .B(n3597), .ZN(n3599)
         );
  OAI21_X1 U4417 ( .B1(n4408), .B2(n4234), .A(n3599), .ZN(n3600) );
  AOI21_X1 U4418 ( .B1(n4339), .B2(n4227), .A(n3600), .ZN(n3601) );
  OAI21_X1 U4419 ( .B1(n3602), .B2(n4237), .A(n3601), .ZN(U3275) );
  NAND3_X1 U4420 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n3603), 
        .ZN(n3605) );
  INV_X1 U4421 ( .A(DATAI_31_), .ZN(n3604) );
  OAI22_X1 U4422 ( .A1(n2169), .A2(n3605), .B1(STATE_REG_SCAN_IN), .B2(n3604), 
        .ZN(U3321) );
  INV_X1 U4423 ( .A(n3607), .ZN(n3609) );
  NOR2_X1 U4424 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  XNOR2_X1 U4425 ( .A(n3606), .B(n3610), .ZN(n3615) );
  AOI22_X1 U4426 ( .A1(n4202), .A2(n3781), .B1(n3780), .B2(n4203), .ZN(n3614)
         );
  NOR2_X1 U4427 ( .A1(n3784), .A2(n4208), .ZN(n3611) );
  AOI211_X1 U4428 ( .C1(n3787), .C2(n3958), .A(n3612), .B(n3611), .ZN(n3613)
         );
  OAI211_X1 U4429 ( .C1(n3615), .C2(n3740), .A(n3614), .B(n3613), .ZN(U3235)
         );
  XNOR2_X1 U4430 ( .A(n3617), .B(n3616), .ZN(n3618) );
  XNOR2_X1 U4431 ( .A(n3619), .B(n3618), .ZN(n3626) );
  AOI22_X1 U4432 ( .A1(n3620), .A2(n3781), .B1(n3690), .B2(n3959), .ZN(n3625)
         );
  NAND2_X1 U4433 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4521) );
  OAI21_X1 U4434 ( .B1(n3770), .B2(n3621), .A(n4521), .ZN(n3622) );
  AOI21_X1 U4435 ( .B1(n3623), .B2(n3772), .A(n3622), .ZN(n3624) );
  OAI211_X1 U4436 ( .C1(n3626), .C2(n3740), .A(n3625), .B(n3624), .ZN(U3221)
         );
  INV_X1 U4437 ( .A(n3628), .ZN(n3630) );
  NOR2_X1 U4438 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  XNOR2_X1 U4439 ( .A(n3627), .B(n3631), .ZN(n3639) );
  AOI22_X1 U4440 ( .A1(n3633), .A2(n3781), .B1(n3780), .B2(n3632), .ZN(n3638)
         );
  NOR2_X1 U4441 ( .A1(STATE_REG_SCAN_IN), .A2(n3634), .ZN(n4515) );
  NOR2_X1 U4442 ( .A1(n3784), .A2(n3635), .ZN(n3636) );
  AOI211_X1 U4443 ( .C1(n3787), .C2(n3962), .A(n4515), .B(n3636), .ZN(n3637)
         );
  OAI211_X1 U4444 ( .C1(n3639), .C2(n3740), .A(n3638), .B(n3637), .ZN(U3233)
         );
  XNOR2_X1 U4445 ( .A(n3640), .B(n3641), .ZN(n3647) );
  AOI22_X1 U4446 ( .A1(n4041), .A2(n3780), .B1(n4049), .B2(n3733), .ZN(n3646)
         );
  INV_X1 U4447 ( .A(n3642), .ZN(n4046) );
  INV_X1 U4448 ( .A(n3955), .ZN(n4270) );
  INV_X1 U4449 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3643) );
  OAI22_X1 U4450 ( .A1(n3770), .A2(n4270), .B1(STATE_REG_SCAN_IN), .B2(n3643), 
        .ZN(n3644) );
  AOI21_X1 U4451 ( .B1(n4046), .B2(n3772), .A(n3644), .ZN(n3645) );
  OAI211_X1 U4452 ( .C1(n3647), .C2(n3740), .A(n3646), .B(n3645), .ZN(U3211)
         );
  NAND2_X1 U4453 ( .A1(n3648), .A2(n3710), .ZN(n3658) );
  AOI21_X1 U4454 ( .B1(n3649), .B2(n3651), .A(n3650), .ZN(n3657) );
  AOI22_X1 U4455 ( .A1(n4110), .A2(n3781), .B1(n3690), .B2(n3956), .ZN(n3656)
         );
  INV_X1 U4456 ( .A(n4106), .ZN(n3654) );
  OAI22_X1 U4457 ( .A1(n3770), .A2(n4292), .B1(STATE_REG_SCAN_IN), .B2(n3652), 
        .ZN(n3653) );
  AOI21_X1 U4458 ( .B1(n3654), .B2(n3772), .A(n3653), .ZN(n3655) );
  OAI211_X1 U4459 ( .C1(n3658), .C2(n3657), .A(n3656), .B(n3655), .ZN(U3213)
         );
  XOR2_X1 U4460 ( .A(n3661), .B(n3660), .Z(n3666) );
  AOI22_X1 U4461 ( .A1(n4187), .A2(n3781), .B1(n3690), .B2(n4188), .ZN(n3665)
         );
  INV_X1 U4462 ( .A(n4192), .ZN(n3663) );
  NAND2_X1 U4463 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4002) );
  OAI21_X1 U4464 ( .B1(n3770), .B2(n4220), .A(n4002), .ZN(n3662) );
  AOI21_X1 U4465 ( .B1(n3663), .B2(n3772), .A(n3662), .ZN(n3664) );
  OAI211_X1 U4466 ( .C1(n3666), .C2(n3740), .A(n3665), .B(n3664), .ZN(U3216)
         );
  OAI211_X1 U4467 ( .C1(n3667), .C2(n3669), .A(n3668), .B(n3710), .ZN(n3674)
         );
  AOI22_X1 U4468 ( .A1(n3787), .A2(n2697), .B1(n3690), .B2(n3169), .ZN(n3673)
         );
  AOI22_X1 U4469 ( .A1(n3671), .A2(n3781), .B1(n3670), .B2(REG3_REG_1__SCAN_IN), .ZN(n3672) );
  NAND3_X1 U4470 ( .A1(n3674), .A2(n3673), .A3(n3672), .ZN(U3219) );
  INV_X1 U4471 ( .A(n3742), .ZN(n3676) );
  OAI21_X1 U4472 ( .B1(n3675), .B2(n3676), .A(n3743), .ZN(n3680) );
  XNOR2_X1 U4473 ( .A(n3678), .B(n3677), .ZN(n3679) );
  XNOR2_X1 U4474 ( .A(n3680), .B(n3679), .ZN(n3686) );
  AOI22_X1 U4475 ( .A1(n4147), .A2(n3781), .B1(n3690), .B2(n4139), .ZN(n3685)
         );
  INV_X1 U4476 ( .A(n3681), .ZN(n4144) );
  INV_X1 U4477 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3682) );
  OAI22_X1 U4478 ( .A1(n3770), .A2(n4304), .B1(STATE_REG_SCAN_IN), .B2(n3682), 
        .ZN(n3683) );
  AOI21_X1 U4479 ( .B1(n4144), .B2(n3772), .A(n3683), .ZN(n3684) );
  OAI211_X1 U4480 ( .C1(n3686), .C2(n3740), .A(n3685), .B(n3684), .ZN(U3220)
         );
  NAND2_X1 U4481 ( .A1(n3762), .A2(n3687), .ZN(n3689) );
  XOR2_X1 U4482 ( .A(n3689), .B(n3688), .Z(n3696) );
  AOI22_X1 U4483 ( .A1(n4078), .A2(n3781), .B1(n3690), .B2(n3955), .ZN(n3695)
         );
  INV_X1 U4484 ( .A(n4074), .ZN(n3693) );
  OAI22_X1 U4485 ( .A1(n3770), .A2(n4281), .B1(STATE_REG_SCAN_IN), .B2(n3691), 
        .ZN(n3692) );
  AOI21_X1 U4486 ( .B1(n3693), .B2(n3772), .A(n3692), .ZN(n3694) );
  OAI211_X1 U4487 ( .C1(n3696), .C2(n3740), .A(n3695), .B(n3694), .ZN(U3222)
         );
  INV_X1 U4488 ( .A(n3776), .ZN(n3698) );
  OAI21_X1 U4489 ( .B1(n3698), .B2(n3777), .A(n3697), .ZN(n3699) );
  XOR2_X1 U4490 ( .A(n3700), .B(n3699), .Z(n3707) );
  AOI22_X1 U4491 ( .A1(n3701), .A2(n3781), .B1(n3780), .B2(n3958), .ZN(n3706)
         );
  INV_X1 U4492 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3702) );
  NOR2_X1 U4493 ( .A1(STATE_REG_SCAN_IN), .A2(n3702), .ZN(n4553) );
  NOR2_X1 U4494 ( .A1(n3784), .A2(n3703), .ZN(n3704) );
  AOI211_X1 U4495 ( .C1(n3787), .C2(n4242), .A(n4553), .B(n3704), .ZN(n3705)
         );
  OAI211_X1 U4496 ( .C1(n3707), .C2(n3740), .A(n3706), .B(n3705), .ZN(U3223)
         );
  NAND2_X1 U4497 ( .A1(n3709), .A2(n3708), .ZN(n3712) );
  OAI211_X1 U4498 ( .C1(n3712), .C2(n2735), .A(n3711), .B(n3710), .ZN(n3720)
         );
  AOI22_X1 U4499 ( .A1(n3714), .A2(n3781), .B1(n3780), .B2(n3713), .ZN(n3719)
         );
  AND2_X1 U4500 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4444) );
  NOR2_X1 U4501 ( .A1(n3784), .A2(n3715), .ZN(n3716) );
  AOI211_X1 U4502 ( .C1(n3787), .C2(n3717), .A(n4444), .B(n3716), .ZN(n3718)
         );
  NAND3_X1 U4503 ( .A1(n3720), .A2(n3719), .A3(n3718), .ZN(U3224) );
  XNOR2_X1 U4504 ( .A(n3723), .B(n3722), .ZN(n3724) );
  XNOR2_X1 U4505 ( .A(n3721), .B(n3724), .ZN(n3728) );
  AOI22_X1 U4506 ( .A1(n4231), .A2(n3781), .B1(n3780), .B2(n3957), .ZN(n3727)
         );
  AND2_X1 U4507 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3988) );
  NOR2_X1 U4508 ( .A1(n3784), .A2(n4226), .ZN(n3725) );
  AOI211_X1 U4509 ( .C1(n3787), .C2(n3779), .A(n3988), .B(n3725), .ZN(n3726)
         );
  OAI211_X1 U4510 ( .C1(n3728), .C2(n3740), .A(n3727), .B(n3726), .ZN(U3225)
         );
  NAND2_X1 U4511 ( .A1(n3729), .A2(n3730), .ZN(n3731) );
  XOR2_X1 U4512 ( .A(n3732), .B(n3731), .Z(n3741) );
  AOI22_X1 U4513 ( .A1(n3734), .A2(n3733), .B1(n3780), .B2(n4087), .ZN(n3739)
         );
  OAI22_X1 U4514 ( .A1(n3770), .A2(n3736), .B1(STATE_REG_SCAN_IN), .B2(n3735), 
        .ZN(n3737) );
  AOI21_X1 U4515 ( .B1(n4093), .B2(n3772), .A(n3737), .ZN(n3738) );
  OAI211_X1 U4516 ( .C1(n3741), .C2(n3740), .A(n3739), .B(n3738), .ZN(U3226)
         );
  NAND2_X1 U4517 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  XNOR2_X1 U4518 ( .A(n3675), .B(n3744), .ZN(n3750) );
  AOI22_X1 U4519 ( .A1(n4172), .A2(n3781), .B1(n3780), .B2(n4156), .ZN(n3749)
         );
  INV_X1 U4520 ( .A(n3745), .ZN(n4171) );
  INV_X1 U4521 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3746) );
  OAI22_X1 U4522 ( .A1(n3770), .A2(n4158), .B1(STATE_REG_SCAN_IN), .B2(n3746), 
        .ZN(n3747) );
  AOI21_X1 U4523 ( .B1(n4171), .B2(n3772), .A(n3747), .ZN(n3748) );
  OAI211_X1 U4524 ( .C1(n3750), .C2(n3740), .A(n3749), .B(n3748), .ZN(U3230)
         );
  INV_X1 U4525 ( .A(n3649), .ZN(n3751) );
  AOI21_X1 U4526 ( .B1(n3753), .B2(n3752), .A(n3751), .ZN(n3760) );
  AOI22_X1 U4527 ( .A1(n4118), .A2(n3781), .B1(n3780), .B2(n4127), .ZN(n3759)
         );
  INV_X1 U4528 ( .A(n4121), .ZN(n3757) );
  INV_X1 U4529 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3754) );
  OAI22_X1 U4530 ( .A1(n3770), .A2(n3755), .B1(STATE_REG_SCAN_IN), .B2(n3754), 
        .ZN(n3756) );
  AOI21_X1 U4531 ( .B1(n3757), .B2(n3772), .A(n3756), .ZN(n3758) );
  OAI211_X1 U4532 ( .C1(n3760), .C2(n3740), .A(n3759), .B(n3758), .ZN(U3232)
         );
  NAND2_X1 U4533 ( .A1(n3761), .A2(n3762), .ZN(n3766) );
  NOR2_X1 U4534 ( .A1(n2150), .A2(n3764), .ZN(n3765) );
  XNOR2_X1 U4535 ( .A(n3766), .B(n3765), .ZN(n3775) );
  AOI22_X1 U4536 ( .A1(n3954), .A2(n3780), .B1(n3781), .B2(n4061), .ZN(n3774)
         );
  INV_X1 U4537 ( .A(n3767), .ZN(n4064) );
  INV_X1 U4538 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3768) );
  OAI22_X1 U4539 ( .A1(n3770), .A2(n3769), .B1(STATE_REG_SCAN_IN), .B2(n3768), 
        .ZN(n3771) );
  AOI21_X1 U4540 ( .B1(n4064), .B2(n3772), .A(n3771), .ZN(n3773) );
  OAI211_X1 U4541 ( .C1(n3775), .C2(n3740), .A(n3774), .B(n3773), .ZN(U3237)
         );
  NAND2_X1 U4542 ( .A1(n3697), .A2(n3776), .ZN(n3778) );
  XOR2_X1 U4543 ( .A(n3778), .B(n3777), .Z(n3790) );
  AOI22_X1 U4544 ( .A1(n3782), .A2(n3781), .B1(n3780), .B2(n3779), .ZN(n3789)
         );
  AND2_X1 U4545 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U4546 ( .A1(n3784), .A2(n3783), .ZN(n3785) );
  AOI211_X1 U4547 ( .C1(n3787), .C2(n3786), .A(n4541), .B(n3785), .ZN(n3788)
         );
  OAI211_X1 U4548 ( .C1(n3790), .C2(n3740), .A(n3789), .B(n3788), .ZN(U3238)
         );
  INV_X1 U4549 ( .A(n3871), .ZN(n3791) );
  NOR2_X1 U4550 ( .A1(n3792), .A2(n3791), .ZN(n3925) );
  NAND2_X1 U4551 ( .A1(n2697), .A2(n4562), .ZN(n3882) );
  OAI211_X1 U4552 ( .C1(n3794), .C2(n4418), .A(n3882), .B(n3793), .ZN(n3797)
         );
  NAND3_X1 U4553 ( .A1(n3797), .A2(n3796), .A3(n3795), .ZN(n3799) );
  OAI211_X1 U4554 ( .C1(n4643), .C2(n3800), .A(n3799), .B(n3798), .ZN(n3803)
         );
  NAND3_X1 U4555 ( .A1(n3803), .A2(n3802), .A3(n3801), .ZN(n3806) );
  NAND3_X1 U4556 ( .A1(n3806), .A2(n3805), .A3(n3804), .ZN(n3810) );
  INV_X1 U4557 ( .A(n3807), .ZN(n3808) );
  AOI21_X1 U4558 ( .B1(n3810), .B2(n3809), .A(n3808), .ZN(n3816) );
  NAND2_X1 U4559 ( .A1(n3812), .A2(n3811), .ZN(n3815) );
  OAI211_X1 U4560 ( .C1(n3816), .C2(n3815), .A(n3814), .B(n3813), .ZN(n3819)
         );
  AND3_X1 U4561 ( .A1(n3819), .A2(n3818), .A3(n3817), .ZN(n3822) );
  OAI21_X1 U4562 ( .B1(n3822), .B2(n3821), .A(n3820), .ZN(n3825) );
  NAND3_X1 U4563 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(n3831) );
  NAND2_X1 U4564 ( .A1(n3827), .A2(n3826), .ZN(n3832) );
  OR2_X1 U4565 ( .A1(n3832), .A2(n3828), .ZN(n3917) );
  INV_X1 U4566 ( .A(n3917), .ZN(n3830) );
  NAND3_X1 U4567 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(n3840) );
  AOI21_X1 U4568 ( .B1(n3834), .B2(n3833), .A(n3832), .ZN(n3839) );
  INV_X1 U4569 ( .A(n3835), .ZN(n3837) );
  NOR4_X1 U4570 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3916)
         );
  NAND2_X1 U4571 ( .A1(n3840), .A2(n3916), .ZN(n3842) );
  INV_X1 U4572 ( .A(n3924), .ZN(n3841) );
  AOI21_X1 U4573 ( .B1(n3842), .B2(n3918), .A(n3841), .ZN(n3848) );
  INV_X1 U4574 ( .A(n3880), .ZN(n3843) );
  AND2_X1 U4575 ( .A1(n3843), .A2(n3891), .ZN(n3844) );
  NAND3_X1 U4576 ( .A1(n3844), .A2(n4099), .A3(n3919), .ZN(n3847) );
  INV_X1 U4577 ( .A(n3844), .ZN(n3921) );
  OAI211_X1 U4578 ( .C1(n3845), .C2(n3921), .A(n3870), .B(n3879), .ZN(n3926)
         );
  INV_X1 U4579 ( .A(n3926), .ZN(n3846) );
  OAI21_X1 U4580 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3855) );
  INV_X1 U4581 ( .A(n3849), .ZN(n4016) );
  INV_X1 U4582 ( .A(n3953), .ZN(n3859) );
  INV_X1 U4583 ( .A(n3850), .ZN(n3851) );
  OAI21_X1 U4584 ( .B1(n4016), .B2(n3859), .A(n3851), .ZN(n3860) );
  NOR2_X1 U4585 ( .A1(n3852), .A2(n3860), .ZN(n3934) );
  INV_X1 U4586 ( .A(n3934), .ZN(n3853) );
  AOI211_X1 U4587 ( .C1(n3925), .C2(n3855), .A(n3854), .B(n3853), .ZN(n3866)
         );
  NOR2_X1 U4588 ( .A1(n3931), .A2(n3930), .ZN(n3861) );
  NAND2_X1 U4589 ( .A1(n3856), .A2(DATAI_30_), .ZN(n3935) );
  AOI222_X1 U4590 ( .A1(n2525), .A2(REG2_REG_31__SCAN_IN), .B1(n2051), .B2(
        REG1_REG_31__SCAN_IN), .C1(n2432), .C2(REG0_REG_31__SCAN_IN), .ZN(
        n3914) );
  INV_X1 U4591 ( .A(n3914), .ZN(n4009) );
  NAND2_X1 U4592 ( .A1(n3857), .A2(DATAI_31_), .ZN(n4010) );
  NAND2_X1 U4593 ( .A1(n4009), .A2(n4010), .ZN(n3862) );
  OAI21_X1 U4594 ( .B1(n3858), .B2(n3935), .A(n3862), .ZN(n3887) );
  AOI21_X1 U4595 ( .B1(n4016), .B2(n3859), .A(n3887), .ZN(n3928) );
  OAI21_X1 U4596 ( .B1(n3861), .B2(n3860), .A(n3928), .ZN(n3933) );
  INV_X1 U4597 ( .A(n3862), .ZN(n3865) );
  INV_X1 U4598 ( .A(n4010), .ZN(n3864) );
  NOR2_X1 U4599 ( .A1(n3863), .A2(n4266), .ZN(n3915) );
  AOI21_X1 U4600 ( .B1(n3864), .B2(n3914), .A(n3915), .ZN(n3896) );
  OAI22_X1 U4601 ( .A1(n3866), .A2(n3933), .B1(n3865), .B2(n3896), .ZN(n3943)
         );
  INV_X1 U4602 ( .A(n3867), .ZN(n3868) );
  OR2_X1 U4603 ( .A1(n3869), .A2(n3868), .ZN(n4055) );
  NAND2_X1 U4604 ( .A1(n3871), .A2(n3870), .ZN(n4071) );
  INV_X1 U4605 ( .A(n4071), .ZN(n3872) );
  NAND4_X1 U4606 ( .A1(n3874), .A2(n3873), .A3(n4055), .A4(n3872), .ZN(n3876)
         );
  NOR2_X1 U4607 ( .A1(n3876), .A2(n3875), .ZN(n3913) );
  XNOR2_X1 U4608 ( .A(n4203), .B(n4191), .ZN(n4184) );
  NOR2_X1 U4609 ( .A1(n3878), .A2(n3877), .ZN(n3885) );
  INV_X1 U4610 ( .A(n3879), .ZN(n3881) );
  OR2_X1 U4611 ( .A1(n3881), .A2(n3880), .ZN(n4085) );
  NAND2_X1 U4612 ( .A1(n3919), .A2(n3924), .ZN(n4136) );
  NAND2_X1 U4613 ( .A1(n3300), .A2(n3882), .ZN(n4628) );
  NOR4_X1 U4614 ( .A1(n3883), .A2(n4085), .A3(n4136), .A4(n4628), .ZN(n3884)
         );
  NAND4_X1 U4615 ( .A1(n4212), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3899)
         );
  INV_X1 U4616 ( .A(n4125), .ZN(n3897) );
  INV_X1 U4617 ( .A(n3887), .ZN(n3895) );
  NAND2_X1 U4618 ( .A1(n3889), .A2(n3888), .ZN(n4166) );
  INV_X1 U4619 ( .A(n4166), .ZN(n3893) );
  NAND2_X1 U4620 ( .A1(n3891), .A2(n3890), .ZN(n4100) );
  NAND2_X1 U4621 ( .A1(n4179), .A2(n4178), .ZN(n4219) );
  NOR4_X1 U4622 ( .A1(n3893), .A2(n4100), .A3(n4219), .A4(n3892), .ZN(n3894)
         );
  NAND4_X1 U4623 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3898)
         );
  NOR3_X1 U4624 ( .A1(n4184), .A2(n3899), .A3(n3898), .ZN(n3900) );
  NAND4_X1 U4625 ( .A1(n3902), .A2(n3901), .A3(n4038), .A4(n3900), .ZN(n3903)
         );
  NOR4_X1 U4626 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3911)
         );
  NOR4_X1 U4627 ( .A1(n2480), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3910)
         );
  NAND4_X1 U4628 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3941)
         );
  NOR2_X1 U4629 ( .A1(n3915), .A2(n3914), .ZN(n3939) );
  OAI21_X1 U4630 ( .B1(n4240), .B2(n3917), .A(n3916), .ZN(n3920) );
  NAND3_X1 U4631 ( .A1(n3920), .A2(n3919), .A3(n3918), .ZN(n3923) );
  INV_X1 U4632 ( .A(n4099), .ZN(n3922) );
  AOI211_X1 U4633 ( .C1(n3924), .C2(n3923), .A(n3922), .B(n3921), .ZN(n3927)
         );
  OAI21_X1 U4634 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n3932) );
  INV_X1 U4635 ( .A(n3928), .ZN(n3929) );
  NOR4_X1 U4636 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3937)
         );
  AOI21_X1 U4637 ( .B1(n4038), .B2(n3934), .A(n3933), .ZN(n3936) );
  OAI22_X1 U4638 ( .A1(n3937), .A2(n3936), .B1(n4009), .B2(n3935), .ZN(n3938)
         );
  OAI21_X1 U4639 ( .B1(n3939), .B2(n4010), .A(n3938), .ZN(n3940) );
  MUX2_X1 U4640 ( .A(n3941), .B(n3940), .S(n4418), .Z(n3942) );
  MUX2_X1 U4641 ( .A(n3943), .B(n3942), .S(n4419), .Z(n3944) );
  XNOR2_X1 U4642 ( .A(n3944), .B(n4003), .ZN(n3952) );
  NAND2_X1 U4643 ( .A1(n3946), .A2(n3945), .ZN(n3947) );
  OAI211_X1 U4644 ( .C1(n3949), .C2(n3948), .A(B_REG_SCAN_IN), .B(n3947), .ZN(
        n3950) );
  OAI21_X1 U4645 ( .B1(n3952), .B2(n3951), .A(n3950), .ZN(U3239) );
  MUX2_X1 U4646 ( .A(DATAO_REG_31__SCAN_IN), .B(n4009), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4647 ( .A(n3953), .B(DATAO_REG_29__SCAN_IN), .S(n3967), .Z(U3579)
         );
  MUX2_X1 U4648 ( .A(n4041), .B(DATAO_REG_28__SCAN_IN), .S(n3967), .Z(U3578)
         );
  MUX2_X1 U4649 ( .A(DATAO_REG_27__SCAN_IN), .B(n3954), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4650 ( .A(n3955), .B(DATAO_REG_26__SCAN_IN), .S(n3967), .Z(U3576)
         );
  MUX2_X1 U4651 ( .A(n4087), .B(DATAO_REG_25__SCAN_IN), .S(n3967), .Z(U3575)
         );
  MUX2_X1 U4652 ( .A(n3956), .B(DATAO_REG_24__SCAN_IN), .S(n3967), .Z(U3574)
         );
  MUX2_X1 U4653 ( .A(n4127), .B(DATAO_REG_23__SCAN_IN), .S(n3967), .Z(U3573)
         );
  MUX2_X1 U4654 ( .A(DATAO_REG_22__SCAN_IN), .B(n4139), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4655 ( .A(n4188), .B(DATAO_REG_20__SCAN_IN), .S(n3967), .Z(U3570)
         );
  MUX2_X1 U4656 ( .A(n4203), .B(DATAO_REG_19__SCAN_IN), .S(n3967), .Z(U3569)
         );
  MUX2_X1 U4657 ( .A(DATAO_REG_18__SCAN_IN), .B(n3957), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4658 ( .A(DATAO_REG_17__SCAN_IN), .B(n3958), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4659 ( .A(n4242), .B(DATAO_REG_15__SCAN_IN), .S(n3967), .Z(U3565)
         );
  MUX2_X1 U4660 ( .A(DATAO_REG_13__SCAN_IN), .B(n3959), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4661 ( .A(DATAO_REG_11__SCAN_IN), .B(n3961), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4662 ( .A(n3962), .B(DATAO_REG_10__SCAN_IN), .S(n3967), .Z(U3560)
         );
  MUX2_X1 U4663 ( .A(n3963), .B(DATAO_REG_8__SCAN_IN), .S(n3967), .Z(U3558) );
  MUX2_X1 U4664 ( .A(DATAO_REG_7__SCAN_IN), .B(n3964), .S(U4043), .Z(U3557) );
  MUX2_X1 U4665 ( .A(n3965), .B(DATAO_REG_5__SCAN_IN), .S(n3967), .Z(U3555) );
  MUX2_X1 U4666 ( .A(n3966), .B(DATAO_REG_3__SCAN_IN), .S(n3967), .Z(U3553) );
  MUX2_X1 U4667 ( .A(n2697), .B(DATAO_REG_0__SCAN_IN), .S(n3967), .Z(U3550) );
  NAND2_X1 U4668 ( .A1(n3989), .A2(n4425), .ZN(n3980) );
  OAI211_X1 U4669 ( .C1(n3970), .C2(n3969), .A(n4555), .B(n3968), .ZN(n3979)
         );
  INV_X1 U4670 ( .A(n3971), .ZN(n3974) );
  OAI211_X1 U4671 ( .C1(n3974), .C2(n3973), .A(n4519), .B(n3972), .ZN(n3978)
         );
  NOR2_X1 U4672 ( .A1(STATE_REG_SCAN_IN), .A2(n3975), .ZN(n3976) );
  AOI21_X1 U4673 ( .B1(n4554), .B2(ADDR_REG_1__SCAN_IN), .A(n3976), .ZN(n3977)
         );
  NAND4_X1 U4674 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(U3241)
         );
  AOI21_X1 U4675 ( .B1(n3983), .B2(n3982), .A(n3981), .ZN(n3992) );
  INV_X1 U4676 ( .A(n4555), .ZN(n4451) );
  AOI221_X1 U4677 ( .B1(n3986), .B2(n3985), .C1(n3984), .C2(n3985), .A(n4548), 
        .ZN(n3987) );
  AOI211_X1 U4678 ( .C1(n4554), .C2(ADDR_REG_17__SCAN_IN), .A(n3988), .B(n3987), .ZN(n3991) );
  NAND2_X1 U4679 ( .A1(n3989), .A2(n4421), .ZN(n3990) );
  OAI211_X1 U4680 ( .C1(n3992), .C2(n4451), .A(n3991), .B(n3990), .ZN(U3257)
         );
  INV_X1 U4681 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3993) );
  MUX2_X1 U4682 ( .A(REG2_REG_19__SCAN_IN), .B(n3993), .S(n4420), .Z(n3996) );
  MUX2_X1 U4683 ( .A(n4317), .B(REG1_REG_19__SCAN_IN), .S(n4420), .Z(n3999) );
  XNOR2_X1 U4684 ( .A(n4000), .B(n3999), .ZN(n4005) );
  NAND2_X1 U4685 ( .A1(n4554), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4001) );
  OAI211_X1 U4686 ( .C1(n4560), .C2(n4003), .A(n4002), .B(n4001), .ZN(n4004)
         );
  AOI21_X1 U4687 ( .B1(n4005), .B2(n4555), .A(n4004), .ZN(n4006) );
  OAI21_X1 U4688 ( .B1(n4007), .B2(n4548), .A(n4006), .ZN(U3259) );
  XNOR2_X1 U4689 ( .A(n4262), .B(n4010), .ZN(n4362) );
  NAND2_X1 U4690 ( .A1(n4009), .A2(n4008), .ZN(n4264) );
  OAI21_X1 U4691 ( .B1(n4010), .B2(n4334), .A(n4264), .ZN(n4359) );
  NAND2_X1 U4692 ( .A1(n4359), .A2(n4227), .ZN(n4012) );
  NAND2_X1 U4693 ( .A1(n4259), .A2(REG2_REG_31__SCAN_IN), .ZN(n4011) );
  OAI211_X1 U4694 ( .C1(n4362), .C2(n4234), .A(n4012), .B(n4011), .ZN(U3260)
         );
  INV_X1 U4695 ( .A(n4013), .ZN(n4025) );
  OAI22_X1 U4696 ( .A1(n4014), .A2(n4228), .B1(n2990), .B2(n4227), .ZN(n4015)
         );
  AOI21_X1 U4697 ( .B1(n4016), .B2(n4232), .A(n4015), .ZN(n4024) );
  INV_X1 U4698 ( .A(n4018), .ZN(n4022) );
  OAI22_X1 U4699 ( .A1(n4020), .A2(n4234), .B1(n4019), .B2(n4225), .ZN(n4021)
         );
  OAI21_X1 U4700 ( .B1(n4022), .B2(n4021), .A(n4227), .ZN(n4023) );
  OAI211_X1 U4701 ( .C1(n4025), .C2(n4237), .A(n4024), .B(n4023), .ZN(U3354)
         );
  INV_X1 U4702 ( .A(n4027), .ZN(n4035) );
  AOI22_X1 U4703 ( .A1(n4028), .A2(n4569), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4428), .ZN(n4031) );
  NAND2_X1 U4704 ( .A1(n4232), .A2(n4029), .ZN(n4030) );
  OAI211_X1 U4705 ( .C1(n4060), .C2(n4228), .A(n4031), .B(n4030), .ZN(n4034)
         );
  NOR2_X1 U4706 ( .A1(n4032), .A2(n4259), .ZN(n4033) );
  OAI21_X1 U4707 ( .B1(n4026), .B2(n4237), .A(n4036), .ZN(U3262) );
  XNOR2_X1 U4708 ( .A(n4037), .B(n4038), .ZN(n4273) );
  INV_X1 U4709 ( .A(n4273), .ZN(n4053) );
  XNOR2_X1 U4710 ( .A(n4039), .B(n4038), .ZN(n4040) );
  NAND2_X1 U4711 ( .A1(n4040), .A2(n4564), .ZN(n4043) );
  NAND2_X1 U4712 ( .A1(n4041), .A2(n4241), .ZN(n4042) );
  NAND2_X1 U4713 ( .A1(n4043), .A2(n4042), .ZN(n4272) );
  INV_X1 U4714 ( .A(n4044), .ZN(n4045) );
  OAI21_X1 U4715 ( .B1(n4062), .B2(n4269), .A(n4045), .ZN(n4369) );
  AOI22_X1 U4716 ( .A1(n4046), .A2(n4569), .B1(n4259), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4047) );
  OAI21_X1 U4717 ( .B1(n4270), .B2(n4228), .A(n4047), .ZN(n4048) );
  AOI21_X1 U4718 ( .B1(n4049), .B2(n4232), .A(n4048), .ZN(n4050) );
  OAI21_X1 U4719 ( .B1(n4369), .B2(n4234), .A(n4050), .ZN(n4051) );
  AOI21_X1 U4720 ( .B1(n4272), .B2(n4227), .A(n4051), .ZN(n4052) );
  OAI21_X1 U4721 ( .B1(n4053), .B2(n4237), .A(n4052), .ZN(U3263) );
  XOR2_X1 U4722 ( .A(n4055), .B(n4054), .Z(n4277) );
  INV_X1 U4723 ( .A(n4277), .ZN(n4068) );
  XNOR2_X1 U4724 ( .A(n4056), .B(n4055), .ZN(n4057) );
  NAND2_X1 U4725 ( .A1(n4057), .A2(n4564), .ZN(n4059) );
  AOI22_X1 U4726 ( .A1(n4087), .A2(n4644), .B1(n4061), .B2(n4642), .ZN(n4058)
         );
  OAI211_X1 U4727 ( .C1(n4060), .C2(n4567), .A(n4059), .B(n4058), .ZN(n4276)
         );
  AND2_X1 U4728 ( .A1(n2074), .A2(n4061), .ZN(n4063) );
  OR2_X1 U4729 ( .A1(n4063), .A2(n4062), .ZN(n4373) );
  AOI22_X1 U4730 ( .A1(n4259), .A2(REG2_REG_26__SCAN_IN), .B1(n4064), .B2(
        n4569), .ZN(n4065) );
  OAI21_X1 U4731 ( .B1(n4373), .B2(n4234), .A(n4065), .ZN(n4066) );
  AOI21_X1 U4732 ( .B1(n4276), .B2(n4227), .A(n4066), .ZN(n4067) );
  OAI21_X1 U4733 ( .B1(n4068), .B2(n4237), .A(n4067), .ZN(U3264) );
  XOR2_X1 U4734 ( .A(n4071), .B(n4069), .Z(n4284) );
  INV_X1 U4735 ( .A(n4284), .ZN(n4082) );
  XOR2_X1 U4736 ( .A(n4071), .B(n4070), .Z(n4072) );
  OAI22_X1 U4737 ( .A1(n4072), .A2(n4221), .B1(n4270), .B2(n4567), .ZN(n4283)
         );
  NAND2_X1 U4738 ( .A1(n4091), .A2(n4078), .ZN(n4073) );
  NAND2_X1 U4739 ( .A1(n2074), .A2(n4073), .ZN(n4377) );
  INV_X1 U4740 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4075) );
  OAI22_X1 U4741 ( .A1(n4227), .A2(n4075), .B1(n4074), .B2(n4225), .ZN(n4077)
         );
  NOR2_X1 U4742 ( .A1(n4228), .A2(n4281), .ZN(n4076) );
  AOI211_X1 U4743 ( .C1(n4232), .C2(n4078), .A(n4077), .B(n4076), .ZN(n4079)
         );
  OAI21_X1 U4744 ( .B1(n4377), .B2(n4234), .A(n4079), .ZN(n4080) );
  AOI21_X1 U4745 ( .B1(n4283), .B2(n4227), .A(n4080), .ZN(n4081) );
  OAI21_X1 U4746 ( .B1(n4082), .B2(n4237), .A(n4081), .ZN(U3265) );
  XOR2_X1 U4747 ( .A(n4083), .B(n4085), .Z(n4288) );
  INV_X1 U4748 ( .A(n4288), .ZN(n4097) );
  XNOR2_X1 U4749 ( .A(n4084), .B(n4085), .ZN(n4090) );
  NOR2_X1 U4750 ( .A1(n4092), .A2(n4334), .ZN(n4086) );
  AOI21_X1 U4751 ( .B1(n4087), .B2(n4241), .A(n4086), .ZN(n4089) );
  NAND2_X1 U4752 ( .A1(n4127), .A2(n4644), .ZN(n4088) );
  OAI211_X1 U4753 ( .C1(n4090), .C2(n4221), .A(n4089), .B(n4088), .ZN(n4287)
         );
  OAI21_X1 U4754 ( .B1(n4103), .B2(n4092), .A(n4091), .ZN(n4381) );
  AOI22_X1 U4755 ( .A1(n4259), .A2(REG2_REG_24__SCAN_IN), .B1(n4093), .B2(
        n4569), .ZN(n4094) );
  OAI21_X1 U4756 ( .B1(n4381), .B2(n4234), .A(n4094), .ZN(n4095) );
  AOI21_X1 U4757 ( .B1(n4287), .B2(n4227), .A(n4095), .ZN(n4096) );
  OAI21_X1 U4758 ( .B1(n4097), .B2(n4237), .A(n4096), .ZN(U3266) );
  XNOR2_X1 U4759 ( .A(n4098), .B(n4100), .ZN(n4295) );
  INV_X1 U4760 ( .A(n4295), .ZN(n4114) );
  OAI21_X1 U4761 ( .B1(n4126), .B2(n4125), .A(n4099), .ZN(n4101) );
  XNOR2_X1 U4762 ( .A(n4101), .B(n4100), .ZN(n4102) );
  OAI22_X1 U4763 ( .A1(n4102), .A2(n4221), .B1(n4281), .B2(n4567), .ZN(n4294)
         );
  INV_X1 U4764 ( .A(n4103), .ZN(n4105) );
  NAND2_X1 U4765 ( .A1(n4120), .A2(n4110), .ZN(n4104) );
  NAND2_X1 U4766 ( .A1(n4105), .A2(n4104), .ZN(n4385) );
  INV_X1 U4767 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4107) );
  OAI22_X1 U4768 ( .A1(n4227), .A2(n4107), .B1(n4106), .B2(n4225), .ZN(n4109)
         );
  NOR2_X1 U4769 ( .A1(n4228), .A2(n4292), .ZN(n4108) );
  AOI211_X1 U4770 ( .C1(n4232), .C2(n4110), .A(n4109), .B(n4108), .ZN(n4111)
         );
  OAI21_X1 U4771 ( .B1(n4385), .B2(n4234), .A(n4111), .ZN(n4112) );
  AOI21_X1 U4772 ( .B1(n4294), .B2(n4227), .A(n4112), .ZN(n4113) );
  OAI21_X1 U4773 ( .B1(n4114), .B2(n4237), .A(n4113), .ZN(U3267) );
  NOR2_X1 U4774 ( .A1(n4115), .A2(n4125), .ZN(n4116) );
  OR2_X1 U4775 ( .A1(n4117), .A2(n4116), .ZN(n4298) );
  NAND2_X1 U4776 ( .A1(n4142), .A2(n4118), .ZN(n4119) );
  NAND2_X1 U4777 ( .A1(n4120), .A2(n4119), .ZN(n4389) );
  INV_X1 U4778 ( .A(n4389), .ZN(n4124) );
  INV_X1 U4779 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4122) );
  OAI22_X1 U4780 ( .A1(n4227), .A2(n4122), .B1(n4121), .B2(n4225), .ZN(n4123)
         );
  AOI21_X1 U4781 ( .B1(n4124), .B2(n4429), .A(n4123), .ZN(n4134) );
  XNOR2_X1 U4782 ( .A(n4126), .B(n4125), .ZN(n4132) );
  NAND2_X1 U4783 ( .A1(n4156), .A2(n4644), .ZN(n4129) );
  NAND2_X1 U4784 ( .A1(n4127), .A2(n4241), .ZN(n4128) );
  OAI211_X1 U4785 ( .C1(n4334), .C2(n4130), .A(n4129), .B(n4128), .ZN(n4131)
         );
  AOI21_X1 U4786 ( .B1(n4132), .B2(n4564), .A(n4131), .ZN(n4299) );
  OR2_X1 U4787 ( .A1(n4299), .A2(n4259), .ZN(n4133) );
  OAI211_X1 U4788 ( .C1(n4298), .C2(n4237), .A(n4134), .B(n4133), .ZN(U3268)
         );
  XNOR2_X1 U4789 ( .A(n4135), .B(n4136), .ZN(n4307) );
  INV_X1 U4790 ( .A(n4307), .ZN(n4151) );
  XNOR2_X1 U4791 ( .A(n4137), .B(n4136), .ZN(n4138) );
  NAND2_X1 U4792 ( .A1(n4138), .A2(n4564), .ZN(n4141) );
  NAND2_X1 U4793 ( .A1(n4139), .A2(n4241), .ZN(n4140) );
  NAND2_X1 U4794 ( .A1(n4141), .A2(n4140), .ZN(n4306) );
  INV_X1 U4795 ( .A(n4310), .ZN(n4143) );
  OAI21_X1 U4796 ( .B1(n4143), .B2(n4303), .A(n4142), .ZN(n4393) );
  AOI22_X1 U4797 ( .A1(n4259), .A2(REG2_REG_21__SCAN_IN), .B1(n4144), .B2(
        n4569), .ZN(n4145) );
  OAI21_X1 U4798 ( .B1(n4304), .B2(n4228), .A(n4145), .ZN(n4146) );
  AOI21_X1 U4799 ( .B1(n4147), .B2(n4232), .A(n4146), .ZN(n4148) );
  OAI21_X1 U4800 ( .B1(n4393), .B2(n4234), .A(n4148), .ZN(n4149) );
  AOI21_X1 U4801 ( .B1(n4306), .B2(n4227), .A(n4149), .ZN(n4150) );
  OAI21_X1 U4802 ( .B1(n4151), .B2(n4237), .A(n4150), .ZN(U3269) );
  INV_X1 U4803 ( .A(n4152), .ZN(n4153) );
  NAND2_X1 U4804 ( .A1(n4154), .A2(n4153), .ZN(n4155) );
  XNOR2_X1 U4805 ( .A(n4155), .B(n4166), .ZN(n4170) );
  AOI22_X1 U4806 ( .A1(n4156), .A2(n4241), .B1(n4172), .B2(n4642), .ZN(n4157)
         );
  OAI21_X1 U4807 ( .B1(n4158), .B2(n4336), .A(n4157), .ZN(n4169) );
  NAND2_X1 U4808 ( .A1(n4217), .A2(n4159), .ZN(n4161) );
  NAND2_X1 U4809 ( .A1(n4161), .A2(n4160), .ZN(n4211) );
  NAND2_X1 U4810 ( .A1(n4209), .A2(n4162), .ZN(n4177) );
  NAND2_X1 U4811 ( .A1(n4177), .A2(n4163), .ZN(n4165) );
  NAND2_X1 U4812 ( .A1(n4165), .A2(n4164), .ZN(n4167) );
  XNOR2_X1 U4813 ( .A(n4167), .B(n4166), .ZN(n4314) );
  NOR2_X1 U4814 ( .A1(n4314), .A2(n4248), .ZN(n4168) );
  AOI211_X1 U4815 ( .C1(n4564), .C2(n4170), .A(n4169), .B(n4168), .ZN(n4313)
         );
  AOI22_X1 U4816 ( .A1(n4259), .A2(REG2_REG_20__SCAN_IN), .B1(n4171), .B2(
        n4569), .ZN(n4174) );
  NAND2_X1 U4817 ( .A1(n2071), .A2(n4172), .ZN(n4311) );
  NAND3_X1 U4818 ( .A1(n4311), .A2(n4429), .A3(n4310), .ZN(n4173) );
  OAI211_X1 U4819 ( .C1(n4314), .C2(n4256), .A(n4174), .B(n4173), .ZN(n4175)
         );
  INV_X1 U4820 ( .A(n4175), .ZN(n4176) );
  OAI21_X1 U4821 ( .B1(n4313), .B2(n4259), .A(n4176), .ZN(U3270) );
  XNOR2_X1 U4822 ( .A(n4177), .B(n4184), .ZN(n4316) );
  INV_X1 U4823 ( .A(n4316), .ZN(n4196) );
  INV_X1 U4824 ( .A(n4178), .ZN(n4180) );
  OAI21_X1 U4825 ( .B1(n4218), .B2(n4180), .A(n4179), .ZN(n4201) );
  INV_X1 U4826 ( .A(n4181), .ZN(n4183) );
  OAI21_X1 U4827 ( .B1(n4201), .B2(n4183), .A(n4182), .ZN(n4185) );
  XNOR2_X1 U4828 ( .A(n4185), .B(n4184), .ZN(n4186) );
  NAND2_X1 U4829 ( .A1(n4186), .A2(n4564), .ZN(n4190) );
  AOI22_X1 U4830 ( .A1(n4188), .A2(n4241), .B1(n4642), .B2(n4187), .ZN(n4189)
         );
  OAI211_X1 U4831 ( .C1(n4220), .C2(n4336), .A(n4190), .B(n4189), .ZN(n4315)
         );
  OAI21_X1 U4832 ( .B1(n4197), .B2(n4191), .A(n2071), .ZN(n4398) );
  NOR2_X1 U4833 ( .A1(n4398), .A2(n4234), .ZN(n4194) );
  OAI22_X1 U4834 ( .A1(n4227), .A2(n3993), .B1(n4192), .B2(n4225), .ZN(n4193)
         );
  AOI211_X1 U4835 ( .C1(n4315), .C2(n4227), .A(n4194), .B(n4193), .ZN(n4195)
         );
  OAI21_X1 U4836 ( .B1(n4196), .B2(n4237), .A(n4195), .ZN(U3271) );
  INV_X1 U4837 ( .A(n4197), .ZN(n4198) );
  OAI211_X1 U4838 ( .C1(n4200), .C2(n4199), .A(n4198), .B(n4674), .ZN(n4319)
         );
  XNOR2_X1 U4839 ( .A(n4201), .B(n4212), .ZN(n4207) );
  AOI22_X1 U4840 ( .A1(n4203), .A2(n4241), .B1(n4202), .B2(n4642), .ZN(n4204)
         );
  OAI21_X1 U4841 ( .B1(n4205), .B2(n4336), .A(n4204), .ZN(n4206) );
  AOI21_X1 U4842 ( .B1(n4207), .B2(n4564), .A(n4206), .ZN(n4320) );
  OAI21_X1 U4843 ( .B1(n4420), .B2(n4319), .A(n4320), .ZN(n4215) );
  OAI22_X1 U4844 ( .A1(n4227), .A2(n2191), .B1(n4208), .B2(n4225), .ZN(n4214)
         );
  INV_X1 U4845 ( .A(n4209), .ZN(n4210) );
  AOI21_X1 U4846 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4321) );
  NOR2_X1 U4847 ( .A1(n4321), .A2(n4237), .ZN(n4213) );
  AOI211_X1 U4848 ( .C1(n4227), .C2(n4215), .A(n4214), .B(n4213), .ZN(n4216)
         );
  INV_X1 U4849 ( .A(n4216), .ZN(U3272) );
  XOR2_X1 U4850 ( .A(n4217), .B(n4219), .Z(n4326) );
  INV_X1 U4851 ( .A(n4326), .ZN(n4238) );
  XOR2_X1 U4852 ( .A(n4219), .B(n4218), .Z(n4222) );
  OAI22_X1 U4853 ( .A1(n4222), .A2(n4221), .B1(n4220), .B2(n4567), .ZN(n4325)
         );
  INV_X1 U4854 ( .A(n4328), .ZN(n4224) );
  OAI21_X1 U4855 ( .B1(n4224), .B2(n4322), .A(n4223), .ZN(n4403) );
  OAI22_X1 U4856 ( .A1(n4227), .A2(n2109), .B1(n4226), .B2(n4225), .ZN(n4230)
         );
  NOR2_X1 U4857 ( .A1(n4228), .A2(n4323), .ZN(n4229) );
  AOI211_X1 U4858 ( .C1(n4232), .C2(n4231), .A(n4230), .B(n4229), .ZN(n4233)
         );
  OAI21_X1 U4859 ( .B1(n4403), .B2(n4234), .A(n4233), .ZN(n4235) );
  AOI21_X1 U4860 ( .B1(n4325), .B2(n4227), .A(n4235), .ZN(n4236) );
  OAI21_X1 U4861 ( .B1(n4238), .B2(n4237), .A(n4236), .ZN(U3273) );
  OAI21_X1 U4862 ( .B1(n4247), .B2(n4240), .A(n4239), .ZN(n4251) );
  AOI22_X1 U4863 ( .A1(n4242), .A2(n4241), .B1(n4642), .B2(n4253), .ZN(n4243)
         );
  OAI21_X1 U4864 ( .B1(n4244), .B2(n4336), .A(n4243), .ZN(n4250) );
  AOI21_X1 U4865 ( .B1(n4247), .B2(n4245), .A(n4246), .ZN(n4348) );
  NOR2_X1 U4866 ( .A1(n4348), .A2(n4248), .ZN(n4249) );
  AOI211_X1 U4867 ( .C1(n4564), .C2(n4251), .A(n4250), .B(n4249), .ZN(n4346)
         );
  AOI22_X1 U4868 ( .A1(n4259), .A2(REG2_REG_14__SCAN_IN), .B1(n4252), .B2(
        n4569), .ZN(n4255) );
  NAND2_X1 U4869 ( .A1(n2061), .A2(n4253), .ZN(n4343) );
  NAND3_X1 U4870 ( .A1(n4344), .A2(n4429), .A3(n4343), .ZN(n4254) );
  OAI211_X1 U4871 ( .C1(n4348), .C2(n4256), .A(n4255), .B(n4254), .ZN(n4257)
         );
  INV_X1 U4872 ( .A(n4257), .ZN(n4258) );
  OAI21_X1 U4873 ( .B1(n4346), .B2(n4259), .A(n4258), .ZN(U3276) );
  NAND2_X1 U4874 ( .A1(n4359), .A2(n4704), .ZN(n4261) );
  NAND2_X1 U4875 ( .A1(n4702), .A2(REG1_REG_31__SCAN_IN), .ZN(n4260) );
  OAI211_X1 U4876 ( .C1(n4362), .C2(n4690), .A(n4261), .B(n4260), .ZN(U3549)
         );
  AOI21_X1 U4877 ( .B1(n4266), .B2(n4263), .A(n4262), .ZN(n4430) );
  INV_X1 U4878 ( .A(n4430), .ZN(n4365) );
  INV_X1 U4879 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4267) );
  INV_X1 U4880 ( .A(n4264), .ZN(n4265) );
  AOI21_X1 U4881 ( .B1(n4266), .B2(n4642), .A(n4265), .ZN(n4432) );
  MUX2_X1 U4882 ( .A(n4267), .B(n4432), .S(n4704), .Z(n4268) );
  OAI21_X1 U4883 ( .B1(n4365), .B2(n4690), .A(n4268), .ZN(U3548) );
  OAI22_X1 U4884 ( .A1(n4270), .A2(n4336), .B1(n4269), .B2(n4334), .ZN(n4271)
         );
  AOI211_X1 U4885 ( .C1(n4273), .C2(n4664), .A(n4272), .B(n4271), .ZN(n4366)
         );
  MUX2_X1 U4886 ( .A(n4274), .B(n4366), .S(n4704), .Z(n4275) );
  OAI21_X1 U4887 ( .B1(n4690), .B2(n4369), .A(n4275), .ZN(U3545) );
  INV_X1 U4888 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4278) );
  AOI21_X1 U4889 ( .B1(n4277), .B2(n4664), .A(n4276), .ZN(n4370) );
  MUX2_X1 U4890 ( .A(n4278), .B(n4370), .S(n4704), .Z(n4279) );
  OAI21_X1 U4891 ( .B1(n4690), .B2(n4373), .A(n4279), .ZN(U3544) );
  INV_X1 U4892 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4285) );
  OAI22_X1 U4893 ( .A1(n4281), .A2(n4336), .B1(n4280), .B2(n4334), .ZN(n4282)
         );
  AOI211_X1 U4894 ( .C1(n4284), .C2(n4664), .A(n4283), .B(n4282), .ZN(n4374)
         );
  MUX2_X1 U4895 ( .A(n4285), .B(n4374), .S(n4704), .Z(n4286) );
  OAI21_X1 U4896 ( .B1(n4690), .B2(n4377), .A(n4286), .ZN(U3543) );
  AOI21_X1 U4897 ( .B1(n4288), .B2(n4664), .A(n4287), .ZN(n4378) );
  MUX2_X1 U4898 ( .A(n4289), .B(n4378), .S(n4704), .Z(n4290) );
  OAI21_X1 U4899 ( .B1(n4690), .B2(n4381), .A(n4290), .ZN(U3542) );
  OAI22_X1 U4900 ( .A1(n4292), .A2(n4336), .B1(n4334), .B2(n4291), .ZN(n4293)
         );
  AOI211_X1 U4901 ( .C1(n4295), .C2(n4664), .A(n4294), .B(n4293), .ZN(n4382)
         );
  MUX2_X1 U4902 ( .A(n4296), .B(n4382), .S(n4704), .Z(n4297) );
  OAI21_X1 U4903 ( .B1(n4690), .B2(n4385), .A(n4297), .ZN(U3541) );
  OR2_X1 U4904 ( .A1(n4298), .A2(n4332), .ZN(n4300) );
  NAND2_X1 U4905 ( .A1(n4300), .A2(n4299), .ZN(n4386) );
  MUX2_X1 U4906 ( .A(REG1_REG_22__SCAN_IN), .B(n4386), .S(n4704), .Z(n4301) );
  INV_X1 U4907 ( .A(n4301), .ZN(n4302) );
  OAI21_X1 U4908 ( .B1(n4690), .B2(n4389), .A(n4302), .ZN(U3540) );
  OAI22_X1 U4909 ( .A1(n4304), .A2(n4336), .B1(n4334), .B2(n4303), .ZN(n4305)
         );
  AOI211_X1 U4910 ( .C1(n4307), .C2(n4664), .A(n4306), .B(n4305), .ZN(n4390)
         );
  MUX2_X1 U4911 ( .A(n4308), .B(n4390), .S(n4704), .Z(n4309) );
  OAI21_X1 U4912 ( .B1(n4690), .B2(n4393), .A(n4309), .ZN(U3539) );
  NAND3_X1 U4913 ( .A1(n4311), .A2(n4674), .A3(n4310), .ZN(n4312) );
  OAI211_X1 U4914 ( .C1(n4314), .C2(n4347), .A(n4313), .B(n4312), .ZN(n4394)
         );
  MUX2_X1 U4915 ( .A(REG1_REG_20__SCAN_IN), .B(n4394), .S(n4704), .Z(U3538) );
  AOI21_X1 U4916 ( .B1(n4316), .B2(n4664), .A(n4315), .ZN(n4395) );
  MUX2_X1 U4917 ( .A(n4317), .B(n4395), .S(n4704), .Z(n4318) );
  OAI21_X1 U4918 ( .B1(n4690), .B2(n4398), .A(n4318), .ZN(U3537) );
  OAI211_X1 U4919 ( .C1(n4321), .C2(n4332), .A(n4320), .B(n4319), .ZN(n4399)
         );
  MUX2_X1 U4920 ( .A(REG1_REG_18__SCAN_IN), .B(n4399), .S(n4704), .Z(U3536) );
  OAI22_X1 U4921 ( .A1(n4323), .A2(n4336), .B1(n4334), .B2(n4322), .ZN(n4324)
         );
  AOI211_X1 U4922 ( .C1(n4326), .C2(n4664), .A(n4325), .B(n4324), .ZN(n4400)
         );
  MUX2_X1 U4923 ( .A(n2315), .B(n4400), .S(n4704), .Z(n4327) );
  OAI21_X1 U4924 ( .B1(n4690), .B2(n4403), .A(n4327), .ZN(U3535) );
  NAND3_X1 U4925 ( .A1(n4329), .A2(n4674), .A3(n4328), .ZN(n4330) );
  OAI211_X1 U4926 ( .C1(n4333), .C2(n4332), .A(n4331), .B(n4330), .ZN(n4404)
         );
  MUX2_X1 U4927 ( .A(n4404), .B(REG1_REG_16__SCAN_IN), .S(n4702), .Z(U3534) );
  OAI22_X1 U4928 ( .A1(n4337), .A2(n4336), .B1(n4335), .B2(n4334), .ZN(n4338)
         );
  AOI211_X1 U4929 ( .C1(n4340), .C2(n4664), .A(n4339), .B(n4338), .ZN(n4405)
         );
  MUX2_X1 U4930 ( .A(n4341), .B(n4405), .S(n4704), .Z(n4342) );
  OAI21_X1 U4931 ( .B1(n4690), .B2(n4408), .A(n4342), .ZN(U3533) );
  NAND3_X1 U4932 ( .A1(n4344), .A2(n4674), .A3(n4343), .ZN(n4345) );
  OAI211_X1 U4933 ( .C1(n4348), .C2(n4347), .A(n4346), .B(n4345), .ZN(n4409)
         );
  MUX2_X1 U4934 ( .A(REG1_REG_14__SCAN_IN), .B(n4409), .S(n4704), .Z(U3532) );
  INV_X1 U4935 ( .A(n4349), .ZN(n4351) );
  AOI21_X1 U4936 ( .B1(n4679), .B2(n4351), .A(n4350), .ZN(n4410) );
  MUX2_X1 U4937 ( .A(n4352), .B(n4410), .S(n4704), .Z(n4353) );
  OAI21_X1 U4938 ( .B1(n4690), .B2(n4413), .A(n4353), .ZN(U3531) );
  INV_X1 U4939 ( .A(n4354), .ZN(n4356) );
  AOI22_X1 U4940 ( .A1(n4356), .A2(n4679), .B1(n4674), .B2(n4355), .ZN(n4357)
         );
  NAND2_X1 U4941 ( .A1(n4358), .A2(n4357), .ZN(n4414) );
  MUX2_X1 U4942 ( .A(REG1_REG_11__SCAN_IN), .B(n4414), .S(n4704), .Z(U3529) );
  NAND2_X1 U4943 ( .A1(n4359), .A2(n4685), .ZN(n4361) );
  NAND2_X1 U4944 ( .A1(n4683), .A2(REG0_REG_31__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U4945 ( .C1(n4362), .C2(n4633), .A(n4361), .B(n4360), .ZN(U3517)
         );
  INV_X1 U4946 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4947 ( .A(n4363), .B(n4432), .S(n4685), .Z(n4364) );
  OAI21_X1 U4948 ( .B1(n4365), .B2(n4633), .A(n4364), .ZN(U3516) );
  INV_X1 U4949 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4367) );
  MUX2_X1 U4950 ( .A(n4367), .B(n4366), .S(n4685), .Z(n4368) );
  OAI21_X1 U4951 ( .B1(n4369), .B2(n4633), .A(n4368), .ZN(U3513) );
  MUX2_X1 U4952 ( .A(n4371), .B(n4370), .S(n4685), .Z(n4372) );
  OAI21_X1 U4953 ( .B1(n4373), .B2(n4633), .A(n4372), .ZN(U3512) );
  INV_X1 U4954 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U4955 ( .A(n4375), .B(n4374), .S(n4685), .Z(n4376) );
  OAI21_X1 U4956 ( .B1(n4377), .B2(n4633), .A(n4376), .ZN(U3511) );
  INV_X1 U4957 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4379) );
  MUX2_X1 U4958 ( .A(n4379), .B(n4378), .S(n4685), .Z(n4380) );
  OAI21_X1 U4959 ( .B1(n4381), .B2(n4633), .A(n4380), .ZN(U3510) );
  INV_X1 U4960 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4383) );
  MUX2_X1 U4961 ( .A(n4383), .B(n4382), .S(n4685), .Z(n4384) );
  OAI21_X1 U4962 ( .B1(n4385), .B2(n4633), .A(n4384), .ZN(U3509) );
  MUX2_X1 U4963 ( .A(REG0_REG_22__SCAN_IN), .B(n4386), .S(n4685), .Z(n4387) );
  INV_X1 U4964 ( .A(n4387), .ZN(n4388) );
  OAI21_X1 U4965 ( .B1(n4389), .B2(n4633), .A(n4388), .ZN(U3508) );
  INV_X1 U4966 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4391) );
  MUX2_X1 U4967 ( .A(n4391), .B(n4390), .S(n4685), .Z(n4392) );
  OAI21_X1 U4968 ( .B1(n4393), .B2(n4633), .A(n4392), .ZN(U3507) );
  MUX2_X1 U4969 ( .A(REG0_REG_20__SCAN_IN), .B(n4394), .S(n4685), .Z(U3506) );
  INV_X1 U4970 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4396) );
  MUX2_X1 U4971 ( .A(n4396), .B(n4395), .S(n4685), .Z(n4397) );
  OAI21_X1 U4972 ( .B1(n4398), .B2(n4633), .A(n4397), .ZN(U3505) );
  MUX2_X1 U4973 ( .A(REG0_REG_18__SCAN_IN), .B(n4399), .S(n4685), .Z(U3503) );
  INV_X1 U4974 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4401) );
  MUX2_X1 U4975 ( .A(n4401), .B(n4400), .S(n4685), .Z(n4402) );
  OAI21_X1 U4976 ( .B1(n4403), .B2(n4633), .A(n4402), .ZN(U3501) );
  MUX2_X1 U4977 ( .A(n4404), .B(REG0_REG_16__SCAN_IN), .S(n4683), .Z(U3499) );
  INV_X1 U4978 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4406) );
  MUX2_X1 U4979 ( .A(n4406), .B(n4405), .S(n4685), .Z(n4407) );
  OAI21_X1 U4980 ( .B1(n4408), .B2(n4633), .A(n4407), .ZN(U3497) );
  MUX2_X1 U4981 ( .A(REG0_REG_14__SCAN_IN), .B(n4409), .S(n4685), .Z(U3495) );
  MUX2_X1 U4982 ( .A(n4411), .B(n4410), .S(n4685), .Z(n4412) );
  OAI21_X1 U4983 ( .B1(n4413), .B2(n4633), .A(n4412), .ZN(U3493) );
  MUX2_X1 U4984 ( .A(REG0_REG_11__SCAN_IN), .B(n4414), .S(n4685), .Z(U3489) );
  MUX2_X1 U4985 ( .A(n2334), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4986 ( .A(n4415), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4987 ( .A(n4416), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4988 ( .A(DATAI_22_), .B(n4417), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4989 ( .A(DATAI_21_), .B(n4418), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4990 ( .A(DATAI_20_), .B(n4419), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4991 ( .A(n4420), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4992 ( .A(DATAI_17_), .B(n4421), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U4993 ( .A(n4422), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4994 ( .A(DATAI_3_), .B(n4423), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4995 ( .A(n4424), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4996 ( .A(n4425), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U4997 ( .A1(U3149), .A2(n4426), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4427) );
  INV_X1 U4998 ( .A(n4427), .ZN(U3324) );
  AOI22_X1 U4999 ( .A1(n4430), .A2(n4429), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4428), .ZN(n4431) );
  OAI21_X1 U5000 ( .B1(n4259), .B2(n4432), .A(n4431), .ZN(U3261) );
  INV_X1 U5001 ( .A(n4435), .ZN(n4433) );
  OAI211_X1 U5002 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4434), .A(n4436), .B(n4433), 
        .ZN(n4439) );
  AOI22_X1 U5003 ( .A1(n4436), .A2(n4435), .B1(n4555), .B2(n4686), .ZN(n4438)
         );
  AOI22_X1 U5004 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4554), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4437) );
  OAI221_X1 U5005 ( .B1(IR_REG_0__SCAN_IN), .B2(n4439), .C1(n2099), .C2(n4438), 
        .A(n4437), .ZN(U3240) );
  AOI211_X1 U5006 ( .C1(n4442), .C2(n4441), .A(n4440), .B(n4451), .ZN(n4443)
         );
  AOI211_X1 U5007 ( .C1(n4554), .C2(ADDR_REG_5__SCAN_IN), .A(n4444), .B(n4443), 
        .ZN(n4449) );
  OAI211_X1 U5008 ( .C1(n4447), .C2(n4446), .A(n4519), .B(n4445), .ZN(n4448)
         );
  OAI211_X1 U5009 ( .C1(n4560), .C2(n4450), .A(n4449), .B(n4448), .ZN(U3245)
         );
  AOI211_X1 U5010 ( .C1(n4698), .C2(n4453), .A(n4452), .B(n4451), .ZN(n4455)
         );
  AOI211_X1 U5011 ( .C1(n4554), .C2(ADDR_REG_6__SCAN_IN), .A(n4455), .B(n4454), 
        .ZN(n4459) );
  OAI211_X1 U5012 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4457), .A(n4519), .B(n4456), 
        .ZN(n4458) );
  OAI211_X1 U5013 ( .C1(n4560), .C2(n4622), .A(n4459), .B(n4458), .ZN(U3246)
         );
  INV_X1 U5014 ( .A(n4460), .ZN(n4462) );
  NAND2_X1 U5015 ( .A1(n4462), .A2(n4461), .ZN(n4464) );
  OAI21_X1 U5016 ( .B1(n4465), .B2(n4464), .A(n4555), .ZN(n4463) );
  AOI21_X1 U5017 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n4467) );
  AOI211_X1 U5018 ( .C1(n4554), .C2(ADDR_REG_7__SCAN_IN), .A(n4467), .B(n4466), 
        .ZN(n4472) );
  OAI211_X1 U5019 ( .C1(n4470), .C2(n4469), .A(n4519), .B(n4468), .ZN(n4471)
         );
  OAI211_X1 U5020 ( .C1(n4560), .C2(n4620), .A(n4472), .B(n4471), .ZN(U3247)
         );
  OAI211_X1 U5021 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4475), .A(n4555), .B(n4474), 
        .ZN(n4479) );
  OAI211_X1 U5022 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4477), .A(n4519), .B(n4476), 
        .ZN(n4478) );
  OAI211_X1 U5023 ( .C1(n4560), .C2(n2114), .A(n4479), .B(n4478), .ZN(n4480)
         );
  AOI211_X1 U5024 ( .C1(n4554), .C2(ADDR_REG_8__SCAN_IN), .A(n4481), .B(n4480), 
        .ZN(n4482) );
  INV_X1 U5025 ( .A(n4482), .ZN(U3248) );
  OAI211_X1 U5026 ( .C1(n4485), .C2(n4484), .A(n4555), .B(n4483), .ZN(n4490)
         );
  OAI211_X1 U5027 ( .C1(n4488), .C2(n4487), .A(n4519), .B(n4486), .ZN(n4489)
         );
  OAI211_X1 U5028 ( .C1(n4560), .C2(n4491), .A(n4490), .B(n4489), .ZN(n4492)
         );
  AOI211_X1 U5029 ( .C1(n4554), .C2(ADDR_REG_9__SCAN_IN), .A(n4493), .B(n4492), 
        .ZN(n4494) );
  INV_X1 U5030 ( .A(n4494), .ZN(U3249) );
  OAI211_X1 U5031 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4497), .A(n4555), .B(n4496), .ZN(n4501) );
  OAI211_X1 U5032 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4499), .A(n4519), .B(n4498), .ZN(n4500) );
  OAI211_X1 U5033 ( .C1(n4560), .C2(n2115), .A(n4501), .B(n4500), .ZN(n4502)
         );
  AOI211_X1 U5034 ( .C1(n4554), .C2(ADDR_REG_10__SCAN_IN), .A(n4503), .B(n4502), .ZN(n4504) );
  INV_X1 U5035 ( .A(n4504), .ZN(U3250) );
  OAI211_X1 U5036 ( .C1(n4507), .C2(n4506), .A(n4555), .B(n4505), .ZN(n4512)
         );
  OAI211_X1 U5037 ( .C1(n4510), .C2(n4509), .A(n4519), .B(n4508), .ZN(n4511)
         );
  OAI211_X1 U5038 ( .C1(n4560), .C2(n4513), .A(n4512), .B(n4511), .ZN(n4514)
         );
  AOI211_X1 U5039 ( .C1(n4554), .C2(ADDR_REG_11__SCAN_IN), .A(n4515), .B(n4514), .ZN(n4516) );
  INV_X1 U5040 ( .A(n4516), .ZN(U3251) );
  OAI211_X1 U5041 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4520), .A(n4519), .B(n4518), .ZN(n4522) );
  NAND2_X1 U5042 ( .A1(n4522), .A2(n4521), .ZN(n4523) );
  AOI21_X1 U5043 ( .B1(n4554), .B2(ADDR_REG_12__SCAN_IN), .A(n4523), .ZN(n4527) );
  OAI211_X1 U5044 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4525), .A(n4555), .B(n4524), .ZN(n4526) );
  OAI211_X1 U5045 ( .C1(n4560), .C2(n2119), .A(n4527), .B(n4526), .ZN(U3252)
         );
  AOI211_X1 U5046 ( .C1(n4530), .C2(n4529), .A(n4528), .B(n4548), .ZN(n4533)
         );
  INV_X1 U5047 ( .A(n4531), .ZN(n4532) );
  AOI211_X1 U5048 ( .C1(n4554), .C2(ADDR_REG_14__SCAN_IN), .A(n4533), .B(n4532), .ZN(n4537) );
  OAI211_X1 U5049 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4535), .A(n4555), .B(n4534), .ZN(n4536) );
  OAI211_X1 U5050 ( .C1(n4560), .C2(n2125), .A(n4537), .B(n4536), .ZN(U3254)
         );
  AOI211_X1 U5051 ( .C1(n2065), .C2(n4539), .A(n4538), .B(n4548), .ZN(n4540)
         );
  AOI211_X1 U5052 ( .C1(n4554), .C2(ADDR_REG_15__SCAN_IN), .A(n4541), .B(n4540), .ZN(n4546) );
  OAI211_X1 U5053 ( .C1(n4544), .C2(n4543), .A(n4555), .B(n4542), .ZN(n4545)
         );
  OAI211_X1 U5054 ( .C1(n4560), .C2(n4547), .A(n4546), .B(n4545), .ZN(U3255)
         );
  AOI221_X1 U5055 ( .B1(n4551), .B2(n4550), .C1(n4549), .C2(n4550), .A(n4548), 
        .ZN(n4552) );
  AOI211_X1 U5056 ( .C1(ADDR_REG_16__SCAN_IN), .C2(n4554), .A(n4553), .B(n4552), .ZN(n4559) );
  OAI221_X1 U5057 ( .B1(n4557), .B2(REG1_REG_16__SCAN_IN), .C1(n4557), .C2(
        n4556), .A(n4555), .ZN(n4558) );
  OAI211_X1 U5058 ( .C1(n4560), .C2(n4610), .A(n4559), .B(n4558), .ZN(U3256)
         );
  NOR2_X1 U5059 ( .A1(n4562), .A2(n4561), .ZN(n4627) );
  INV_X1 U5060 ( .A(n4563), .ZN(n4568) );
  OAI21_X1 U5061 ( .B1(n4565), .B2(n4564), .A(n4628), .ZN(n4566) );
  OAI21_X1 U5062 ( .B1(n2705), .B2(n4567), .A(n4566), .ZN(n4626) );
  AOI21_X1 U5063 ( .B1(n4627), .B2(n4568), .A(n4626), .ZN(n4573) );
  AOI22_X1 U5064 ( .A1(n4570), .A2(n4628), .B1(REG3_REG_0__SCAN_IN), .B2(n4569), .ZN(n4571) );
  OAI221_X1 U5065 ( .B1(n4259), .B2(n4573), .C1(n4227), .C2(n4572), .A(n4571), 
        .ZN(U3290) );
  NOR2_X1 U5066 ( .A1(n4604), .A2(n4574), .ZN(U3291) );
  INV_X1 U5067 ( .A(D_REG_30__SCAN_IN), .ZN(n4575) );
  NOR2_X1 U5068 ( .A1(n4604), .A2(n4575), .ZN(U3292) );
  INV_X1 U5069 ( .A(D_REG_29__SCAN_IN), .ZN(n4576) );
  NOR2_X1 U5070 ( .A1(n4604), .A2(n4576), .ZN(U3293) );
  INV_X1 U5071 ( .A(D_REG_28__SCAN_IN), .ZN(n4577) );
  NOR2_X1 U5072 ( .A1(n4604), .A2(n4577), .ZN(U3294) );
  INV_X1 U5073 ( .A(D_REG_27__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U5074 ( .A1(n4604), .A2(n4578), .ZN(U3295) );
  INV_X1 U5075 ( .A(D_REG_26__SCAN_IN), .ZN(n4579) );
  NOR2_X1 U5076 ( .A1(n4604), .A2(n4579), .ZN(U3296) );
  INV_X1 U5077 ( .A(D_REG_25__SCAN_IN), .ZN(n4580) );
  NOR2_X1 U5078 ( .A1(n4604), .A2(n4580), .ZN(U3297) );
  INV_X1 U5079 ( .A(D_REG_24__SCAN_IN), .ZN(n4581) );
  NOR2_X1 U5080 ( .A1(n4604), .A2(n4581), .ZN(U3298) );
  INV_X1 U5081 ( .A(D_REG_23__SCAN_IN), .ZN(n4582) );
  NOR2_X1 U5082 ( .A1(n4604), .A2(n4582), .ZN(U3299) );
  INV_X1 U5083 ( .A(D_REG_22__SCAN_IN), .ZN(n4583) );
  NOR2_X1 U5084 ( .A1(n4604), .A2(n4583), .ZN(U3300) );
  NOR2_X1 U5085 ( .A1(n4604), .A2(n4584), .ZN(U3301) );
  INV_X1 U5086 ( .A(D_REG_20__SCAN_IN), .ZN(n4585) );
  NOR2_X1 U5087 ( .A1(n4604), .A2(n4585), .ZN(U3302) );
  INV_X1 U5088 ( .A(D_REG_19__SCAN_IN), .ZN(n4586) );
  NOR2_X1 U5089 ( .A1(n4604), .A2(n4586), .ZN(U3303) );
  INV_X1 U5090 ( .A(D_REG_18__SCAN_IN), .ZN(n4587) );
  NOR2_X1 U5091 ( .A1(n4604), .A2(n4587), .ZN(U3304) );
  INV_X1 U5092 ( .A(D_REG_17__SCAN_IN), .ZN(n4588) );
  NOR2_X1 U5093 ( .A1(n4604), .A2(n4588), .ZN(U3305) );
  INV_X1 U5094 ( .A(D_REG_16__SCAN_IN), .ZN(n4589) );
  NOR2_X1 U5095 ( .A1(n4604), .A2(n4589), .ZN(U3306) );
  INV_X1 U5096 ( .A(D_REG_15__SCAN_IN), .ZN(n4590) );
  NOR2_X1 U5097 ( .A1(n4604), .A2(n4590), .ZN(U3307) );
  INV_X1 U5098 ( .A(D_REG_14__SCAN_IN), .ZN(n4591) );
  NOR2_X1 U5099 ( .A1(n4604), .A2(n4591), .ZN(U3308) );
  INV_X1 U5100 ( .A(D_REG_13__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U5101 ( .A1(n4604), .A2(n4592), .ZN(U3309) );
  INV_X1 U5102 ( .A(D_REG_12__SCAN_IN), .ZN(n4593) );
  NOR2_X1 U5103 ( .A1(n4604), .A2(n4593), .ZN(U3310) );
  INV_X1 U5104 ( .A(D_REG_11__SCAN_IN), .ZN(n4594) );
  NOR2_X1 U5105 ( .A1(n4604), .A2(n4594), .ZN(U3311) );
  NOR2_X1 U5106 ( .A1(n4604), .A2(n4595), .ZN(U3312) );
  INV_X1 U5107 ( .A(D_REG_9__SCAN_IN), .ZN(n4596) );
  NOR2_X1 U5108 ( .A1(n4604), .A2(n4596), .ZN(U3313) );
  NOR2_X1 U5109 ( .A1(n4604), .A2(n4597), .ZN(U3314) );
  INV_X1 U5110 ( .A(D_REG_7__SCAN_IN), .ZN(n4598) );
  NOR2_X1 U5111 ( .A1(n4604), .A2(n4598), .ZN(U3315) );
  INV_X1 U5112 ( .A(D_REG_6__SCAN_IN), .ZN(n4599) );
  NOR2_X1 U5113 ( .A1(n4604), .A2(n4599), .ZN(U3316) );
  INV_X1 U5114 ( .A(D_REG_5__SCAN_IN), .ZN(n4600) );
  NOR2_X1 U5115 ( .A1(n4604), .A2(n4600), .ZN(U3317) );
  INV_X1 U5116 ( .A(D_REG_4__SCAN_IN), .ZN(n4601) );
  NOR2_X1 U5117 ( .A1(n4604), .A2(n4601), .ZN(U3318) );
  INV_X1 U5118 ( .A(D_REG_3__SCAN_IN), .ZN(n4602) );
  NOR2_X1 U5119 ( .A1(n4604), .A2(n4602), .ZN(U3319) );
  INV_X1 U5120 ( .A(D_REG_2__SCAN_IN), .ZN(n4603) );
  NOR2_X1 U5121 ( .A1(n4604), .A2(n4603), .ZN(U3320) );
  AOI21_X1 U5122 ( .B1(U3149), .B2(n4606), .A(n4605), .ZN(U3329) );
  AOI22_X1 U5123 ( .A1(STATE_REG_SCAN_IN), .A2(n4608), .B1(n4607), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5124 ( .A1(STATE_REG_SCAN_IN), .A2(n4610), .B1(n4609), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5125 ( .A1(U3149), .A2(n4611), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4612) );
  INV_X1 U5126 ( .A(n4612), .ZN(U3337) );
  INV_X1 U5127 ( .A(DATAI_14_), .ZN(n4613) );
  AOI22_X1 U5128 ( .A1(STATE_REG_SCAN_IN), .A2(n2125), .B1(n4613), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5129 ( .A(DATAI_12_), .ZN(n4614) );
  AOI22_X1 U5130 ( .A1(STATE_REG_SCAN_IN), .A2(n2119), .B1(n4614), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5131 ( .A1(U3149), .A2(n4615), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4616) );
  INV_X1 U5132 ( .A(n4616), .ZN(U3341) );
  INV_X1 U5133 ( .A(DATAI_10_), .ZN(n4617) );
  AOI22_X1 U5134 ( .A1(STATE_REG_SCAN_IN), .A2(n2115), .B1(n4617), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5135 ( .A(DATAI_8_), .ZN(n4618) );
  AOI22_X1 U5136 ( .A1(STATE_REG_SCAN_IN), .A2(n2114), .B1(n4618), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5137 ( .A(DATAI_7_), .ZN(n4619) );
  AOI22_X1 U5138 ( .A1(STATE_REG_SCAN_IN), .A2(n4620), .B1(n4619), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5139 ( .A(DATAI_6_), .ZN(n4621) );
  AOI22_X1 U5140 ( .A1(STATE_REG_SCAN_IN), .A2(n4622), .B1(n4621), .B2(U3149), 
        .ZN(U3346) );
  OAI22_X1 U5141 ( .A1(U3149), .A2(n4623), .B1(DATAI_5_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4624) );
  INV_X1 U5142 ( .A(n4624), .ZN(U3347) );
  OAI22_X1 U5143 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4625) );
  INV_X1 U5144 ( .A(n4625), .ZN(U3352) );
  AOI211_X1 U5145 ( .C1(n4679), .C2(n4628), .A(n4627), .B(n4626), .ZN(n4687)
         );
  INV_X1 U5146 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5147 ( .A1(n4685), .A2(n4687), .B1(n4629), .B2(n4683), .ZN(U3467)
         );
  AOI21_X1 U5148 ( .B1(n4679), .B2(n4631), .A(n4630), .ZN(n4693) );
  INV_X1 U5149 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5150 ( .A1(n4633), .A2(n4689), .B1(n4685), .B2(n4632), .ZN(n4634)
         );
  INV_X1 U5151 ( .A(n4634), .ZN(n4635) );
  OAI21_X1 U5152 ( .B1(n4693), .B2(n4683), .A(n4635), .ZN(U3469) );
  NOR3_X1 U5153 ( .A1(n4637), .A2(n4636), .A3(n4667), .ZN(n4639) );
  AOI211_X1 U5154 ( .C1(n4679), .C2(n4640), .A(n4639), .B(n4638), .ZN(n4695)
         );
  INV_X1 U5155 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5156 ( .A1(n4685), .A2(n4695), .B1(n4641), .B2(n4683), .ZN(U3471)
         );
  AOI22_X1 U5157 ( .A1(n3169), .A2(n4644), .B1(n4643), .B2(n4642), .ZN(n4645)
         );
  OAI21_X1 U5158 ( .B1(n4646), .B2(n4667), .A(n4645), .ZN(n4648) );
  AOI211_X1 U5159 ( .C1(n4679), .C2(n4649), .A(n4648), .B(n4647), .ZN(n4696)
         );
  AOI22_X1 U5160 ( .A1(n4685), .A2(n4696), .B1(n4650), .B2(n4683), .ZN(U3473)
         );
  INV_X1 U5161 ( .A(n4651), .ZN(n4653) );
  AOI211_X1 U5162 ( .C1(n4654), .C2(n4679), .A(n4653), .B(n4652), .ZN(n4697)
         );
  INV_X1 U5163 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5164 ( .A1(n4685), .A2(n4697), .B1(n4655), .B2(n4683), .ZN(U3475)
         );
  NOR3_X1 U5165 ( .A1(n4657), .A2(n4656), .A3(n4667), .ZN(n4659) );
  AOI211_X1 U5166 ( .C1(n4679), .C2(n4660), .A(n4659), .B(n4658), .ZN(n4699)
         );
  AOI22_X1 U5167 ( .A1(n4685), .A2(n4699), .B1(n4661), .B2(n4683), .ZN(U3479)
         );
  AOI211_X1 U5168 ( .C1(n4665), .C2(n4664), .A(n4663), .B(n4662), .ZN(n4700)
         );
  INV_X1 U5169 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5170 ( .A1(n4685), .A2(n4700), .B1(n4666), .B2(n4683), .ZN(U3481)
         );
  NOR3_X1 U5171 ( .A1(n4669), .A2(n4668), .A3(n4667), .ZN(n4671) );
  AOI211_X1 U5172 ( .C1(n4672), .C2(n4679), .A(n4671), .B(n4670), .ZN(n4701)
         );
  INV_X1 U5173 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5174 ( .A1(n4685), .A2(n4701), .B1(n4673), .B2(n4683), .ZN(U3483)
         );
  NAND2_X1 U5175 ( .A1(n4675), .A2(n4674), .ZN(n4676) );
  NOR2_X1 U5176 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  AOI21_X1 U5177 ( .B1(n4680), .B2(n4679), .A(n4678), .ZN(n4681) );
  INV_X1 U5178 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5179 ( .A1(n4685), .A2(n4703), .B1(n4684), .B2(n4683), .ZN(U3487)
         );
  AOI22_X1 U5180 ( .A1(n4704), .A2(n4687), .B1(n4686), .B2(n4702), .ZN(U3518)
         );
  OAI22_X1 U5181 ( .A1(n4690), .A2(n4689), .B1(n4704), .B2(n4688), .ZN(n4691)
         );
  INV_X1 U5182 ( .A(n4691), .ZN(n4692) );
  OAI21_X1 U5183 ( .B1(n4693), .B2(n4702), .A(n4692), .ZN(U3519) );
  AOI22_X1 U5184 ( .A1(n4704), .A2(n4695), .B1(n4694), .B2(n4702), .ZN(U3520)
         );
  AOI22_X1 U5185 ( .A1(n4704), .A2(n4696), .B1(n2374), .B2(n4702), .ZN(U3521)
         );
  AOI22_X1 U5186 ( .A1(n4704), .A2(n4697), .B1(n2378), .B2(n4702), .ZN(U3522)
         );
  AOI22_X1 U5187 ( .A1(n4704), .A2(n4699), .B1(n4698), .B2(n4702), .ZN(U3524)
         );
  AOI22_X1 U5188 ( .A1(n4704), .A2(n4700), .B1(n2409), .B2(n4702), .ZN(U3525)
         );
  AOI22_X1 U5189 ( .A1(n4704), .A2(n4701), .B1(n2420), .B2(n4702), .ZN(U3526)
         );
  AOI22_X1 U5190 ( .A1(n4704), .A2(n4703), .B1(n2439), .B2(n4702), .ZN(U3528)
         );
  AOI21_X1 U2358 ( .B1(n3734), .B2(n3956), .A(n4083), .ZN(n2559) );
  CLKBUF_X1 U2316 ( .A(n2720), .Z(n2825) );
  AND2_X1 U2368 ( .A1(n2939), .A2(n3132), .ZN(n2909) );
  CLKBUF_X1 U35070 ( .A(n3857), .Z(n3856) );
  NOR2_X1 U35350 ( .A1(n4223), .A2(n4202), .ZN(n4197) );
  AND2_X1 U35470 ( .A1(n2671), .A2(n2670), .ZN(n4674) );
endmodule

