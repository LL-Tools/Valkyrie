

module b20_C_gen_AntiSAT_k_256_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4502, n4503, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537;

  NOR2_X2 U5008 ( .A1(n9741), .A2(n9578), .ZN(n9577) );
  AOI22_X1 U5009 ( .A1(n9609), .A2(n5806), .B1(n9806), .B2(n9630), .ZN(n9595)
         );
  NAND2_X1 U5010 ( .A1(n5057), .A2(n4539), .ZN(n9656) );
  INV_X1 U5011 ( .A(n8957), .ZN(n8940) );
  NAND2_X1 U5012 ( .A1(n7566), .A2(n7568), .ZN(n7567) );
  INV_X1 U5013 ( .A(n5574), .ZN(n5867) );
  INV_X1 U5014 ( .A(n6163), .ZN(n6125) );
  CLKBUF_X2 U5015 ( .A(n4542), .Z(n5594) );
  INV_X2 U5016 ( .A(n6966), .ZN(n5571) );
  NAND4_X1 U5017 ( .A1(n5536), .A2(n5535), .A3(n5534), .A4(n5533), .ZN(n5964)
         );
  AND3_X2 U5018 ( .A1(n5544), .A2(n4792), .A3(n4791), .ZN(n8454) );
  AND2_X4 U5019 ( .A1(n5497), .A2(n9824), .ZN(n5547) );
  INV_X1 U5020 ( .A(n5982), .ZN(n6157) );
  INV_X1 U5021 ( .A(n6161), .ZN(n6131) );
  NAND2_X1 U5022 ( .A1(n9595), .A2(n5807), .ZN(n5808) );
  INV_X1 U5023 ( .A(n9366), .ZN(n5559) );
  NOR2_X1 U5024 ( .A1(n4873), .A2(n5490), .ZN(n5493) );
  OR2_X1 U5025 ( .A1(n9140), .A2(n8640), .ZN(n6571) );
  AND2_X1 U5026 ( .A1(n9140), .A2(n8640), .ZN(n6743) );
  INV_X1 U5027 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5128) );
  INV_X1 U5028 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6233) );
  OR2_X1 U5029 ( .A1(n9493), .A2(n9503), .ZN(n9482) );
  NAND2_X1 U5030 ( .A1(n8130), .A2(n8129), .ZN(n8542) );
  XNOR2_X1 U5031 ( .A(n5189), .B(n6410), .ZN(n8805) );
  OAI21_X1 U5032 ( .B1(n8805), .B2(n4859), .A(n4858), .ZN(n8820) );
  NAND2_X1 U5033 ( .A1(n5414), .A2(n5410), .ZN(n5411) );
  OAI21_X2 U5034 ( .B1(n8118), .B2(n5000), .A(n4999), .ZN(n4998) );
  NAND2_X2 U5035 ( .A1(n7980), .A2(n7979), .ZN(n8118) );
  OAI21_X2 U5036 ( .B1(n6851), .B2(P2_D_REG_0__SCAN_IN), .A(n7102), .ZN(n6852)
         );
  NAND2_X2 U5037 ( .A1(n6848), .A2(n6847), .ZN(n6851) );
  NAND2_X2 U5038 ( .A1(n5150), .A2(n5158), .ZN(n9937) );
  NAND4_X2 U5039 ( .A1(n5539), .A2(n5540), .A3(n4793), .A4(n4794), .ZN(n5545)
         );
  XNOR2_X2 U5040 ( .A(n6232), .B(n9209), .ZN(n6239) );
  NAND2_X2 U5041 ( .A1(n9208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6232) );
  NAND2_X2 U5042 ( .A1(n5412), .A2(n5411), .ZN(n5922) );
  AOI21_X2 U5043 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(n8128) );
  NAND2_X2 U5044 ( .A1(n4998), .A2(n4997), .ZN(n8063) );
  NAND2_X2 U5045 ( .A1(n5257), .A2(n5154), .ZN(n7150) );
  AOI22_X2 U5046 ( .A1(n9656), .A2(n5771), .B1(n9766), .B2(n9415), .ZN(n9641)
         );
  XNOR2_X2 U5047 ( .A(n5202), .B(n5201), .ZN(n8838) );
  OAI21_X2 U5048 ( .B1(n9972), .B2(n4864), .A(n4863), .ZN(n9996) );
  XNOR2_X2 U5049 ( .A(n5187), .B(n6388), .ZN(n9972) );
  INV_X4 U5050 ( .A(n6158), .ZN(n5972) );
  OAI21_X1 U5051 ( .B1(n9259), .B2(n6056), .A(n6055), .ZN(n6061) );
  NAND2_X2 U5052 ( .A1(n6609), .A2(n6613), .ZN(n6776) );
  NAND2_X4 U5053 ( .A1(n7345), .A2(n5951), .ZN(n6158) );
  NAND4_X1 U5054 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n8780)
         );
  INV_X8 U5055 ( .A(n6881), .ZN(n6837) );
  BUF_X2 U5056 ( .A(n5585), .Z(n8393) );
  BUF_X4 U5057 ( .A(n6265), .Z(n4502) );
  INV_X2 U5058 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U5059 ( .B1(n4804), .B2(n4805), .A(n4592), .ZN(n4661) );
  AND2_X1 U5060 ( .A1(n4892), .A2(n4608), .ZN(n5942) );
  AND2_X1 U5061 ( .A1(n9513), .A2(n9512), .ZN(n9722) );
  OR2_X1 U5062 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  AND2_X1 U5063 ( .A1(n4778), .A2(n4777), .ZN(n8610) );
  NOR2_X1 U5064 ( .A1(n4811), .A2(n4817), .ZN(n4810) );
  NAND2_X1 U5065 ( .A1(n8533), .A2(n4808), .ZN(n4805) );
  OAI21_X1 U5066 ( .B1(n4634), .B2(n4633), .A(n4630), .ZN(n5019) );
  NAND2_X1 U5067 ( .A1(n4611), .A2(n4616), .ZN(n9236) );
  NAND2_X1 U5068 ( .A1(n9233), .A2(n6081), .ZN(n9239) );
  AND2_X1 U5069 ( .A1(n9400), .A2(n9399), .ZN(n9404) );
  NAND2_X1 U5070 ( .A1(n9041), .A2(n6806), .ZN(n9038) );
  OAI21_X1 U5071 ( .B1(n7963), .B2(n4751), .A(n4747), .ZN(n8084) );
  NAND2_X1 U5072 ( .A1(n7879), .A2(n6336), .ZN(n7963) );
  NAND2_X1 U5073 ( .A1(n4526), .A2(n6001), .ZN(n7528) );
  AND2_X1 U5074 ( .A1(n8465), .A2(n8462), .ZN(n7600) );
  AND2_X1 U5075 ( .A1(n4851), .A2(n5181), .ZN(n5182) );
  NAND2_X1 U5076 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  INV_X2 U5077 ( .A(n10061), .ZN(n10052) );
  NOR2_X1 U5078 ( .A1(n7507), .A2(n5083), .ZN(n5175) );
  AND2_X1 U5079 ( .A1(n5965), .A2(n5030), .ZN(n5968) );
  INV_X1 U5080 ( .A(n9490), .ZN(n9856) );
  AND2_X1 U5081 ( .A1(n5573), .A2(n4720), .ZN(n9860) );
  NAND4_X1 U5082 ( .A1(n6288), .A2(n6287), .A3(n6286), .A4(n6285), .ZN(n8778)
         );
  NAND2_X2 U5083 ( .A1(n5949), .A2(n5951), .ZN(n6161) );
  NAND4_X1 U5084 ( .A1(n6271), .A2(n6270), .A3(n6269), .A4(n6268), .ZN(n8781)
         );
  AND3_X2 U5085 ( .A1(n6264), .A2(n6263), .A3(n6262), .ZN(n7953) );
  OAI211_X1 U5086 ( .C1(n5574), .C2(n6937), .A(n5554), .B(n5553), .ZN(n9366)
         );
  AND2_X1 U5087 ( .A1(n5162), .A2(n6902), .ZN(n9949) );
  AND2_X1 U5088 ( .A1(n6966), .A2(n6272), .ZN(n5585) );
  MUX2_X1 U5089 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5422), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5424) );
  INV_X2 U5090 ( .A(n6834), .ZN(n8864) );
  AND2_X1 U5091 ( .A1(n9824), .A2(n5499), .ZN(n5538) );
  INV_X1 U5092 ( .A(n5498), .ZN(n9824) );
  INV_X1 U5093 ( .A(n5428), .ZN(n4503) );
  NAND2_X1 U5094 ( .A1(n4525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5119) );
  NAND3_X1 U5095 ( .A1(n5496), .A2(n9817), .A3(n5495), .ZN(n5498) );
  OR2_X1 U5096 ( .A1(n6234), .A2(n6233), .ZN(n6236) );
  OR2_X1 U5097 ( .A1(n5493), .A2(n5625), .ZN(n5491) );
  MUX2_X1 U5098 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5413), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5415) );
  AND2_X1 U5099 ( .A1(n5114), .A2(n4754), .ZN(n6234) );
  INV_X2 U5100 ( .A(n9213), .ZN(n8665) );
  AND2_X1 U5101 ( .A1(n4512), .A2(n5059), .ZN(n5463) );
  NOR3_X1 U5102 ( .A1(n4505), .A2(P2_IR_REG_28__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .ZN(n4754) );
  OR2_X1 U5103 ( .A1(n5005), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5104 ( .A1(n5291), .A2(n5292), .ZN(n5313) );
  NAND2_X1 U5105 ( .A1(n5259), .A2(n5094), .ZN(n5163) );
  AND2_X2 U5106 ( .A1(n7147), .A2(n4857), .ZN(n5259) );
  AND4_X1 U5107 ( .A1(n5087), .A2(n5133), .A3(n5126), .A4(n5164), .ZN(n5093)
         );
  AND4_X1 U5108 ( .A1(n5168), .A2(n5128), .A3(n5089), .A4(n5088), .ZN(n5090)
         );
  AND2_X1 U5109 ( .A1(n5401), .A2(n10408), .ZN(n5453) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4610) );
  INV_X1 U5111 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5094) );
  INV_X1 U5113 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5126) );
  NOR3_X1 U5114 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5103) );
  INV_X1 U5115 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4788) );
  INV_X1 U5116 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5133) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5449) );
  INV_X4 U5118 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5119 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4857) );
  INV_X1 U5120 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5168) );
  INV_X1 U5121 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U5122 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5092) );
  INV_X1 U5123 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5164) );
  NOR2_X1 U5124 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5091) );
  OAI22_X1 U5125 ( .A1(n8956), .A2(n8955), .B1(n8969), .B2(n9161), .ZN(n8601)
         );
  AOI21_X2 U5126 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9984), .A(n9996), .ZN(
        n5189) );
  AOI22_X2 U5127 ( .A1(n9641), .A2(n5781), .B1(n9653), .B2(n9663), .ZN(n9626)
         );
  NOR2_X2 U5128 ( .A1(n8820), .A2(n5196), .ZN(n5202) );
  NAND2_X2 U5129 ( .A1(n6238), .A2(n6241), .ZN(n6283) );
  AND2_X1 U5130 ( .A1(n6239), .A2(n6240), .ZN(n6265) );
  AOI21_X1 U5131 ( .B1(n4828), .B2(n4830), .A(n8376), .ZN(n4827) );
  INV_X1 U5132 ( .A(n4831), .ZN(n4830) );
  AND2_X1 U5133 ( .A1(n5099), .A2(n4698), .ZN(n4697) );
  AND2_X1 U5134 ( .A1(n5021), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5135 ( .A1(n4632), .A2(n6104), .ZN(n4631) );
  INV_X1 U5136 ( .A(n5009), .ZN(n4632) );
  NAND2_X1 U5137 ( .A1(n5383), .A2(n5382), .ZN(n5849) );
  XNOR2_X1 U5138 ( .A(n5465), .B(n5419), .ZN(n8525) );
  AOI21_X1 U5139 ( .B1(n4939), .B2(n4649), .A(n4648), .ZN(n4647) );
  INV_X1 U5140 ( .A(n5346), .ZN(n4649) );
  NAND2_X1 U5141 ( .A1(n4650), .A2(n5346), .ZN(n5732) );
  AOI21_X1 U5142 ( .B1(n5610), .B2(n4952), .A(n4951), .ZN(n4950) );
  INV_X1 U5143 ( .A(n5322), .ZN(n4952) );
  INV_X1 U5144 ( .A(n5325), .ZN(n4951) );
  AOI21_X1 U5145 ( .B1(n9317), .B2(n9318), .A(n4628), .ZN(n4627) );
  INV_X1 U5146 ( .A(n6137), .ZN(n4628) );
  AND2_X1 U5147 ( .A1(n8495), .A2(n8290), .ZN(n9509) );
  OAI211_X1 U5148 ( .C1(n4800), .C2(n5906), .A(n4803), .B(n4798), .ZN(n8300)
         );
  NAND2_X1 U5149 ( .A1(n8294), .A2(n4976), .ZN(n4803) );
  MUX2_X1 U5150 ( .A(n8331), .B(n8330), .S(n8398), .Z(n8337) );
  OR2_X1 U5151 ( .A1(n8368), .A2(n4826), .ZN(n4822) );
  INV_X1 U5152 ( .A(n4827), .ZN(n4826) );
  NAND2_X1 U5153 ( .A1(n8290), .A2(n8289), .ZN(n8389) );
  OR2_X1 U5154 ( .A1(n9741), .A2(n9553), .ZN(n8438) );
  NOR2_X1 U5155 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5401) );
  INV_X1 U5156 ( .A(n5506), .ZN(n5348) );
  OR2_X1 U5157 ( .A1(n5654), .A2(n4598), .ZN(n4597) );
  NAND2_X1 U5158 ( .A1(n4967), .A2(n4599), .ZN(n4598) );
  INV_X1 U5159 ( .A(n5653), .ZN(n4599) );
  AOI21_X1 U5160 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(n6760) );
  NOR2_X1 U5161 ( .A1(n8902), .A2(n6742), .ZN(n6746) );
  OAI21_X1 U5162 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n6747) );
  INV_X1 U5163 ( .A(n6240), .ZN(n6241) );
  INV_X1 U5164 ( .A(n6795), .ZN(n4762) );
  OR2_X1 U5165 ( .A1(n8780), .A2(n10024), .ZN(n6617) );
  INV_X1 U5166 ( .A(n8914), .ZN(n6820) );
  OR2_X1 U5167 ( .A1(n8618), .A2(n8939), .ZN(n6735) );
  OR2_X1 U5168 ( .A1(n9178), .A2(n9003), .ZN(n8595) );
  OR2_X1 U5169 ( .A1(n9201), .A2(n8211), .ZN(n6683) );
  INV_X1 U5170 ( .A(n6801), .ZN(n4779) );
  INV_X1 U5171 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5118) );
  INV_X1 U5172 ( .A(n5080), .ZN(n5016) );
  AOI21_X1 U5173 ( .B1(n4552), .B2(n8495), .A(n4517), .ZN(n4818) );
  OR2_X1 U5174 ( .A1(n9730), .A2(n9554), .ZN(n8490) );
  NAND2_X1 U5175 ( .A1(n9601), .A2(n4603), .ZN(n4897) );
  NOR2_X1 U5176 ( .A1(n4901), .A2(n4604), .ZN(n4603) );
  INV_X1 U5177 ( .A(n8369), .ZN(n4604) );
  INV_X1 U5178 ( .A(n5920), .ZN(n4901) );
  NAND2_X1 U5179 ( .A1(n9590), .A2(n4954), .ZN(n8374) );
  INV_X1 U5180 ( .A(n4707), .ZN(n4706) );
  OAI21_X1 U5181 ( .B1(n5047), .B2(n4708), .A(n5081), .ZN(n4707) );
  NAND2_X1 U5182 ( .A1(n5056), .A2(n5743), .ZN(n5055) );
  INV_X1 U5183 ( .A(n9704), .ZN(n5056) );
  INV_X1 U5184 ( .A(n7107), .ZN(n8410) );
  NAND2_X1 U5185 ( .A1(n5922), .A2(n5926), .ZN(n6966) );
  XNOR2_X1 U5186 ( .A(n6199), .B(n6198), .ZN(n6201) );
  AND2_X1 U5187 ( .A1(n5862), .A2(n5387), .ZN(n5848) );
  NAND2_X1 U5188 ( .A1(n5377), .A2(n5376), .ZN(n4930) );
  NAND2_X1 U5189 ( .A1(n4956), .A2(n4957), .ZN(n5484) );
  AOI21_X1 U5190 ( .B1(n4958), .B2(n4960), .A(n4577), .ZN(n4957) );
  NAND2_X1 U5191 ( .A1(n5773), .A2(n4958), .ZN(n4956) );
  INV_X1 U5192 ( .A(SI_11_), .ZN(n10263) );
  NAND2_X1 U5193 ( .A1(n5338), .A2(SI_12_), .ZN(n5339) );
  OR2_X1 U5194 ( .A1(n5660), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U5195 ( .A1(n4904), .A2(n4950), .ZN(n5638) );
  NAND2_X1 U5196 ( .A1(n4516), .A2(n4902), .ZN(n4904) );
  XNOR2_X1 U5197 ( .A(n5123), .B(n5122), .ZN(n5209) );
  NAND2_X1 U5198 ( .A1(n4511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5123) );
  INV_X1 U5199 ( .A(n6283), .ZN(n6550) );
  NOR2_X1 U5200 ( .A1(n8233), .A2(n6844), .ZN(n5110) );
  OAI21_X1 U5201 ( .B1(n5289), .B2(n8863), .A(n4685), .ZN(n4684) );
  INV_X1 U5202 ( .A(n5287), .ZN(n4685) );
  NAND2_X1 U5203 ( .A1(n4868), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5204 ( .A1(n5203), .A2(n4868), .ZN(n4866) );
  INV_X1 U5205 ( .A(n5206), .ZN(n4868) );
  NAND2_X1 U5206 ( .A1(n9145), .A2(n8939), .ZN(n4777) );
  NAND2_X1 U5207 ( .A1(n9178), .A2(n8977), .ZN(n4786) );
  AND2_X1 U5208 ( .A1(n8980), .A2(n4786), .ZN(n4785) );
  OR2_X1 U5209 ( .A1(n9188), .A2(n9037), .ZN(n6696) );
  OAI21_X1 U5210 ( .B1(n8084), .B2(n6655), .A(n6664), .ZN(n8163) );
  NAND2_X1 U5211 ( .A1(n6399), .A2(n6398), .ZN(n9052) );
  NOR2_X1 U5212 ( .A1(n4584), .A2(n4740), .ZN(n4739) );
  NOR2_X1 U5213 ( .A1(n5112), .A2(n4505), .ZN(n6231) );
  XNOR2_X1 U5214 ( .A(n5119), .B(n5118), .ZN(n6772) );
  INV_X1 U5215 ( .A(n5313), .ZN(n6272) );
  NOR2_X1 U5216 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  NAND2_X1 U5217 ( .A1(n4627), .A2(n4624), .ZN(n4623) );
  INV_X1 U5218 ( .A(n9317), .ZN(n4624) );
  INV_X1 U5219 ( .A(n4627), .ZN(n4625) );
  OAI21_X1 U5220 ( .B1(n8053), .B2(n4614), .A(n4612), .ZN(n9400) );
  NOR2_X1 U5221 ( .A1(n4510), .A2(n4616), .ZN(n4614) );
  AOI22_X1 U5222 ( .A1(n4510), .A2(n4547), .B1(n4616), .B2(n4613), .ZN(n4612)
         );
  INV_X1 U5223 ( .A(n8001), .ZN(n8537) );
  AOI211_X1 U5224 ( .C1(n8531), .C2(n8530), .A(n8529), .B(n8528), .ZN(n8532)
         );
  AND4_X1 U5225 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n6150)
         );
  INV_X1 U5226 ( .A(n5538), .ZN(n5803) );
  NOR2_X1 U5227 ( .A1(n9525), .A2(n5045), .ZN(n5044) );
  INV_X1 U5228 ( .A(n5860), .ZN(n5045) );
  AOI21_X1 U5229 ( .B1(n5036), .B2(n5034), .A(n4573), .ZN(n5033) );
  AOI21_X1 U5230 ( .B1(n4927), .B2(n4926), .A(n4925), .ZN(n4924) );
  INV_X1 U5231 ( .A(n8366), .ZN(n4925) );
  INV_X1 U5232 ( .A(n9627), .ZN(n4926) );
  OAI21_X1 U5233 ( .B1(n7894), .B2(n4708), .A(n4706), .ZN(n5744) );
  OR2_X1 U5234 ( .A1(n7863), .A2(n7873), .ZN(n8314) );
  OR2_X1 U5235 ( .A1(n9422), .A2(n7863), .ZN(n5635) );
  NAND2_X1 U5236 ( .A1(n7342), .A2(n9860), .ZN(n5575) );
  NOR2_X1 U5237 ( .A1(n5472), .A2(n5471), .ZN(n5474) );
  NAND2_X1 U5238 ( .A1(n4959), .A2(n4961), .ZN(n5794) );
  OR2_X1 U5239 ( .A1(n5773), .A2(n4960), .ZN(n4959) );
  OAI21_X1 U5240 ( .B1(n5732), .B2(n4944), .A(n4942), .ZN(n5746) );
  INV_X1 U5241 ( .A(n9590), .ZN(n9256) );
  XNOR2_X1 U5242 ( .A(n4595), .B(n8434), .ZN(n5929) );
  NAND2_X1 U5243 ( .A1(n9507), .A2(n8290), .ZN(n4595) );
  NAND2_X1 U5244 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  NAND2_X1 U5245 ( .A1(n6652), .A2(n6651), .ZN(n6657) );
  NAND2_X1 U5246 ( .A1(n4845), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U5247 ( .A1(n8306), .A2(n8398), .ZN(n4845) );
  AOI21_X1 U5248 ( .B1(n8308), .B2(n8309), .A(n4844), .ZN(n4843) );
  INV_X1 U5249 ( .A(n8313), .ZN(n4841) );
  NAND2_X1 U5250 ( .A1(n8321), .A2(n4837), .ZN(n8323) );
  NOR2_X1 U5251 ( .A1(n4839), .A2(n4838), .ZN(n4837) );
  INV_X1 U5252 ( .A(n8319), .ZN(n4838) );
  NAND2_X1 U5253 ( .A1(n8342), .A2(n4849), .ZN(n4848) );
  AND2_X1 U5254 ( .A1(n4850), .A2(n8341), .ZN(n4849) );
  OR2_X1 U5255 ( .A1(n8343), .A2(n9408), .ZN(n4850) );
  AND2_X1 U5256 ( .A1(n4834), .A2(n4829), .ZN(n4828) );
  INV_X1 U5257 ( .A(n8372), .ZN(n4834) );
  NAND2_X1 U5258 ( .A1(n4831), .A2(n4836), .ZN(n4829) );
  INV_X1 U5259 ( .A(n9558), .ZN(n4655) );
  AND2_X1 U5260 ( .A1(n9611), .A2(n4531), .ZN(n4654) );
  OR2_X1 U5261 ( .A1(n9483), .A2(n8432), .ZN(n8516) );
  INV_X1 U5262 ( .A(n4936), .ZN(n4648) );
  AOI21_X1 U5263 ( .B1(n4938), .B2(n4942), .A(n4937), .ZN(n4936) );
  INV_X1 U5264 ( .A(n5353), .ZN(n4937) );
  AND2_X1 U5265 ( .A1(n4944), .A2(n4941), .ZN(n4938) );
  NOR2_X1 U5266 ( .A1(n5349), .A2(n4946), .ZN(n4945) );
  INV_X1 U5267 ( .A(n4948), .ZN(n4946) );
  INV_X1 U5268 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10230) );
  AND2_X1 U5269 ( .A1(n7683), .A2(n7681), .ZN(n7750) );
  OAI21_X1 U5270 ( .B1(n7150), .B2(n5155), .A(n5156), .ZN(n7157) );
  NAND2_X1 U5271 ( .A1(n8797), .A2(n5270), .ZN(n5271) );
  NAND2_X1 U5272 ( .A1(n8043), .A2(n4663), .ZN(n5276) );
  OR2_X1 U5273 ( .A1(n6377), .A2(n6380), .ZN(n4663) );
  OR2_X1 U5274 ( .A1(n8727), .A2(n8992), .ZN(n6716) );
  INV_X1 U5275 ( .A(n4761), .ZN(n4760) );
  OAI21_X1 U5276 ( .B1(n6794), .B2(n4762), .A(n6796), .ZN(n4761) );
  NAND2_X1 U5277 ( .A1(n8030), .A2(n4688), .ZN(n6651) );
  OR2_X1 U5278 ( .A1(n8775), .A2(n7710), .ZN(n6789) );
  OR2_X1 U5279 ( .A1(n9161), .A2(n8603), .ZN(n6721) );
  INV_X1 U5280 ( .A(n5103), .ZN(n5004) );
  NOR2_X1 U5281 ( .A1(n5005), .A2(n4696), .ZN(n4695) );
  INV_X1 U5282 ( .A(n4697), .ZN(n4696) );
  AND2_X1 U5283 ( .A1(n5096), .A2(n5097), .ZN(n5003) );
  INV_X1 U5284 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5097) );
  INV_X1 U5285 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5096) );
  OR2_X1 U5286 ( .A1(n5141), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5129) );
  NOR2_X1 U5287 ( .A1(n6088), .A2(n4618), .ZN(n4617) );
  INV_X1 U5288 ( .A(n8054), .ZN(n4618) );
  NAND2_X1 U5289 ( .A1(n5028), .A2(n5027), .ZN(n5029) );
  INV_X1 U5290 ( .A(n5949), .ZN(n5027) );
  INV_X1 U5291 ( .A(n5947), .ZN(n5028) );
  NAND3_X1 U5292 ( .A1(n4636), .A2(n4635), .A3(n4629), .ZN(n4634) );
  NOR2_X1 U5293 ( .A1(n9311), .A2(n5013), .ZN(n4635) );
  INV_X1 U5294 ( .A(n9404), .ZN(n4629) );
  INV_X1 U5295 ( .A(n6104), .ZN(n4633) );
  AND2_X1 U5296 ( .A1(n5022), .A2(n4560), .ZN(n5021) );
  OR2_X1 U5297 ( .A1(n6116), .A2(n9327), .ZN(n5022) );
  NAND2_X1 U5298 ( .A1(n6087), .A2(n4576), .ZN(n4616) );
  AND2_X1 U5299 ( .A1(n4822), .A2(n4555), .ZN(n8378) );
  NOR2_X1 U5300 ( .A1(n4833), .A2(n8389), .ZN(n4821) );
  NAND2_X1 U5301 ( .A1(n8434), .A2(n8495), .ZN(n4819) );
  NOR3_X1 U5302 ( .A1(n8386), .A2(n9483), .A3(n4819), .ZN(n4809) );
  OAI21_X1 U5303 ( .B1(n4816), .B2(n9483), .A(n4820), .ZN(n4813) );
  INV_X1 U5304 ( .A(n7845), .ZN(n4680) );
  OR2_X1 U5305 ( .A1(n9720), .A2(n9520), .ZN(n8495) );
  NOR2_X1 U5306 ( .A1(n9529), .A2(n4877), .ZN(n4876) );
  INV_X1 U5307 ( .A(n4878), .ZN(n4877) );
  NOR2_X1 U5308 ( .A1(n9730), .A2(n9562), .ZN(n4878) );
  INV_X1 U5309 ( .A(n5039), .ZN(n5034) );
  AOI21_X1 U5310 ( .B1(n5920), .B2(n4900), .A(n4899), .ZN(n4898) );
  INV_X1 U5311 ( .A(n8438), .ZN(n4899) );
  INV_X1 U5312 ( .A(n8430), .ZN(n4900) );
  NOR2_X1 U5313 ( .A1(n9618), .A2(n4881), .ZN(n4880) );
  INV_X1 U5314 ( .A(n4882), .ZN(n4881) );
  NOR2_X1 U5315 ( .A1(n9408), .A2(n4886), .ZN(n4885) );
  INV_X1 U5316 ( .A(n4887), .ZN(n4886) );
  AND2_X1 U5317 ( .A1(n7818), .A2(n9907), .ZN(n7817) );
  NOR2_X1 U5318 ( .A1(n8419), .A2(n5916), .ZN(n4910) );
  NOR2_X1 U5319 ( .A1(n5678), .A2(n5677), .ZN(n5695) );
  OR2_X1 U5320 ( .A1(n5646), .A2(n5645), .ZN(n5664) );
  NAND2_X1 U5321 ( .A1(n5913), .A2(n5912), .ZN(n8465) );
  INV_X1 U5322 ( .A(n8418), .ZN(n5912) );
  OR2_X1 U5323 ( .A1(n7480), .A2(n9265), .ZN(n8416) );
  OR2_X1 U5324 ( .A1(n9256), .A2(n9596), .ZN(n9578) );
  NOR2_X2 U5325 ( .A1(n9766), .A2(n9673), .ZN(n9664) );
  AND2_X1 U5326 ( .A1(n7609), .A2(n7717), .ZN(n7818) );
  INV_X1 U5327 ( .A(n5848), .ZN(n4933) );
  INV_X1 U5328 ( .A(n5879), .ZN(n4932) );
  INV_X1 U5329 ( .A(n5388), .ZN(n4934) );
  AND2_X1 U5330 ( .A1(n5599), .A2(n5060), .ZN(n5059) );
  NOR2_X1 U5331 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5060) );
  NOR2_X1 U5332 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5429) );
  AND2_X1 U5333 ( .A1(n5382), .A2(n5381), .ZN(n5834) );
  AND2_X1 U5334 ( .A1(n5376), .A2(n5375), .ZN(n5822) );
  INV_X1 U5335 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5476) );
  AOI21_X1 U5336 ( .B1(n4580), .B2(n5362), .A(n4962), .ZN(n4961) );
  NOR2_X1 U5337 ( .A1(n5361), .A2(SI_20_), .ZN(n4962) );
  NOR2_X1 U5338 ( .A1(n4545), .A2(n5025), .ZN(n5024) );
  INV_X1 U5339 ( .A(n5452), .ZN(n5025) );
  NAND2_X1 U5340 ( .A1(n4597), .A2(n4964), .ZN(n5704) );
  NOR2_X1 U5341 ( .A1(n5671), .A2(n4971), .ZN(n4970) );
  INV_X1 U5342 ( .A(n5334), .ZN(n4971) );
  OR2_X1 U5343 ( .A1(n5688), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5689) );
  NOR2_X1 U5344 ( .A1(n5330), .A2(n5637), .ZN(n4646) );
  NOR2_X1 U5345 ( .A1(n5061), .A2(n5062), .ZN(n5332) );
  OAI21_X1 U5346 ( .B1(n6272), .B2(n4602), .A(n4601), .ZN(n5319) );
  NAND2_X1 U5347 ( .A1(n6272), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4601) );
  OR2_X1 U5348 ( .A1(n5603), .A2(n4789), .ZN(n4903) );
  NAND3_X1 U5349 ( .A1(n5584), .A2(n5312), .A3(n5318), .ZN(n4902) );
  INV_X1 U5350 ( .A(n5291), .ZN(n4709) );
  AOI21_X1 U5351 ( .B1(n8556), .B2(n8688), .A(n8693), .ZN(n4995) );
  NAND2_X1 U5352 ( .A1(n4994), .A2(n8692), .ZN(n4993) );
  NAND2_X1 U5353 ( .A1(n4995), .A2(n4996), .ZN(n4994) );
  INV_X1 U5354 ( .A(n8556), .ZN(n4996) );
  INV_X1 U5355 ( .A(n8719), .ZN(n4986) );
  INV_X1 U5356 ( .A(n8574), .ZN(n4981) );
  NOR2_X1 U5357 ( .A1(n8728), .A2(n8729), .ZN(n8556) );
  INV_X1 U5358 ( .A(n7987), .ZN(n4999) );
  NAND2_X1 U5359 ( .A1(n6751), .A2(n6881), .ZN(n6758) );
  NAND2_X1 U5360 ( .A1(n6750), .A2(n5073), .ZN(n6751) );
  AND2_X1 U5361 ( .A1(n4731), .A2(n4729), .ZN(n4728) );
  INV_X1 U5362 ( .A(n5074), .ZN(n4732) );
  AND4_X1 U5363 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n8558)
         );
  INV_X1 U5364 ( .A(n8790), .ZN(n4852) );
  XNOR2_X1 U5365 ( .A(n5271), .B(n6353), .ZN(n7780) );
  NAND2_X1 U5366 ( .A1(n7780), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U5367 ( .A1(n4872), .A2(n4871), .ZN(n4870) );
  INV_X1 U5368 ( .A(n7824), .ZN(n4871) );
  NAND2_X1 U5369 ( .A1(n8044), .A2(n8045), .ZN(n8043) );
  XNOR2_X1 U5370 ( .A(n5276), .B(n6388), .ZN(n9966) );
  NAND2_X1 U5371 ( .A1(n9987), .A2(n9988), .ZN(n9986) );
  XNOR2_X1 U5372 ( .A(n5278), .B(n6410), .ZN(n8815) );
  NAND2_X1 U5373 ( .A1(n9986), .A2(n4668), .ZN(n5278) );
  NAND2_X1 U5374 ( .A1(n9984), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4668) );
  OR2_X1 U5375 ( .A1(n8805), .A2(n9048), .ZN(n4861) );
  NAND2_X1 U5376 ( .A1(n6753), .A2(n6749), .ZN(n6829) );
  NAND2_X1 U5377 ( .A1(n6226), .A2(n10254), .ZN(n6476) );
  INV_X1 U5378 ( .A(n6469), .ZN(n6226) );
  OR2_X1 U5379 ( .A1(n6443), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6454) );
  AOI21_X1 U5380 ( .B1(n9038), .B2(n6810), .A(n4524), .ZN(n9014) );
  OR2_X1 U5381 ( .A1(n6371), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6381) );
  OR2_X1 U5382 ( .A1(n6315), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U5383 ( .A1(n6304), .A2(n6624), .ZN(n7632) );
  AND2_X1 U5384 ( .A1(n6547), .A2(n6546), .ZN(n6825) );
  AOI21_X1 U5385 ( .B1(n4765), .B2(n6823), .A(n6822), .ZN(n4764) );
  NAND2_X1 U5386 ( .A1(n8890), .A2(n9057), .ZN(n8893) );
  XNOR2_X1 U5387 ( .A(n9134), .B(n8905), .ZN(n8888) );
  NOR2_X1 U5388 ( .A1(n4734), .A2(n6740), .ZN(n4733) );
  INV_X1 U5389 ( .A(n6520), .ZN(n4734) );
  INV_X1 U5390 ( .A(n4770), .ZN(n4767) );
  AND2_X1 U5391 ( .A1(n6483), .A2(n6482), .ZN(n8939) );
  OR2_X1 U5392 ( .A1(n9167), .A2(n8558), .ZN(n8952) );
  AOI21_X1 U5393 ( .B1(n4785), .B2(n8991), .A(n4549), .ZN(n4784) );
  OR2_X1 U5394 ( .A1(n8990), .A2(n8991), .ZN(n4787) );
  AND2_X1 U5395 ( .A1(n8595), .A2(n6711), .ZN(n8991) );
  NOR2_X1 U5396 ( .A1(n6576), .A2(n4743), .ZN(n4742) );
  INV_X1 U5397 ( .A(n6684), .ZN(n4743) );
  AND4_X1 U5398 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n9037)
         );
  NAND2_X1 U5399 ( .A1(n9052), .A2(n6683), .ZN(n4744) );
  AND2_X1 U5400 ( .A1(n7288), .A2(n6837), .ZN(n9057) );
  AND2_X1 U5401 ( .A1(n6836), .A2(n6837), .ZN(n9055) );
  NAND2_X1 U5402 ( .A1(n6864), .A2(n6828), .ZN(n9060) );
  INV_X1 U5403 ( .A(n6558), .ZN(n6451) );
  INV_X1 U5404 ( .A(n6261), .ZN(n6450) );
  NAND2_X1 U5405 ( .A1(n6798), .A2(n4781), .ZN(n4780) );
  NOR2_X1 U5406 ( .A1(n6800), .A2(n4782), .ZN(n4781) );
  INV_X1 U5407 ( .A(n6797), .ZN(n4782) );
  INV_X1 U5408 ( .A(n9055), .ZN(n9004) );
  INV_X1 U5409 ( .A(n9057), .ZN(n9036) );
  NAND2_X1 U5410 ( .A1(n8169), .A2(n6387), .ZN(n4741) );
  NAND2_X1 U5411 ( .A1(n7998), .A2(n6604), .ZN(n10054) );
  OR2_X1 U5412 ( .A1(n7251), .A2(n9206), .ZN(n7261) );
  INV_X1 U5413 ( .A(n9060), .ZN(n8989) );
  AND2_X1 U5414 ( .A1(n7245), .A2(n7254), .ZN(n7258) );
  NAND2_X1 U5415 ( .A1(n5100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U5416 ( .A1(n5107), .A2(n5106), .ZN(n5108) );
  XNOR2_X1 U5417 ( .A(n5113), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6831) );
  AND2_X1 U5418 ( .A1(n5117), .A2(n5112), .ZN(n6865) );
  AND2_X1 U5419 ( .A1(n4528), .A2(n5098), .ZN(n4509) );
  INV_X1 U5420 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U5421 ( .A1(n6030), .A2(n6033), .ZN(n5018) );
  NAND2_X1 U5422 ( .A1(n7567), .A2(n4642), .ZN(n6030) );
  AND2_X1 U5423 ( .A1(n4643), .A2(n6024), .ZN(n4642) );
  INV_X1 U5424 ( .A(n6028), .ZN(n4643) );
  NOR2_X1 U5425 ( .A1(n4640), .A2(n4641), .ZN(n4639) );
  INV_X1 U5426 ( .A(n5999), .ZN(n4641) );
  NOR2_X1 U5427 ( .A1(n5016), .A2(n5015), .ZN(n5010) );
  INV_X1 U5428 ( .A(n9398), .ZN(n4636) );
  NAND2_X1 U5429 ( .A1(n4621), .A2(n4620), .ZN(n9382) );
  AOI21_X1 U5430 ( .B1(n4507), .B2(n4625), .A(n4578), .ZN(n4620) );
  AND4_X1 U5431 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n6182)
         );
  NAND2_X1 U5432 ( .A1(n5800), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5433 ( .A1(n6980), .A2(n9432), .ZN(n7092) );
  NAND2_X1 U5434 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5435 ( .A1(n7004), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4675) );
  AND2_X1 U5436 ( .A1(n4674), .A2(n4673), .ZN(n7017) );
  INV_X1 U5437 ( .A(n6989), .ZN(n4673) );
  NOR2_X1 U5438 ( .A1(n7017), .A2(n4672), .ZN(n7019) );
  AND2_X1 U5439 ( .A1(n7020), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5440 ( .A1(n7218), .A2(n4590), .ZN(n7221) );
  OR2_X1 U5441 ( .A1(n7735), .A2(n7734), .ZN(n7846) );
  NAND2_X1 U5442 ( .A1(n9517), .A2(n8289), .ZN(n9508) );
  NAND2_X1 U5443 ( .A1(n9508), .A2(n9509), .ZN(n9507) );
  NAND2_X1 U5444 ( .A1(n5043), .A2(n4543), .ZN(n9501) );
  AND2_X1 U5445 ( .A1(n5887), .A2(n5874), .ZN(n9530) );
  AND4_X1 U5446 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(n9553)
         );
  AND4_X1 U5447 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n9554)
         );
  NAND2_X1 U5448 ( .A1(n4897), .A2(n4898), .ZN(n9550) );
  NAND2_X1 U5449 ( .A1(n4897), .A2(n4895), .ZN(n9552) );
  NOR2_X1 U5450 ( .A1(n9558), .A2(n4896), .ZN(n4895) );
  INV_X1 U5451 ( .A(n4898), .ZN(n4896) );
  OR2_X1 U5452 ( .A1(n9745), .A2(n9614), .ZN(n5807) );
  AND2_X1 U5453 ( .A1(n8374), .A2(n9570), .ZN(n8430) );
  AOI21_X1 U5454 ( .B1(n4924), .B2(n4928), .A(n4832), .ZN(n4923) );
  AND2_X1 U5455 ( .A1(n8442), .A2(n8366), .ZN(n9611) );
  NAND2_X1 U5456 ( .A1(n5919), .A2(n8354), .ZN(n9628) );
  NAND2_X1 U5457 ( .A1(n9657), .A2(n4905), .ZN(n5919) );
  AND2_X1 U5458 ( .A1(n9640), .A2(n8349), .ZN(n4905) );
  INV_X1 U5459 ( .A(n9699), .ZN(n9662) );
  NAND2_X1 U5460 ( .A1(n9679), .A2(n4906), .ZN(n9657) );
  NOR2_X1 U5461 ( .A1(n9660), .A2(n4907), .ZN(n4906) );
  AND2_X1 U5462 ( .A1(n8341), .A2(n9678), .ZN(n9704) );
  OR2_X1 U5463 ( .A1(n5054), .A2(n5055), .ZN(n5053) );
  AOI21_X1 U5464 ( .B1(n4919), .B2(n8423), .A(n4918), .ZN(n4917) );
  INV_X1 U5465 ( .A(n8338), .ZN(n4918) );
  INV_X1 U5466 ( .A(n5716), .ZN(n5050) );
  NOR2_X1 U5467 ( .A1(n5049), .A2(n5048), .ZN(n5047) );
  INV_X1 U5468 ( .A(n4551), .ZN(n5049) );
  NOR2_X1 U5469 ( .A1(n8336), .A2(n4920), .ZN(n4919) );
  OR2_X1 U5470 ( .A1(n7895), .A2(n8423), .ZN(n4921) );
  XNOR2_X1 U5471 ( .A(n9783), .B(n9397), .ZN(n8336) );
  OR2_X1 U5472 ( .A1(n8147), .A2(n9418), .ZN(n5716) );
  NAND2_X1 U5473 ( .A1(n7894), .A2(n8423), .ZN(n7893) );
  OR2_X1 U5474 ( .A1(n9358), .A2(n9420), .ZN(n5683) );
  AND2_X1 U5475 ( .A1(n8419), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5476 ( .A1(n4718), .A2(n5652), .ZN(n4717) );
  INV_X1 U5477 ( .A(n7472), .ZN(n4718) );
  INV_X1 U5478 ( .A(n5652), .ZN(n4719) );
  NAND2_X1 U5479 ( .A1(n7473), .A2(n7472), .ZN(n7471) );
  NAND2_X1 U5480 ( .A1(n7360), .A2(n7433), .ZN(n5608) );
  OR2_X1 U5481 ( .A1(n8295), .A2(n5908), .ZN(n5909) );
  NAND2_X1 U5482 ( .A1(n8523), .A2(n7081), .ZN(n9684) );
  INV_X1 U5483 ( .A(n9684), .ZN(n9696) );
  NAND2_X1 U5484 ( .A1(n5921), .A2(n8505), .ZN(n9701) );
  NAND2_X1 U5485 ( .A1(n7331), .A2(n8525), .ZN(n9707) );
  INV_X1 U5486 ( .A(n9698), .ZN(n9686) );
  NAND2_X1 U5487 ( .A1(n5418), .A2(n5417), .ZN(n9493) );
  INV_X1 U5488 ( .A(n9701), .ZN(n9681) );
  OAI211_X1 U5489 ( .C1(P1_B_REG_SCAN_IN), .C2(n5471), .A(n5432), .B(n5473), 
        .ZN(n9867) );
  OAI21_X1 U5490 ( .B1(n6201), .B2(n10441), .A(n6200), .ZN(n6247) );
  OR2_X1 U5491 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  XNOR2_X1 U5492 ( .A(n6247), .B(n6246), .ZN(n8664) );
  XNOR2_X1 U5493 ( .A(n6201), .B(SI_29_), .ZN(n9215) );
  XNOR2_X1 U5494 ( .A(n5866), .B(n5865), .ZN(n8236) );
  NAND2_X1 U5495 ( .A1(n5863), .A2(n5862), .ZN(n5866) );
  XNOR2_X1 U5496 ( .A(n5849), .B(n5848), .ZN(n8231) );
  NAND2_X1 U5497 ( .A1(n4503), .A2(n5423), .ZN(n5427) );
  INV_X1 U5498 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5467) );
  OAI21_X1 U5499 ( .B1(n5758), .B2(n4656), .A(n5356), .ZN(n5773) );
  INV_X1 U5500 ( .A(n5757), .ZN(n4656) );
  AND2_X1 U5501 ( .A1(n5024), .A2(n5760), .ZN(n5023) );
  NAND2_X1 U5502 ( .A1(n4947), .A2(n4948), .ZN(n5508) );
  INV_X1 U5503 ( .A(n5337), .ZN(n4968) );
  NAND2_X1 U5504 ( .A1(n5656), .A2(n4970), .ZN(n4969) );
  NAND2_X1 U5505 ( .A1(n5656), .A2(n5334), .ZN(n5672) );
  OR2_X1 U5506 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  NAND2_X1 U5507 ( .A1(n5319), .A2(SI_6_), .ZN(n5322) );
  NAND2_X1 U5508 ( .A1(n4662), .A2(n10217), .ZN(n5324) );
  INV_X1 U5509 ( .A(n5323), .ZN(n4662) );
  NAND3_X1 U5510 ( .A1(n4902), .A2(n5519), .A3(n4903), .ZN(n5518) );
  NAND2_X1 U5511 ( .A1(n4989), .A2(n8993), .ZN(n4988) );
  INV_X1 U5512 ( .A(n8550), .ZN(n4989) );
  AND4_X1 U5513 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n9003)
         );
  INV_X1 U5514 ( .A(n8891), .ZN(n8640) );
  AND2_X1 U5515 ( .A1(n8125), .A2(n8211), .ZN(n8126) );
  INV_X1 U5516 ( .A(n8558), .ZN(n8978) );
  NAND4_X1 U5517 ( .A1(n6310), .A2(n6309), .A3(n6308), .A4(n6307), .ZN(n8776)
         );
  OR2_X1 U5518 ( .A1(n7245), .A2(n5249), .ZN(n8779) );
  NAND2_X1 U5519 ( .A1(n8823), .A2(n8824), .ZN(n8822) );
  INV_X1 U5520 ( .A(n8876), .ZN(n9994) );
  NOR2_X1 U5521 ( .A1(n8837), .A2(n5203), .ZN(n5207) );
  NAND2_X1 U5522 ( .A1(n5290), .A2(n4683), .ZN(n4682) );
  OR2_X1 U5523 ( .A1(n5255), .A2(n8858), .ZN(n5290) );
  INV_X1 U5524 ( .A(n4684), .ZN(n4683) );
  AND3_X1 U5525 ( .A1(n6282), .A2(n6281), .A3(n6280), .ZN(n10024) );
  INV_X1 U5526 ( .A(n10054), .ZN(n10047) );
  NAND2_X1 U5527 ( .A1(n6212), .A2(n6211), .ZN(n9070) );
  NAND2_X1 U5528 ( .A1(n9132), .A2(n10065), .ZN(n9078) );
  INV_X1 U5529 ( .A(n6825), .ZN(n9134) );
  AND3_X1 U5530 ( .A1(n6291), .A2(n6290), .A3(n6289), .ZN(n7958) );
  OR2_X1 U5531 ( .A1(n6558), .A2(n5293), .ZN(n6264) );
  AND2_X1 U5532 ( .A1(n6850), .A2(n6849), .ZN(n9207) );
  OR2_X1 U5533 ( .A1(n6851), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6850) );
  INV_X1 U5534 ( .A(n9614), .ZN(n9290) );
  NAND2_X1 U5535 ( .A1(n4894), .A2(n5628), .ZN(n7863) );
  NAND2_X1 U5536 ( .A1(n6950), .A2(n5867), .ZN(n4894) );
  AND4_X1 U5537 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n9242)
         );
  AND2_X1 U5538 ( .A1(n6054), .A2(n9349), .ZN(n6055) );
  NAND2_X1 U5539 ( .A1(n5751), .A2(n5750), .ZN(n9770) );
  INV_X1 U5540 ( .A(n9637), .ZN(n9756) );
  AND2_X1 U5541 ( .A1(n6101), .A2(n6100), .ZN(n9373) );
  INV_X1 U5542 ( .A(n9668), .ZN(n9766) );
  INV_X1 U5543 ( .A(n9386), .ZN(n9396) );
  INV_X1 U5544 ( .A(n9299), .ZN(n9407) );
  AOI21_X1 U5545 ( .B1(n8532), .B2(n4515), .A(n8540), .ZN(n4806) );
  INV_X1 U5546 ( .A(n8532), .ZN(n4807) );
  OAI21_X1 U5547 ( .B1(n9428), .B2(n6979), .A(n4681), .ZN(n9434) );
  NAND2_X1 U5548 ( .A1(n9428), .A2(n6979), .ZN(n4681) );
  NOR2_X1 U5549 ( .A1(n7056), .A2(n4671), .ZN(n7034) );
  AND2_X1 U5550 ( .A1(n7062), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4671) );
  INV_X1 U5551 ( .A(n5901), .ZN(n5457) );
  OR2_X1 U5552 ( .A1(n9866), .A2(n5457), .ZN(n9495) );
  INV_X1 U5553 ( .A(n9859), .ZN(n9492) );
  AND2_X1 U5554 ( .A1(n8284), .A2(n8283), .ZN(n8592) );
  AOI21_X1 U5555 ( .B1(n9498), .B2(n9909), .A(n4553), .ZN(n4608) );
  AND2_X1 U5556 ( .A1(n4955), .A2(n5813), .ZN(n9590) );
  NAND2_X1 U5557 ( .A1(n8013), .A2(n5867), .ZN(n4955) );
  INV_X1 U5558 ( .A(n4721), .ZN(n4720) );
  OAI21_X1 U5559 ( .B1(n5574), .B2(n6932), .A(n5572), .ZN(n4721) );
  NAND2_X1 U5560 ( .A1(n5585), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5561 ( .A1(n5409), .A2(n5625), .ZN(n5410) );
  NAND2_X1 U5562 ( .A1(n6608), .A2(n6609), .ZN(n6612) );
  INV_X1 U5563 ( .A(n5907), .ZN(n4802) );
  NAND2_X1 U5564 ( .A1(n4689), .A2(n4687), .ZN(n6654) );
  NAND2_X1 U5565 ( .A1(n6646), .A2(n6837), .ZN(n4689) );
  NAND2_X1 U5566 ( .A1(n6657), .A2(n6881), .ZN(n4687) );
  AND2_X1 U5567 ( .A1(n8307), .A2(n4976), .ZN(n4844) );
  AND2_X1 U5568 ( .A1(n6674), .A2(n6881), .ZN(n4694) );
  INV_X1 U5569 ( .A(n8320), .ZN(n4839) );
  NAND2_X1 U5570 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  AOI21_X1 U5571 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6705) );
  AOI22_X1 U5572 ( .A1(n8344), .A2(n4976), .B1(n8346), .B2(n8345), .ZN(n4846)
         );
  NAND2_X1 U5573 ( .A1(n4848), .A2(n8398), .ZN(n4847) );
  AOI21_X1 U5574 ( .B1(n8367), .B2(n4835), .A(n4832), .ZN(n4831) );
  INV_X1 U5575 ( .A(n5745), .ZN(n4941) );
  NOR2_X1 U5576 ( .A1(n6728), .A2(n5064), .ZN(n4701) );
  NOR2_X1 U5577 ( .A1(n8609), .A2(n6738), .ZN(n4699) );
  NAND2_X1 U5578 ( .A1(n6739), .A2(n4775), .ZN(n4700) );
  NAND2_X1 U5579 ( .A1(n5103), .A2(n5006), .ZN(n5005) );
  NOR2_X1 U5580 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5006) );
  OR2_X1 U5581 ( .A1(n8379), .A2(n8377), .ZN(n4833) );
  AOI21_X1 U5582 ( .B1(n4827), .B2(n4825), .A(n4824), .ZN(n4823) );
  INV_X1 U5583 ( .A(n8375), .ZN(n4824) );
  INV_X1 U5584 ( .A(n4828), .ZN(n4825) );
  NAND2_X1 U5585 ( .A1(n5944), .A2(n8525), .ZN(n5950) );
  NOR2_X1 U5586 ( .A1(n9756), .A2(n9761), .ZN(n4882) );
  NOR2_X1 U5587 ( .A1(n9783), .A2(n8147), .ZN(n4887) );
  NOR2_X1 U5588 ( .A1(n7608), .A2(n7613), .ZN(n7609) );
  INV_X1 U5589 ( .A(n5792), .ZN(n5363) );
  NAND2_X1 U5590 ( .A1(n5350), .A2(n10411), .ZN(n5353) );
  AND2_X1 U5591 ( .A1(n5340), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U5592 ( .A1(n5343), .A2(n5342), .ZN(n5346) );
  NAND3_X1 U5593 ( .A1(n4712), .A2(n4711), .A3(n4710), .ZN(n5291) );
  INV_X1 U5594 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5595 ( .A1(n7292), .A2(n7291), .ZN(n7295) );
  NOR2_X1 U5596 ( .A1(n6829), .A2(n8905), .ZN(n6748) );
  INV_X1 U5597 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10204) );
  INV_X1 U5598 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U5599 ( .A1(n6216), .A2(n6215), .ZN(n6360) );
  INV_X1 U5600 ( .A(n6347), .ZN(n6216) );
  NAND2_X1 U5601 ( .A1(n10008), .A2(n4756), .ZN(n6650) );
  NAND2_X1 U5602 ( .A1(n8778), .A2(n7958), .ZN(n6632) );
  AND2_X1 U5603 ( .A1(n7805), .A2(n8869), .ZN(n7293) );
  OR2_X1 U5604 ( .A1(n6851), .A2(n6863), .ZN(n6882) );
  INV_X1 U5605 ( .A(n6823), .ZN(n4766) );
  INV_X1 U5606 ( .A(n4768), .ZN(n4765) );
  NOR2_X1 U5607 ( .A1(n4522), .A2(n4775), .ZN(n4774) );
  NOR2_X1 U5608 ( .A1(n6818), .A2(n8769), .ZN(n4770) );
  AND2_X1 U5609 ( .A1(n9155), .A2(n8957), .ZN(n6730) );
  OR2_X1 U5610 ( .A1(n6813), .A2(n8993), .ZN(n6708) );
  INV_X1 U5611 ( .A(n6676), .ZN(n4740) );
  AND2_X1 U5612 ( .A1(n6865), .A2(n7805), .ZN(n7463) );
  INV_X1 U5613 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5089) );
  INV_X1 U5614 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5088) );
  OR2_X1 U5615 ( .A1(n6071), .A2(n8142), .ZN(n6085) );
  AND2_X1 U5616 ( .A1(n5948), .A2(n5950), .ZN(n5949) );
  AOI21_X1 U5617 ( .B1(n5012), .B2(n5010), .A(n4569), .ZN(n5009) );
  INV_X1 U5618 ( .A(n6089), .ZN(n4615) );
  INV_X1 U5619 ( .A(n4617), .ZN(n4613) );
  AND2_X1 U5620 ( .A1(n8520), .A2(n8435), .ZN(n8522) );
  NOR2_X1 U5621 ( .A1(n9536), .A2(n4653), .ZN(n8431) );
  OR2_X1 U5622 ( .A1(n9529), .A2(n6150), .ZN(n8513) );
  NAND2_X1 U5623 ( .A1(n9628), .A2(n9627), .ZN(n4929) );
  AOI21_X1 U5624 ( .B1(n5055), .B2(n5052), .A(n5756), .ZN(n5051) );
  NAND2_X1 U5625 ( .A1(n4706), .A2(n4704), .ZN(n4703) );
  NOR2_X1 U5626 ( .A1(n5058), .A2(n5046), .ZN(n4704) );
  INV_X1 U5627 ( .A(n7895), .ZN(n4607) );
  INV_X1 U5628 ( .A(n8426), .ZN(n4915) );
  INV_X1 U5629 ( .A(n4919), .ZN(n4916) );
  INV_X1 U5630 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5709) );
  INV_X1 U5631 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5677) );
  OR2_X1 U5632 ( .A1(n5664), .A2(n7123), .ZN(n5678) );
  INV_X1 U5633 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5617) );
  INV_X1 U5634 ( .A(n5950), .ZN(n7345) );
  NAND2_X1 U5635 ( .A1(n9664), .A2(n4882), .ZN(n9631) );
  NAND2_X1 U5636 ( .A1(n9664), .A2(n9653), .ZN(n9646) );
  NAND2_X1 U5637 ( .A1(n7817), .A2(n8024), .ZN(n8005) );
  NAND2_X1 U5638 ( .A1(n4874), .A2(n7443), .ZN(n7275) );
  NAND2_X1 U5639 ( .A1(n5396), .A2(n5395), .ZN(n6199) );
  NOR2_X1 U5640 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5400) );
  NAND2_X1 U5641 ( .A1(n5463), .A2(n5419), .ZN(n5458) );
  INV_X1 U5642 ( .A(n5772), .ZN(n4963) );
  INV_X1 U5643 ( .A(n4945), .ZN(n4944) );
  AOI21_X1 U5644 ( .B1(n4943), .B2(n4945), .A(n4550), .ZN(n4942) );
  INV_X1 U5645 ( .A(n4949), .ZN(n4943) );
  NAND2_X1 U5646 ( .A1(n5347), .A2(n5729), .ZN(n4948) );
  OR2_X1 U5647 ( .A1(n5347), .A2(n5729), .ZN(n4949) );
  INV_X1 U5648 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U5649 ( .A1(n4600), .A2(n5702), .ZN(n5341) );
  NAND2_X1 U5650 ( .A1(n4597), .A2(n4596), .ZN(n4600) );
  NOR2_X1 U5651 ( .A1(n4965), .A2(SI_13_), .ZN(n4596) );
  NAND2_X1 U5652 ( .A1(n5522), .A2(n5399), .ZN(n5613) );
  INV_X1 U5653 ( .A(n8668), .ZN(n8641) );
  INV_X1 U5654 ( .A(n9058), .ZN(n8544) );
  AND2_X1 U5655 ( .A1(n8700), .A2(n8571), .ZN(n8574) );
  INV_X1 U5656 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U5657 ( .A1(n8552), .A2(n8551), .ZN(n8686) );
  AND2_X1 U5658 ( .A1(n8120), .A2(n8772), .ZN(n5001) );
  INV_X1 U5659 ( .A(n4992), .ZN(n4991) );
  OAI21_X1 U5660 ( .B1(n4993), .B2(n4995), .A(n8739), .ZN(n4992) );
  NAND2_X1 U5661 ( .A1(n8751), .A2(n8752), .ZN(n4985) );
  AND2_X1 U5662 ( .A1(n8751), .A2(n4986), .ZN(n4984) );
  XNOR2_X1 U5663 ( .A(n6835), .B(n6834), .ZN(n7288) );
  OR2_X1 U5664 ( .A1(n6524), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6535) );
  INV_X1 U5665 ( .A(n8014), .ZN(n4730) );
  OR2_X1 U5666 ( .A1(n7157), .A2(n7156), .ZN(n7159) );
  NAND2_X1 U5667 ( .A1(n7159), .A2(n5156), .ZN(n9932) );
  OAI21_X1 U5668 ( .B1(n9949), .B2(n4856), .A(n4854), .ZN(n6905) );
  INV_X1 U5669 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5670 ( .A(n6902), .ZN(n4856) );
  NAND2_X1 U5671 ( .A1(n9949), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9948) );
  AND2_X1 U5672 ( .A1(n5171), .A2(n7503), .ZN(n6920) );
  OR2_X1 U5673 ( .A1(n5170), .A2(n6945), .ZN(n5171) );
  NAND2_X1 U5674 ( .A1(n6920), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7505) );
  OR2_X1 U5675 ( .A1(n7590), .A2(n5084), .ZN(n4853) );
  OR2_X1 U5676 ( .A1(n7773), .A2(n5183), .ZN(n4872) );
  NAND2_X1 U5677 ( .A1(n7779), .A2(n5272), .ZN(n7832) );
  XNOR2_X1 U5678 ( .A(n5185), .B(n6367), .ZN(n7930) );
  AND2_X1 U5679 ( .A1(n4870), .A2(n4869), .ZN(n5185) );
  NAND2_X1 U5680 ( .A1(n7835), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5681 ( .A1(n7925), .A2(n5275), .ZN(n8044) );
  NAND2_X1 U5682 ( .A1(n9965), .A2(n5277), .ZN(n9987) );
  NAND2_X1 U5683 ( .A1(n4865), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4864) );
  NAND2_X1 U5684 ( .A1(n5188), .A2(n4865), .ZN(n4863) );
  INV_X1 U5685 ( .A(n9997), .ZN(n4865) );
  XNOR2_X1 U5686 ( .A(n5280), .B(n5201), .ZN(n8849) );
  NAND2_X1 U5687 ( .A1(n8822), .A2(n4669), .ZN(n5280) );
  OR2_X1 U5688 ( .A1(n6421), .A2(n9114), .ZN(n4669) );
  INV_X1 U5689 ( .A(n5209), .ZN(n6834) );
  AND2_X1 U5690 ( .A1(n6519), .A2(n6735), .ZN(n6520) );
  NAND2_X1 U5691 ( .A1(n6227), .A2(n10231), .ZN(n6524) );
  INV_X1 U5692 ( .A(n6476), .ZN(n6227) );
  OR2_X1 U5693 ( .A1(n6496), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U5694 ( .A1(n6225), .A2(n6224), .ZN(n6494) );
  INV_X1 U5695 ( .A(n6505), .ZN(n6225) );
  OR2_X1 U5696 ( .A1(n6494), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6496) );
  OR2_X1 U5697 ( .A1(n6503), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U5698 ( .A1(n6223), .A2(n10204), .ZN(n6503) );
  INV_X1 U5699 ( .A(n6454), .ZN(n6223) );
  AND4_X1 U5700 ( .A1(n6440), .A2(n6439), .A3(n6438), .A4(n6437), .ZN(n9005)
         );
  NAND2_X1 U5701 ( .A1(n4738), .A2(n4737), .ZN(n9009) );
  AND2_X1 U5702 ( .A1(n9010), .A2(n6693), .ZN(n4737) );
  AND2_X1 U5703 ( .A1(n6708), .A2(n6692), .ZN(n9010) );
  NAND2_X1 U5704 ( .A1(n6222), .A2(n6221), .ZN(n6443) );
  INV_X1 U5705 ( .A(n6434), .ZN(n6222) );
  NAND2_X1 U5706 ( .A1(n6220), .A2(n10459), .ZN(n6424) );
  INV_X1 U5707 ( .A(n6413), .ZN(n6220) );
  OR2_X1 U5708 ( .A1(n6424), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6434) );
  OR2_X1 U5709 ( .A1(n6403), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U5710 ( .A1(n6219), .A2(n6218), .ZN(n6403) );
  INV_X1 U5711 ( .A(n6391), .ZN(n6219) );
  NAND2_X1 U5712 ( .A1(n6217), .A2(n10460), .ZN(n6391) );
  INV_X1 U5713 ( .A(n6381), .ZN(n6217) );
  OR2_X1 U5714 ( .A1(n6360), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6371) );
  AOI21_X1 U5715 ( .B1(n4760), .B2(n4762), .A(n4532), .ZN(n4758) );
  INV_X1 U5716 ( .A(n7982), .ZN(n8162) );
  AOI21_X1 U5717 ( .B1(n4750), .B2(n4749), .A(n4748), .ZN(n4747) );
  INV_X1 U5718 ( .A(n6656), .ZN(n4748) );
  INV_X1 U5719 ( .A(n6658), .ZN(n4749) );
  NAND2_X1 U5720 ( .A1(n4759), .A2(n6795), .ZN(n8086) );
  NAND2_X1 U5721 ( .A1(n8098), .A2(n6794), .ZN(n4759) );
  NAND2_X1 U5722 ( .A1(n4753), .A2(n6651), .ZN(n8097) );
  NAND2_X1 U5723 ( .A1(n7963), .A2(n6658), .ZN(n4753) );
  OR2_X1 U5724 ( .A1(n6337), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U5725 ( .A1(n7948), .A2(n8774), .ZN(n7962) );
  NAND2_X1 U5726 ( .A1(n4755), .A2(n6788), .ZN(n7965) );
  INV_X1 U5727 ( .A(n7882), .ZN(n4755) );
  AND2_X1 U5728 ( .A1(n7880), .A2(n6788), .ZN(n6786) );
  AND2_X1 U5729 ( .A1(n7885), .A2(n6789), .ZN(n7882) );
  NAND2_X1 U5730 ( .A1(n6650), .A2(n7962), .ZN(n7885) );
  NOR2_X1 U5731 ( .A1(n6633), .A2(n4746), .ZN(n4745) );
  INV_X1 U5732 ( .A(n6635), .ZN(n4746) );
  OR2_X1 U5733 ( .A1(n8778), .A2(n7958), .ZN(n7629) );
  AND2_X1 U5734 ( .A1(n7692), .A2(n6783), .ZN(n7636) );
  INV_X1 U5735 ( .A(n6779), .ZN(n7618) );
  OR3_X1 U5736 ( .A1(n7450), .A2(n7449), .A3(n7448), .ZN(n7455) );
  AND2_X1 U5737 ( .A1(n10040), .A2(n6604), .ZN(n7257) );
  AND2_X1 U5738 ( .A1(n6543), .A2(n6572), .ZN(n4735) );
  AND2_X1 U5739 ( .A1(n4769), .A2(n4773), .ZN(n4768) );
  OR2_X1 U5740 ( .A1(n4522), .A2(n4776), .ZN(n4773) );
  NAND2_X1 U5741 ( .A1(n4774), .A2(n4770), .ZN(n4769) );
  AND2_X1 U5742 ( .A1(n6821), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U5743 ( .A1(n4774), .A2(n4772), .ZN(n4771) );
  INV_X1 U5744 ( .A(n6819), .ZN(n4772) );
  NAND2_X1 U5745 ( .A1(n6475), .A2(n6474), .ZN(n8618) );
  AND2_X1 U5746 ( .A1(n8928), .A2(n8927), .ZN(n8944) );
  AND4_X1 U5747 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n8603)
         );
  AND2_X1 U5748 ( .A1(n6721), .A2(n6722), .ZN(n8955) );
  OR2_X1 U5749 ( .A1(n8981), .A2(n8950), .ZN(n8964) );
  NAND2_X1 U5750 ( .A1(n6502), .A2(n6501), .ZN(n8727) );
  AND2_X1 U5751 ( .A1(n6683), .A2(n6684), .ZN(n9053) );
  AND2_X1 U5752 ( .A1(n7262), .A2(n9063), .ZN(n7242) );
  INV_X1 U5753 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6235) );
  AND2_X1 U5754 ( .A1(n5105), .A2(n4511), .ZN(n6847) );
  INV_X1 U5755 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5002) );
  INV_X1 U5756 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5098) );
  INV_X1 U5757 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5177) );
  NOR2_X1 U5758 ( .A1(n5167), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5172) );
  INV_X1 U5759 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U5760 ( .A1(n8053), .A2(n6074), .ZN(n9233) );
  NAND2_X1 U5761 ( .A1(n8053), .A2(n4617), .ZN(n4611) );
  NAND2_X1 U5762 ( .A1(n5029), .A2(n4544), .ZN(n5030) );
  NAND2_X1 U5763 ( .A1(n4634), .A2(n5009), .ZN(n9271) );
  NAND2_X1 U5764 ( .A1(n7870), .A2(n6042), .ZN(n9259) );
  NAND2_X1 U5765 ( .A1(n7869), .A2(n7871), .ZN(n7870) );
  NOR2_X1 U5766 ( .A1(n5777), .A2(n8272), .ZN(n5786) );
  AND2_X1 U5767 ( .A1(n5786), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U5768 ( .A1(n5019), .A2(n5020), .ZN(n6121) );
  AOI21_X1 U5769 ( .B1(n5021), .B2(n9327), .A(n4579), .ZN(n5020) );
  NAND2_X1 U5770 ( .A1(n5981), .A2(n7183), .ZN(n9363) );
  AND2_X1 U5771 ( .A1(n8592), .A2(n9410), .ZN(n8402) );
  OAI21_X1 U5772 ( .B1(n8388), .B2(n4819), .A(n4810), .ZN(n8396) );
  NOR2_X1 U5773 ( .A1(n4974), .A2(n8592), .ZN(n4973) );
  OAI21_X1 U5774 ( .B1(n9483), .B2(n4976), .A(n4975), .ZN(n4974) );
  OAI21_X1 U5775 ( .B1(n8388), .B2(n4814), .A(n4812), .ZN(n8399) );
  NAND2_X1 U5776 ( .A1(n4815), .A2(n9790), .ZN(n4814) );
  INV_X1 U5777 ( .A(n4819), .ZN(n4815) );
  NOR2_X1 U5778 ( .A1(n7033), .A2(n4567), .ZN(n7058) );
  NOR2_X1 U5779 ( .A1(n7058), .A2(n7057), .ZN(n7056) );
  NOR2_X1 U5780 ( .A1(n7221), .A2(n7220), .ZN(n7374) );
  NOR2_X1 U5781 ( .A1(n4680), .A2(n7848), .ZN(n4679) );
  NOR2_X1 U5782 ( .A1(n7915), .A2(n7914), .ZN(n8075) );
  NAND2_X1 U5783 ( .A1(n8252), .A2(n4664), .ZN(n9474) );
  NAND2_X1 U5784 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  INV_X1 U5785 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5786 ( .A1(n9577), .A2(n4513), .ZN(n9503) );
  AND4_X1 U5787 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5889), .ZN(n9520)
         );
  NAND2_X1 U5788 ( .A1(n9577), .A2(n4876), .ZN(n9527) );
  INV_X1 U5789 ( .A(n9557), .ZN(n5847) );
  NAND2_X1 U5790 ( .A1(n9577), .A2(n9800), .ZN(n9559) );
  NOR2_X1 U5791 ( .A1(n8373), .A2(n5037), .ZN(n5036) );
  INV_X1 U5792 ( .A(n5040), .ZN(n5037) );
  NOR2_X1 U5793 ( .A1(n5821), .A2(n5042), .ZN(n5039) );
  OR2_X1 U5794 ( .A1(n9256), .A2(n4954), .ZN(n5040) );
  NAND2_X1 U5795 ( .A1(n9601), .A2(n8369), .ZN(n8243) );
  NAND2_X1 U5796 ( .A1(n8243), .A2(n8430), .ZN(n9571) );
  NAND2_X1 U5797 ( .A1(n9664), .A2(n4537), .ZN(n9596) );
  NAND2_X1 U5798 ( .A1(n4929), .A2(n4927), .ZN(n9610) );
  AND2_X1 U5799 ( .A1(n8359), .A2(n8360), .ZN(n9627) );
  NAND2_X1 U5800 ( .A1(n5738), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U5801 ( .A1(n4605), .A2(n8339), .ZN(n9695) );
  NAND2_X1 U5802 ( .A1(n4914), .A2(n4606), .ZN(n4605) );
  AOI21_X1 U5803 ( .B1(n4917), .B2(n4916), .A(n4915), .ZN(n4914) );
  NAND2_X1 U5804 ( .A1(n4607), .A2(n4917), .ZN(n4606) );
  NAND2_X1 U5805 ( .A1(n7817), .A2(n4514), .ZN(n9705) );
  NAND2_X1 U5806 ( .A1(n7817), .A2(n4885), .ZN(n9708) );
  OR2_X1 U5807 ( .A1(n5710), .A2(n5709), .ZN(n5722) );
  NOR2_X1 U5808 ( .A1(n5722), .A2(n7729), .ZN(n5736) );
  NAND2_X1 U5809 ( .A1(n4909), .A2(n4908), .ZN(n7808) );
  OR2_X1 U5810 ( .A1(n4911), .A2(n5916), .ZN(n4908) );
  NOR2_X1 U5811 ( .A1(n7657), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U5812 ( .A1(n7599), .A2(n8322), .ZN(n7658) );
  AOI21_X1 U5813 ( .B1(n4716), .B2(n4719), .A(n4548), .ZN(n4715) );
  AND4_X1 U5814 ( .A1(n5682), .A2(n5681), .A3(n5680), .A4(n5679), .ZN(n7809)
         );
  NAND2_X1 U5815 ( .A1(n7600), .A2(n7601), .ZN(n7599) );
  NAND2_X1 U5816 ( .A1(n7577), .A2(n7489), .ZN(n7491) );
  OR2_X1 U5817 ( .A1(n7491), .A2(n7863), .ZN(n7474) );
  NOR2_X1 U5818 ( .A1(n7275), .A2(n7283), .ZN(n7367) );
  AND2_X1 U5819 ( .A1(n7367), .A2(n9882), .ZN(n7489) );
  AND4_X1 U5820 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n7858)
         );
  NAND2_X1 U5821 ( .A1(n7365), .A2(n8412), .ZN(n7364) );
  NAND2_X1 U5822 ( .A1(n7279), .A2(n7443), .ZN(n5591) );
  NAND2_X1 U5823 ( .A1(n7232), .A2(n8460), .ZN(n8293) );
  NAND2_X1 U5824 ( .A1(n5984), .A2(n5559), .ZN(n5561) );
  NAND2_X1 U5825 ( .A1(n4790), .A2(n5905), .ZN(n7340) );
  XNOR2_X1 U5826 ( .A(n5545), .B(n8454), .ZN(n7107) );
  NOR2_X1 U5827 ( .A1(n7185), .A2(n7108), .ZN(n7351) );
  OR2_X1 U5828 ( .A1(n9867), .A2(n5445), .ZN(n7324) );
  AND2_X1 U5829 ( .A1(n9410), .A2(n8582), .ZN(n9715) );
  INV_X1 U5830 ( .A(n9909), .ZN(n9786) );
  AND2_X1 U5831 ( .A1(n5470), .A2(n5469), .ZN(n7326) );
  INV_X1 U5832 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5494) );
  NOR2_X1 U5833 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5407) );
  NOR2_X1 U5834 ( .A1(n4873), .A2(n5489), .ZN(n5492) );
  XNOR2_X1 U5835 ( .A(n4935), .B(n5882), .ZN(n8593) );
  INV_X1 U5836 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U5837 ( .A1(n5421), .A2(n5420), .ZN(n5428) );
  AND3_X1 U5838 ( .A1(n5460), .A2(n5476), .A3(n5467), .ZN(n5420) );
  INV_X1 U5839 ( .A(n5458), .ZN(n5421) );
  XNOR2_X1 U5840 ( .A(n5477), .B(n5476), .ZN(n8011) );
  OAI21_X1 U5841 ( .B1(n5484), .B2(n5483), .A(n5367), .ZN(n5810) );
  AND2_X1 U5842 ( .A1(n5372), .A2(n5371), .ZN(n5809) );
  INV_X1 U5843 ( .A(SI_19_), .ZN(n5357) );
  INV_X1 U5844 ( .A(n8525), .ZN(n8503) );
  AND2_X1 U5845 ( .A1(n5705), .A2(n5692), .ZN(n7381) );
  NAND2_X1 U5846 ( .A1(n4645), .A2(n4541), .ZN(n5654) );
  NAND2_X1 U5847 ( .A1(n5518), .A2(n4535), .ZN(n4645) );
  AND2_X1 U5848 ( .A1(n5661), .A2(n5688), .ZN(n7219) );
  OAI21_X1 U5849 ( .B1(n5638), .B2(n5637), .A(n5636), .ZN(n5640) );
  INV_X1 U5850 ( .A(n5613), .ZN(n5524) );
  NAND2_X1 U5851 ( .A1(n4610), .A2(n4609), .ZN(n5586) );
  INV_X1 U5852 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4609) );
  OR2_X1 U5853 ( .A1(n4891), .A2(SI_1_), .ZN(n4890) );
  AND4_X1 U5854 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n8175)
         );
  INV_X1 U5855 ( .A(n7397), .ZN(n7398) );
  AND2_X1 U5856 ( .A1(n6566), .A2(n6565), .ZN(n8767) );
  CLKBUF_X1 U5857 ( .A(n7314), .Z(n7315) );
  AND4_X1 U5858 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n8992)
         );
  AND3_X1 U5859 ( .A1(n6465), .A2(n6464), .A3(n6463), .ZN(n8921) );
  AND3_X1 U5860 ( .A1(n4987), .A2(n8545), .A3(n4986), .ZN(n8753) );
  NAND2_X1 U5861 ( .A1(n4987), .A2(n8545), .ZN(n8718) );
  OR2_X1 U5862 ( .A1(n7986), .A2(n8210), .ZN(n4997) );
  OR2_X1 U5863 ( .A1(n8191), .A2(n5001), .ZN(n5000) );
  AND2_X1 U5864 ( .A1(n7266), .A2(n7265), .ZN(n8725) );
  AND2_X1 U5865 ( .A1(n6442), .A2(n6441), .ZN(n8765) );
  NAND2_X1 U5866 ( .A1(n7259), .A2(n9061), .ZN(n8723) );
  INV_X1 U5867 ( .A(n8747), .ZN(n8758) );
  NAND2_X1 U5868 ( .A1(n7390), .A2(n8014), .ZN(n8747) );
  AOI21_X1 U5869 ( .B1(n6599), .B2(n4728), .A(n4594), .ZN(n4726) );
  AOI21_X1 U5870 ( .B1(n6764), .B2(n6881), .A(n6596), .ZN(n6767) );
  AND3_X1 U5871 ( .A1(n6758), .A2(n6757), .A3(n4529), .ZN(n6764) );
  NAND2_X1 U5872 ( .A1(n4520), .A2(n7805), .ZN(n4723) );
  INV_X1 U5873 ( .A(n8603), .ZN(n8969) );
  NAND4_X1 U5874 ( .A1(n6321), .A2(n6320), .A3(n6319), .A4(n6318), .ZN(n8775)
         );
  NAND2_X1 U5875 ( .A1(n6550), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6279) );
  OR2_X1 U5876 ( .A1(n6436), .A2(n7156), .ZN(n6260) );
  NAND2_X1 U5877 ( .A1(n6267), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6269) );
  OR2_X1 U5878 ( .A1(P2_U3150), .A2(n5286), .ZN(n9982) );
  INV_X1 U5879 ( .A(n4870), .ZN(n7823) );
  INV_X1 U5880 ( .A(n4872), .ZN(n7825) );
  MUX2_X1 U5881 ( .A(n5253), .B(n8779), .S(n6835), .Z(n9983) );
  NOR2_X1 U5882 ( .A1(n9972), .A2(n6393), .ZN(n9975) );
  INV_X1 U5883 ( .A(n4861), .ZN(n8804) );
  NAND2_X1 U5884 ( .A1(n8814), .A2(n5279), .ZN(n8823) );
  NAND2_X1 U5885 ( .A1(n4862), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U5886 ( .A1(n5190), .A2(n4862), .ZN(n4858) );
  INV_X1 U5887 ( .A(n8821), .ZN(n4862) );
  INV_X1 U5888 ( .A(n5190), .ZN(n4860) );
  NOR2_X1 U5889 ( .A1(n8838), .A2(n9019), .ZN(n8837) );
  AND2_X1 U5890 ( .A1(n7143), .A2(n6834), .ZN(n9974) );
  NAND2_X1 U5891 ( .A1(n6560), .A2(n6559), .ZN(n8659) );
  NAND2_X1 U5892 ( .A1(n8919), .A2(n8933), .ZN(n4778) );
  NAND2_X1 U5893 ( .A1(n6467), .A2(n6466), .ZN(n8681) );
  NAND2_X1 U5894 ( .A1(n4787), .A2(n4785), .ZN(n8976) );
  NAND2_X1 U5895 ( .A1(n6430), .A2(n6696), .ZN(n9022) );
  NAND2_X1 U5896 ( .A1(n6432), .A2(n6431), .ZN(n9110) );
  NAND2_X1 U5897 ( .A1(n4686), .A2(n6950), .ZN(n6345) );
  NAND2_X1 U5898 ( .A1(n7632), .A2(n6635), .ZN(n7691) );
  INV_X1 U5899 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7560) );
  OR2_X1 U5900 ( .A1(n10054), .A2(n6868), .ZN(n9063) );
  NAND2_X1 U5901 ( .A1(n7258), .A2(n7257), .ZN(n9061) );
  INV_X1 U5902 ( .A(n9061), .ZN(n10019) );
  NAND2_X1 U5903 ( .A1(n6249), .A2(n6248), .ZN(n9128) );
  NAND2_X1 U5904 ( .A1(n8661), .A2(n10040), .ZN(n6843) );
  AOI21_X1 U5905 ( .B1(n8895), .B2(n9060), .A(n8894), .ZN(n9132) );
  NAND2_X1 U5906 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U5907 ( .A1(n8891), .A2(n9055), .ZN(n8892) );
  NAND2_X1 U5908 ( .A1(n6534), .A2(n6533), .ZN(n9140) );
  OR2_X1 U5909 ( .A1(n6558), .A2(n6532), .ZN(n6533) );
  NAND2_X1 U5910 ( .A1(n4736), .A2(n6572), .ZN(n8900) );
  AND2_X1 U5911 ( .A1(n6523), .A2(n6522), .ZN(n8914) );
  AND2_X1 U5912 ( .A1(n6461), .A2(n6460), .ZN(n9150) );
  INV_X1 U5913 ( .A(n8681), .ZN(n9155) );
  NAND2_X1 U5914 ( .A1(n6493), .A2(n6492), .ZN(n9161) );
  NAND2_X1 U5915 ( .A1(n6485), .A2(n6484), .ZN(n9167) );
  INV_X1 U5916 ( .A(n8727), .ZN(n9175) );
  NAND2_X1 U5917 ( .A1(n6453), .A2(n6452), .ZN(n9178) );
  INV_X1 U5918 ( .A(n8765), .ZN(n6813) );
  NAND2_X1 U5919 ( .A1(n6423), .A2(n6422), .ZN(n9188) );
  NAND2_X1 U5920 ( .A1(n6412), .A2(n6411), .ZN(n9194) );
  NAND2_X1 U5921 ( .A1(n4744), .A2(n6684), .ZN(n9035) );
  NAND2_X1 U5922 ( .A1(n6402), .A2(n6401), .ZN(n9201) );
  NAND2_X1 U5923 ( .A1(n6390), .A2(n6389), .ZN(n8227) );
  INV_X1 U5924 ( .A(n9174), .ZN(n9200) );
  NAND2_X1 U5925 ( .A1(n4780), .A2(n6799), .ZN(n8208) );
  NAND2_X1 U5926 ( .A1(n4741), .A2(n6676), .ZN(n8205) );
  AND3_X1 U5927 ( .A1(n10051), .A2(n10050), .A3(n10049), .ZN(n10067) );
  INV_X1 U5928 ( .A(n8030), .ZN(n7973) );
  INV_X1 U5929 ( .A(n6578), .ZN(n7939) );
  AND2_X1 U5930 ( .A1(n6772), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7254) );
  INV_X1 U5931 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9209) );
  INV_X1 U5932 ( .A(n6847), .ZN(n8233) );
  INV_X1 U5933 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U5934 ( .A1(n5108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  OR2_X1 U5935 ( .A1(n5107), .A2(n5106), .ZN(n5109) );
  INV_X1 U5936 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8016) );
  INV_X1 U5937 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7999) );
  INV_X1 U5938 ( .A(n6831), .ZN(n7998) );
  INV_X1 U5939 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7651) );
  INV_X1 U5940 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7565) );
  INV_X1 U5941 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7413) );
  INV_X1 U5942 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7287) );
  INV_X1 U5943 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7178) );
  INV_X1 U5944 ( .A(n6356), .ZN(n7835) );
  INV_X1 U5945 ( .A(n8795), .ZN(n6952) );
  OAI21_X1 U5946 ( .B1(n5149), .B2(n5148), .A(n5147), .ZN(n5150) );
  NOR2_X1 U5947 ( .A1(n5259), .A2(n6233), .ZN(n5149) );
  AND2_X1 U5948 ( .A1(n8011), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6890) );
  AND4_X1 U5949 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n7571)
         );
  AND4_X1 U5950 ( .A1(n5651), .A2(n5650), .A3(n5649), .A4(n5648), .ZN(n9265)
         );
  OR2_X1 U5951 ( .A1(n6173), .A2(n9402), .ZN(n5068) );
  INV_X1 U5952 ( .A(n5018), .ZN(n5017) );
  AOI21_X1 U5953 ( .B1(n6117), .B2(n6116), .A(n9327), .ZN(n9288) );
  NAND2_X1 U5954 ( .A1(n9271), .A2(n6104), .ZN(n6117) );
  NAND2_X1 U5955 ( .A1(n5796), .A2(n5795), .ZN(n9618) );
  NAND2_X1 U5956 ( .A1(n4622), .A2(n4627), .ZN(n9295) );
  NAND2_X1 U5957 ( .A1(n9249), .A2(n9317), .ZN(n4622) );
  NAND2_X1 U5958 ( .A1(n4619), .A2(n4507), .ZN(n9381) );
  INV_X1 U5959 ( .A(n5010), .ZN(n5007) );
  OR2_X1 U5960 ( .A1(n5011), .A2(n9404), .ZN(n5008) );
  NAND2_X1 U5961 ( .A1(n4636), .A2(n5014), .ZN(n5011) );
  NAND2_X1 U5962 ( .A1(n5825), .A2(n5824), .ZN(n9741) );
  OR2_X1 U5963 ( .A1(n9249), .A2(n9318), .ZN(n4626) );
  AND4_X1 U5964 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n7873)
         );
  INV_X1 U5965 ( .A(n5545), .ZN(n7190) );
  NAND2_X1 U5966 ( .A1(n8053), .A2(n8054), .ZN(n8140) );
  INV_X1 U5967 ( .A(n5032), .ZN(n5031) );
  AND2_X1 U5968 ( .A1(n6181), .A2(n5922), .ZN(n9391) );
  NAND2_X1 U5969 ( .A1(n5851), .A2(n5850), .ZN(n9730) );
  NAND2_X1 U5970 ( .A1(n9434), .A2(n9433), .ZN(n9432) );
  INV_X1 U5971 ( .A(n4674), .ZN(n6990) );
  NAND2_X1 U5972 ( .A1(n7034), .A2(n7035), .ZN(n7116) );
  NOR2_X1 U5973 ( .A1(n4670), .A2(n7374), .ZN(n9838) );
  AND2_X1 U5974 ( .A1(n7375), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4670) );
  NAND2_X1 U5975 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
  NOR2_X1 U5976 ( .A1(n8075), .A2(n4667), .ZN(n8079) );
  AND2_X1 U5977 ( .A1(n8076), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U5978 ( .A1(n8079), .A2(n8078), .ZN(n8252) );
  INV_X1 U5979 ( .A(n9849), .ZN(n9471) );
  NOR2_X1 U5980 ( .A1(n8580), .A2(n9707), .ZN(n8588) );
  NAND2_X1 U5981 ( .A1(n9510), .A2(n9701), .ZN(n9513) );
  AND2_X1 U5982 ( .A1(n5043), .A2(n4527), .ZN(n9502) );
  OR2_X1 U5983 ( .A1(n9556), .A2(n9555), .ZN(n9734) );
  NAND2_X1 U5984 ( .A1(n5808), .A2(n5041), .ZN(n8241) );
  OAI21_X1 U5985 ( .B1(n9628), .B2(n4928), .A(n4924), .ZN(n9602) );
  AND2_X1 U5986 ( .A1(n4657), .A2(n5785), .ZN(n9637) );
  NAND2_X1 U5987 ( .A1(n7802), .A2(n5867), .ZN(n4657) );
  NAND2_X1 U5988 ( .A1(n9657), .A2(n8349), .ZN(n9643) );
  AND2_X1 U5989 ( .A1(n5762), .A2(n5761), .ZN(n9668) );
  NAND2_X1 U5990 ( .A1(n9679), .A2(n8480), .ZN(n9659) );
  AND2_X1 U5991 ( .A1(n5053), .A2(n5052), .ZN(n9672) );
  INV_X1 U5992 ( .A(n5053), .ZN(n9702) );
  NAND2_X1 U5993 ( .A1(n4913), .A2(n4917), .ZN(n8196) );
  NAND2_X1 U5994 ( .A1(n7895), .A2(n4919), .ZN(n4913) );
  NAND2_X1 U5995 ( .A1(n4705), .A2(n5046), .ZN(n8198) );
  NAND2_X1 U5996 ( .A1(n7894), .A2(n5047), .ZN(n4705) );
  NAND2_X1 U5997 ( .A1(n4921), .A2(n8335), .ZN(n8003) );
  NAND2_X1 U5998 ( .A1(n7893), .A2(n5716), .ZN(n8002) );
  NAND2_X1 U5999 ( .A1(n6177), .A2(n9874), .ZN(n9490) );
  OAI21_X1 U6000 ( .B1(n7473), .B2(n4719), .A(n4716), .ZN(n7604) );
  NAND2_X1 U6001 ( .A1(n7471), .A2(n5652), .ZN(n7605) );
  INV_X1 U6002 ( .A(n9495), .ZN(n9853) );
  NAND2_X1 U6003 ( .A1(n5675), .A2(n5674), .ZN(n9358) );
  INV_X1 U6004 ( .A(n9860), .ZN(n7235) );
  INV_X1 U6005 ( .A(n8454), .ZN(n7185) );
  INV_X1 U6006 ( .A(n9618), .ZN(n9806) );
  AND2_X1 U6007 ( .A1(n5951), .A2(n6890), .ZN(n9874) );
  XNOR2_X1 U6008 ( .A(n6210), .B(n6209), .ZN(n9816) );
  OAI21_X1 U6009 ( .B1(n6247), .B2(n6246), .A(n6207), .ZN(n6210) );
  INV_X1 U6010 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10409) );
  INV_X1 U6011 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10494) );
  NOR2_X1 U6012 ( .A1(n5425), .A2(n5625), .ZN(n5426) );
  INV_X1 U6013 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10414) );
  INV_X1 U6014 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U6015 ( .A1(n5475), .A2(n5462), .ZN(n8001) );
  INV_X1 U6016 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U6017 ( .A1(n5026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5456) );
  INV_X1 U6018 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10214) );
  INV_X1 U6019 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10422) );
  INV_X1 U6020 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7321) );
  NAND2_X1 U6021 ( .A1(n4969), .A2(n4967), .ZN(n5687) );
  NAND2_X1 U6022 ( .A1(n4969), .A2(n5337), .ZN(n5685) );
  INV_X1 U6023 ( .A(n7381), .ZN(n9844) );
  AND2_X1 U6024 ( .A1(n5641), .A2(n5627), .ZN(n7062) );
  NAND2_X1 U6025 ( .A1(n5611), .A2(n5610), .ZN(n5609) );
  NAND2_X1 U6026 ( .A1(n5602), .A2(n5318), .ZN(n5520) );
  NAND2_X1 U6027 ( .A1(n5568), .A2(n5569), .ZN(n6932) );
  NAND2_X1 U6028 ( .A1(n4797), .A2(n4796), .ZN(n4795) );
  INV_X1 U6029 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4797) );
  NOR2_X1 U6030 ( .A1(n6931), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U6031 ( .A(n5543), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9428) );
  AOI21_X1 U6032 ( .B1(n5288), .B2(n9994), .A(n4682), .ZN(n5071) );
  OR2_X1 U6033 ( .A1(n5210), .A2(n9998), .ZN(n5086) );
  OAI21_X1 U6034 ( .B1(n9227), .B2(n9226), .A(n9383), .ZN(n9231) );
  AOI211_X1 U6035 ( .C1(n9256), .C2(n9407), .A(n9255), .B(n9254), .ZN(n9257)
         );
  NAND2_X1 U6036 ( .A1(n4806), .A2(n4807), .ZN(n4659) );
  NAND2_X1 U6037 ( .A1(n4806), .A2(n8401), .ZN(n4658) );
  INV_X1 U6038 ( .A(n4661), .ZN(n4660) );
  AND2_X1 U6039 ( .A1(n4892), .A2(n4893), .ZN(n9500) );
  NOR2_X1 U6040 ( .A1(n5480), .A2(n5482), .ZN(n5932) );
  OAI21_X1 U6041 ( .B1(n5942), .B2(n9911), .A(n5943), .ZN(P1_U3519) );
  NOR2_X1 U6042 ( .A1(n5939), .A2(n5941), .ZN(n5943) );
  AND4_X1 U6043 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(n5984)
         );
  AND2_X1 U6044 ( .A1(n4728), .A2(n4520), .ZN(n4506) );
  INV_X2 U6045 ( .A(n6322), .ZN(n4686) );
  AND2_X1 U6046 ( .A1(n4623), .A2(n9296), .ZN(n4507) );
  AND2_X1 U6047 ( .A1(n4982), .A2(n8940), .ZN(n4508) );
  OAI211_X1 U6048 ( .C1(n5574), .C2(n6934), .A(n5590), .B(n5589), .ZN(n7198)
         );
  INV_X1 U6049 ( .A(n7198), .ZN(n7443) );
  OR2_X1 U6050 ( .A1(n6081), .A2(n4615), .ZN(n4510) );
  NAND2_X1 U6051 ( .A1(n6521), .A2(n6520), .ZN(n8608) );
  NAND3_X1 U6052 ( .A1(n5191), .A2(n4509), .A3(n4695), .ZN(n4511) );
  AND3_X1 U6053 ( .A1(n4534), .A2(n5070), .A3(n5453), .ZN(n4512) );
  AND2_X1 U6054 ( .A1(n4876), .A2(n4875), .ZN(n4513) );
  AND2_X1 U6055 ( .A1(n4885), .A2(n4884), .ZN(n4514) );
  NAND4_X1 U6056 ( .A1(n8507), .A2(n5457), .A3(n8537), .A4(n8503), .ZN(n4515)
         );
  AND3_X1 U6057 ( .A1(n4903), .A2(n5519), .A3(n5610), .ZN(n4516) );
  AND2_X1 U6058 ( .A1(n8390), .A2(n4976), .ZN(n4517) );
  INV_X1 U6059 ( .A(n9907), .ZN(n8058) );
  AND2_X1 U6060 ( .A1(n5694), .A2(n5693), .ZN(n9907) );
  INV_X1 U6061 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6230) );
  AND3_X1 U6062 ( .A1(n6335), .A2(n6334), .A3(n6333), .ZN(n7948) );
  OAI21_X1 U6063 ( .B1(n4650), .B2(n4940), .A(n4647), .ZN(n5758) );
  AND3_X1 U6064 ( .A1(n8430), .A2(n9627), .A3(n4654), .ZN(n4518) );
  OR2_X1 U6065 ( .A1(n5728), .A2(n5050), .ZN(n4519) );
  NAND2_X1 U6066 ( .A1(n5719), .A2(n5452), .ZN(n5509) );
  XNOR2_X1 U6067 ( .A(n4637), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6068 ( .A1(n6030), .A2(n6034), .ZN(n7855) );
  NAND2_X1 U6069 ( .A1(n4963), .A2(n4572), .ZN(n4960) );
  AND2_X1 U6070 ( .A1(n4961), .A2(n4583), .ZN(n4958) );
  NAND2_X1 U6071 ( .A1(n5031), .A2(n7528), .ZN(n7404) );
  AND2_X1 U6072 ( .A1(n5136), .A2(n5135), .ZN(n6400) );
  AND2_X1 U6073 ( .A1(n4730), .A2(n8869), .ZN(n4520) );
  NAND2_X1 U6074 ( .A1(n5474), .A2(n5473), .ZN(n5951) );
  XNOR2_X1 U6075 ( .A(n5456), .B(n5455), .ZN(n5901) );
  NAND2_X1 U6076 ( .A1(n5208), .A2(n5209), .ZN(n6261) );
  NAND3_X1 U6077 ( .A1(n6260), .A2(n6259), .A3(n5076), .ZN(n7298) );
  INV_X1 U6078 ( .A(n8773), .ZN(n4688) );
  AOI21_X1 U6079 ( .B1(n8552), .B2(n4995), .A(n4993), .ZN(n4990) );
  AND2_X1 U6080 ( .A1(n8686), .A2(n8556), .ZN(n4521) );
  AND2_X2 U6081 ( .A1(n5457), .A2(n8001), .ZN(n8398) );
  AND2_X1 U6082 ( .A1(n6238), .A2(n6240), .ZN(n6267) );
  AND2_X1 U6083 ( .A1(n8904), .A2(n6820), .ZN(n4522) );
  XNOR2_X1 U6084 ( .A(n6236), .B(n6235), .ZN(n6240) );
  INV_X1 U6085 ( .A(n4928), .ZN(n4927) );
  NAND2_X1 U6086 ( .A1(n8359), .A2(n9611), .ZN(n4928) );
  OR2_X1 U6087 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4523) );
  NAND2_X1 U6088 ( .A1(n9637), .A2(n9613), .ZN(n8359) );
  AND2_X1 U6089 ( .A1(n5599), .A2(n5398), .ZN(n5522) );
  NOR2_X1 U6090 ( .A1(n6809), .A2(n6808), .ZN(n4524) );
  INV_X1 U6091 ( .A(n8933), .ZN(n4775) );
  OR2_X1 U6092 ( .A1(n5112), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4525) );
  AND2_X1 U6093 ( .A1(n7167), .A2(n5999), .ZN(n4526) );
  NAND4_X1 U6094 ( .A1(n6299), .A2(n6298), .A3(n6297), .A4(n6296), .ZN(n8777)
         );
  INV_X1 U6095 ( .A(n8777), .ZN(n6303) );
  INV_X1 U6096 ( .A(n8322), .ZN(n4912) );
  NAND2_X1 U6097 ( .A1(n5029), .A2(n5951), .ZN(n5982) );
  NAND2_X1 U6098 ( .A1(n9795), .A2(n6150), .ZN(n4527) );
  NAND2_X1 U6099 ( .A1(n8395), .A2(n8394), .ZN(n9483) );
  INV_X1 U6100 ( .A(n9483), .ZN(n9790) );
  OR2_X1 U6101 ( .A1(n6741), .A2(n6740), .ZN(n8609) );
  AND2_X1 U6102 ( .A1(n5003), .A2(n5002), .ZN(n4528) );
  OR3_X1 U6103 ( .A1(n6760), .A2(n6759), .A3(n6829), .ZN(n4529) );
  NAND2_X1 U6104 ( .A1(n5486), .A2(n5485), .ZN(n9745) );
  INV_X1 U6105 ( .A(n9603), .ZN(n4832) );
  INV_X1 U6106 ( .A(n8335), .ZN(n4920) );
  AND2_X1 U6107 ( .A1(n5914), .A2(n8314), .ZN(n4530) );
  XNOR2_X1 U6108 ( .A(n5491), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5497) );
  NOR2_X1 U6109 ( .A1(n5586), .A2(n4523), .ZN(n5599) );
  AND4_X1 U6110 ( .A1(n9603), .A2(n9640), .A3(n8429), .A4(n8428), .ZN(n4531)
         );
  AND2_X1 U6111 ( .A1(n10039), .A2(n8772), .ZN(n4532) );
  NAND2_X1 U6112 ( .A1(n5191), .A2(n4528), .ZN(n4533) );
  INV_X1 U6113 ( .A(n9783), .ZN(n9248) );
  NAND2_X1 U6114 ( .A1(n5721), .A2(n5720), .ZN(n9783) );
  NOR2_X1 U6115 ( .A1(n9250), .A2(n9251), .ZN(n9249) );
  AOI21_X1 U6116 ( .B1(n6842), .B2(n9060), .A(n6841), .ZN(n8655) );
  AND4_X1 U6117 ( .A1(n5449), .A2(n5402), .A3(n5690), .A4(n5760), .ZN(n4534)
         );
  AND2_X1 U6118 ( .A1(n4950), .A2(n4646), .ZN(n4535) );
  AND2_X1 U6119 ( .A1(n4626), .A2(n9317), .ZN(n4536) );
  NAND2_X1 U6120 ( .A1(n5191), .A2(n4509), .ZN(n6769) );
  AND4_X1 U6121 ( .A1(n5669), .A2(n5668), .A3(n5667), .A4(n5666), .ZN(n9353)
         );
  AND2_X1 U6122 ( .A1(n4880), .A2(n9600), .ZN(n4537) );
  AND2_X1 U6123 ( .A1(n5735), .A2(n5734), .ZN(n9832) );
  AND2_X1 U6124 ( .A1(n5038), .A2(n5040), .ZN(n4538) );
  INV_X1 U6125 ( .A(n9529), .ZN(n9795) );
  NAND2_X1 U6126 ( .A1(n5869), .A2(n5868), .ZN(n9529) );
  INV_X1 U6127 ( .A(n9761), .ZN(n9653) );
  NAND2_X1 U6128 ( .A1(n5776), .A2(n5775), .ZN(n9761) );
  NAND2_X1 U6129 ( .A1(n9577), .A2(n4878), .ZN(n4879) );
  INV_X1 U6130 ( .A(n9562), .ZN(n9800) );
  NAND2_X1 U6131 ( .A1(n5836), .A2(n5835), .ZN(n9562) );
  INV_X1 U6132 ( .A(n8147), .ZN(n8024) );
  NAND2_X1 U6133 ( .A1(n5708), .A2(n5707), .ZN(n8147) );
  AND2_X1 U6134 ( .A1(n9709), .A2(n9416), .ZN(n5058) );
  INV_X1 U6135 ( .A(n5058), .ZN(n5052) );
  NAND2_X1 U6136 ( .A1(n5458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5466) );
  OR2_X1 U6137 ( .A1(n9677), .A2(n9662), .ZN(n4539) );
  OR2_X1 U6138 ( .A1(n7751), .A2(n7750), .ZN(n4540) );
  OR2_X1 U6139 ( .A1(n8659), .A2(n8767), .ZN(n6753) );
  AND2_X1 U6140 ( .A1(n5332), .A2(n4644), .ZN(n4541) );
  NOR2_X2 U6141 ( .A1(n5499), .A2(n9824), .ZN(n4542) );
  AND2_X1 U6142 ( .A1(n5893), .A2(n4527), .ZN(n4543) );
  OR2_X1 U6143 ( .A1(n8781), .A2(n7301), .ZN(n7461) );
  INV_X1 U6144 ( .A(n4965), .ZN(n4964) );
  OAI21_X1 U6145 ( .B1(n4970), .B2(n4966), .A(n5339), .ZN(n4965) );
  AND2_X1 U6146 ( .A1(n7108), .A2(n5951), .ZN(n4544) );
  AND2_X1 U6147 ( .A1(n5454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4545) );
  INV_X1 U6148 ( .A(n4836), .ZN(n4835) );
  NOR2_X1 U6149 ( .A1(n8366), .A2(n8398), .ZN(n4836) );
  AND2_X1 U6150 ( .A1(n4861), .A2(n4860), .ZN(n4546) );
  NAND2_X1 U6151 ( .A1(n6074), .A2(n6089), .ZN(n4547) );
  AND2_X1 U6152 ( .A1(n8513), .A2(n8289), .ZN(n9525) );
  INV_X1 U6153 ( .A(n4817), .ZN(n4816) );
  OAI21_X1 U6154 ( .B1(n8392), .B2(n4818), .A(n8391), .ZN(n4817) );
  INV_X1 U6155 ( .A(n5046), .ZN(n4708) );
  NAND2_X1 U6156 ( .A1(n4551), .A2(n4519), .ZN(n5046) );
  AND2_X1 U6157 ( .A1(n5670), .A2(n9353), .ZN(n4548) );
  INV_X1 U6158 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U6159 ( .A1(n8727), .A2(n8970), .ZN(n4549) );
  NAND2_X1 U6160 ( .A1(n9427), .A2(n9860), .ZN(n8460) );
  AND3_X1 U6161 ( .A1(n5191), .A2(n4509), .A3(n4698), .ZN(n5114) );
  INV_X1 U6162 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U6163 ( .A1(n4752), .A2(n6651), .ZN(n4751) );
  INV_X1 U6164 ( .A(n4967), .ZN(n4966) );
  NOR2_X1 U6165 ( .A1(n5684), .A2(n4968), .ZN(n4967) );
  AND2_X1 U6166 ( .A1(n5348), .A2(SI_16_), .ZN(n4550) );
  INV_X1 U6167 ( .A(n7342), .ZN(n9427) );
  AND4_X1 U6168 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n7342)
         );
  NAND2_X1 U6169 ( .A1(n9783), .A2(n9417), .ZN(n4551) );
  INV_X1 U6170 ( .A(n4940), .ZN(n4939) );
  NAND2_X1 U6171 ( .A1(n4942), .A2(n4941), .ZN(n4940) );
  INV_X1 U6172 ( .A(n7360), .ZN(n9425) );
  AND4_X1 U6173 ( .A1(n5598), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n7360)
         );
  NAND2_X1 U6174 ( .A1(n8387), .A2(n8385), .ZN(n4552) );
  INV_X1 U6175 ( .A(n7279), .ZN(n9426) );
  AND4_X1 U6176 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n7279)
         );
  NAND2_X1 U6177 ( .A1(n9496), .A2(n4893), .ZN(n4553) );
  INV_X1 U6178 ( .A(n8434), .ZN(n8392) );
  AND2_X1 U6179 ( .A1(n8496), .A2(n8499), .ZN(n8434) );
  AND2_X1 U6180 ( .A1(n6674), .A2(n6837), .ZN(n4554) );
  AND2_X1 U6181 ( .A1(n4823), .A2(n4821), .ZN(n4555) );
  AND2_X1 U6182 ( .A1(n5051), .A2(n4703), .ZN(n4556) );
  AND2_X1 U6183 ( .A1(n4779), .A2(n6799), .ZN(n4557) );
  AND2_X1 U6184 ( .A1(n4706), .A2(n5052), .ZN(n4558) );
  AND2_X1 U6185 ( .A1(n4787), .A2(n4786), .ZN(n4559) );
  NAND2_X1 U6186 ( .A1(n9286), .A2(n9285), .ZN(n4560) );
  AND2_X1 U6187 ( .A1(n8641), .A2(n8637), .ZN(n4561) );
  INV_X1 U6188 ( .A(n5610), .ZN(n4953) );
  AND2_X1 U6189 ( .A1(n5325), .A2(n5324), .ZN(n5610) );
  NAND2_X1 U6190 ( .A1(n5604), .A2(n5603), .ZN(n5602) );
  OR3_X1 U6191 ( .A1(n5112), .A2(n5004), .A3(P2_IR_REG_22__SCAN_IN), .ZN(n4562) );
  INV_X1 U6192 ( .A(n8373), .ZN(n9572) );
  AND2_X1 U6193 ( .A1(n8438), .A2(n8447), .ZN(n8373) );
  AND2_X1 U6194 ( .A1(n4929), .A2(n8359), .ZN(n4563) );
  INV_X1 U6195 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6196 ( .A1(n4771), .A2(n4766), .ZN(n4564) );
  INV_X1 U6197 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4713) );
  INV_X1 U6198 ( .A(n4502), .ZN(n6506) );
  AND4_X1 U6199 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n9576)
         );
  INV_X1 U6200 ( .A(n9576), .ZN(n4954) );
  NAND2_X1 U6201 ( .A1(n5884), .A2(n5883), .ZN(n9720) );
  INV_X1 U6202 ( .A(n9720), .ZN(n4875) );
  AND2_X1 U6203 ( .A1(n7817), .A2(n4887), .ZN(n4565) );
  AND2_X1 U6204 ( .A1(n5191), .A2(n5096), .ZN(n5193) );
  OR3_X1 U6205 ( .A1(n6173), .A2(n6172), .A3(n9402), .ZN(n4566) );
  AND2_X1 U6206 ( .A1(n7036), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U6207 ( .A1(n5719), .A2(n5024), .ZN(n5759) );
  NOR2_X1 U6208 ( .A1(n9404), .A2(n9398), .ZN(n4568) );
  INV_X1 U6209 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4698) );
  INV_X1 U6210 ( .A(n8099), .ZN(n4752) );
  XNOR2_X1 U6211 ( .A(n5102), .B(n5101), .ZN(n6845) );
  INV_X1 U6212 ( .A(n8480), .ZN(n4907) );
  AND2_X1 U6213 ( .A1(n6091), .A2(n6093), .ZN(n4569) );
  NOR2_X1 U6214 ( .A1(n9975), .A2(n5188), .ZN(n4570) );
  AND2_X1 U6215 ( .A1(n4921), .A2(n4919), .ZN(n4571) );
  NAND2_X1 U6216 ( .A1(n9664), .A2(n4880), .ZN(n4883) );
  OR2_X1 U6217 ( .A1(n5362), .A2(n10483), .ZN(n4572) );
  AND2_X1 U6218 ( .A1(n9741), .A2(n9413), .ZN(n4573) );
  NOR2_X1 U6219 ( .A1(n5460), .A2(n5625), .ZN(n4574) );
  NAND2_X1 U6220 ( .A1(n4983), .A2(n4985), .ZN(n4575) );
  NAND2_X1 U6221 ( .A1(n6084), .A2(n6083), .ZN(n4576) );
  INV_X1 U6222 ( .A(n5014), .ZN(n5013) );
  NAND2_X1 U6223 ( .A1(n5016), .A2(n5015), .ZN(n5014) );
  INV_X1 U6224 ( .A(n9311), .ZN(n5012) );
  INV_X1 U6225 ( .A(n5042), .ZN(n5041) );
  NOR2_X1 U6226 ( .A1(n9600), .A2(n9290), .ZN(n5042) );
  AND2_X1 U6227 ( .A1(n5363), .A2(SI_21_), .ZN(n4577) );
  NAND2_X1 U6228 ( .A1(n9384), .A2(n9380), .ZN(n4578) );
  AND2_X1 U6229 ( .A1(n6119), .A2(n6118), .ZN(n4579) );
  NAND2_X1 U6230 ( .A1(n5361), .A2(SI_20_), .ZN(n4580) );
  INV_X1 U6231 ( .A(n6802), .ZN(n4691) );
  AND3_X1 U6232 ( .A1(n9228), .A2(n9229), .A3(n9230), .ZN(n4581) );
  AND2_X1 U6233 ( .A1(n5008), .A2(n5007), .ZN(n4582) );
  OR2_X1 U6234 ( .A1(n5363), .A2(SI_21_), .ZN(n4583) );
  NOR2_X1 U6235 ( .A1(n8227), .A2(n8174), .ZN(n4584) );
  AND2_X1 U6236 ( .A1(n9015), .A2(n6696), .ZN(n4585) );
  NAND2_X1 U6237 ( .A1(n5451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5719) );
  AND2_X1 U6238 ( .A1(n4738), .A2(n6693), .ZN(n4586) );
  NOR2_X1 U6239 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4587) );
  AND2_X1 U6240 ( .A1(n4985), .A2(n4988), .ZN(n4588) );
  NAND2_X1 U6241 ( .A1(n5512), .A2(n5511), .ZN(n9709) );
  INV_X1 U6242 ( .A(n9709), .ZN(n4884) );
  INV_X1 U6243 ( .A(n7848), .ZN(n4678) );
  XNOR2_X1 U6244 ( .A(n5466), .B(n5467), .ZN(n8406) );
  INV_X1 U6245 ( .A(n8406), .ZN(n5944) );
  INV_X1 U6246 ( .A(n8423), .ZN(n5048) );
  NAND2_X1 U6247 ( .A1(n5191), .A2(n5003), .ZN(n5198) );
  AND2_X1 U6248 ( .A1(n7543), .A2(n7542), .ZN(n7670) );
  INV_X1 U6249 ( .A(n8398), .ZN(n4976) );
  NAND2_X1 U6250 ( .A1(n7528), .A2(n6003), .ZN(n7403) );
  NAND2_X1 U6251 ( .A1(n5018), .A2(n6034), .ZN(n7869) );
  AND2_X1 U6252 ( .A1(n5017), .A2(n6034), .ZN(n4589) );
  AND2_X1 U6253 ( .A1(n7219), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4590) );
  AND2_X1 U6254 ( .A1(n4753), .A2(n4750), .ZN(n4591) );
  INV_X1 U6255 ( .A(SI_20_), .ZN(n10483) );
  INV_X1 U6256 ( .A(n9926), .ZN(n9923) );
  XNOR2_X1 U6257 ( .A(n5121), .B(n6230), .ZN(n5208) );
  NAND4_X1 U6258 ( .A1(n6332), .A2(n6331), .A3(n6330), .A4(n6329), .ZN(n8774)
         );
  INV_X1 U6259 ( .A(n8774), .ZN(n4756) );
  AND2_X1 U6260 ( .A1(n5971), .A2(n7078), .ZN(n7181) );
  INV_X1 U6261 ( .A(n7230), .ZN(n4874) );
  INV_X1 U6262 ( .A(n8432), .ZN(n4975) );
  OR2_X1 U6263 ( .A1(n8539), .A2(n8538), .ZN(n4592) );
  NOR2_X1 U6264 ( .A1(n6775), .A2(n6774), .ZN(n4593) );
  INV_X1 U6265 ( .A(n8261), .ZN(n4666) );
  XNOR2_X1 U6266 ( .A(n6449), .B(n5098), .ZN(n8869) );
  INV_X1 U6267 ( .A(n8869), .ZN(n7462) );
  INV_X1 U6268 ( .A(n7805), .ZN(n4729) );
  XNOR2_X1 U6269 ( .A(n6770), .B(n4698), .ZN(n7805) );
  NAND2_X1 U6270 ( .A1(n9456), .A2(n9457), .ZN(n4676) );
  NAND2_X1 U6271 ( .A1(n4730), .A2(n7462), .ZN(n4594) );
  INV_X1 U6272 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4796) );
  INV_X1 U6273 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4711) );
  INV_X1 U6274 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4602) );
  INV_X1 U6275 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U6276 ( .A1(n5341), .A2(n5340), .ZN(n5718) );
  NAND2_X1 U6277 ( .A1(n9552), .A2(n8448), .ZN(n9542) );
  NAND2_X1 U6278 ( .A1(n9231), .A2(n4581), .ZN(P1_U3214) );
  OR2_X1 U6279 ( .A1(n9249), .A2(n4625), .ZN(n4619) );
  NAND2_X1 U6280 ( .A1(n9249), .A2(n4507), .ZN(n4621) );
  NAND2_X1 U6281 ( .A1(n5431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U6282 ( .A1(n7204), .A2(n7205), .ZN(n7168) );
  OAI211_X1 U6283 ( .C1(n5995), .C2(n4641), .A(n4638), .B(n6002), .ZN(n6003)
         );
  NAND2_X1 U6284 ( .A1(n7204), .A2(n4639), .ZN(n4638) );
  INV_X1 U6285 ( .A(n7205), .ZN(n4640) );
  NAND2_X1 U6286 ( .A1(n7168), .A2(n5995), .ZN(n7167) );
  NAND2_X1 U6287 ( .A1(n7567), .A2(n6024), .ZN(n6029) );
  NAND3_X1 U6288 ( .A1(n4950), .A2(n4646), .A3(n4953), .ZN(n4644) );
  NAND2_X1 U6289 ( .A1(n4651), .A2(n5341), .ZN(n4650) );
  INV_X1 U6290 ( .A(n5717), .ZN(n4652) );
  NAND3_X1 U6291 ( .A1(n8373), .A2(n4655), .A3(n4518), .ZN(n4653) );
  OAI21_X1 U6292 ( .B1(n5773), .B2(n5772), .A(n5361), .ZN(n5782) );
  NAND3_X1 U6293 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(P1_U3242) );
  INV_X2 U6294 ( .A(n6272), .ZN(n5416) );
  MUX2_X1 U6295 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6272), .Z(n5323) );
  AOI21_X1 U6296 ( .B1(n7846), .B2(n7845), .A(n4678), .ZN(n7912) );
  NAND2_X1 U6297 ( .A1(n7847), .A2(n4677), .ZN(n7849) );
  NAND2_X1 U6298 ( .A1(n7846), .A2(n4679), .ZN(n4677) );
  NAND2_X1 U6299 ( .A1(n6958), .A2(n4686), .ZN(n6355) );
  NAND2_X1 U6300 ( .A1(n6976), .A2(n4686), .ZN(n6369) );
  NAND2_X1 U6301 ( .A1(n7137), .A2(n4686), .ZN(n6390) );
  NAND2_X1 U6302 ( .A1(n7177), .A2(n4686), .ZN(n6402) );
  NAND2_X1 U6303 ( .A1(n7226), .A2(n4686), .ZN(n6412) );
  NAND2_X1 U6304 ( .A1(n7411), .A2(n4686), .ZN(n6432) );
  NAND2_X1 U6305 ( .A1(n7286), .A2(n4686), .ZN(n6423) );
  NAND2_X1 U6306 ( .A1(n7564), .A2(n4686), .ZN(n6442) );
  NAND2_X1 U6307 ( .A1(n7650), .A2(n4686), .ZN(n6453) );
  NAND2_X1 U6308 ( .A1(n7997), .A2(n4686), .ZN(n6493) );
  NAND2_X1 U6309 ( .A1(n7867), .A2(n4686), .ZN(n6485) );
  NAND2_X1 U6310 ( .A1(n7802), .A2(n4686), .ZN(n6502) );
  NAND2_X1 U6311 ( .A1(n8013), .A2(n4686), .ZN(n6467) );
  NAND2_X1 U6312 ( .A1(n8137), .A2(n4686), .ZN(n6461) );
  NAND2_X1 U6313 ( .A1(n8223), .A2(n4686), .ZN(n6475) );
  NAND2_X1 U6314 ( .A1(n8231), .A2(n4686), .ZN(n6523) );
  NAND2_X1 U6315 ( .A1(n8593), .A2(n4686), .ZN(n6547) );
  NAND2_X1 U6316 ( .A1(n8236), .A2(n4686), .ZN(n6534) );
  NAND2_X1 U6317 ( .A1(n9215), .A2(n4686), .ZN(n6560) );
  NAND2_X1 U6318 ( .A1(n8664), .A2(n4686), .ZN(n6249) );
  NAND2_X1 U6319 ( .A1(n9816), .A2(n4686), .ZN(n6212) );
  NAND4_X1 U6320 ( .A1(n4693), .A2(n4692), .A3(n6677), .A4(n4691), .ZN(n4690)
         );
  NAND2_X1 U6321 ( .A1(n6672), .A2(n4554), .ZN(n4692) );
  NAND2_X1 U6322 ( .A1(n6673), .A2(n4694), .ZN(n4693) );
  NAND3_X1 U6323 ( .A1(n4692), .A2(n4693), .A3(n6677), .ZN(n6679) );
  NAND2_X1 U6324 ( .A1(n4690), .A2(n6678), .ZN(n6681) );
  NAND3_X1 U6325 ( .A1(n5191), .A2(n4697), .A3(n4509), .ZN(n5112) );
  NAND2_X1 U6326 ( .A1(n7894), .A2(n4558), .ZN(n4702) );
  NAND2_X1 U6327 ( .A1(n4556), .A2(n4702), .ZN(n5057) );
  NAND2_X1 U6328 ( .A1(n4709), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U6329 ( .A1(n7473), .A2(n4716), .ZN(n4714) );
  NAND2_X1 U6330 ( .A1(n4714), .A2(n4715), .ZN(n7656) );
  NAND2_X2 U6331 ( .A1(n6966), .A2(n6931), .ZN(n5574) );
  OAI21_X2 U6332 ( .B1(n5808), .B2(n5035), .A(n5033), .ZN(n9557) );
  NAND3_X1 U6333 ( .A1(n4725), .A2(n4724), .A3(n4722), .ZN(P2_U3296) );
  OR2_X1 U6334 ( .A1(n6771), .A2(n4723), .ZN(n4722) );
  AOI21_X1 U6335 ( .B1(n6599), .B2(n4506), .A(n4593), .ZN(n4724) );
  NAND2_X1 U6336 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  OR2_X1 U6337 ( .A1(n6771), .A2(n4729), .ZN(n4727) );
  NAND2_X1 U6338 ( .A1(n6597), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U6339 ( .A1(n6521), .A2(n4733), .ZN(n4736) );
  NAND2_X1 U6340 ( .A1(n4736), .A2(n4735), .ZN(n6544) );
  NAND2_X1 U6341 ( .A1(n6430), .A2(n4585), .ZN(n4738) );
  NAND2_X1 U6342 ( .A1(n4741), .A2(n4739), .ZN(n6399) );
  NAND2_X1 U6343 ( .A1(n4744), .A2(n4742), .ZN(n6420) );
  NAND2_X1 U6344 ( .A1(n7632), .A2(n4745), .ZN(n6313) );
  NAND2_X1 U6345 ( .A1(n8098), .A2(n4760), .ZN(n4757) );
  NAND2_X1 U6346 ( .A1(n4757), .A2(n4758), .ZN(n8158) );
  OAI21_X1 U6347 ( .B1(n8937), .B2(n4771), .A(n4768), .ZN(n8903) );
  INV_X1 U6348 ( .A(n4763), .ZN(n8889) );
  OAI21_X1 U6349 ( .B1(n8937), .B2(n4564), .A(n4764), .ZN(n4763) );
  OAI21_X2 U6350 ( .B1(n8937), .B2(n6819), .A(n4767), .ZN(n8919) );
  NAND2_X1 U6351 ( .A1(n4780), .A2(n4557), .ZN(n8206) );
  NAND2_X1 U6352 ( .A1(n6798), .A2(n6797), .ZN(n8172) );
  NAND2_X1 U6353 ( .A1(n8990), .A2(n4785), .ZN(n4783) );
  NAND2_X1 U6354 ( .A1(n4783), .A2(n4784), .ZN(n8968) );
  INV_X1 U6355 ( .A(n4787), .ZN(n8988) );
  MUX2_X1 U6356 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6272), .Z(n5314) );
  MUX2_X1 U6357 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6272), .Z(n5328) );
  NAND3_X1 U6358 ( .A1(n4788), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6359 ( .A1(n5584), .A2(n5312), .ZN(n5604) );
  INV_X1 U6360 ( .A(n5318), .ZN(n4789) );
  OAI21_X1 U6361 ( .B1(n8410), .B2(n7109), .A(n4790), .ZN(n7110) );
  NAND2_X1 U6362 ( .A1(n8410), .A2(n7109), .ZN(n4790) );
  NAND2_X1 U6363 ( .A1(n5538), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4794) );
  OR2_X1 U6364 ( .A1(n5574), .A2(n6943), .ZN(n4792) );
  NAND2_X1 U6365 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4795), .ZN(n5552) );
  NAND2_X1 U6366 ( .A1(n8460), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U6367 ( .A1(n4799), .A2(n8398), .ZN(n4798) );
  NAND2_X1 U6368 ( .A1(n4801), .A2(n8296), .ZN(n4799) );
  NAND2_X1 U6369 ( .A1(n8460), .A2(n8398), .ZN(n4800) );
  NAND2_X1 U6370 ( .A1(n5906), .A2(n5907), .ZN(n7232) );
  INV_X1 U6371 ( .A(n8534), .ZN(n4804) );
  INV_X1 U6372 ( .A(n8540), .ZN(n4808) );
  NAND3_X1 U6373 ( .A1(n4512), .A2(n5059), .A3(n5405), .ZN(n4873) );
  NOR2_X1 U6374 ( .A1(n8386), .A2(n4819), .ZN(n4811) );
  NOR2_X1 U6375 ( .A1(n4809), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6376 ( .A1(n9483), .A2(n8398), .ZN(n4820) );
  NAND2_X1 U6377 ( .A1(n4822), .A2(n4823), .ZN(n8382) );
  NAND2_X1 U6378 ( .A1(n4840), .A2(n8312), .ZN(n8321) );
  AOI21_X1 U6379 ( .B1(n4847), .B2(n4846), .A(n9683), .ZN(n8351) );
  OR3_X1 U6380 ( .A1(n8340), .A2(n8477), .A3(n8478), .ZN(n8342) );
  AOI21_X1 U6381 ( .B1(n8365), .B2(n8398), .A(n8364), .ZN(n8368) );
  NOR2_X4 U6382 ( .A1(n5095), .A2(n5163), .ZN(n5191) );
  OAI21_X1 U6383 ( .B1(n8318), .B2(n8467), .A(n8470), .ZN(n8331) );
  AOI211_X1 U6384 ( .C1(n8337), .C2(n8474), .A(n4920), .B(n8336), .ZN(n8340)
         );
  NAND2_X1 U6385 ( .A1(n8399), .A2(n8400), .ZN(n4978) );
  OAI211_X1 U6386 ( .C1(n8300), .C2(n8299), .A(n8458), .B(n8459), .ZN(n8303)
         );
  NAND2_X1 U6387 ( .A1(n4978), .A2(n4972), .ZN(n8401) );
  NAND2_X1 U6388 ( .A1(n8397), .A2(n9483), .ZN(n4977) );
  AOI21_X1 U6389 ( .B1(n4977), .B2(n4973), .A(n8526), .ZN(n4972) );
  MUX2_X1 U6390 ( .A(n8353), .B(n8352), .S(n8398), .Z(n8363) );
  AOI21_X1 U6391 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8364) );
  INV_X1 U6392 ( .A(n4853), .ZN(n8791) );
  INV_X1 U6393 ( .A(n4851), .ZN(n8789) );
  NOR2_X1 U6394 ( .A1(n7589), .A2(n10012), .ZN(n7590) );
  OAI21_X1 U6395 ( .B1(n4856), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6901), .ZN(
        n4855) );
  OAI21_X1 U6396 ( .B1(n8838), .B2(n4867), .A(n4866), .ZN(n8857) );
  NAND2_X1 U6397 ( .A1(n4873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5413) );
  INV_X1 U6398 ( .A(n4879), .ZN(n9526) );
  INV_X1 U6399 ( .A(n4883), .ZN(n9617) );
  OAI211_X1 U6400 ( .C1(n5292), .C2(n4713), .A(n4889), .B(n4888), .ZN(n4891)
         );
  NAND3_X1 U6401 ( .A1(n5292), .A2(n5291), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4889) );
  NAND2_X1 U6402 ( .A1(n5295), .A2(n4890), .ZN(n5541) );
  NAND2_X1 U6403 ( .A1(n4891), .A2(SI_1_), .ZN(n5295) );
  NAND2_X1 U6404 ( .A1(n5929), .A2(n9701), .ZN(n4892) );
  OR2_X2 U6405 ( .A1(n5942), .A2(n9923), .ZN(n5931) );
  INV_X1 U6406 ( .A(n5928), .ZN(n4893) );
  NAND2_X1 U6407 ( .A1(n7600), .A2(n4910), .ZN(n4909) );
  NAND2_X1 U6408 ( .A1(n9628), .A2(n4924), .ZN(n4922) );
  NAND2_X1 U6409 ( .A1(n4922), .A2(n4923), .ZN(n9601) );
  NAND2_X1 U6410 ( .A1(n4930), .A2(n5834), .ZN(n5383) );
  XNOR2_X1 U6411 ( .A(n4930), .B(n5834), .ZN(n8223) );
  NAND2_X1 U6412 ( .A1(n5849), .A2(n5848), .ZN(n5863) );
  NAND2_X1 U6413 ( .A1(n5863), .A2(n5388), .ZN(n5880) );
  OAI21_X1 U6414 ( .B1(n5849), .B2(n4934), .A(n4931), .ZN(n4935) );
  AOI21_X1 U6415 ( .B1(n4933), .B2(n5388), .A(n4932), .ZN(n4931) );
  NAND2_X1 U6416 ( .A1(n5732), .A2(n4949), .ZN(n4947) );
  NAND2_X1 U6417 ( .A1(n5518), .A2(n5322), .ZN(n5611) );
  NAND2_X1 U6418 ( .A1(n4980), .A2(n4979), .ZN(n8617) );
  AOI21_X1 U6419 ( .B1(n8573), .B2(n8957), .A(n4981), .ZN(n4979) );
  NAND2_X1 U6420 ( .A1(n8676), .A2(n8573), .ZN(n4980) );
  INV_X1 U6421 ( .A(n8676), .ZN(n4982) );
  NAND2_X1 U6422 ( .A1(n4983), .A2(n4588), .ZN(n8687) );
  NAND3_X1 U6423 ( .A1(n4987), .A2(n4984), .A3(n8545), .ZN(n4983) );
  OR2_X2 U6424 ( .A1(n8547), .A2(n8546), .ZN(n4987) );
  OAI21_X2 U6425 ( .B1(n8552), .B2(n4993), .A(n4991), .ZN(n8562) );
  NAND2_X1 U6426 ( .A1(n8638), .A2(n8637), .ZN(n8667) );
  NAND2_X2 U6427 ( .A1(n8628), .A2(n8627), .ZN(n8638) );
  NAND2_X1 U6428 ( .A1(n8638), .A2(n4561), .ZN(n8669) );
  NAND2_X2 U6429 ( .A1(n7792), .A2(n7791), .ZN(n7980) );
  INV_X1 U6430 ( .A(n9303), .ZN(n5015) );
  INV_X1 U6431 ( .A(n6121), .ZN(n9338) );
  NAND2_X1 U6432 ( .A1(n5719), .A2(n5023), .ZN(n5026) );
  NAND2_X2 U6433 ( .A1(n5947), .A2(n5951), .ZN(n6163) );
  NAND2_X1 U6434 ( .A1(n6003), .A2(n6006), .ZN(n5032) );
  NAND2_X1 U6435 ( .A1(n5032), .A2(n7528), .ZN(n6016) );
  INV_X1 U6436 ( .A(n5036), .ZN(n5035) );
  NAND2_X1 U6437 ( .A1(n5038), .A2(n5036), .ZN(n9569) );
  NAND2_X1 U6438 ( .A1(n5808), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U6439 ( .A1(n5861), .A2(n5044), .ZN(n5043) );
  NAND2_X1 U6440 ( .A1(n5861), .A2(n5860), .ZN(n9524) );
  INV_X1 U6441 ( .A(n5744), .ZN(n5054) );
  NAND2_X1 U6442 ( .A1(n5744), .A2(n5743), .ZN(n9703) );
  XNOR2_X1 U6443 ( .A(n5704), .B(n5703), .ZN(n7137) );
  OAI21_X1 U6444 ( .B1(n5313), .B2(n5297), .A(n5296), .ZN(n5300) );
  NAND2_X1 U6445 ( .A1(n5313), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5296) );
  NAND2_X2 U6446 ( .A1(n7295), .A2(n7294), .ZN(n7678) );
  OR2_X1 U6447 ( .A1(n6231), .A2(n6233), .ZN(n5121) );
  INV_X1 U6448 ( .A(n7461), .ZN(n6605) );
  NAND2_X1 U6449 ( .A1(n8566), .A2(n8565), .ZN(n8573) );
  INV_X1 U6450 ( .A(n8686), .ZN(n8730) );
  NAND2_X1 U6451 ( .A1(n5463), .A2(n5079), .ZN(n5414) );
  OR2_X1 U6452 ( .A1(n6507), .A2(n6266), .ZN(n6270) );
  NAND2_X1 U6453 ( .A1(n9382), .A2(n6156), .ZN(n9223) );
  NOR2_X1 U6454 ( .A1(n9223), .A2(n5068), .ZN(n6195) );
  NAND2_X1 U6455 ( .A1(n9223), .A2(n6169), .ZN(n6197) );
  AND2_X1 U6456 ( .A1(n8001), .A2(n8406), .ZN(n7331) );
  NAND2_X1 U6457 ( .A1(n5415), .A2(n5414), .ZN(n5926) );
  OAI21_X1 U6458 ( .B1(n5982), .B2(n8454), .A(n5973), .ZN(n5974) );
  INV_X1 U6459 ( .A(n5497), .ZN(n5499) );
  OR3_X1 U6460 ( .A1(n5492), .A2(n5494), .A3(n5625), .ZN(n5496) );
  AOI21_X2 U6461 ( .B1(n8128), .B2(n8127), .A(n8126), .ZN(n8130) );
  NAND2_X2 U6463 ( .A1(n7455), .A2(n9061), .ZN(n10023) );
  NAND3_X1 U6464 ( .A1(n7450), .A2(n6884), .A3(n6883), .ZN(n10068) );
  AND2_X1 U6465 ( .A1(n6872), .A2(n6871), .ZN(n10061) );
  NOR2_X1 U6466 ( .A1(n5330), .A2(n5636), .ZN(n5061) );
  INV_X1 U6467 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5152) );
  AND2_X1 U6468 ( .A1(n7998), .A2(n6868), .ZN(n10040) );
  INV_X1 U6469 ( .A(n8922), .ZN(n8904) );
  OR2_X1 U6470 ( .A1(n5200), .A2(n5199), .ZN(n8845) );
  AND2_X1 U6471 ( .A1(n5331), .A2(n10454), .ZN(n5062) );
  OR2_X1 U6472 ( .A1(n6888), .A2(n9174), .ZN(n5063) );
  NAND2_X1 U6473 ( .A1(n6727), .A2(n6726), .ZN(n5064) );
  OR3_X1 U6474 ( .A1(n8699), .A2(n8978), .A3(n6881), .ZN(n5065) );
  AND2_X1 U6475 ( .A1(n9027), .A2(n6688), .ZN(n5066) );
  NOR2_X1 U6476 ( .A1(n6517), .A2(n8925), .ZN(n5067) );
  OR2_X1 U6477 ( .A1(n6888), .A2(n9101), .ZN(n5069) );
  AND3_X1 U6478 ( .A1(n5400), .A2(n5446), .A3(n10230), .ZN(n5070) );
  AND2_X1 U6479 ( .A1(n6754), .A2(n6753), .ZN(n5072) );
  AND2_X1 U6480 ( .A1(n6762), .A2(n6749), .ZN(n5073) );
  NOR2_X1 U6481 ( .A1(n5938), .A2(n9814), .ZN(n5939) );
  AND2_X1 U6482 ( .A1(n6254), .A2(n6762), .ZN(n5074) );
  NOR2_X1 U6483 ( .A1(n8596), .A2(n6730), .ZN(n5075) );
  INV_X1 U6484 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5297) );
  AND4_X1 U6485 ( .A1(n5727), .A2(n5726), .A3(n5725), .A4(n5724), .ZN(n9397)
         );
  INV_X1 U6486 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6215) );
  AND2_X1 U6487 ( .A1(n6258), .A2(n6257), .ZN(n5076) );
  INV_X1 U6488 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5293) );
  AND2_X1 U6489 ( .A1(n5678), .A2(n5677), .ZN(n5077) );
  AND2_X1 U6490 ( .A1(n6786), .A2(n7762), .ZN(n5078) );
  INV_X1 U6491 ( .A(n7298), .ZN(n7297) );
  AND2_X1 U6492 ( .A1(n6555), .A2(n6554), .ZN(n6824) );
  INV_X1 U6493 ( .A(n6824), .ZN(n8905) );
  INV_X1 U6494 ( .A(n9307), .ZN(n9697) );
  AND4_X1 U6495 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n9307)
         );
  AND4_X1 U6496 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n8993)
         );
  INV_X1 U6497 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5419) );
  NOR2_X1 U6498 ( .A1(n5408), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5079) );
  INV_X1 U6499 ( .A(n7657), .ZN(n5917) );
  XNOR2_X1 U6500 ( .A(n6161), .B(n5956), .ZN(n5080) );
  OR2_X1 U6501 ( .A1(n9832), .A2(n9307), .ZN(n5081) );
  INV_X1 U6502 ( .A(n9832), .ZN(n9408) );
  NAND2_X1 U6503 ( .A1(n8952), .A2(n6721), .ZN(n5082) );
  INV_X1 U6504 ( .A(n7613), .ZN(n5670) );
  NAND2_X1 U6505 ( .A1(n7329), .A2(n9490), .ZN(n9670) );
  AND2_X2 U6506 ( .A1(n5937), .A2(n5936), .ZN(n9913) );
  INV_X1 U6507 ( .A(n9509), .ZN(n5893) );
  AND2_X1 U6508 ( .A1(n6941), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5083) );
  AND2_X1 U6509 ( .A1(n5176), .A2(n6948), .ZN(n5084) );
  AND2_X1 U6510 ( .A1(n5207), .A2(n5206), .ZN(n5085) );
  INV_X1 U6511 ( .A(n6865), .ZN(n6604) );
  NAND2_X1 U6512 ( .A1(n6605), .A2(n6604), .ZN(n6606) );
  INV_X1 U6513 ( .A(n6609), .ZN(n6610) );
  NAND2_X1 U6514 ( .A1(n6610), .A2(n6881), .ZN(n6611) );
  NAND2_X1 U6515 ( .A1(n6612), .A2(n6611), .ZN(n6616) );
  INV_X1 U6516 ( .A(n8945), .ZN(n6726) );
  NOR2_X1 U6517 ( .A1(n6725), .A2(n6730), .ZN(n6727) );
  INV_X1 U6518 ( .A(n8993), .ZN(n6812) );
  INV_X1 U6519 ( .A(SI_9_), .ZN(n10454) );
  NAND2_X1 U6520 ( .A1(n5074), .A2(n6568), .ZN(n6569) );
  NAND2_X1 U6521 ( .A1(n9937), .A2(n5152), .ZN(n5151) );
  INV_X1 U6522 ( .A(n6092), .ZN(n6093) );
  INV_X1 U6523 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6524 ( .A1(n5901), .A2(n8537), .ZN(n5948) );
  INV_X1 U6525 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6526 ( .A1(n8636), .A2(n8922), .ZN(n8637) );
  OAI21_X1 U6527 ( .B1(n9937), .B2(n5152), .A(n5151), .ZN(n9933) );
  INV_X1 U6528 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5195) );
  INV_X1 U6529 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10460) );
  AND2_X1 U6530 ( .A1(n7692), .A2(n6786), .ZN(n6787) );
  INV_X1 U6531 ( .A(n7885), .ZN(n6336) );
  NOR2_X1 U6532 ( .A1(n9274), .A2(n9373), .ZN(n6102) );
  INV_X1 U6533 ( .A(n7406), .ZN(n6006) );
  NOR2_X1 U6534 ( .A1(n9783), .A2(n9417), .ZN(n5728) );
  NAND2_X1 U6535 ( .A1(n7358), .A2(n8301), .ZN(n7414) );
  OR2_X1 U6536 ( .A1(n5489), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6537 ( .A1(n5427), .A2(n5426), .ZN(n5430) );
  INV_X1 U6538 ( .A(SI_22_), .ZN(n10241) );
  INV_X1 U6539 ( .A(SI_17_), .ZN(n10411) );
  INV_X1 U6540 ( .A(SI_14_), .ZN(n5342) );
  INV_X1 U6541 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5399) );
  INV_X1 U6542 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6543 ( .A1(n6261), .A2(n6272), .ZN(n6322) );
  INV_X1 U6544 ( .A(n6507), .ZN(n6561) );
  NOR2_X1 U6545 ( .A1(n6421), .A2(n5195), .ZN(n5196) );
  INV_X1 U6546 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5122) );
  AOI21_X1 U6547 ( .B1(n7693), .B2(n6787), .A(n5078), .ZN(n7966) );
  AOI22_X1 U6548 ( .A1(n8968), .A2(n8967), .B1(n8558), .B2(n8699), .ZN(n8956)
         );
  INV_X1 U6549 ( .A(n9047), .ZN(n8211) );
  INV_X1 U6550 ( .A(n6087), .ZN(n6088) );
  INV_X1 U6551 ( .A(n7856), .ZN(n6033) );
  XNOR2_X1 U6552 ( .A(n5974), .B(n6161), .ZN(n5977) );
  OR2_X1 U6553 ( .A1(n5765), .A2(n5487), .ZN(n5777) );
  AND2_X1 U6554 ( .A1(n9489), .A2(n5888), .ZN(n9505) );
  AND2_X1 U6555 ( .A1(n5736), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U6556 ( .A1(n9907), .A2(n6063), .ZN(n5701) );
  NAND2_X1 U6557 ( .A1(n5907), .A2(n8457), .ZN(n8403) );
  NOR2_X1 U6558 ( .A1(n5938), .A2(n9780), .ZN(n5480) );
  NAND2_X1 U6559 ( .A1(n5901), .A2(n8525), .ZN(n5945) );
  OR2_X1 U6560 ( .A1(n7480), .A2(n7862), .ZN(n5652) );
  OR2_X1 U6561 ( .A1(n9423), .A2(n7525), .ZN(n5624) );
  NAND2_X1 U6562 ( .A1(n5909), .A2(n8459), .ZN(n7277) );
  INV_X1 U6563 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5455) );
  INV_X1 U6564 ( .A(SI_15_), .ZN(n5729) );
  INV_X1 U6565 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5690) );
  INV_X1 U6566 ( .A(n8780), .ZN(n7391) );
  AND2_X1 U6567 ( .A1(n8625), .A2(n8621), .ZN(n8701) );
  INV_X1 U6568 ( .A(n8761), .ZN(n8735) );
  NAND2_X1 U6569 ( .A1(n7256), .A2(n7288), .ZN(n8757) );
  INV_X1 U6570 ( .A(n8845), .ZN(n5201) );
  OR2_X1 U6571 ( .A1(n6548), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8657) );
  NOR2_X1 U6572 ( .A1(n9207), .A2(n7292), .ZN(n7449) );
  OR2_X1 U6573 ( .A1(n7455), .A2(n9063), .ZN(n8984) );
  AND2_X1 U6574 ( .A1(n6566), .A2(n6245), .ZN(n8880) );
  OR2_X1 U6575 ( .A1(n9194), .A2(n8544), .ZN(n6688) );
  INV_X1 U6576 ( .A(n9056), .ZN(n8174) );
  AND2_X1 U6577 ( .A1(n7243), .A2(n7258), .ZN(n7264) );
  INV_X1 U6578 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7729) );
  INV_X1 U6579 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7123) );
  AND2_X1 U6580 ( .A1(n9224), .A2(n9225), .ZN(n6156) );
  AND3_X1 U6581 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5592) );
  INV_X1 U6582 ( .A(n9393), .ZN(n9355) );
  INV_X1 U6583 ( .A(n9391), .ZN(n9376) );
  AND2_X1 U6584 ( .A1(n5797), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5799) );
  INV_X1 U6585 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8272) );
  NOR2_X1 U6586 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  NOR2_X1 U6587 ( .A1(n9562), .A2(n9544), .ZN(n5846) );
  INV_X1 U6588 ( .A(n9745), .ZN(n9600) );
  INV_X1 U6589 ( .A(n9414), .ZN(n9663) );
  AND2_X1 U6590 ( .A1(n8537), .A2(n5944), .ZN(n8523) );
  AOI22_X1 U6591 ( .A1(n9511), .A2(n9698), .B1(n9696), .B2(n9545), .ZN(n9512)
         );
  AND2_X1 U6592 ( .A1(n8479), .A2(n8339), .ZN(n8426) );
  INV_X1 U6593 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5460) );
  INV_X1 U6594 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5760) );
  INV_X1 U6595 ( .A(n6272), .ZN(n6931) );
  INV_X1 U6596 ( .A(n8757), .ZN(n8733) );
  INV_X1 U6597 ( .A(n8725), .ZN(n8754) );
  AND2_X1 U6598 ( .A1(n6531), .A2(n6530), .ZN(n8922) );
  NAND2_X1 U6599 ( .A1(n5111), .A2(n5110), .ZN(n7245) );
  AND3_X1 U6600 ( .A1(n7255), .A2(n10054), .A3(n6833), .ZN(n8102) );
  INV_X1 U6601 ( .A(n9069), .ZN(n9023) );
  OR2_X1 U6602 ( .A1(n8102), .A2(n7624), .ZN(n10004) );
  INV_X1 U6603 ( .A(n8984), .ZN(n10017) );
  INV_X1 U6604 ( .A(n9101), .ZN(n9121) );
  AND2_X1 U6605 ( .A1(n6419), .A2(n6688), .ZN(n9039) );
  OR2_X1 U6606 ( .A1(n8102), .A2(n10040), .ZN(n10045) );
  OR2_X1 U6607 ( .A1(n7261), .A2(n7242), .ZN(n6872) );
  AND3_X1 U6608 ( .A1(n6955), .A2(n7326), .A3(n7324), .ZN(n6183) );
  INV_X1 U6609 ( .A(n9402), .ZN(n9383) );
  AND3_X1 U6610 ( .A1(n5925), .A2(n5924), .A3(n5923), .ZN(n8432) );
  AND4_X1 U6611 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n9687)
         );
  AND4_X1 U6612 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n9685)
         );
  INV_X1 U6613 ( .A(n9852), .ZN(n9455) );
  AND2_X1 U6614 ( .A1(n6988), .A2(n7083), .ZN(n9849) );
  AND2_X1 U6615 ( .A1(n6988), .A2(n5926), .ZN(n9459) );
  NOR2_X1 U6616 ( .A1(n9722), .A2(n9866), .ZN(n9514) );
  AND2_X1 U6617 ( .A1(n8370), .A2(n8369), .ZN(n9603) );
  AND2_X1 U6618 ( .A1(n8523), .A2(n5922), .ZN(n9698) );
  INV_X1 U6619 ( .A(n9693), .ZN(n9863) );
  AND2_X1 U6620 ( .A1(n5945), .A2(n7331), .ZN(n9829) );
  NAND2_X1 U6621 ( .A1(n7346), .A2(n5904), .ZN(n9909) );
  AND2_X1 U6622 ( .A1(n8398), .A2(n8525), .ZN(n7114) );
  NAND2_X1 U6623 ( .A1(n5424), .A2(n5427), .ZN(n5471) );
  INV_X1 U6624 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10084) );
  INV_X1 U6625 ( .A(n8618), .ZN(n9145) );
  INV_X1 U6626 ( .A(n8109), .ZN(n10033) );
  INV_X1 U6627 ( .A(n8921), .ZN(n8769) );
  INV_X1 U6628 ( .A(n9037), .ZN(n9016) );
  INV_X1 U6629 ( .A(n9974), .ZN(n9998) );
  INV_X1 U6630 ( .A(n10023), .ZN(n8033) );
  NAND2_X1 U6631 ( .A1(n10023), .A2(n10004), .ZN(n9069) );
  NAND2_X1 U6632 ( .A1(n9078), .A2(n9077), .ZN(n9080) );
  NAND2_X1 U6633 ( .A1(n10065), .A2(n10047), .ZN(n9101) );
  NAND2_X1 U6634 ( .A1(n10065), .A2(n10045), .ZN(n9124) );
  NAND2_X1 U6635 ( .A1(n10052), .A2(n10047), .ZN(n9174) );
  NAND2_X1 U6636 ( .A1(n10052), .A2(n10045), .ZN(n9204) );
  NAND2_X1 U6637 ( .A1(n6851), .A2(n7258), .ZN(n7101) );
  INV_X1 U6638 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7868) );
  INV_X1 U6639 ( .A(n6400), .ZN(n9984) );
  AND2_X1 U6640 ( .A1(n6178), .A2(n9490), .ZN(n9299) );
  NAND2_X1 U6641 ( .A1(n6183), .A2(n6168), .ZN(n9402) );
  INV_X1 U6642 ( .A(n6150), .ZN(n9545) );
  INV_X1 U6643 ( .A(n9685), .ZN(n9416) );
  INV_X1 U6644 ( .A(n9397), .ZN(n9417) );
  INV_X1 U6645 ( .A(n9459), .ZN(n9845) );
  OR2_X1 U6646 ( .A1(n6970), .A2(n6968), .ZN(n9852) );
  OR2_X1 U6647 ( .A1(n9866), .A2(n7347), .ZN(n9693) );
  OR2_X1 U6648 ( .A1(n9866), .A2(n7330), .ZN(n9859) );
  NAND2_X1 U6649 ( .A1(n9926), .A2(n9829), .ZN(n9780) );
  AND2_X2 U6650 ( .A1(n5479), .A2(n5478), .ZN(n9926) );
  NAND2_X1 U6651 ( .A1(n9913), .A2(n9829), .ZN(n9814) );
  INV_X1 U6652 ( .A(n9913), .ZN(n9911) );
  INV_X1 U6653 ( .A(n9871), .ZN(n9868) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10415) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10206) );
  INV_X2 U6656 ( .A(n8779), .ZN(P2_U3893) );
  NAND2_X1 U6657 ( .A1(n5086), .A2(n5071), .ZN(P2_U3200) );
  AND2_X2 U6658 ( .A1(n6891), .A2(n6890), .ZN(P1_U3973) );
  NAND4_X1 U6659 ( .A1(n5093), .A2(n5090), .A3(n5092), .A4(n5091), .ZN(n5095)
         );
  NAND2_X1 U6660 ( .A1(n5119), .A2(n5118), .ZN(n5100) );
  INV_X1 U6661 ( .A(n6845), .ZN(n5111) );
  NAND2_X1 U6662 ( .A1(n4562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5104) );
  MUX2_X1 U6663 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5104), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5105) );
  INV_X1 U6664 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6665 ( .A1(n5109), .A2(n5108), .ZN(n6844) );
  NAND2_X1 U6666 ( .A1(n5112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5113) );
  INV_X1 U6667 ( .A(n5114), .ZN(n5115) );
  NAND2_X1 U6668 ( .A1(n5115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6669 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5116), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5117) );
  NAND2_X2 U6670 ( .A1(n6831), .A2(n6865), .ZN(n6881) );
  NAND2_X1 U6671 ( .A1(n7245), .A2(n6881), .ZN(n5120) );
  NAND2_X1 U6672 ( .A1(n5120), .A2(n6772), .ZN(n5252) );
  NAND2_X1 U6673 ( .A1(n5252), .A2(n6261), .ZN(n5124) );
  NAND2_X1 U6674 ( .A1(n5124), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  OR2_X1 U6675 ( .A1(n5163), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6676 ( .A1(n5172), .A2(n5173), .ZN(n5143) );
  INV_X1 U6677 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5125) );
  NAND4_X1 U6678 ( .A1(n5177), .A2(n5126), .A3(n5087), .A4(n5125), .ZN(n5127)
         );
  NOR2_X1 U6679 ( .A1(n5143), .A2(n5127), .ZN(n5139) );
  NAND2_X1 U6680 ( .A1(n5139), .A2(n5128), .ZN(n5141) );
  NAND2_X1 U6681 ( .A1(n5129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5137) );
  INV_X1 U6682 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6683 ( .A1(n5137), .A2(n5130), .ZN(n5131) );
  NAND2_X1 U6684 ( .A1(n5131), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6685 ( .A1(n5134), .A2(n5133), .ZN(n5136) );
  NAND2_X1 U6686 ( .A1(n5136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U6687 ( .A(n5132), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6410) );
  OR2_X1 U6688 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  XNOR2_X1 U6689 ( .A(n5137), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U6690 ( .A1(n5141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  XNOR2_X1 U6691 ( .A(n5138), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6377) );
  INV_X1 U6692 ( .A(n6377), .ZN(n8047) );
  OR2_X1 U6693 ( .A1(n5139), .A2(n6233), .ZN(n5140) );
  MUX2_X1 U6694 ( .A(n5140), .B(P2_IR_REG_31__SCAN_IN), .S(n5128), .Z(n5142)
         );
  NAND2_X1 U6695 ( .A1(n5142), .A2(n5141), .ZN(n7928) );
  INV_X1 U6696 ( .A(n7928), .ZN(n6367) );
  NAND2_X1 U6697 ( .A1(n5143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5178) );
  OAI21_X1 U6698 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6699 ( .A1(n5178), .A2(n5144), .ZN(n5146) );
  OAI21_X1 U6700 ( .B1(n5146), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5145) );
  XNOR2_X1 U6701 ( .A(n5145), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6356) );
  XNOR2_X1 U6702 ( .A(n5146), .B(n5087), .ZN(n6353) );
  NAND2_X1 U6703 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5148), .ZN(n5147) );
  NAND2_X1 U6704 ( .A1(n5259), .A2(n5148), .ZN(n5158) );
  NAND2_X1 U6705 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5153) );
  MUX2_X1 U6706 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5153), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5154) );
  INV_X1 U6707 ( .A(n5259), .ZN(n5257) );
  INV_X1 U6708 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5214) );
  NOR2_X1 U6709 ( .A1(n5214), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6710 ( .A1(n5259), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5156) );
  INV_X1 U6711 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U6712 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  NAND2_X1 U6713 ( .A1(n9937), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6714 ( .A1(n9931), .A2(n5157), .ZN(n5161) );
  NAND2_X1 U6715 ( .A1(n5158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5159) );
  MUX2_X1 U6716 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5159), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5160) );
  NAND2_X1 U6717 ( .A1(n5160), .A2(n5163), .ZN(n9953) );
  OR2_X1 U6718 ( .A1(n5161), .A2(n9953), .ZN(n5162) );
  NAND2_X1 U6719 ( .A1(n5161), .A2(n9953), .ZN(n6902) );
  NAND2_X1 U6720 ( .A1(n5163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6721 ( .A(n5165), .B(n5164), .ZN(n6935) );
  INV_X1 U6722 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U6723 ( .A(n6935), .B(n6293), .ZN(n6901) );
  NAND2_X1 U6724 ( .A1(n6935), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6725 ( .A1(n6905), .A2(n5166), .ZN(n5170) );
  NAND2_X1 U6726 ( .A1(n5167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6727 ( .A(n5169), .B(n5168), .ZN(n6945) );
  NAND2_X1 U6728 ( .A1(n5170), .A2(n6945), .ZN(n7503) );
  OR2_X1 U6729 ( .A1(n5172), .A2(n6233), .ZN(n5174) );
  XNOR2_X1 U6730 ( .A(n5174), .B(n5173), .ZN(n6941) );
  XNOR2_X1 U6731 ( .A(n6941), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7504) );
  AOI21_X1 U6732 ( .B1(n7505), .B2(n7503), .A(n7504), .ZN(n7507) );
  XNOR2_X1 U6733 ( .A(n5178), .B(n5177), .ZN(n6948) );
  INV_X1 U6734 ( .A(n6948), .ZN(n7594) );
  XNOR2_X1 U6735 ( .A(n5175), .B(n7594), .ZN(n7589) );
  INV_X1 U6736 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10012) );
  INV_X1 U6737 ( .A(n5175), .ZN(n5176) );
  NAND2_X1 U6738 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6739 ( .A1(n5179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5180) );
  XNOR2_X1 U6740 ( .A(n5180), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U6741 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6952), .ZN(n5181) );
  OAI21_X1 U6742 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6952), .A(n5181), .ZN(
        n8790) );
  NOR2_X1 U6743 ( .A1(n6353), .A2(n5182), .ZN(n5183) );
  INV_X1 U6744 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8107) );
  XNOR2_X1 U6745 ( .A(n5182), .B(n6353), .ZN(n7774) );
  NOR2_X1 U6746 ( .A1(n8107), .A2(n7774), .ZN(n7773) );
  NAND2_X1 U6747 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7835), .ZN(n5184) );
  OAI21_X1 U6748 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7835), .A(n5184), .ZN(
        n7824) );
  NOR2_X1 U6749 ( .A1(n6367), .A2(n5185), .ZN(n5186) );
  INV_X1 U6750 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7931) );
  NOR2_X1 U6751 ( .A1(n7931), .A2(n7930), .ZN(n7929) );
  NOR2_X1 U6752 ( .A1(n5186), .A2(n7929), .ZN(n8036) );
  INV_X1 U6753 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8177) );
  AOI22_X1 U6754 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6377), .B1(n8047), .B2(
        n8177), .ZN(n8035) );
  NOR2_X1 U6755 ( .A1(n8036), .A2(n8035), .ZN(n8034) );
  AOI21_X2 U6756 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8047), .A(n8034), .ZN(
        n5187) );
  NOR2_X1 U6757 ( .A1(n6388), .A2(n5187), .ZN(n5188) );
  INV_X1 U6758 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6393) );
  INV_X1 U6759 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6405) );
  XNOR2_X1 U6760 ( .A(n6400), .B(n6405), .ZN(n9997) );
  NOR2_X1 U6761 ( .A1(n6410), .A2(n5189), .ZN(n5190) );
  INV_X1 U6762 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9048) );
  NOR2_X1 U6763 ( .A1(n5191), .A2(n6233), .ZN(n5192) );
  MUX2_X1 U6764 ( .A(n6233), .B(n5192), .S(P2_IR_REG_16__SCAN_IN), .Z(n5194)
         );
  OR2_X1 U6765 ( .A1(n5194), .A2(n5193), .ZN(n8832) );
  INV_X1 U6766 ( .A(n8832), .ZN(n6421) );
  AOI22_X1 U6767 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n6421), .B1(n8832), .B2(
        n5195), .ZN(n8821) );
  NOR2_X1 U6768 ( .A1(n5193), .A2(n6233), .ZN(n5197) );
  MUX2_X1 U6769 ( .A(n6233), .B(n5197), .S(P2_IR_REG_17__SCAN_IN), .Z(n5200)
         );
  INV_X1 U6770 ( .A(n5198), .ZN(n5199) );
  INV_X1 U6771 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9019) );
  NOR2_X1 U6772 ( .A1(n5201), .A2(n5202), .ZN(n5203) );
  NAND2_X1 U6773 ( .A1(n5198), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6774 ( .A(n5204), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8863) );
  INV_X1 U6775 ( .A(n8863), .ZN(n8858) );
  INV_X1 U6776 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5205) );
  AOI22_X1 U6777 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8863), .B1(n8858), .B2(
        n5205), .ZN(n5206) );
  NOR2_X1 U6778 ( .A1(n8857), .A2(n5085), .ZN(n5210) );
  NOR2_X1 U6779 ( .A1(n5208), .A2(P2_U3151), .ZN(n9218) );
  AND2_X1 U6780 ( .A1(n5252), .A2(n9218), .ZN(n7143) );
  INV_X1 U6781 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6433) );
  MUX2_X1 U6782 ( .A(n9019), .B(n6433), .S(n8864), .Z(n5248) );
  XNOR2_X1 U6783 ( .A(n5248), .B(n8845), .ZN(n8841) );
  MUX2_X1 U6784 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8864), .Z(n5211) );
  OR2_X1 U6785 ( .A1(n5211), .A2(n8832), .ZN(n5246) );
  XNOR2_X1 U6786 ( .A(n5211), .B(n6421), .ZN(n8828) );
  MUX2_X1 U6787 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8864), .Z(n5212) );
  INV_X1 U6788 ( .A(n6410), .ZN(n8811) );
  OR2_X1 U6789 ( .A1(n5212), .A2(n8811), .ZN(n5245) );
  XNOR2_X1 U6790 ( .A(n5212), .B(n6410), .ZN(n8808) );
  MUX2_X1 U6791 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8864), .Z(n5213) );
  OR2_X1 U6792 ( .A1(n5213), .A2(n9984), .ZN(n5244) );
  XNOR2_X1 U6793 ( .A(n5213), .B(n6400), .ZN(n9991) );
  MUX2_X1 U6794 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8864), .Z(n5242) );
  INV_X1 U6795 ( .A(n6388), .ZN(n9963) );
  OR2_X1 U6796 ( .A1(n5242), .A2(n9963), .ZN(n5243) );
  MUX2_X1 U6797 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8864), .Z(n5239) );
  INV_X1 U6798 ( .A(n5239), .ZN(n5240) );
  MUX2_X1 U6799 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8864), .Z(n5220) );
  MUX2_X1 U6800 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8864), .Z(n5215) );
  XOR2_X1 U6801 ( .A(n7150), .B(n5215), .Z(n7149) );
  INV_X1 U6802 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6266) );
  MUX2_X1 U6803 ( .A(n5214), .B(n6266), .S(n8864), .Z(n7141) );
  NAND2_X1 U6804 ( .A1(n7141), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7148) );
  AOI22_X1 U6805 ( .A1(n7149), .A2(n7148), .B1(n5215), .B2(n7150), .ZN(n9940)
         );
  MUX2_X1 U6806 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8864), .Z(n5216) );
  XNOR2_X1 U6807 ( .A(n5216), .B(n9937), .ZN(n9941) );
  INV_X1 U6808 ( .A(n9937), .ZN(n5218) );
  INV_X1 U6809 ( .A(n5216), .ZN(n5217) );
  OAI22_X1 U6810 ( .A1(n9940), .A2(n9941), .B1(n5218), .B2(n5217), .ZN(n9956)
         );
  MUX2_X1 U6811 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8864), .Z(n5219) );
  XNOR2_X1 U6812 ( .A(n5219), .B(n9953), .ZN(n9957) );
  NOR2_X1 U6813 ( .A1(n9956), .A2(n9957), .ZN(n9955) );
  NOR2_X1 U6814 ( .A1(n5219), .A2(n9953), .ZN(n6892) );
  XNOR2_X1 U6815 ( .A(n5220), .B(n6935), .ZN(n6895) );
  NOR3_X1 U6816 ( .A1(n9955), .A2(n6892), .A3(n6895), .ZN(n6893) );
  AOI21_X1 U6817 ( .B1(n5220), .B2(n6935), .A(n6893), .ZN(n6915) );
  MUX2_X1 U6818 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8864), .Z(n5221) );
  XNOR2_X1 U6819 ( .A(n5221), .B(n6945), .ZN(n6914) );
  INV_X1 U6820 ( .A(n6945), .ZN(n5267) );
  INV_X1 U6821 ( .A(n5221), .ZN(n5222) );
  OAI22_X1 U6822 ( .A1(n6915), .A2(n6914), .B1(n5267), .B2(n5222), .ZN(n7498)
         );
  INV_X1 U6823 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6314) );
  INV_X1 U6824 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6317) );
  MUX2_X1 U6825 ( .A(n6314), .B(n6317), .S(n8864), .Z(n5223) );
  INV_X1 U6826 ( .A(n6941), .ZN(n7512) );
  NAND2_X1 U6827 ( .A1(n5223), .A2(n7512), .ZN(n5224) );
  OAI21_X1 U6828 ( .B1(n5223), .B2(n7512), .A(n5224), .ZN(n7497) );
  NOR2_X1 U6829 ( .A1(n7498), .A2(n7497), .ZN(n7585) );
  INV_X1 U6830 ( .A(n5224), .ZN(n7584) );
  MUX2_X1 U6831 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8864), .Z(n5225) );
  NOR2_X1 U6832 ( .A1(n5225), .A2(n6948), .ZN(n5226) );
  AOI21_X1 U6833 ( .B1(n5225), .B2(n6948), .A(n5226), .ZN(n7583) );
  OAI21_X1 U6834 ( .B1(n7585), .B2(n7584), .A(n7583), .ZN(n8784) );
  INV_X1 U6835 ( .A(n5226), .ZN(n8783) );
  INV_X1 U6836 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8026) );
  INV_X1 U6837 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6339) );
  MUX2_X1 U6838 ( .A(n8026), .B(n6339), .S(n8864), .Z(n5227) );
  NAND2_X1 U6839 ( .A1(n5227), .A2(n8795), .ZN(n5230) );
  INV_X1 U6840 ( .A(n5227), .ZN(n5228) );
  NAND2_X1 U6841 ( .A1(n5228), .A2(n6952), .ZN(n5229) );
  NAND2_X1 U6842 ( .A1(n5230), .A2(n5229), .ZN(n8782) );
  AOI21_X1 U6843 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n8786) );
  INV_X1 U6844 ( .A(n5230), .ZN(n7776) );
  INV_X1 U6845 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6346) );
  MUX2_X1 U6846 ( .A(n8107), .B(n6346), .S(n8864), .Z(n5231) );
  NAND2_X1 U6847 ( .A1(n5231), .A2(n6353), .ZN(n7827) );
  INV_X1 U6848 ( .A(n5231), .ZN(n5232) );
  INV_X1 U6849 ( .A(n6353), .ZN(n7782) );
  NAND2_X1 U6850 ( .A1(n5232), .A2(n7782), .ZN(n5233) );
  AND2_X1 U6851 ( .A1(n7827), .A2(n5233), .ZN(n7775) );
  OAI21_X1 U6852 ( .B1(n8786), .B2(n7776), .A(n7775), .ZN(n7828) );
  INV_X1 U6853 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6362) );
  INV_X1 U6854 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6359) );
  MUX2_X1 U6855 ( .A(n6362), .B(n6359), .S(n8864), .Z(n5234) );
  NAND2_X1 U6856 ( .A1(n5234), .A2(n6356), .ZN(n5237) );
  INV_X1 U6857 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6858 ( .A1(n5235), .A2(n7835), .ZN(n5236) );
  NAND2_X1 U6859 ( .A1(n5237), .A2(n5236), .ZN(n7826) );
  AOI21_X1 U6860 ( .B1(n7828), .B2(n7827), .A(n7826), .ZN(n7830) );
  INV_X1 U6861 ( .A(n5237), .ZN(n5238) );
  NOR2_X1 U6862 ( .A1(n7830), .A2(n5238), .ZN(n7924) );
  XNOR2_X1 U6863 ( .A(n5239), .B(n7928), .ZN(n7923) );
  NOR2_X1 U6864 ( .A1(n7924), .A2(n7923), .ZN(n7922) );
  AOI21_X1 U6865 ( .B1(n6367), .B2(n5240), .A(n7922), .ZN(n8042) );
  INV_X1 U6866 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6380) );
  MUX2_X1 U6867 ( .A(n8177), .B(n6380), .S(n8864), .Z(n5241) );
  NAND2_X1 U6868 ( .A1(n5241), .A2(n6377), .ZN(n8037) );
  NOR2_X1 U6869 ( .A1(n5241), .A2(n6377), .ZN(n8039) );
  AOI21_X1 U6870 ( .B1(n8042), .B2(n8037), .A(n8039), .ZN(n9968) );
  XNOR2_X1 U6871 ( .A(n5242), .B(n6388), .ZN(n9969) );
  NAND2_X1 U6872 ( .A1(n9968), .A2(n9969), .ZN(n9967) );
  NAND2_X1 U6873 ( .A1(n5243), .A2(n9967), .ZN(n9990) );
  NAND2_X1 U6874 ( .A1(n9991), .A2(n9990), .ZN(n9989) );
  NAND2_X1 U6875 ( .A1(n5244), .A2(n9989), .ZN(n8807) );
  NAND2_X1 U6876 ( .A1(n8808), .A2(n8807), .ZN(n8806) );
  NAND2_X1 U6877 ( .A1(n5245), .A2(n8806), .ZN(n8827) );
  NAND2_X1 U6878 ( .A1(n8828), .A2(n8827), .ZN(n8826) );
  NAND2_X1 U6879 ( .A1(n5246), .A2(n8826), .ZN(n8840) );
  NAND2_X1 U6880 ( .A1(n8841), .A2(n8840), .ZN(n8839) );
  INV_X1 U6881 ( .A(n8839), .ZN(n5247) );
  AOI21_X1 U6882 ( .B1(n5248), .B2(n5201), .A(n5247), .ZN(n5251) );
  MUX2_X1 U6883 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8864), .Z(n5250) );
  NOR2_X1 U6884 ( .A1(n5251), .A2(n5250), .ZN(n8861) );
  INV_X1 U6885 ( .A(n7254), .ZN(n5249) );
  NOR2_X1 U6886 ( .A1(n8861), .A2(n8779), .ZN(n5254) );
  NAND2_X1 U6887 ( .A1(n5251), .A2(n5250), .ZN(n8862) );
  NOR2_X1 U6888 ( .A1(n8864), .A2(P2_U3151), .ZN(n8237) );
  NAND2_X1 U6889 ( .A1(n5252), .A2(n8237), .ZN(n5253) );
  INV_X1 U6890 ( .A(n5208), .ZN(n6835) );
  INV_X1 U6891 ( .A(n9983), .ZN(n8796) );
  AOI21_X1 U6892 ( .B1(n5254), .B2(n8862), .A(n8796), .ZN(n5255) );
  INV_X1 U6893 ( .A(n8862), .ZN(n5256) );
  NOR2_X2 U6894 ( .A1(n8779), .A2(n6835), .ZN(n9993) );
  OAI21_X1 U6895 ( .B1(n8861), .B2(n5256), .A(n9993), .ZN(n5289) );
  INV_X1 U6896 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8855) );
  AOI22_X1 U6897 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8858), .B1(n8863), .B2(
        n8855), .ZN(n5283) );
  INV_X1 U6898 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9114) );
  AOI22_X1 U6899 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8832), .B1(n6421), .B2(
        n9114), .ZN(n8824) );
  INV_X1 U6900 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9120) );
  AOI22_X1 U6901 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9984), .B1(n6400), .B2(
        n9120), .ZN(n9988) );
  AOI22_X1 U6902 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8047), .B1(n6377), .B2(
        n6380), .ZN(n8045) );
  NAND2_X1 U6903 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7835), .ZN(n5273) );
  AOI22_X1 U6904 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7835), .B1(n6356), .B2(
        n6359), .ZN(n7833) );
  NAND2_X1 U6905 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6952), .ZN(n5270) );
  AOI22_X1 U6906 ( .A1(n8795), .A2(n6339), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n6952), .ZN(n8798) );
  INV_X1 U6907 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6275) );
  MUX2_X1 U6908 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6275), .S(n9937), .Z(n9929)
         );
  INV_X1 U6909 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7147) );
  AND2_X1 U6910 ( .A1(n7147), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5258) );
  OAI22_X1 U6911 ( .A1(n7150), .A2(n5258), .B1(n5257), .B2(n6266), .ZN(n7152)
         );
  INV_X1 U6912 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7151) );
  OR2_X1 U6913 ( .A1(n7152), .A2(n7151), .ZN(n7154) );
  NAND2_X1 U6914 ( .A1(n5259), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6915 ( .A1(n7154), .A2(n5260), .ZN(n9928) );
  NAND2_X1 U6916 ( .A1(n9929), .A2(n9928), .ZN(n9927) );
  NAND2_X1 U6917 ( .A1(n9937), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6918 ( .A1(n9927), .A2(n5261), .ZN(n5263) );
  INV_X1 U6919 ( .A(n9953), .ZN(n5262) );
  XNOR2_X1 U6920 ( .A(n5263), .B(n5262), .ZN(n9945) );
  NAND2_X1 U6921 ( .A1(n9945), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6922 ( .A1(n5263), .A2(n9953), .ZN(n5264) );
  NAND2_X1 U6923 ( .A1(n5265), .A2(n5264), .ZN(n6898) );
  INV_X1 U6924 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6295) );
  MUX2_X1 U6925 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6295), .S(n6935), .Z(n6899)
         );
  NAND2_X1 U6926 ( .A1(n6898), .A2(n6899), .ZN(n6897) );
  NAND2_X1 U6927 ( .A1(n6935), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6928 ( .A1(n6897), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6929 ( .A(n5268), .B(n5267), .ZN(n6918) );
  AOI22_X1 U6930 ( .A1(n6918), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n6945), .B2(
        n5268), .ZN(n7500) );
  MUX2_X1 U6931 ( .A(n6317), .B(P2_REG1_REG_6__SCAN_IN), .S(n6941), .Z(n7501)
         );
  NOR2_X1 U6932 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  AOI21_X1 U6933 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6941), .A(n7499), .ZN(
        n5269) );
  XOR2_X1 U6934 ( .A(n6948), .B(n5269), .Z(n7582) );
  INV_X1 U6935 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6328) );
  OAI22_X1 U6936 ( .A1(n7582), .A2(n6328), .B1(n7594), .B2(n5269), .ZN(n8799)
         );
  NAND2_X1 U6937 ( .A1(n8798), .A2(n8799), .ZN(n8797) );
  NAND2_X1 U6938 ( .A1(n7782), .A2(n5271), .ZN(n5272) );
  NAND2_X1 U6939 ( .A1(n7833), .A2(n7832), .ZN(n7831) );
  NAND2_X1 U6940 ( .A1(n5273), .A2(n7831), .ZN(n5274) );
  NAND2_X1 U6941 ( .A1(n7928), .A2(n5274), .ZN(n5275) );
  XNOR2_X1 U6942 ( .A(n6367), .B(n5274), .ZN(n7926) );
  NAND2_X1 U6943 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7926), .ZN(n7925) );
  NAND2_X1 U6944 ( .A1(n9963), .A2(n5276), .ZN(n5277) );
  NAND2_X1 U6945 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U6946 ( .A1(n8811), .A2(n5278), .ZN(n5279) );
  NAND2_X1 U6947 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8815), .ZN(n8814) );
  NAND2_X1 U6948 ( .A1(n8845), .A2(n5280), .ZN(n5281) );
  NAND2_X1 U6949 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8849), .ZN(n8848) );
  NAND2_X1 U6950 ( .A1(n5281), .A2(n8848), .ZN(n5282) );
  NAND2_X1 U6951 ( .A1(n5283), .A2(n5282), .ZN(n8854) );
  OAI21_X1 U6952 ( .B1(n5283), .B2(n5282), .A(n8854), .ZN(n5288) );
  INV_X1 U6953 ( .A(n7143), .ZN(n5284) );
  OR2_X1 U6954 ( .A1(n5284), .A2(n6834), .ZN(n8876) );
  INV_X1 U6955 ( .A(n6772), .ZN(n5285) );
  NOR2_X1 U6956 ( .A1(n7245), .A2(n5285), .ZN(n5286) );
  INV_X1 U6957 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U6958 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8756) );
  OAI21_X1 U6959 ( .B1(n9982), .B2(n10144), .A(n8756), .ZN(n5287) );
  MUX2_X1 U6960 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5313), .Z(n5294) );
  NAND2_X1 U6961 ( .A1(n5294), .A2(SI_0_), .ZN(n5542) );
  OAI21_X1 U6962 ( .B1(n5541), .B2(n5542), .A(n5295), .ZN(n5550) );
  INV_X1 U6963 ( .A(n5300), .ZN(n5299) );
  INV_X1 U6964 ( .A(SI_2_), .ZN(n5298) );
  NAND2_X1 U6965 ( .A1(n5299), .A2(n5298), .ZN(n5301) );
  NAND2_X1 U6966 ( .A1(n5300), .A2(SI_2_), .ZN(n5302) );
  AND2_X1 U6967 ( .A1(n5301), .A2(n5302), .ZN(n5549) );
  NAND2_X1 U6968 ( .A1(n5550), .A2(n5549), .ZN(n5548) );
  NAND2_X1 U6969 ( .A1(n5548), .A2(n5302), .ZN(n5567) );
  MUX2_X1 U6970 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5313), .Z(n5305) );
  INV_X1 U6971 ( .A(n5305), .ZN(n5304) );
  INV_X1 U6972 ( .A(SI_3_), .ZN(n5303) );
  NAND2_X1 U6973 ( .A1(n5304), .A2(n5303), .ZN(n5306) );
  NAND2_X1 U6974 ( .A1(n5305), .A2(SI_3_), .ZN(n5307) );
  AND2_X1 U6975 ( .A1(n5306), .A2(n5307), .ZN(n5566) );
  NAND2_X1 U6976 ( .A1(n5567), .A2(n5566), .ZN(n5569) );
  NAND2_X1 U6977 ( .A1(n5569), .A2(n5307), .ZN(n5582) );
  MUX2_X1 U6978 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5313), .Z(n5308) );
  NAND2_X1 U6979 ( .A1(n5308), .A2(SI_4_), .ZN(n5312) );
  INV_X1 U6980 ( .A(n5308), .ZN(n5310) );
  INV_X1 U6981 ( .A(SI_4_), .ZN(n5309) );
  NAND2_X1 U6982 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  AND2_X1 U6983 ( .A1(n5312), .A2(n5311), .ZN(n5581) );
  NAND2_X1 U6984 ( .A1(n5582), .A2(n5581), .ZN(n5584) );
  NAND2_X1 U6985 ( .A1(n5314), .A2(SI_5_), .ZN(n5318) );
  INV_X1 U6986 ( .A(n5314), .ZN(n5316) );
  INV_X1 U6987 ( .A(SI_5_), .ZN(n5315) );
  NAND2_X1 U6988 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  AND2_X1 U6989 ( .A1(n5318), .A2(n5317), .ZN(n5603) );
  INV_X1 U6990 ( .A(n5319), .ZN(n5320) );
  INV_X1 U6991 ( .A(SI_6_), .ZN(n10434) );
  NAND2_X1 U6992 ( .A1(n5320), .A2(n10434), .ZN(n5321) );
  AND2_X1 U6993 ( .A1(n5322), .A2(n5321), .ZN(n5519) );
  NAND2_X1 U6994 ( .A1(n5323), .A2(SI_7_), .ZN(n5325) );
  INV_X1 U6995 ( .A(SI_7_), .ZN(n10217) );
  XNOR2_X1 U6996 ( .A(n5328), .B(SI_8_), .ZN(n5637) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5327) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5326) );
  MUX2_X1 U6999 ( .A(n5327), .B(n5326), .S(n5416), .Z(n5331) );
  XNOR2_X1 U7000 ( .A(n5331), .B(SI_9_), .ZN(n5639) );
  INV_X1 U7001 ( .A(n5639), .ZN(n5330) );
  INV_X1 U7002 ( .A(n5328), .ZN(n5329) );
  INV_X1 U7003 ( .A(SI_8_), .ZN(n10245) );
  NAND2_X1 U7004 ( .A1(n5329), .A2(n10245), .ZN(n5636) );
  MUX2_X1 U7005 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n5416), .Z(n5333) );
  NAND2_X1 U7006 ( .A1(n5333), .A2(SI_10_), .ZN(n5334) );
  OAI21_X1 U7007 ( .B1(n5333), .B2(SI_10_), .A(n5334), .ZN(n5653) );
  MUX2_X1 U7008 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5416), .Z(n5335) );
  XNOR2_X1 U7009 ( .A(n5335), .B(SI_11_), .ZN(n5671) );
  INV_X1 U7010 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U7011 ( .A1(n5336), .A2(n10263), .ZN(n5337) );
  MUX2_X1 U7012 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5416), .Z(n5338) );
  OAI21_X1 U7013 ( .B1(n5338), .B2(SI_12_), .A(n5339), .ZN(n5684) );
  MUX2_X1 U7014 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5416), .Z(n5702) );
  NAND2_X1 U7015 ( .A1(n5704), .A2(SI_13_), .ZN(n5340) );
  MUX2_X1 U7016 ( .A(n7178), .B(n10206), .S(n5416), .Z(n5343) );
  INV_X1 U7017 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U7018 ( .A1(n5344), .A2(SI_14_), .ZN(n5345) );
  NAND2_X1 U7019 ( .A1(n5346), .A2(n5345), .ZN(n5717) );
  MUX2_X1 U7020 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5416), .Z(n5730) );
  INV_X1 U7021 ( .A(n5730), .ZN(n5347) );
  MUX2_X1 U7022 ( .A(n7287), .B(n7321), .S(n5416), .Z(n5506) );
  NOR2_X1 U7023 ( .A1(n5348), .A2(SI_16_), .ZN(n5349) );
  MUX2_X1 U7024 ( .A(n7413), .B(n10422), .S(n5416), .Z(n5350) );
  INV_X1 U7025 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U7026 ( .A1(n5351), .A2(SI_17_), .ZN(n5352) );
  NAND2_X1 U7027 ( .A1(n5353), .A2(n5352), .ZN(n5745) );
  MUX2_X1 U7028 ( .A(n7565), .B(n10214), .S(n6931), .Z(n5354) );
  XNOR2_X1 U7029 ( .A(n5354), .B(SI_18_), .ZN(n5757) );
  INV_X1 U7030 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U7031 ( .A1(n5355), .A2(SI_18_), .ZN(n5356) );
  MUX2_X1 U7032 ( .A(n7651), .B(n10415), .S(n6931), .Z(n5358) );
  NAND2_X1 U7033 ( .A1(n5358), .A2(n5357), .ZN(n5361) );
  INV_X1 U7034 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U7035 ( .A1(n5359), .A2(SI_19_), .ZN(n5360) );
  NAND2_X1 U7036 ( .A1(n5361), .A2(n5360), .ZN(n5772) );
  MUX2_X1 U7037 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5416), .Z(n5783) );
  INV_X1 U7038 ( .A(n5783), .ZN(n5362) );
  MUX2_X1 U7039 ( .A(n7868), .B(n7891), .S(n5416), .Z(n5792) );
  MUX2_X1 U7040 ( .A(n7999), .B(n10469), .S(n6931), .Z(n5364) );
  NAND2_X1 U7041 ( .A1(n5364), .A2(n10241), .ZN(n5367) );
  INV_X1 U7042 ( .A(n5364), .ZN(n5365) );
  NAND2_X1 U7043 ( .A1(n5365), .A2(SI_22_), .ZN(n5366) );
  NAND2_X1 U7044 ( .A1(n5367), .A2(n5366), .ZN(n5483) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5368) );
  MUX2_X1 U7046 ( .A(n8016), .B(n5368), .S(n5416), .Z(n5369) );
  INV_X1 U7047 ( .A(SI_23_), .ZN(n10265) );
  NAND2_X1 U7048 ( .A1(n5369), .A2(n10265), .ZN(n5372) );
  INV_X1 U7049 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U7050 ( .A1(n5370), .A2(SI_23_), .ZN(n5371) );
  NAND2_X1 U7051 ( .A1(n5810), .A2(n5809), .ZN(n5812) );
  NAND2_X1 U7052 ( .A1(n5812), .A2(n5372), .ZN(n5823) );
  INV_X1 U7053 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8138) );
  MUX2_X1 U7054 ( .A(n8138), .B(n10414), .S(n5416), .Z(n5373) );
  INV_X1 U7055 ( .A(SI_24_), .ZN(n10397) );
  NAND2_X1 U7056 ( .A1(n5373), .A2(n10397), .ZN(n5376) );
  INV_X1 U7057 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U7058 ( .A1(n5374), .A2(SI_24_), .ZN(n5375) );
  NAND2_X1 U7059 ( .A1(n5823), .A2(n5822), .ZN(n5377) );
  INV_X1 U7060 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8224) );
  MUX2_X1 U7061 ( .A(n8224), .B(n10494), .S(n6931), .Z(n5379) );
  INV_X1 U7062 ( .A(SI_25_), .ZN(n5378) );
  NAND2_X1 U7063 ( .A1(n5379), .A2(n5378), .ZN(n5382) );
  INV_X1 U7064 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U7065 ( .A1(n5380), .A2(SI_25_), .ZN(n5381) );
  INV_X1 U7066 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8232) );
  MUX2_X1 U7067 ( .A(n8232), .B(n10409), .S(n6931), .Z(n5385) );
  INV_X1 U7068 ( .A(SI_26_), .ZN(n5384) );
  NAND2_X1 U7069 ( .A1(n5385), .A2(n5384), .ZN(n5862) );
  INV_X1 U7070 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U7071 ( .A1(n5386), .A2(SI_26_), .ZN(n5387) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6532) );
  INV_X1 U7073 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10182) );
  MUX2_X1 U7074 ( .A(n6532), .B(n10182), .S(n6931), .Z(n5389) );
  INV_X1 U7075 ( .A(SI_27_), .ZN(n10406) );
  NAND2_X1 U7076 ( .A1(n5389), .A2(n10406), .ZN(n5864) );
  AND2_X1 U7077 ( .A1(n5862), .A2(n5864), .ZN(n5388) );
  INV_X1 U7078 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U7079 ( .A1(n5390), .A2(SI_27_), .ZN(n5879) );
  MUX2_X1 U7080 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6931), .Z(n5392) );
  INV_X1 U7081 ( .A(SI_28_), .ZN(n5393) );
  XNOR2_X1 U7082 ( .A(n5392), .B(n5393), .ZN(n5881) );
  AND2_X1 U7083 ( .A1(n5879), .A2(n5881), .ZN(n5391) );
  NAND2_X1 U7084 ( .A1(n5880), .A2(n5391), .ZN(n5396) );
  INV_X1 U7085 ( .A(n5392), .ZN(n5394) );
  NAND2_X1 U7086 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  INV_X1 U7087 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9217) );
  INV_X1 U7088 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5397) );
  MUX2_X1 U7089 ( .A(n9217), .B(n5397), .S(n6931), .Z(n6198) );
  NOR2_X1 U7090 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5402) );
  NOR2_X1 U7091 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5404) );
  NOR2_X1 U7092 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5403) );
  NAND4_X1 U7093 ( .A1(n5429), .A2(n5404), .A3(n5403), .A4(n5460), .ZN(n5408)
         );
  INV_X1 U7094 ( .A(n5408), .ZN(n5405) );
  NAND2_X1 U7095 ( .A1(n5406), .A2(n5409), .ZN(n5489) );
  NOR2_X1 U7096 ( .A1(n5492), .A2(n5407), .ZN(n5412) );
  NAND2_X1 U7097 ( .A1(n9215), .A2(n5867), .ZN(n5418) );
  NAND2_X1 U7098 ( .A1(n8393), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5417) );
  INV_X1 U7099 ( .A(n9493), .ZN(n5938) );
  NAND2_X1 U7100 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5422) );
  INV_X1 U7101 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5423) );
  INV_X1 U7102 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5425) );
  AOI21_X1 U7103 ( .B1(n4503), .B2(n5429), .A(n4587), .ZN(n5431) );
  NAND2_X1 U7104 ( .A1(n5430), .A2(n5431), .ZN(n5472) );
  NAND3_X1 U7105 ( .A1(n5472), .A2(P1_B_REG_SCAN_IN), .A3(n5471), .ZN(n5432)
         );
  OR2_X1 U7106 ( .A1(n9867), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5435) );
  INV_X1 U7107 ( .A(n5472), .ZN(n5433) );
  OR2_X1 U7108 ( .A1(n5473), .A2(n5433), .ZN(n5434) );
  NAND2_X1 U7109 ( .A1(n5435), .A2(n5434), .ZN(n6167) );
  NOR4_X1 U7110 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5444) );
  NOR4_X1 U7111 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5443) );
  INV_X1 U7112 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9869) );
  INV_X1 U7113 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9870) );
  INV_X1 U7114 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10392) );
  INV_X1 U7115 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U7116 ( .A1(n9869), .A2(n9870), .A3(n10392), .A4(n10428), .ZN(n5441) );
  NOR4_X1 U7117 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5439) );
  NOR4_X1 U7118 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5438) );
  NOR4_X1 U7119 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5437) );
  NOR4_X1 U7120 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5436) );
  NAND4_X1 U7121 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(n5440)
         );
  NOR4_X1 U7122 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5441), .A4(n5440), .ZN(n5442) );
  AND3_X1 U7123 ( .A1(n5444), .A2(n5443), .A3(n5442), .ZN(n5445) );
  NOR2_X1 U7124 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5448) );
  NOR2_X1 U7125 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5447) );
  AND4_X1 U7126 ( .A1(n5449), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n5450)
         );
  NAND2_X1 U7127 ( .A1(n5524), .A2(n5450), .ZN(n5451) );
  NAND2_X1 U7128 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n5452) );
  INV_X1 U7129 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U7130 ( .A1(n5466), .A2(n5467), .ZN(n5461) );
  NAND2_X1 U7131 ( .A1(n5461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7132 ( .A1(n5459), .A2(n5460), .ZN(n5475) );
  NAND2_X1 U7133 ( .A1(n4574), .A2(n5461), .ZN(n5462) );
  INV_X1 U7134 ( .A(n5463), .ZN(n5464) );
  NAND2_X1 U7135 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7136 ( .A1(n7114), .A2(n8406), .ZN(n6176) );
  NAND3_X1 U7137 ( .A1(n6167), .A2(n7324), .A3(n6176), .ZN(n5933) );
  AND2_X1 U7138 ( .A1(n8523), .A2(n5945), .ZN(n5934) );
  NOR2_X1 U7139 ( .A1(n5933), .A2(n5934), .ZN(n5479) );
  OR2_X1 U7140 ( .A1(n9867), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5470) );
  INV_X1 U7141 ( .A(n5471), .ZN(n5468) );
  OR2_X1 U7142 ( .A1(n5473), .A2(n5468), .ZN(n5469) );
  NAND2_X1 U7143 ( .A1(n5475), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7144 ( .A1(n7326), .A2(n9874), .ZN(n9872) );
  INV_X1 U7145 ( .A(n9872), .ZN(n5478) );
  INV_X1 U7146 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5481) );
  NOR2_X1 U7147 ( .A1(n9926), .A2(n5481), .ZN(n5482) );
  XNOR2_X1 U7148 ( .A(n5484), .B(n5483), .ZN(n7997) );
  NAND2_X1 U7149 ( .A1(n7997), .A2(n5867), .ZN(n5486) );
  NAND2_X1 U7150 ( .A1(n8393), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7151 ( .A1(n5592), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5618) );
  NOR2_X1 U7152 ( .A1(n5618), .A2(n5617), .ZN(n5629) );
  NAND2_X1 U7153 ( .A1(n5629), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7154 ( .A1(n5695), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7155 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5487) );
  OR2_X1 U7156 ( .A1(n5799), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7157 ( .A1(n5799), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5814) );
  AND2_X1 U7158 ( .A1(n5488), .A2(n5814), .ZN(n9598) );
  INV_X1 U7159 ( .A(n5493), .ZN(n9817) );
  NAND2_X1 U7160 ( .A1(n5494), .A2(n5625), .ZN(n5495) );
  NAND2_X1 U7161 ( .A1(n9598), .A2(n5547), .ZN(n5505) );
  INV_X1 U7162 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5502) );
  AND2_X2 U7163 ( .A1(n5499), .A2(n5498), .ZN(n5800) );
  BUF_X2 U7164 ( .A(n5800), .Z(n8285) );
  NAND2_X1 U7165 ( .A1(n8285), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7166 ( .A1(n5594), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5500) );
  OAI211_X1 U7167 ( .C1(n5502), .C2(n5803), .A(n5501), .B(n5500), .ZN(n5503)
         );
  INV_X1 U7168 ( .A(n5503), .ZN(n5504) );
  NAND2_X1 U7169 ( .A1(n5505), .A2(n5504), .ZN(n9614) );
  XNOR2_X1 U7170 ( .A(n5506), .B(SI_16_), .ZN(n5507) );
  XNOR2_X1 U7171 ( .A(n5508), .B(n5507), .ZN(n7286) );
  NAND2_X1 U7172 ( .A1(n7286), .A2(n5867), .ZN(n5512) );
  OAI21_X1 U7173 ( .B1(n5509), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U7174 ( .A(n5510), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8076) );
  AOI22_X1 U7175 ( .A1(n8393), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5571), .B2(
        n8076), .ZN(n5511) );
  OR2_X1 U7176 ( .A1(n5738), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5513) );
  AND2_X1 U7177 ( .A1(n5765), .A2(n5513), .ZN(n9710) );
  NAND2_X1 U7178 ( .A1(n5547), .A2(n9710), .ZN(n5517) );
  INV_X2 U7179 ( .A(n5803), .ZN(n5870) );
  NAND2_X1 U7180 ( .A1(n5870), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7181 ( .A1(n8285), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7182 ( .A1(n5594), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5514) );
  OR2_X1 U7183 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  NAND2_X1 U7184 ( .A1(n5518), .A2(n5521), .ZN(n6942) );
  OR2_X1 U7185 ( .A1(n6942), .A2(n5574), .ZN(n5527) );
  NOR2_X1 U7186 ( .A1(n5522), .A2(n5625), .ZN(n5523) );
  MUX2_X1 U7187 ( .A(n5625), .B(n5523), .S(P1_IR_REG_6__SCAN_IN), .Z(n5525) );
  OR2_X1 U7188 ( .A1(n5525), .A2(n5524), .ZN(n7016) );
  INV_X1 U7189 ( .A(n7016), .ZN(n7020) );
  AOI22_X1 U7190 ( .A1(n5585), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5571), .B2(
        n7020), .ZN(n5526) );
  NAND2_X1 U7191 ( .A1(n5527), .A2(n5526), .ZN(n7534) );
  NAND2_X1 U7192 ( .A1(n5870), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5532) );
  OAI21_X1 U7193 ( .B1(n5592), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5618), .ZN(
        n5528) );
  INV_X1 U7194 ( .A(n5528), .ZN(n7537) );
  NAND2_X1 U7195 ( .A1(n5547), .A2(n7537), .ZN(n5531) );
  NAND2_X1 U7196 ( .A1(n8285), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7197 ( .A1(n5594), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5529) );
  INV_X1 U7198 ( .A(n7571), .ZN(n9424) );
  NAND2_X1 U7199 ( .A1(n5547), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7200 ( .A1(n5800), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7201 ( .A1(n5538), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7202 ( .A1(n4542), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7203 ( .A1(n5416), .A2(SI_0_), .ZN(n5537) );
  XNOR2_X1 U7204 ( .A(n5537), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9828) );
  MUX2_X1 U7205 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9828), .S(n6966), .Z(n7108) );
  NAND2_X1 U7206 ( .A1(n5964), .A2(n7108), .ZN(n7106) );
  NAND2_X1 U7207 ( .A1(n5547), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7208 ( .A1(n4542), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5540) );
  XNOR2_X1 U7209 ( .A(n5541), .B(n5542), .ZN(n6943) );
  NAND2_X1 U7210 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5543) );
  NAND2_X1 U7211 ( .A1(n5571), .A2(n9428), .ZN(n5544) );
  NAND2_X1 U7212 ( .A1(n7106), .A2(n7107), .ZN(n7105) );
  NAND2_X1 U7213 ( .A1(n7190), .A2(n8454), .ZN(n5546) );
  NAND2_X1 U7214 ( .A1(n7105), .A2(n5546), .ZN(n7348) );
  NAND2_X1 U7215 ( .A1(n5547), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7216 ( .A1(n5800), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7217 ( .A1(n5538), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7218 ( .A1(n4542), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7219 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U7220 ( .A1(n5548), .A2(n5551), .ZN(n6937) );
  NAND2_X1 U7221 ( .A1(n5585), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5554) );
  XNOR2_X1 U7222 ( .A(n5552), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U7223 ( .A1(n5571), .A2(n7098), .ZN(n5553) );
  NAND2_X1 U7224 ( .A1(n5984), .A2(n9366), .ZN(n5907) );
  NAND4_X1 U7225 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(n5560)
         );
  NAND2_X1 U7226 ( .A1(n5560), .A2(n5559), .ZN(n8457) );
  NAND2_X1 U7227 ( .A1(n7348), .A2(n8403), .ZN(n7350) );
  NAND2_X1 U7228 ( .A1(n7350), .A2(n5561), .ZN(n7228) );
  INV_X1 U7229 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U7230 ( .A1(n5547), .A2(n9855), .ZN(n5565) );
  NAND2_X1 U7231 ( .A1(n5538), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7232 ( .A1(n5800), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7233 ( .A1(n4542), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5562) );
  OR2_X1 U7234 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U7235 ( .A1(n5585), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7236 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  XNOR2_X1 U7237 ( .A(n5570), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U7238 ( .A1(n5571), .A2(n9439), .ZN(n5572) );
  NAND2_X1 U7239 ( .A1(n7342), .A2(n7235), .ZN(n8298) );
  NAND2_X1 U7240 ( .A1(n8298), .A2(n8460), .ZN(n8404) );
  NAND2_X1 U7241 ( .A1(n7228), .A2(n8404), .ZN(n7229) );
  NAND2_X1 U7242 ( .A1(n7229), .A2(n5575), .ZN(n7195) );
  NAND2_X1 U7243 ( .A1(n5538), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5580) );
  INV_X1 U7244 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5576) );
  XNOR2_X1 U7245 ( .A(n5576), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U7246 ( .A1(n5547), .A2(n7440), .ZN(n5579) );
  NAND2_X1 U7247 ( .A1(n8285), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7248 ( .A1(n4542), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5577) );
  OR2_X1 U7249 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  NAND2_X1 U7250 ( .A1(n5584), .A2(n5583), .ZN(n6934) );
  NAND2_X1 U7251 ( .A1(n5585), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5590) );
  OR2_X1 U7252 ( .A1(n5586), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7253 ( .A1(n5587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5588) );
  XNOR2_X1 U7254 ( .A(n5588), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U7255 ( .A1(n5571), .A2(n7077), .ZN(n5589) );
  NAND2_X1 U7256 ( .A1(n7279), .A2(n7198), .ZN(n8296) );
  NAND2_X1 U7257 ( .A1(n9426), .A2(n7443), .ZN(n8459) );
  NAND2_X1 U7258 ( .A1(n8296), .A2(n8459), .ZN(n8405) );
  NAND2_X1 U7259 ( .A1(n7195), .A2(n8405), .ZN(n7194) );
  NAND2_X1 U7260 ( .A1(n7194), .A2(n5591), .ZN(n7274) );
  NAND2_X1 U7261 ( .A1(n5870), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5598) );
  AOI21_X1 U7262 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5593) );
  NOR2_X1 U7263 ( .A1(n5593), .A2(n5592), .ZN(n7430) );
  NAND2_X1 U7264 ( .A1(n5547), .A2(n7430), .ZN(n5597) );
  NAND2_X1 U7265 ( .A1(n8285), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7266 ( .A1(n5594), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5595) );
  INV_X1 U7267 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  NOR2_X1 U7268 ( .A1(n5599), .A2(n5625), .ZN(n5600) );
  MUX2_X1 U7269 ( .A(n5625), .B(n5600), .S(P1_IR_REG_5__SCAN_IN), .Z(n5601) );
  OR2_X1 U7270 ( .A1(n5601), .A2(n5522), .ZN(n9452) );
  INV_X1 U7271 ( .A(n9452), .ZN(n7004) );
  AOI22_X1 U7272 ( .A1(n5585), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5571), .B2(
        n7004), .ZN(n5607) );
  OR2_X1 U7273 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U7274 ( .A1(n5602), .A2(n5605), .ZN(n6944) );
  OR2_X1 U7275 ( .A1(n6944), .A2(n5574), .ZN(n5606) );
  NAND2_X1 U7276 ( .A1(n5607), .A2(n5606), .ZN(n7283) );
  NAND2_X1 U7277 ( .A1(n7360), .A2(n7283), .ZN(n8302) );
  INV_X1 U7278 ( .A(n7283), .ZN(n7433) );
  NAND2_X1 U7279 ( .A1(n9425), .A2(n7433), .ZN(n8458) );
  NAND2_X1 U7280 ( .A1(n8302), .A2(n8458), .ZN(n7276) );
  NAND2_X1 U7281 ( .A1(n7274), .A2(n7276), .ZN(n7273) );
  NAND2_X1 U7282 ( .A1(n7273), .A2(n5608), .ZN(n7365) );
  NAND2_X1 U7283 ( .A1(n7571), .A2(n7534), .ZN(n8301) );
  INV_X1 U7284 ( .A(n7534), .ZN(n9882) );
  NAND2_X1 U7285 ( .A1(n9882), .A2(n9424), .ZN(n8304) );
  NAND2_X1 U7286 ( .A1(n8301), .A2(n8304), .ZN(n8412) );
  OAI21_X1 U7287 ( .B1(n7534), .B2(n9424), .A(n7364), .ZN(n7488) );
  OR2_X1 U7288 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U7289 ( .A1(n5609), .A2(n5612), .ZN(n6949) );
  OR2_X1 U7290 ( .A1(n6949), .A2(n5574), .ZN(n5616) );
  NAND2_X1 U7291 ( .A1(n5613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5614) );
  XNOR2_X1 U7292 ( .A(n5614), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7293 ( .A1(n8393), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5571), .B2(
        n7036), .ZN(n5615) );
  NAND2_X1 U7294 ( .A1(n5616), .A2(n5615), .ZN(n7525) );
  NAND2_X1 U7295 ( .A1(n5870), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5623) );
  AND2_X1 U7296 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NOR2_X1 U7297 ( .A1(n5629), .A2(n5619), .ZN(n7570) );
  NAND2_X1 U7298 ( .A1(n5547), .A2(n7570), .ZN(n5622) );
  NAND2_X1 U7299 ( .A1(n8285), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7300 ( .A1(n5594), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5620) );
  OR2_X1 U7301 ( .A1(n7525), .A2(n7858), .ZN(n5914) );
  NAND2_X1 U7302 ( .A1(n7525), .A2(n7858), .ZN(n7415) );
  NAND2_X1 U7303 ( .A1(n5914), .A2(n7415), .ZN(n8313) );
  NAND2_X1 U7304 ( .A1(n7488), .A2(n8313), .ZN(n7487) );
  INV_X1 U7305 ( .A(n7858), .ZN(n9423) );
  NAND2_X1 U7306 ( .A1(n7487), .A2(n5624), .ZN(n7421) );
  XNOR2_X1 U7307 ( .A(n5638), .B(n5637), .ZN(n6950) );
  NOR2_X1 U7308 ( .A1(n5613), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5658) );
  OR2_X1 U7309 ( .A1(n5658), .A2(n5625), .ZN(n5626) );
  INV_X1 U7310 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U7311 ( .A1(n5626), .A2(n10382), .ZN(n5641) );
  OR2_X1 U7312 ( .A1(n5626), .A2(n10382), .ZN(n5627) );
  AOI22_X1 U7313 ( .A1(n8393), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5571), .B2(
        n7062), .ZN(n5628) );
  OR2_X1 U7314 ( .A1(n5629), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5630) );
  AND2_X1 U7315 ( .A1(n5646), .A2(n5630), .ZN(n7857) );
  NAND2_X1 U7316 ( .A1(n5547), .A2(n7857), .ZN(n5634) );
  NAND2_X1 U7317 ( .A1(n5870), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7318 ( .A1(n8285), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7319 ( .A1(n5594), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7320 ( .A1(n7863), .A2(n7873), .ZN(n8319) );
  NAND2_X1 U7321 ( .A1(n8314), .A2(n8319), .ZN(n7420) );
  NAND2_X1 U7322 ( .A1(n7421), .A2(n7420), .ZN(n7419) );
  INV_X1 U7323 ( .A(n7873), .ZN(n9422) );
  NAND2_X1 U7324 ( .A1(n7419), .A2(n5635), .ZN(n7473) );
  XNOR2_X1 U7325 ( .A(n5640), .B(n5639), .ZN(n6958) );
  NAND2_X1 U7326 ( .A1(n6958), .A2(n5867), .ZN(n5644) );
  NAND2_X1 U7327 ( .A1(n5641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5642) );
  XNOR2_X1 U7328 ( .A(n5642), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7120) );
  AOI22_X1 U7329 ( .A1(n8393), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5571), .B2(
        n7120), .ZN(n5643) );
  NAND2_X1 U7330 ( .A1(n5644), .A2(n5643), .ZN(n7480) );
  NAND2_X1 U7331 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  AND2_X1 U7332 ( .A1(n5664), .A2(n5647), .ZN(n7477) );
  NAND2_X1 U7333 ( .A1(n5547), .A2(n7477), .ZN(n5651) );
  NAND2_X1 U7334 ( .A1(n5870), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7335 ( .A1(n8285), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7336 ( .A1(n5594), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7337 ( .A1(n7480), .A2(n9265), .ZN(n8320) );
  NAND2_X1 U7338 ( .A1(n8416), .A2(n8320), .ZN(n7472) );
  INV_X1 U7339 ( .A(n9265), .ZN(n7862) );
  NAND2_X1 U7340 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NAND2_X1 U7341 ( .A1(n5656), .A2(n5655), .ZN(n6962) );
  OR2_X1 U7342 ( .A1(n6962), .A2(n5574), .ZN(n5663) );
  NOR2_X1 U7343 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5657) );
  NAND2_X1 U7344 ( .A1(n5658), .A2(n5657), .ZN(n5660) );
  NAND2_X1 U7345 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5659) );
  MUX2_X1 U7346 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5659), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5661) );
  AOI22_X1 U7347 ( .A1(n8393), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5571), .B2(
        n7219), .ZN(n5662) );
  NAND2_X1 U7348 ( .A1(n5663), .A2(n5662), .ZN(n7613) );
  NAND2_X1 U7349 ( .A1(n5870), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7350 ( .A1(n5664), .A2(n7123), .ZN(n5665) );
  AND2_X1 U7351 ( .A1(n5678), .A2(n5665), .ZN(n7606) );
  NAND2_X1 U7352 ( .A1(n5547), .A2(n7606), .ZN(n5668) );
  NAND2_X1 U7353 ( .A1(n8285), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7354 ( .A1(n5594), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5666) );
  OR2_X1 U7355 ( .A1(n7613), .A2(n9353), .ZN(n8463) );
  NAND2_X1 U7356 ( .A1(n7613), .A2(n9353), .ZN(n8322) );
  NAND2_X1 U7357 ( .A1(n8463), .A2(n8322), .ZN(n8419) );
  INV_X1 U7358 ( .A(n9353), .ZN(n9421) );
  XNOR2_X1 U7359 ( .A(n5672), .B(n5671), .ZN(n6976) );
  NAND2_X1 U7360 ( .A1(n6976), .A2(n5867), .ZN(n5675) );
  NAND2_X1 U7361 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U7362 ( .A(n5673), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7375) );
  AOI22_X1 U7363 ( .A1(n8393), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5571), .B2(
        n7375), .ZN(n5674) );
  NOR2_X1 U7364 ( .A1(n5695), .A2(n5077), .ZN(n9352) );
  NAND2_X1 U7365 ( .A1(n5547), .A2(n9352), .ZN(n5682) );
  NAND2_X1 U7366 ( .A1(n5870), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7367 ( .A1(n8285), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7368 ( .A1(n5594), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5679) );
  OR2_X1 U7369 ( .A1(n9358), .A2(n7809), .ZN(n8324) );
  NAND2_X1 U7370 ( .A1(n9358), .A2(n7809), .ZN(n8325) );
  NAND2_X1 U7371 ( .A1(n8324), .A2(n8325), .ZN(n7657) );
  NAND2_X1 U7372 ( .A1(n7656), .A2(n7657), .ZN(n7655) );
  INV_X1 U7373 ( .A(n7809), .ZN(n9420) );
  NAND2_X1 U7374 ( .A1(n7655), .A2(n5683), .ZN(n7814) );
  NAND2_X1 U7375 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U7376 ( .A1(n5687), .A2(n5686), .ZN(n7048) );
  OR2_X1 U7377 ( .A1(n7048), .A2(n5574), .ZN(n5694) );
  NAND2_X1 U7378 ( .A1(n5689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7379 ( .A1(n5691), .A2(n5690), .ZN(n5705) );
  OR2_X1 U7380 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  AOI22_X1 U7381 ( .A1(n8393), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5571), .B2(
        n7381), .ZN(n5693) );
  NAND2_X1 U7382 ( .A1(n5870), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7383 ( .A1(n8285), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5699) );
  OR2_X1 U7384 ( .A1(n5695), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5696) );
  AND2_X1 U7385 ( .A1(n5696), .A2(n5710), .ZN(n8055) );
  NAND2_X1 U7386 ( .A1(n5547), .A2(n8055), .ZN(n5698) );
  NAND2_X1 U7387 ( .A1(n5594), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5697) );
  NAND4_X1 U7388 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n9419)
         );
  NAND2_X1 U7389 ( .A1(n9907), .A2(n9419), .ZN(n8328) );
  INV_X1 U7390 ( .A(n9419), .ZN(n6063) );
  NAND2_X1 U7391 ( .A1(n8058), .A2(n6063), .ZN(n8470) );
  NAND2_X1 U7392 ( .A1(n8328), .A2(n8470), .ZN(n7813) );
  NAND2_X1 U7393 ( .A1(n7814), .A2(n7813), .ZN(n7812) );
  NAND2_X1 U7394 ( .A1(n7812), .A2(n5701), .ZN(n7894) );
  XNOR2_X1 U7395 ( .A(n5702), .B(SI_13_), .ZN(n5703) );
  NAND2_X1 U7396 ( .A1(n7137), .A2(n5867), .ZN(n5708) );
  NAND2_X1 U7397 ( .A1(n5705), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U7398 ( .A(n5706), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7731) );
  AOI22_X1 U7399 ( .A1(n7731), .A2(n5571), .B1(n8393), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7400 ( .A1(n5710), .A2(n5709), .ZN(n5711) );
  AND2_X1 U7401 ( .A1(n5722), .A2(n5711), .ZN(n8143) );
  NAND2_X1 U7402 ( .A1(n5547), .A2(n8143), .ZN(n5715) );
  NAND2_X1 U7403 ( .A1(n5870), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7404 ( .A1(n8285), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7405 ( .A1(n5594), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5712) );
  OR2_X1 U7406 ( .A1(n8147), .A2(n9242), .ZN(n8335) );
  NAND2_X1 U7407 ( .A1(n8147), .A2(n9242), .ZN(n8474) );
  NAND2_X1 U7408 ( .A1(n8335), .A2(n8474), .ZN(n8423) );
  INV_X1 U7409 ( .A(n9242), .ZN(n9418) );
  XNOR2_X1 U7410 ( .A(n5718), .B(n5717), .ZN(n7177) );
  NAND2_X1 U7411 ( .A1(n7177), .A2(n5867), .ZN(n5721) );
  XNOR2_X1 U7412 ( .A(n5719), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7841) );
  AOI22_X1 U7413 ( .A1(n8393), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5571), .B2(
        n7841), .ZN(n5720) );
  NAND2_X1 U7414 ( .A1(n5870), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5727) );
  AND2_X1 U7415 ( .A1(n5722), .A2(n7729), .ZN(n5723) );
  NOR2_X1 U7416 ( .A1(n5736), .A2(n5723), .ZN(n9241) );
  NAND2_X1 U7417 ( .A1(n5547), .A2(n9241), .ZN(n5726) );
  NAND2_X1 U7418 ( .A1(n8285), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7419 ( .A1(n5594), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5724) );
  XNOR2_X1 U7420 ( .A(n5730), .B(n5729), .ZN(n5731) );
  XNOR2_X1 U7421 ( .A(n5732), .B(n5731), .ZN(n7226) );
  NAND2_X1 U7422 ( .A1(n7226), .A2(n5867), .ZN(n5735) );
  INV_X1 U7423 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U7424 ( .A(n5509), .B(n5733), .ZN(n7848) );
  AOI22_X1 U7425 ( .A1(n8393), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5571), .B2(
        n7848), .ZN(n5734) );
  NOR2_X1 U7426 ( .A1(n5736), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5737) );
  OR2_X1 U7427 ( .A1(n5738), .A2(n5737), .ZN(n8199) );
  INV_X1 U7428 ( .A(n8199), .ZN(n9392) );
  NAND2_X1 U7429 ( .A1(n5547), .A2(n9392), .ZN(n5742) );
  NAND2_X1 U7430 ( .A1(n8285), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7431 ( .A1(n5870), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7432 ( .A1(n5594), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7433 ( .A1(n9832), .A2(n9307), .ZN(n5743) );
  OR2_X1 U7434 ( .A1(n9709), .A2(n9685), .ZN(n8341) );
  NAND2_X1 U7435 ( .A1(n9709), .A2(n9685), .ZN(n9678) );
  XNOR2_X1 U7436 ( .A(n5746), .B(n5745), .ZN(n7411) );
  NAND2_X1 U7437 ( .A1(n7411), .A2(n5867), .ZN(n5751) );
  OR2_X1 U7438 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5747) );
  AND2_X1 U7439 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5747), .ZN(n5748) );
  OR2_X1 U7440 ( .A1(n5509), .A2(n5748), .ZN(n5749) );
  INV_X1 U7441 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10318) );
  XNOR2_X1 U7442 ( .A(n5749), .B(n10318), .ZN(n8261) );
  AOI22_X1 U7443 ( .A1(n8393), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5571), .B2(
        n8261), .ZN(n5750) );
  NAND2_X1 U7444 ( .A1(n5800), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U7445 ( .A(n5765), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U7446 ( .A1(n5547), .A2(n9675), .ZN(n5754) );
  NAND2_X1 U7447 ( .A1(n5870), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7448 ( .A1(n5594), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5752) );
  NAND4_X1 U7449 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n9699)
         );
  NOR2_X1 U7450 ( .A1(n9770), .A2(n9699), .ZN(n5756) );
  INV_X1 U7451 ( .A(n9770), .ZN(n9677) );
  XNOR2_X1 U7452 ( .A(n5758), .B(n5757), .ZN(n7564) );
  NAND2_X1 U7453 ( .A1(n7564), .A2(n5867), .ZN(n5762) );
  XNOR2_X1 U7454 ( .A(n5759), .B(n5760), .ZN(n8262) );
  AOI22_X1 U7455 ( .A1(n8393), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5571), .B2(
        n8262), .ZN(n5761) );
  INV_X1 U7456 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5764) );
  INV_X1 U7457 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5763) );
  OAI21_X1 U7458 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5766) );
  AND2_X1 U7459 ( .A1(n5766), .A2(n5777), .ZN(n9665) );
  NAND2_X1 U7460 ( .A1(n9665), .A2(n5547), .ZN(n5770) );
  NAND2_X1 U7461 ( .A1(n5870), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7462 ( .A1(n8285), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7463 ( .A1(n5594), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7464 ( .A1(n9668), .A2(n9687), .ZN(n5771) );
  INV_X1 U7465 ( .A(n9687), .ZN(n9415) );
  XNOR2_X1 U7466 ( .A(n5773), .B(n5772), .ZN(n7650) );
  NAND2_X1 U7467 ( .A1(n7650), .A2(n5867), .ZN(n5776) );
  AOI22_X1 U7468 ( .A1(n8393), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5457), .B2(
        n5571), .ZN(n5775) );
  AND2_X1 U7469 ( .A1(n5777), .A2(n8272), .ZN(n5778) );
  OR2_X1 U7470 ( .A1(n5778), .A2(n5786), .ZN(n9649) );
  AOI22_X1 U7471 ( .A1(n5870), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8285), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7472 ( .A1(n5594), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5779) );
  OAI211_X1 U7473 ( .C1(n9649), .C2(n5790), .A(n5780), .B(n5779), .ZN(n9414)
         );
  NAND2_X1 U7474 ( .A1(n9761), .A2(n9414), .ZN(n5781) );
  XNOR2_X1 U7475 ( .A(n5783), .B(n10483), .ZN(n5784) );
  XNOR2_X1 U7476 ( .A(n5782), .B(n5784), .ZN(n7802) );
  NAND2_X1 U7477 ( .A1(n8393), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U7478 ( .A1(n5786), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5787) );
  OR2_X1 U7479 ( .A1(n5797), .A2(n5787), .ZN(n9633) );
  INV_X1 U7480 ( .A(n5547), .ZN(n5790) );
  AOI22_X1 U7481 ( .A1(n5870), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n8285), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7482 ( .A1(n5594), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5788) );
  OAI211_X1 U7483 ( .C1(n9633), .C2(n5790), .A(n5789), .B(n5788), .ZN(n9613)
         );
  INV_X1 U7484 ( .A(n9613), .ZN(n9645) );
  NAND2_X1 U7485 ( .A1(n9637), .A2(n9645), .ZN(n5791) );
  XNOR2_X1 U7486 ( .A(n5792), .B(SI_21_), .ZN(n5793) );
  XNOR2_X1 U7487 ( .A(n5794), .B(n5793), .ZN(n7867) );
  NAND2_X1 U7488 ( .A1(n7867), .A2(n5867), .ZN(n5796) );
  NAND2_X1 U7489 ( .A1(n8393), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5795) );
  NOR2_X1 U7490 ( .A1(n5797), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5798) );
  OR2_X1 U7491 ( .A1(n5799), .A2(n5798), .ZN(n9619) );
  INV_X1 U7492 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U7493 ( .A1(n5800), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7494 ( .A1(n5594), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5801) );
  OAI211_X1 U7495 ( .C1(n9752), .C2(n5803), .A(n5802), .B(n5801), .ZN(n5804)
         );
  INV_X1 U7496 ( .A(n5804), .ZN(n5805) );
  OAI21_X1 U7497 ( .B1(n9619), .B2(n5790), .A(n5805), .ZN(n9604) );
  NAND2_X1 U7498 ( .A1(n9618), .A2(n9604), .ZN(n5806) );
  INV_X1 U7499 ( .A(n9604), .ZN(n9630) );
  OR2_X1 U7500 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  NAND2_X1 U7501 ( .A1(n5812), .A2(n5811), .ZN(n8013) );
  NAND2_X1 U7502 ( .A1(n8393), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7503 ( .A1(n5870), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5820) );
  INV_X1 U7504 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U7505 ( .A1(n9252), .A2(n5814), .ZN(n5816) );
  INV_X1 U7506 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U7507 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n5815), .ZN(n5828) );
  AND2_X1 U7508 ( .A1(n5816), .A2(n5828), .ZN(n9587) );
  NAND2_X1 U7509 ( .A1(n5547), .A2(n9587), .ZN(n5819) );
  NAND2_X1 U7510 ( .A1(n8285), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7511 ( .A1(n5594), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5817) );
  NOR2_X1 U7512 ( .A1(n9590), .A2(n9576), .ZN(n5821) );
  XNOR2_X1 U7513 ( .A(n5823), .B(n5822), .ZN(n8137) );
  NAND2_X1 U7514 ( .A1(n8137), .A2(n5867), .ZN(n5825) );
  NAND2_X1 U7515 ( .A1(n8393), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7516 ( .A1(n8285), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7517 ( .A1(n5870), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5832) );
  INV_X1 U7518 ( .A(n5828), .ZN(n5826) );
  NAND2_X1 U7519 ( .A1(n5826), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5839) );
  INV_X1 U7520 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7521 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  AND2_X1 U7522 ( .A1(n5839), .A2(n5829), .ZN(n9579) );
  NAND2_X1 U7523 ( .A1(n5547), .A2(n9579), .ZN(n5831) );
  NAND2_X1 U7524 ( .A1(n5594), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7525 ( .A1(n9741), .A2(n9553), .ZN(n8447) );
  INV_X1 U7526 ( .A(n9553), .ZN(n9413) );
  NAND2_X1 U7527 ( .A1(n8223), .A2(n5867), .ZN(n5836) );
  NAND2_X1 U7528 ( .A1(n8393), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7529 ( .A1(n5870), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7530 ( .A1(n8285), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5843) );
  INV_X1 U7531 ( .A(n5839), .ZN(n5837) );
  NAND2_X1 U7532 ( .A1(n5837), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5854) );
  INV_X1 U7533 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7534 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AND2_X1 U7535 ( .A1(n5854), .A2(n5840), .ZN(n9563) );
  NAND2_X1 U7536 ( .A1(n5547), .A2(n9563), .ZN(n5842) );
  NAND2_X1 U7537 ( .A1(n5594), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5841) );
  NAND4_X1 U7538 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n9544)
         );
  NAND2_X1 U7539 ( .A1(n9562), .A2(n9544), .ZN(n5845) );
  OAI21_X2 U7540 ( .B1(n5847), .B2(n5846), .A(n5845), .ZN(n9537) );
  NAND2_X1 U7541 ( .A1(n8231), .A2(n5867), .ZN(n5851) );
  NAND2_X1 U7542 ( .A1(n8393), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7543 ( .A1(n5870), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7544 ( .A1(n5800), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5858) );
  INV_X1 U7545 ( .A(n5854), .ZN(n5852) );
  NAND2_X1 U7546 ( .A1(n5852), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5873) );
  INV_X1 U7547 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7548 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  AND2_X1 U7549 ( .A1(n5873), .A2(n5855), .ZN(n9538) );
  NAND2_X1 U7550 ( .A1(n5547), .A2(n9538), .ZN(n5857) );
  NAND2_X1 U7551 ( .A1(n5594), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7552 ( .A1(n9730), .A2(n9554), .ZN(n8509) );
  NAND2_X1 U7553 ( .A1(n8490), .A2(n8509), .ZN(n9536) );
  NAND2_X1 U7554 ( .A1(n9537), .A2(n9536), .ZN(n5861) );
  INV_X1 U7555 ( .A(n9554), .ZN(n9412) );
  NAND2_X1 U7556 ( .A1(n9730), .A2(n9412), .ZN(n5860) );
  AND2_X1 U7557 ( .A1(n5864), .A2(n5879), .ZN(n5865) );
  NAND2_X1 U7558 ( .A1(n8236), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U7559 ( .A1(n8393), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7560 ( .A1(n8285), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7561 ( .A1(n5870), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5877) );
  INV_X1 U7562 ( .A(n5873), .ZN(n5871) );
  NAND2_X1 U7563 ( .A1(n5871), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5887) );
  INV_X1 U7564 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7565 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  NAND2_X1 U7566 ( .A1(n5547), .A2(n9530), .ZN(n5876) );
  NAND2_X1 U7567 ( .A1(n5594), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7568 ( .A1(n9529), .A2(n6150), .ZN(n8289) );
  NAND2_X1 U7569 ( .A1(n8593), .A2(n5867), .ZN(n5884) );
  NAND2_X1 U7570 ( .A1(n8393), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7571 ( .A1(n5870), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5892) );
  INV_X1 U7572 ( .A(n5887), .ZN(n5885) );
  NAND2_X1 U7573 ( .A1(n5885), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9489) );
  INV_X1 U7574 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7575 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  NAND2_X1 U7576 ( .A1(n5547), .A2(n9505), .ZN(n5891) );
  NAND2_X1 U7577 ( .A1(n5800), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7578 ( .A1(n5594), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7579 ( .A1(n9720), .A2(n9520), .ZN(n8290) );
  INV_X1 U7580 ( .A(n9520), .ZN(n9411) );
  NAND2_X1 U7581 ( .A1(n9720), .A2(n9411), .ZN(n5894) );
  NAND2_X1 U7582 ( .A1(n9501), .A2(n5894), .ZN(n5900) );
  NAND2_X1 U7583 ( .A1(n5870), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5899) );
  INV_X1 U7584 ( .A(n9489), .ZN(n5895) );
  NAND2_X1 U7585 ( .A1(n5547), .A2(n5895), .ZN(n5898) );
  NAND2_X1 U7586 ( .A1(n5800), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7587 ( .A1(n5594), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5896) );
  OR2_X1 U7588 ( .A1(n9493), .A2(n6182), .ZN(n8496) );
  NAND2_X1 U7589 ( .A1(n9493), .A2(n6182), .ZN(n8499) );
  XNOR2_X1 U7590 ( .A(n5900), .B(n8434), .ZN(n9498) );
  INV_X1 U7591 ( .A(n5945), .ZN(n8530) );
  NAND2_X1 U7592 ( .A1(n8530), .A2(n8523), .ZN(n6179) );
  INV_X1 U7593 ( .A(n7331), .ZN(n5903) );
  NAND2_X1 U7594 ( .A1(n5945), .A2(n5948), .ZN(n5902) );
  NAND3_X1 U7595 ( .A1(n6179), .A2(n5903), .A3(n5902), .ZN(n7346) );
  INV_X1 U7596 ( .A(n7114), .ZN(n5904) );
  INV_X1 U7597 ( .A(n7108), .ZN(n7337) );
  NOR2_X1 U7598 ( .A1(n5964), .A2(n7337), .ZN(n7109) );
  NAND2_X1 U7599 ( .A1(n7190), .A2(n7185), .ZN(n5905) );
  NAND2_X1 U7600 ( .A1(n7340), .A2(n8457), .ZN(n5906) );
  NAND2_X1 U7601 ( .A1(n8293), .A2(n8298), .ZN(n8295) );
  INV_X1 U7602 ( .A(n8296), .ZN(n5908) );
  NAND2_X1 U7603 ( .A1(n7277), .A2(n8302), .ZN(n5910) );
  NAND2_X1 U7604 ( .A1(n5910), .A2(n8458), .ZN(n7358) );
  INV_X1 U7605 ( .A(n7414), .ZN(n5913) );
  NAND2_X1 U7606 ( .A1(n8319), .A2(n7415), .ZN(n8310) );
  NAND3_X1 U7607 ( .A1(n8416), .A2(n8310), .A3(n8314), .ZN(n5911) );
  NAND2_X1 U7608 ( .A1(n5911), .A2(n8320), .ZN(n8418) );
  AND3_X1 U7609 ( .A1(n8416), .A2(n4530), .A3(n8304), .ZN(n5915) );
  OR2_X1 U7610 ( .A1(n8418), .A2(n5915), .ZN(n8462) );
  INV_X1 U7611 ( .A(n8419), .ZN(n7601) );
  INV_X1 U7612 ( .A(n8324), .ZN(n5916) );
  INV_X1 U7613 ( .A(n7813), .ZN(n8421) );
  NAND2_X1 U7614 ( .A1(n7808), .A2(n8421), .ZN(n7807) );
  NAND2_X1 U7615 ( .A1(n7807), .A2(n8470), .ZN(n7895) );
  NAND2_X1 U7616 ( .A1(n9783), .A2(n9397), .ZN(n8338) );
  OR2_X1 U7617 ( .A1(n9408), .A2(n9307), .ZN(n8479) );
  NAND2_X1 U7618 ( .A1(n9408), .A2(n9307), .ZN(n8339) );
  NAND2_X1 U7619 ( .A1(n9695), .A2(n9704), .ZN(n9694) );
  OR2_X1 U7620 ( .A1(n9770), .A2(n9662), .ZN(n8480) );
  NAND2_X1 U7621 ( .A1(n9770), .A2(n9662), .ZN(n8347) );
  NAND2_X1 U7622 ( .A1(n8480), .A2(n8347), .ZN(n9683) );
  INV_X1 U7623 ( .A(n9678), .ZN(n8477) );
  NOR2_X1 U7624 ( .A1(n9683), .A2(n8477), .ZN(n5918) );
  NAND2_X1 U7625 ( .A1(n9694), .A2(n5918), .ZN(n9679) );
  OR2_X1 U7626 ( .A1(n9766), .A2(n9687), .ZN(n8348) );
  NAND2_X1 U7627 ( .A1(n9766), .A2(n9687), .ZN(n8349) );
  NAND2_X1 U7628 ( .A1(n8348), .A2(n8349), .ZN(n9660) );
  OR2_X1 U7629 ( .A1(n9761), .A2(n9663), .ZN(n8354) );
  NAND2_X1 U7630 ( .A1(n9761), .A2(n9663), .ZN(n8492) );
  NAND2_X1 U7631 ( .A1(n8354), .A2(n8492), .ZN(n9642) );
  NAND2_X1 U7632 ( .A1(n9756), .A2(n9645), .ZN(n8360) );
  INV_X1 U7633 ( .A(n8359), .ZN(n8357) );
  OR2_X1 U7634 ( .A1(n9618), .A2(n9630), .ZN(n8442) );
  NAND2_X1 U7635 ( .A1(n9618), .A2(n9630), .ZN(n8366) );
  OR2_X1 U7636 ( .A1(n9745), .A2(n9290), .ZN(n8370) );
  NAND2_X1 U7637 ( .A1(n9745), .A2(n9290), .ZN(n8369) );
  NAND2_X1 U7638 ( .A1(n9256), .A2(n9576), .ZN(n9570) );
  INV_X1 U7639 ( .A(n9570), .ZN(n8367) );
  NOR2_X1 U7640 ( .A1(n9572), .A2(n8367), .ZN(n5920) );
  INV_X1 U7641 ( .A(n9544), .ZN(n9575) );
  OR2_X1 U7642 ( .A1(n9562), .A2(n9575), .ZN(n8441) );
  NAND2_X1 U7643 ( .A1(n9562), .A2(n9575), .ZN(n8448) );
  NAND2_X1 U7644 ( .A1(n8441), .A2(n8448), .ZN(n9558) );
  INV_X1 U7645 ( .A(n9536), .ZN(n9543) );
  NAND2_X1 U7646 ( .A1(n9542), .A2(n9543), .ZN(n9541) );
  NAND2_X1 U7647 ( .A1(n9541), .A2(n8509), .ZN(n9518) );
  NAND2_X1 U7648 ( .A1(n9518), .A2(n9525), .ZN(n9517) );
  NAND2_X1 U7649 ( .A1(n5457), .A2(n8537), .ZN(n5921) );
  NAND2_X1 U7650 ( .A1(n5944), .A2(n8503), .ZN(n8505) );
  INV_X1 U7651 ( .A(n5922), .ZN(n7081) );
  NAND2_X1 U7652 ( .A1(n5870), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7653 ( .A1(n5594), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7654 ( .A1(n8285), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5923) );
  INV_X1 U7655 ( .A(n5926), .ZN(n6987) );
  NAND2_X1 U7656 ( .A1(n6987), .A2(P1_B_REG_SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7657 ( .A1(n9698), .A2(n5927), .ZN(n8581) );
  OAI22_X1 U7658 ( .A1(n9520), .A2(n9684), .B1(n8432), .B2(n8581), .ZN(n5928)
         );
  AND2_X1 U7659 ( .A1(n7351), .A2(n5559), .ZN(n7352) );
  NAND2_X1 U7660 ( .A1(n7352), .A2(n9860), .ZN(n7230) );
  INV_X1 U7661 ( .A(n7525), .ZN(n7577) );
  OR2_X1 U7662 ( .A1(n7474), .A2(n7480), .ZN(n7608) );
  INV_X1 U7663 ( .A(n9358), .ZN(n7717) );
  OR2_X2 U7664 ( .A1(n9770), .A2(n9705), .ZN(n9673) );
  AOI21_X1 U7665 ( .B1(n9493), .B2(n9503), .A(n9707), .ZN(n5930) );
  NAND2_X1 U7666 ( .A1(n5930), .A2(n9482), .ZN(n9496) );
  NAND2_X1 U7667 ( .A1(n5932), .A2(n5931), .ZN(P1_U3551) );
  INV_X1 U7668 ( .A(n5933), .ZN(n5937) );
  INV_X1 U7669 ( .A(n5934), .ZN(n7323) );
  NAND2_X1 U7670 ( .A1(n9874), .A2(n7323), .ZN(n5935) );
  NOR2_X1 U7671 ( .A1(n7326), .A2(n5935), .ZN(n5936) );
  INV_X1 U7672 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5940) );
  NOR2_X1 U7673 ( .A1(n9913), .A2(n5940), .ZN(n5941) );
  NAND2_X1 U7674 ( .A1(n5945), .A2(n5950), .ZN(n5946) );
  NAND2_X1 U7675 ( .A1(n5946), .A2(n5948), .ZN(n5947) );
  NAND2_X1 U7676 ( .A1(n9618), .A2(n6157), .ZN(n5953) );
  NAND2_X1 U7677 ( .A1(n9604), .A2(n5972), .ZN(n5952) );
  NAND2_X1 U7678 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  XNOR2_X1 U7679 ( .A(n5954), .B(n6131), .ZN(n9286) );
  INV_X1 U7680 ( .A(n9286), .ZN(n6119) );
  AND2_X1 U7681 ( .A1(n9604), .A2(n6125), .ZN(n5955) );
  AOI21_X1 U7682 ( .B1(n9618), .B2(n5972), .A(n5955), .ZN(n9285) );
  INV_X1 U7683 ( .A(n9285), .ZN(n6118) );
  AOI22_X1 U7684 ( .A1(n9709), .A2(n6157), .B1(n5972), .B2(n9416), .ZN(n5956)
         );
  OAI22_X1 U7685 ( .A1(n7279), .A2(n6158), .B1(n7443), .B2(n5982), .ZN(n5957)
         );
  XNOR2_X1 U7686 ( .A(n5957), .B(n6131), .ZN(n5996) );
  OR2_X1 U7687 ( .A1(n7279), .A2(n6163), .ZN(n5959) );
  NAND2_X1 U7688 ( .A1(n5972), .A2(n7198), .ZN(n5958) );
  NAND2_X1 U7689 ( .A1(n5959), .A2(n5958), .ZN(n5997) );
  XNOR2_X1 U7690 ( .A(n5996), .B(n5997), .ZN(n7169) );
  OAI22_X1 U7691 ( .A1(n7342), .A2(n6158), .B1(n9860), .B2(n5982), .ZN(n5960)
         );
  XNOR2_X1 U7692 ( .A(n5960), .B(n6131), .ZN(n5994) );
  OR2_X1 U7693 ( .A1(n7342), .A2(n6163), .ZN(n5962) );
  NAND2_X1 U7694 ( .A1(n5972), .A2(n7235), .ZN(n5961) );
  NAND2_X1 U7695 ( .A1(n5962), .A2(n5961), .ZN(n5993) );
  INV_X1 U7696 ( .A(n5993), .ZN(n5963) );
  NAND2_X1 U7697 ( .A1(n5994), .A2(n5963), .ZN(n7170) );
  AND2_X1 U7698 ( .A1(n7169), .A2(n7170), .ZN(n5995) );
  NAND2_X1 U7699 ( .A1(n5964), .A2(n5972), .ZN(n5965) );
  NAND2_X1 U7700 ( .A1(n5968), .A2(n6131), .ZN(n5971) );
  INV_X1 U7701 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5966) );
  OR2_X1 U7702 ( .A1(n5951), .A2(n5966), .ZN(n5967) );
  NAND2_X1 U7703 ( .A1(n5968), .A2(n5967), .ZN(n7080) );
  NAND2_X1 U7704 ( .A1(n5964), .A2(n6125), .ZN(n5970) );
  INV_X1 U7705 ( .A(n5951), .ZN(n6891) );
  AOI22_X1 U7706 ( .A1(n5972), .A2(n7108), .B1(n6891), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7707 ( .A1(n5970), .A2(n5969), .ZN(n7079) );
  NAND2_X1 U7708 ( .A1(n7080), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U7709 ( .A1(n5545), .A2(n5972), .ZN(n5973) );
  NAND2_X1 U7710 ( .A1(n5545), .A2(n6125), .ZN(n5976) );
  OR2_X1 U7711 ( .A1(n8454), .A2(n6158), .ZN(n5975) );
  NAND2_X1 U7712 ( .A1(n5976), .A2(n5975), .ZN(n5978) );
  NAND2_X1 U7713 ( .A1(n5977), .A2(n5978), .ZN(n7182) );
  NAND2_X1 U7714 ( .A1(n7181), .A2(n7182), .ZN(n5981) );
  INV_X1 U7715 ( .A(n5977), .ZN(n5980) );
  INV_X1 U7716 ( .A(n5978), .ZN(n5979) );
  NAND2_X1 U7717 ( .A1(n5980), .A2(n5979), .ZN(n7183) );
  OAI22_X1 U7718 ( .A1(n5982), .A2(n5559), .B1(n5984), .B2(n6158), .ZN(n5983)
         );
  XNOR2_X1 U7719 ( .A(n5983), .B(n6131), .ZN(n5990) );
  INV_X1 U7720 ( .A(n5990), .ZN(n5987) );
  OR2_X1 U7721 ( .A1(n5984), .A2(n6163), .ZN(n5986) );
  NAND2_X1 U7722 ( .A1(n5972), .A2(n9366), .ZN(n5985) );
  NAND2_X1 U7723 ( .A1(n5986), .A2(n5985), .ZN(n5988) );
  NAND2_X1 U7724 ( .A1(n5987), .A2(n5988), .ZN(n5991) );
  INV_X1 U7725 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7726 ( .A1(n5990), .A2(n5989), .ZN(n5992) );
  AND2_X1 U7727 ( .A1(n5991), .A2(n5992), .ZN(n9364) );
  NAND2_X1 U7728 ( .A1(n9363), .A2(n9364), .ZN(n9362) );
  NAND2_X1 U7729 ( .A1(n9362), .A2(n5992), .ZN(n7204) );
  XNOR2_X1 U7730 ( .A(n5994), .B(n5993), .ZN(n7205) );
  INV_X1 U7731 ( .A(n5996), .ZN(n5998) );
  NAND2_X1 U7732 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  OAI22_X1 U7733 ( .A1(n7360), .A2(n6158), .B1(n7433), .B2(n5982), .ZN(n6000)
         );
  XNOR2_X1 U7734 ( .A(n6000), .B(n6161), .ZN(n6002) );
  INV_X1 U7735 ( .A(n6002), .ZN(n6001) );
  OR2_X1 U7736 ( .A1(n7360), .A2(n6163), .ZN(n6005) );
  NAND2_X1 U7737 ( .A1(n7283), .A2(n5972), .ZN(n6004) );
  NAND2_X1 U7738 ( .A1(n6005), .A2(n6004), .ZN(n7406) );
  NAND2_X1 U7739 ( .A1(n7534), .A2(n6157), .ZN(n6007) );
  OAI21_X1 U7740 ( .B1(n7571), .B2(n6158), .A(n6007), .ZN(n6008) );
  XNOR2_X1 U7741 ( .A(n6008), .B(n6131), .ZN(n6011) );
  OR2_X1 U7742 ( .A1(n7571), .A2(n6163), .ZN(n6010) );
  NAND2_X1 U7743 ( .A1(n7534), .A2(n5972), .ZN(n6009) );
  AND2_X1 U7744 ( .A1(n6010), .A2(n6009), .ZN(n6012) );
  NAND2_X1 U7745 ( .A1(n6011), .A2(n6012), .ZN(n6017) );
  INV_X1 U7746 ( .A(n6011), .ZN(n6014) );
  INV_X1 U7747 ( .A(n6012), .ZN(n6013) );
  NAND2_X1 U7748 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  AND2_X1 U7749 ( .A1(n6017), .A2(n6015), .ZN(n7529) );
  NAND2_X1 U7750 ( .A1(n6016), .A2(n7529), .ZN(n7531) );
  NAND2_X1 U7751 ( .A1(n7531), .A2(n6017), .ZN(n7566) );
  NAND2_X1 U7752 ( .A1(n7525), .A2(n6157), .ZN(n6019) );
  OR2_X1 U7753 ( .A1(n7858), .A2(n6158), .ZN(n6018) );
  NAND2_X1 U7754 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  XNOR2_X1 U7755 ( .A(n6020), .B(n6161), .ZN(n6021) );
  AOI22_X1 U7756 ( .A1(n7525), .A2(n5972), .B1(n9423), .B2(n6125), .ZN(n6022)
         );
  XNOR2_X1 U7757 ( .A(n6021), .B(n6022), .ZN(n7568) );
  INV_X1 U7758 ( .A(n6021), .ZN(n6023) );
  NAND2_X1 U7759 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  NAND2_X1 U7760 ( .A1(n7863), .A2(n6157), .ZN(n6026) );
  OR2_X1 U7761 ( .A1(n7873), .A2(n6158), .ZN(n6025) );
  NAND2_X1 U7762 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7763 ( .A(n6027), .B(n6131), .ZN(n6028) );
  NAND2_X1 U7764 ( .A1(n6029), .A2(n6028), .ZN(n6034) );
  NAND2_X1 U7765 ( .A1(n7863), .A2(n5972), .ZN(n6032) );
  OR2_X1 U7766 ( .A1(n7873), .A2(n6163), .ZN(n6031) );
  NAND2_X1 U7767 ( .A1(n6032), .A2(n6031), .ZN(n7856) );
  NAND2_X1 U7768 ( .A1(n7480), .A2(n6157), .ZN(n6036) );
  OR2_X1 U7769 ( .A1(n9265), .A2(n6158), .ZN(n6035) );
  NAND2_X1 U7770 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  XNOR2_X1 U7771 ( .A(n6037), .B(n6161), .ZN(n6039) );
  NOR2_X1 U7772 ( .A1(n9265), .A2(n6163), .ZN(n6038) );
  AOI21_X1 U7773 ( .B1(n7480), .B2(n5972), .A(n6038), .ZN(n6040) );
  XNOR2_X1 U7774 ( .A(n6039), .B(n6040), .ZN(n7871) );
  INV_X1 U7775 ( .A(n6039), .ZN(n6041) );
  NAND2_X1 U7776 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7777 ( .A1(n7613), .A2(n6157), .ZN(n6044) );
  OR2_X1 U7778 ( .A1(n9353), .A2(n6158), .ZN(n6043) );
  NAND2_X1 U7779 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  XNOR2_X1 U7780 ( .A(n6045), .B(n6131), .ZN(n6047) );
  NOR2_X1 U7781 ( .A1(n9353), .A2(n6163), .ZN(n6046) );
  AOI21_X1 U7782 ( .B1(n7613), .B2(n5972), .A(n6046), .ZN(n9263) );
  AND2_X1 U7783 ( .A1(n6047), .A2(n9263), .ZN(n6056) );
  INV_X1 U7784 ( .A(n6047), .ZN(n9260) );
  INV_X1 U7785 ( .A(n9263), .ZN(n6048) );
  NAND2_X1 U7786 ( .A1(n9260), .A2(n6048), .ZN(n6054) );
  NAND2_X1 U7787 ( .A1(n9358), .A2(n6157), .ZN(n6050) );
  OR2_X1 U7788 ( .A1(n7809), .A2(n6158), .ZN(n6049) );
  NAND2_X1 U7789 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7790 ( .A(n6051), .B(n6161), .ZN(n6057) );
  NAND2_X1 U7791 ( .A1(n9358), .A2(n5972), .ZN(n6053) );
  OR2_X1 U7792 ( .A1(n7809), .A2(n6163), .ZN(n6052) );
  NAND2_X1 U7793 ( .A1(n6053), .A2(n6052), .ZN(n6058) );
  NAND2_X1 U7794 ( .A1(n6057), .A2(n6058), .ZN(n9349) );
  INV_X1 U7795 ( .A(n6057), .ZN(n6060) );
  INV_X1 U7796 ( .A(n6058), .ZN(n6059) );
  NAND2_X1 U7797 ( .A1(n6060), .A2(n6059), .ZN(n9348) );
  NAND2_X2 U7798 ( .A1(n6061), .A2(n9348), .ZN(n8053) );
  OAI22_X1 U7799 ( .A1(n9907), .A2(n5982), .B1(n6063), .B2(n6158), .ZN(n6062)
         );
  XNOR2_X1 U7800 ( .A(n6062), .B(n6131), .ZN(n6077) );
  OAI22_X1 U7801 ( .A1(n9907), .A2(n6158), .B1(n6063), .B2(n6163), .ZN(n6075)
         );
  XNOR2_X1 U7802 ( .A(n6077), .B(n6075), .ZN(n8054) );
  NAND2_X1 U7803 ( .A1(n8147), .A2(n6157), .ZN(n6065) );
  OR2_X1 U7804 ( .A1(n9242), .A2(n6158), .ZN(n6064) );
  NAND2_X1 U7805 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  XNOR2_X1 U7806 ( .A(n6066), .B(n6161), .ZN(n6070) );
  INV_X1 U7807 ( .A(n6070), .ZN(n6068) );
  NOR2_X1 U7808 ( .A1(n9242), .A2(n6163), .ZN(n6067) );
  AOI21_X1 U7809 ( .B1(n8147), .B2(n5972), .A(n6067), .ZN(n6069) );
  NAND2_X1 U7810 ( .A1(n6068), .A2(n6069), .ZN(n6078) );
  INV_X1 U7811 ( .A(n6078), .ZN(n6071) );
  XNOR2_X1 U7812 ( .A(n6070), .B(n6069), .ZN(n8142) );
  AND2_X1 U7813 ( .A1(n8054), .A2(n6085), .ZN(n6073) );
  OAI22_X1 U7814 ( .A1(n9248), .A2(n5982), .B1(n9397), .B2(n6158), .ZN(n6072)
         );
  XNOR2_X1 U7815 ( .A(n6072), .B(n6131), .ZN(n6086) );
  AND2_X1 U7816 ( .A1(n6073), .A2(n6086), .ZN(n6074) );
  INV_X1 U7817 ( .A(n6086), .ZN(n6083) );
  INV_X1 U7818 ( .A(n6085), .ZN(n6079) );
  INV_X1 U7819 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7820 ( .A1(n6077), .A2(n6076), .ZN(n8139) );
  AND2_X1 U7821 ( .A1(n8139), .A2(n6078), .ZN(n6084) );
  OR2_X1 U7822 ( .A1(n6079), .A2(n6084), .ZN(n6080) );
  OR2_X1 U7823 ( .A1(n6083), .A2(n6080), .ZN(n9232) );
  OAI22_X1 U7824 ( .A1(n9248), .A2(n6158), .B1(n9397), .B2(n6163), .ZN(n9234)
         );
  AND2_X1 U7825 ( .A1(n9232), .A2(n9234), .ZN(n6081) );
  OAI22_X1 U7826 ( .A1(n9832), .A2(n5982), .B1(n9307), .B2(n6158), .ZN(n6082)
         );
  XNOR2_X1 U7827 ( .A(n6082), .B(n6131), .ZN(n6089) );
  OR2_X1 U7828 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  OAI22_X1 U7829 ( .A1(n9832), .A2(n6158), .B1(n9307), .B2(n6163), .ZN(n9399)
         );
  AOI21_X1 U7830 ( .B1(n9239), .B2(n9236), .A(n6089), .ZN(n9398) );
  AOI22_X1 U7831 ( .A1(n9709), .A2(n5972), .B1(n6125), .B2(n9416), .ZN(n9303)
         );
  OAI22_X1 U7832 ( .A1(n9677), .A2(n6158), .B1(n9662), .B2(n6163), .ZN(n6092)
         );
  AOI22_X1 U7833 ( .A1(n9770), .A2(n6157), .B1(n5972), .B2(n9699), .ZN(n6090)
         );
  XNOR2_X1 U7834 ( .A(n6090), .B(n6161), .ZN(n6091) );
  XOR2_X1 U7835 ( .A(n6092), .B(n6091), .Z(n9311) );
  NAND2_X1 U7836 ( .A1(n9761), .A2(n6157), .ZN(n6095) );
  NAND2_X1 U7837 ( .A1(n9414), .A2(n5972), .ZN(n6094) );
  NAND2_X1 U7838 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  XNOR2_X1 U7839 ( .A(n6096), .B(n6161), .ZN(n9277) );
  NAND2_X1 U7840 ( .A1(n9761), .A2(n5972), .ZN(n6098) );
  NAND2_X1 U7841 ( .A1(n9414), .A2(n6125), .ZN(n6097) );
  NAND2_X1 U7842 ( .A1(n6098), .A2(n6097), .ZN(n9275) );
  NAND2_X1 U7843 ( .A1(n9277), .A2(n9275), .ZN(n9324) );
  INV_X1 U7844 ( .A(n9324), .ZN(n6103) );
  AOI22_X1 U7845 ( .A1(n9766), .A2(n6157), .B1(n5972), .B2(n9415), .ZN(n6099)
         );
  XNOR2_X1 U7846 ( .A(n6099), .B(n6161), .ZN(n9274) );
  OR2_X1 U7847 ( .A1(n9668), .A2(n6158), .ZN(n6101) );
  OR2_X1 U7848 ( .A1(n9687), .A2(n6163), .ZN(n6100) );
  INV_X1 U7849 ( .A(n9277), .ZN(n6111) );
  INV_X1 U7850 ( .A(n9274), .ZN(n9272) );
  INV_X1 U7851 ( .A(n9373), .ZN(n6105) );
  OAI21_X1 U7852 ( .B1(n9272), .B2(n6105), .A(n9275), .ZN(n6110) );
  NOR3_X1 U7853 ( .A1(n9272), .A2(n9275), .A3(n6105), .ZN(n6109) );
  OAI22_X1 U7854 ( .A1(n9637), .A2(n5982), .B1(n9645), .B2(n6158), .ZN(n6106)
         );
  XNOR2_X1 U7855 ( .A(n6106), .B(n6161), .ZN(n6112) );
  OR2_X1 U7856 ( .A1(n9637), .A2(n6158), .ZN(n6108) );
  NAND2_X1 U7857 ( .A1(n9613), .A2(n6125), .ZN(n6107) );
  NAND2_X1 U7858 ( .A1(n6108), .A2(n6107), .ZN(n6113) );
  NOR2_X1 U7859 ( .A1(n6112), .A2(n6113), .ZN(n9326) );
  AOI211_X1 U7860 ( .C1(n6111), .C2(n6110), .A(n6109), .B(n9326), .ZN(n6116)
         );
  INV_X1 U7861 ( .A(n6112), .ZN(n6115) );
  INV_X1 U7862 ( .A(n6113), .ZN(n6114) );
  NOR2_X1 U7863 ( .A1(n6115), .A2(n6114), .ZN(n9327) );
  AOI22_X1 U7864 ( .A1(n9745), .A2(n6157), .B1(n5972), .B2(n9614), .ZN(n6120)
         );
  XOR2_X1 U7865 ( .A(n6161), .B(n6120), .Z(n9336) );
  INV_X1 U7866 ( .A(n9336), .ZN(n6123) );
  OAI22_X1 U7867 ( .A1(n9600), .A2(n6158), .B1(n9290), .B2(n6163), .ZN(n9335)
         );
  OAI21_X1 U7868 ( .B1(n6121), .B2(n9336), .A(n9335), .ZN(n6122) );
  OAI21_X1 U7869 ( .B1(n9338), .B2(n6123), .A(n6122), .ZN(n9250) );
  AOI22_X1 U7870 ( .A1(n9256), .A2(n6157), .B1(n5972), .B2(n4954), .ZN(n6124)
         );
  XNOR2_X1 U7871 ( .A(n6124), .B(n6161), .ZN(n6127) );
  AOI22_X1 U7872 ( .A1(n9256), .A2(n5972), .B1(n6125), .B2(n4954), .ZN(n6126)
         );
  NAND2_X1 U7873 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  OAI21_X1 U7874 ( .B1(n6127), .B2(n6126), .A(n6128), .ZN(n9251) );
  INV_X1 U7875 ( .A(n6128), .ZN(n9318) );
  NAND2_X1 U7876 ( .A1(n9741), .A2(n6157), .ZN(n6130) );
  OR2_X1 U7877 ( .A1(n9553), .A2(n6158), .ZN(n6129) );
  NAND2_X1 U7878 ( .A1(n6130), .A2(n6129), .ZN(n6132) );
  XNOR2_X1 U7879 ( .A(n6132), .B(n6131), .ZN(n6135) );
  NOR2_X1 U7880 ( .A1(n9553), .A2(n6163), .ZN(n6133) );
  AOI21_X1 U7881 ( .B1(n9741), .B2(n5972), .A(n6133), .ZN(n6134) );
  NAND2_X1 U7882 ( .A1(n6135), .A2(n6134), .ZN(n6137) );
  OR2_X1 U7883 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  AND2_X1 U7884 ( .A1(n6137), .A2(n6136), .ZN(n9317) );
  OAI22_X1 U7885 ( .A1(n9800), .A2(n6158), .B1(n9575), .B2(n6163), .ZN(n6146)
         );
  NAND2_X1 U7886 ( .A1(n9562), .A2(n6157), .ZN(n6139) );
  NAND2_X1 U7887 ( .A1(n9544), .A2(n5972), .ZN(n6138) );
  NAND2_X1 U7888 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  XNOR2_X1 U7889 ( .A(n6140), .B(n6161), .ZN(n6145) );
  XOR2_X1 U7890 ( .A(n6146), .B(n6145), .Z(n9296) );
  NAND2_X1 U7891 ( .A1(n9730), .A2(n6157), .ZN(n6142) );
  OR2_X1 U7892 ( .A1(n9554), .A2(n6158), .ZN(n6141) );
  NAND2_X1 U7893 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  XNOR2_X1 U7894 ( .A(n6143), .B(n6161), .ZN(n6155) );
  NOR2_X1 U7895 ( .A1(n9554), .A2(n6163), .ZN(n6144) );
  AOI21_X1 U7896 ( .B1(n9730), .B2(n5972), .A(n6144), .ZN(n6153) );
  XNOR2_X1 U7897 ( .A(n6155), .B(n6153), .ZN(n9384) );
  INV_X1 U7898 ( .A(n6145), .ZN(n6148) );
  INV_X1 U7899 ( .A(n6146), .ZN(n6147) );
  NAND2_X1 U7900 ( .A1(n6148), .A2(n6147), .ZN(n9380) );
  AOI22_X1 U7901 ( .A1(n9529), .A2(n6157), .B1(n5972), .B2(n9545), .ZN(n6149)
         );
  XOR2_X1 U7902 ( .A(n6161), .B(n6149), .Z(n6152) );
  OAI22_X1 U7903 ( .A1(n9795), .A2(n6158), .B1(n6150), .B2(n6163), .ZN(n6151)
         );
  NOR2_X1 U7904 ( .A1(n6152), .A2(n6151), .ZN(n6171) );
  AOI21_X1 U7905 ( .B1(n6152), .B2(n6151), .A(n6171), .ZN(n9224) );
  INV_X1 U7906 ( .A(n6153), .ZN(n6154) );
  NAND2_X1 U7907 ( .A1(n6155), .A2(n6154), .ZN(n9225) );
  NAND2_X1 U7908 ( .A1(n9720), .A2(n6157), .ZN(n6160) );
  OR2_X1 U7909 ( .A1(n9520), .A2(n6158), .ZN(n6159) );
  NAND2_X1 U7910 ( .A1(n6160), .A2(n6159), .ZN(n6162) );
  XNOR2_X1 U7911 ( .A(n6162), .B(n6161), .ZN(n6166) );
  NOR2_X1 U7912 ( .A1(n9520), .A2(n6163), .ZN(n6164) );
  AOI21_X1 U7913 ( .B1(n9720), .B2(n5972), .A(n6164), .ZN(n6165) );
  XNOR2_X1 U7914 ( .A(n6166), .B(n6165), .ZN(n6170) );
  INV_X1 U7915 ( .A(n6167), .ZN(n6955) );
  NOR2_X1 U7916 ( .A1(n9829), .A2(n8523), .ZN(n6184) );
  AND2_X1 U7917 ( .A1(n9874), .A2(n6184), .ZN(n6168) );
  NOR3_X1 U7918 ( .A1(n6171), .A2(n6170), .A3(n9402), .ZN(n6169) );
  INV_X1 U7919 ( .A(n6170), .ZN(n6173) );
  INV_X1 U7920 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U7921 ( .A1(n7331), .A2(n8503), .ZN(n7330) );
  INV_X1 U7922 ( .A(n7330), .ZN(n6174) );
  AND2_X1 U7923 ( .A1(n9874), .A2(n6174), .ZN(n6175) );
  NAND2_X1 U7924 ( .A1(n6183), .A2(n6175), .ZN(n6178) );
  INV_X1 U7925 ( .A(n6176), .ZN(n6177) );
  INV_X1 U7926 ( .A(n6179), .ZN(n7332) );
  NAND2_X1 U7927 ( .A1(n9874), .A2(n7332), .ZN(n8536) );
  INV_X1 U7928 ( .A(n8536), .ZN(n6180) );
  NAND2_X1 U7929 ( .A1(n6183), .A2(n6180), .ZN(n6189) );
  INV_X1 U7930 ( .A(n6189), .ZN(n6181) );
  INV_X1 U7931 ( .A(n6182), .ZN(n9511) );
  AOI22_X1 U7932 ( .A1(n9391), .A2(n9511), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6191) );
  INV_X1 U7933 ( .A(n6183), .ZN(n6188) );
  INV_X1 U7934 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7935 ( .A1(n8503), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7800) );
  NAND3_X1 U7936 ( .A1(n8536), .A2(n6185), .A3(n7800), .ZN(n6187) );
  NAND3_X1 U7937 ( .A1(n7323), .A2(n5951), .A3(n8011), .ZN(n6186) );
  AOI21_X1 U7938 ( .B1(n6188), .B2(n6187), .A(n6186), .ZN(n7186) );
  NOR2_X2 U7939 ( .A1(n7186), .A2(P1_U3086), .ZN(n9393) );
  NOR2_X2 U7940 ( .A1(n6189), .A2(n5922), .ZN(n9386) );
  AOI22_X1 U7941 ( .A1(n9393), .A2(n9505), .B1(n9386), .B2(n9545), .ZN(n6190)
         );
  OAI211_X1 U7942 ( .C1(n4875), .C2(n9299), .A(n6191), .B(n6190), .ZN(n6192)
         );
  INV_X1 U7943 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7944 ( .A1(n4566), .A2(n6193), .ZN(n6194) );
  NOR2_X1 U7945 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  NAND2_X1 U7946 ( .A1(n6197), .A2(n6196), .ZN(P1_U3220) );
  INV_X1 U7947 ( .A(SI_29_), .ZN(n10441) );
  INV_X1 U7948 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8666) );
  INV_X1 U7949 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6202) );
  MUX2_X1 U7950 ( .A(n8666), .B(n6202), .S(n6931), .Z(n6204) );
  INV_X1 U7951 ( .A(SI_30_), .ZN(n6203) );
  NAND2_X1 U7952 ( .A1(n6204), .A2(n6203), .ZN(n6207) );
  INV_X1 U7953 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U7954 ( .A1(n6205), .A2(SI_30_), .ZN(n6206) );
  NAND2_X1 U7955 ( .A1(n6207), .A2(n6206), .ZN(n6246) );
  MUX2_X1 U7956 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6931), .Z(n6208) );
  INV_X1 U7957 ( .A(SI_31_), .ZN(n10229) );
  XNOR2_X1 U7958 ( .A(n6208), .B(n10229), .ZN(n6209) );
  NAND2_X2 U7959 ( .A1(n6261), .A2(n5416), .ZN(n6558) );
  INV_X1 U7960 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9210) );
  OR2_X1 U7961 ( .A1(n6558), .A2(n9210), .ZN(n6211) );
  NAND2_X1 U7962 ( .A1(n10159), .A2(n7560), .ZN(n6305) );
  INV_X1 U7963 ( .A(n6305), .ZN(n6213) );
  NAND2_X1 U7964 ( .A1(n6213), .A2(n10435), .ZN(n6315) );
  INV_X1 U7965 ( .A(n6326), .ZN(n6214) );
  NAND2_X1 U7966 ( .A1(n6214), .A2(n10457), .ZN(n6337) );
  INV_X1 U7967 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6218) );
  INV_X1 U7968 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6221) );
  INV_X1 U7969 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6224) );
  INV_X1 U7970 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10254) );
  INV_X1 U7971 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10231) );
  INV_X1 U7972 ( .A(n6535), .ZN(n6229) );
  INV_X1 U7973 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7974 ( .A1(n6229), .A2(n6228), .ZN(n6548) );
  INV_X1 U7975 ( .A(n8657), .ZN(n6237) );
  NAND2_X1 U7976 ( .A1(n6234), .A2(n6235), .ZN(n9208) );
  INV_X1 U7977 ( .A(n6239), .ZN(n6238) );
  NAND2_X1 U7978 ( .A1(n6237), .A2(n6550), .ZN(n6566) );
  INV_X1 U7979 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U7980 ( .A1(n4502), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6243) );
  NAND2_X2 U7981 ( .A1(n6239), .A2(n6241), .ZN(n6507) );
  INV_X1 U7982 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9072) );
  OR2_X1 U7983 ( .A1(n6507), .A2(n9072), .ZN(n6242) );
  OAI211_X1 U7984 ( .C1(n8883), .C2(n6436), .A(n6243), .B(n6242), .ZN(n6244)
         );
  INV_X1 U7985 ( .A(n6244), .ZN(n6245) );
  NOR2_X1 U7986 ( .A1(n9070), .A2(n8880), .ZN(n6766) );
  INV_X1 U7987 ( .A(n6766), .ZN(n6254) );
  OR2_X1 U7988 ( .A1(n6558), .A2(n8666), .ZN(n6248) );
  INV_X1 U7989 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U7990 ( .A1(n6561), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7991 ( .A1(n4502), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6250) );
  OAI211_X1 U7992 ( .C1(n8886), .C2(n6436), .A(n6251), .B(n6250), .ZN(n6252)
         );
  INV_X1 U7993 ( .A(n6252), .ZN(n6253) );
  NAND2_X1 U7994 ( .A1(n6566), .A2(n6253), .ZN(n8766) );
  INV_X1 U7995 ( .A(n8766), .ZN(n6255) );
  NAND2_X1 U7996 ( .A1(n9128), .A2(n6255), .ZN(n6762) );
  OR2_X1 U7997 ( .A1(n9128), .A2(n6255), .ZN(n6754) );
  INV_X1 U7998 ( .A(n6754), .ZN(n6761) );
  NAND2_X1 U7999 ( .A1(n6761), .A2(n9070), .ZN(n6256) );
  NAND2_X1 U8000 ( .A1(n9070), .A2(n8880), .ZN(n6765) );
  NAND3_X1 U8001 ( .A1(n6256), .A2(n6765), .A3(n6865), .ZN(n6597) );
  INV_X4 U8002 ( .A(n6267), .ZN(n6436) );
  OR2_X1 U8003 ( .A1(n6507), .A2(n7151), .ZN(n6259) );
  NAND2_X1 U8004 ( .A1(n6265), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6258) );
  INV_X1 U8005 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7319) );
  OR2_X1 U8006 ( .A1(n6283), .A2(n7319), .ZN(n6257) );
  OR2_X1 U8007 ( .A1(n6322), .A2(n6943), .ZN(n6263) );
  OR2_X1 U8008 ( .A1(n6261), .A2(n7150), .ZN(n6262) );
  OR2_X2 U8009 ( .A1(n7298), .A2(n7953), .ZN(n6609) );
  NAND2_X1 U8010 ( .A1(n7298), .A2(n7953), .ZN(n6613) );
  INV_X1 U8011 ( .A(n6776), .ZN(n6577) );
  NAND2_X1 U8012 ( .A1(n4502), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6271) );
  INV_X1 U8013 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7269) );
  OR2_X1 U8014 ( .A1(n6283), .A2(n7269), .ZN(n6268) );
  NAND2_X1 U8015 ( .A1(n6272), .A2(SI_0_), .ZN(n6273) );
  XNOR2_X1 U8016 ( .A(n6273), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9222) );
  MUX2_X1 U8017 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9222), .S(n6261), .Z(n7456) );
  INV_X1 U8018 ( .A(n7456), .ZN(n7301) );
  NAND2_X1 U8019 ( .A1(n6577), .A2(n6605), .ZN(n7459) );
  NAND2_X1 U8020 ( .A1(n7459), .A2(n6609), .ZN(n7617) );
  INV_X1 U8021 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6274) );
  OR2_X1 U8022 ( .A1(n6506), .A2(n6274), .ZN(n6278) );
  OR2_X1 U8023 ( .A1(n6436), .A2(n5152), .ZN(n6277) );
  OR2_X1 U8024 ( .A1(n6507), .A2(n6275), .ZN(n6276) );
  OR2_X1 U8025 ( .A1(n6558), .A2(n5297), .ZN(n6282) );
  OR2_X1 U8026 ( .A1(n6322), .A2(n6937), .ZN(n6281) );
  OR2_X1 U8027 ( .A1(n6261), .A2(n9937), .ZN(n6280) );
  NAND2_X1 U8028 ( .A1(n8780), .A2(n10024), .ZN(n6618) );
  NAND2_X1 U8029 ( .A1(n6617), .A2(n6618), .ZN(n6779) );
  NAND2_X1 U8030 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  NAND2_X1 U8031 ( .A1(n7616), .A2(n6617), .ZN(n7553) );
  NAND2_X1 U8032 ( .A1(n4502), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6288) );
  OR2_X1 U8033 ( .A1(n6283), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6287) );
  INV_X1 U8034 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7559) );
  OR2_X1 U8035 ( .A1(n6436), .A2(n7559), .ZN(n6286) );
  INV_X1 U8036 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6284) );
  OR2_X1 U8037 ( .A1(n6507), .A2(n6284), .ZN(n6285) );
  INV_X1 U8038 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6933) );
  OR2_X1 U8039 ( .A1(n6558), .A2(n6933), .ZN(n6291) );
  OR2_X1 U8040 ( .A1(n6322), .A2(n6932), .ZN(n6290) );
  OR2_X1 U8041 ( .A1(n6261), .A2(n9953), .ZN(n6289) );
  NAND2_X1 U8042 ( .A1(n7629), .A2(n6632), .ZN(n7556) );
  INV_X1 U8043 ( .A(n7556), .ZN(n6292) );
  NAND2_X1 U8044 ( .A1(n7553), .A2(n6292), .ZN(n7630) );
  NAND2_X1 U8045 ( .A1(n7630), .A2(n7629), .ZN(n6304) );
  NAND2_X1 U8046 ( .A1(n4502), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6299) );
  OR2_X1 U8047 ( .A1(n6436), .A2(n6293), .ZN(n6298) );
  NAND2_X1 U8048 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6294) );
  AND2_X1 U8049 ( .A1(n6305), .A2(n6294), .ZN(n10016) );
  OR2_X1 U8050 ( .A1(n6283), .A2(n10016), .ZN(n6297) );
  OR2_X1 U8051 ( .A1(n6507), .A2(n6295), .ZN(n6296) );
  INV_X1 U8052 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6936) );
  OR2_X1 U8053 ( .A1(n6558), .A2(n6936), .ZN(n6301) );
  OR2_X1 U8054 ( .A1(n6322), .A2(n6934), .ZN(n6300) );
  OAI211_X1 U8055 ( .C1(n6261), .C2(n6935), .A(n6301), .B(n6300), .ZN(n10018)
         );
  NAND2_X1 U8056 ( .A1(n8777), .A2(n10018), .ZN(n7692) );
  INV_X1 U8057 ( .A(n10018), .ZN(n6302) );
  NAND2_X1 U8058 ( .A1(n6303), .A2(n6302), .ZN(n6783) );
  INV_X1 U8059 ( .A(n7636), .ZN(n6624) );
  OR2_X1 U8060 ( .A1(n8777), .A2(n6302), .ZN(n6635) );
  NAND2_X1 U8061 ( .A1(n4502), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6310) );
  INV_X1 U8062 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7696) );
  OR2_X1 U8063 ( .A1(n6436), .A2(n7696), .ZN(n6309) );
  NAND2_X1 U8064 ( .A1(n6305), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6306) );
  AND2_X1 U8065 ( .A1(n6315), .A2(n6306), .ZN(n7697) );
  OR2_X1 U8066 ( .A1(n6283), .A2(n7697), .ZN(n6308) );
  INV_X1 U8067 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6917) );
  OR2_X1 U8068 ( .A1(n6507), .A2(n6917), .ZN(n6307) );
  INV_X1 U8069 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6946) );
  OR2_X1 U8070 ( .A1(n6558), .A2(n6946), .ZN(n6312) );
  OR2_X1 U8071 ( .A1(n6322), .A2(n6944), .ZN(n6311) );
  OAI211_X1 U8072 ( .C1(n6261), .C2(n6945), .A(n6312), .B(n6311), .ZN(n6578)
         );
  NOR2_X1 U8073 ( .A1(n8776), .A2(n7939), .ZN(n6633) );
  NAND2_X1 U8074 ( .A1(n8776), .A2(n7939), .ZN(n6638) );
  NAND2_X1 U8075 ( .A1(n6313), .A2(n6638), .ZN(n7767) );
  NAND2_X1 U8076 ( .A1(n4502), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6321) );
  OR2_X1 U8077 ( .A1(n6436), .A2(n6314), .ZN(n6320) );
  NAND2_X1 U8078 ( .A1(n6315), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6316) );
  AND2_X1 U8079 ( .A1(n6326), .A2(n6316), .ZN(n7769) );
  OR2_X1 U8080 ( .A1(n6283), .A2(n7769), .ZN(n6319) );
  OR2_X1 U8081 ( .A1(n6507), .A2(n6317), .ZN(n6318) );
  OR2_X1 U8082 ( .A1(n6322), .A2(n6942), .ZN(n6324) );
  INV_X1 U8083 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6940) );
  OR2_X1 U8084 ( .A1(n6558), .A2(n6940), .ZN(n6323) );
  OAI211_X1 U8085 ( .C1(n6261), .C2(n6941), .A(n6324), .B(n6323), .ZN(n7710)
         );
  INV_X1 U8086 ( .A(n7710), .ZN(n10029) );
  AND2_X1 U8087 ( .A1(n8775), .A2(n10029), .ZN(n6639) );
  OR2_X1 U8088 ( .A1(n8775), .A2(n10029), .ZN(n6628) );
  OAI21_X1 U8089 ( .B1(n7767), .B2(n6639), .A(n6628), .ZN(n6325) );
  INV_X1 U8090 ( .A(n6325), .ZN(n7879) );
  OR2_X1 U8091 ( .A1(n6436), .A2(n10012), .ZN(n6332) );
  NAND2_X1 U8092 ( .A1(n6326), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6327) );
  AND2_X1 U8093 ( .A1(n6337), .A2(n6327), .ZN(n10007) );
  OR2_X1 U8094 ( .A1(n6283), .A2(n10007), .ZN(n6331) );
  NAND2_X1 U8095 ( .A1(n4502), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6330) );
  OR2_X1 U8096 ( .A1(n6507), .A2(n6328), .ZN(n6329) );
  OR2_X1 U8097 ( .A1(n6322), .A2(n6949), .ZN(n6335) );
  INV_X1 U8098 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6947) );
  OR2_X1 U8099 ( .A1(n6558), .A2(n6947), .ZN(n6334) );
  OR2_X1 U8100 ( .A1(n6261), .A2(n6948), .ZN(n6333) );
  NAND2_X1 U8101 ( .A1(n4502), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6343) );
  OR2_X1 U8102 ( .A1(n6436), .A2(n8026), .ZN(n6342) );
  NAND2_X1 U8103 ( .A1(n6337), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6338) );
  AND2_X1 U8104 ( .A1(n6347), .A2(n6338), .ZN(n8025) );
  OR2_X1 U8105 ( .A1(n6283), .A2(n8025), .ZN(n6341) );
  OR2_X1 U8106 ( .A1(n6507), .A2(n6339), .ZN(n6340) );
  NAND4_X1 U8107 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n8773)
         );
  INV_X1 U8108 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6954) );
  OR2_X1 U8109 ( .A1(n6558), .A2(n6954), .ZN(n6344) );
  OAI211_X1 U8110 ( .C1(n6261), .C2(n6952), .A(n6345), .B(n6344), .ZN(n8030)
         );
  NAND2_X1 U8111 ( .A1(n8773), .A2(n7973), .ZN(n6645) );
  AND2_X1 U8112 ( .A1(n7962), .A2(n6645), .ZN(n6658) );
  NAND2_X1 U8113 ( .A1(n4502), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6352) );
  OR2_X1 U8114 ( .A1(n6507), .A2(n6346), .ZN(n6351) );
  NAND2_X1 U8115 ( .A1(n6347), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6348) );
  AND2_X1 U8116 ( .A1(n6360), .A2(n6348), .ZN(n8106) );
  OR2_X1 U8117 ( .A1(n6283), .A2(n8106), .ZN(n6350) );
  OR2_X1 U8118 ( .A1(n6436), .A2(n8107), .ZN(n6349) );
  NAND4_X1 U8119 ( .A1(n6352), .A2(n6351), .A3(n6350), .A4(n6349), .ZN(n8114)
         );
  AOI22_X1 U8120 ( .A1(n6451), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6450), .B2(
        n6353), .ZN(n6354) );
  NAND2_X1 U8121 ( .A1(n6355), .A2(n6354), .ZN(n8109) );
  OR2_X1 U8122 ( .A1(n8114), .A2(n10033), .ZN(n6652) );
  NAND2_X1 U8123 ( .A1(n10033), .A2(n8114), .ZN(n6656) );
  NAND2_X1 U8124 ( .A1(n6652), .A2(n6656), .ZN(n8099) );
  OR2_X1 U8125 ( .A1(n6962), .A2(n6322), .ZN(n6358) );
  AOI22_X1 U8126 ( .A1(n6451), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6450), .B2(
        n6356), .ZN(n6357) );
  NAND2_X1 U8127 ( .A1(n6358), .A2(n6357), .ZN(n10039) );
  INV_X1 U8128 ( .A(n10039), .ZN(n8094) );
  NAND2_X1 U8129 ( .A1(n4502), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6366) );
  OR2_X1 U8130 ( .A1(n6507), .A2(n6359), .ZN(n6365) );
  NAND2_X1 U8131 ( .A1(n6360), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6361) );
  AND2_X1 U8132 ( .A1(n6371), .A2(n6361), .ZN(n8092) );
  OR2_X1 U8133 ( .A1(n6283), .A2(n8092), .ZN(n6364) );
  OR2_X1 U8134 ( .A1(n6436), .A2(n6362), .ZN(n6363) );
  NAND4_X1 U8135 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n8772)
         );
  AND2_X1 U8136 ( .A1(n8094), .A2(n8772), .ZN(n6655) );
  INV_X1 U8137 ( .A(n8772), .ZN(n8100) );
  NAND2_X1 U8138 ( .A1(n10039), .A2(n8100), .ZN(n6664) );
  AOI22_X1 U8139 ( .A1(n6451), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6450), .B2(
        n6367), .ZN(n6368) );
  NAND2_X1 U8140 ( .A1(n6369), .A2(n6368), .ZN(n10048) );
  NAND2_X1 U8141 ( .A1(n4502), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6376) );
  INV_X1 U8142 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6370) );
  OR2_X1 U8143 ( .A1(n6507), .A2(n6370), .ZN(n6375) );
  NAND2_X1 U8144 ( .A1(n6371), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6372) );
  AND2_X1 U8145 ( .A1(n6381), .A2(n6372), .ZN(n8183) );
  OR2_X1 U8146 ( .A1(n6283), .A2(n8183), .ZN(n6374) );
  OR2_X1 U8147 ( .A1(n6436), .A2(n7931), .ZN(n6373) );
  OR2_X1 U8148 ( .A1(n10048), .A2(n8175), .ZN(n6668) );
  NAND2_X1 U8149 ( .A1(n10048), .A2(n8175), .ZN(n8168) );
  NAND2_X1 U8150 ( .A1(n6668), .A2(n8168), .ZN(n7982) );
  NAND2_X1 U8151 ( .A1(n8163), .A2(n8162), .ZN(n8169) );
  OR2_X1 U8152 ( .A1(n7048), .A2(n6322), .ZN(n6379) );
  AOI22_X1 U8153 ( .A1(n6451), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6450), .B2(
        n6377), .ZN(n6378) );
  NAND2_X1 U8154 ( .A1(n6379), .A2(n6378), .ZN(n8179) );
  INV_X1 U8155 ( .A(n8179), .ZN(n10055) );
  NAND2_X1 U8156 ( .A1(n4502), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6386) );
  OR2_X1 U8157 ( .A1(n6507), .A2(n6380), .ZN(n6385) );
  NAND2_X1 U8158 ( .A1(n6381), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6382) );
  AND2_X1 U8159 ( .A1(n6391), .A2(n6382), .ZN(n8176) );
  OR2_X1 U8160 ( .A1(n6283), .A2(n8176), .ZN(n6384) );
  OR2_X1 U8161 ( .A1(n6436), .A2(n8177), .ZN(n6383) );
  NAND4_X1 U8162 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n8770)
         );
  NAND2_X1 U8163 ( .A1(n10055), .A2(n8770), .ZN(n6676) );
  INV_X1 U8164 ( .A(n8770), .ZN(n8210) );
  NAND2_X1 U8165 ( .A1(n8179), .A2(n8210), .ZN(n6675) );
  NAND2_X1 U8166 ( .A1(n6676), .A2(n6675), .ZN(n8171) );
  INV_X1 U8167 ( .A(n8168), .ZN(n6669) );
  NOR2_X1 U8168 ( .A1(n8171), .A2(n6669), .ZN(n6387) );
  AOI22_X1 U8169 ( .A1(n6451), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6450), .B2(
        n6388), .ZN(n6389) );
  NAND2_X1 U8170 ( .A1(n4502), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6397) );
  INV_X1 U8171 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8226) );
  OR2_X1 U8172 ( .A1(n6507), .A2(n8226), .ZN(n6396) );
  NAND2_X1 U8173 ( .A1(n6391), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6392) );
  AND2_X1 U8174 ( .A1(n6403), .A2(n6392), .ZN(n8219) );
  OR2_X1 U8175 ( .A1(n6283), .A2(n8219), .ZN(n6395) );
  OR2_X1 U8176 ( .A1(n6436), .A2(n6393), .ZN(n6394) );
  NAND4_X1 U8177 ( .A1(n6397), .A2(n6396), .A3(n6395), .A4(n6394), .ZN(n9056)
         );
  NAND2_X1 U8178 ( .A1(n8227), .A2(n8174), .ZN(n6398) );
  AOI22_X1 U8179 ( .A1(n6451), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6450), .B2(
        n6400), .ZN(n6401) );
  NAND2_X1 U8180 ( .A1(n4502), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6409) );
  OR2_X1 U8181 ( .A1(n6507), .A2(n9120), .ZN(n6408) );
  NAND2_X1 U8182 ( .A1(n6403), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6404) );
  AND2_X1 U8183 ( .A1(n6413), .A2(n6404), .ZN(n9062) );
  OR2_X1 U8184 ( .A1(n6283), .A2(n9062), .ZN(n6407) );
  OR2_X1 U8185 ( .A1(n6436), .A2(n6405), .ZN(n6406) );
  NAND4_X1 U8186 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n9047)
         );
  NAND2_X1 U8187 ( .A1(n9201), .A2(n8211), .ZN(n6684) );
  AOI22_X1 U8188 ( .A1(n6451), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6450), .B2(
        n6410), .ZN(n6411) );
  NAND2_X1 U8189 ( .A1(n4502), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6418) );
  INV_X1 U8190 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9117) );
  OR2_X1 U8191 ( .A1(n6507), .A2(n9117), .ZN(n6417) );
  NAND2_X1 U8192 ( .A1(n6413), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6414) );
  AND2_X1 U8193 ( .A1(n6424), .A2(n6414), .ZN(n8131) );
  OR2_X1 U8194 ( .A1(n6283), .A2(n8131), .ZN(n6416) );
  OR2_X1 U8195 ( .A1(n6436), .A2(n9048), .ZN(n6415) );
  NAND4_X1 U8196 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n9058)
         );
  AND2_X1 U8197 ( .A1(n9194), .A2(n8544), .ZN(n6576) );
  INV_X1 U8198 ( .A(n6576), .ZN(n6419) );
  NAND2_X1 U8199 ( .A1(n6420), .A2(n6688), .ZN(n9026) );
  AOI22_X1 U8200 ( .A1(n6451), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6450), .B2(
        n6421), .ZN(n6422) );
  NAND2_X1 U8201 ( .A1(n4502), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6429) );
  OR2_X1 U8202 ( .A1(n6507), .A2(n9114), .ZN(n6428) );
  NAND2_X1 U8203 ( .A1(n6424), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6425) );
  AND2_X1 U8204 ( .A1(n6434), .A2(n6425), .ZN(n9031) );
  OR2_X1 U8205 ( .A1(n6283), .A2(n9031), .ZN(n6427) );
  OR2_X1 U8206 ( .A1(n6436), .A2(n5195), .ZN(n6426) );
  NAND2_X1 U8207 ( .A1(n9188), .A2(n9037), .ZN(n6694) );
  NAND2_X1 U8208 ( .A1(n9026), .A2(n6694), .ZN(n6430) );
  AOI22_X1 U8209 ( .A1(n6451), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6450), .B2(
        n5201), .ZN(n6431) );
  NAND2_X1 U8210 ( .A1(n4502), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6440) );
  OR2_X1 U8211 ( .A1(n6507), .A2(n6433), .ZN(n6439) );
  NAND2_X1 U8212 ( .A1(n6434), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6435) );
  AND2_X1 U8213 ( .A1(n6443), .A2(n6435), .ZN(n9018) );
  OR2_X1 U8214 ( .A1(n6283), .A2(n9018), .ZN(n6438) );
  OR2_X1 U8215 ( .A1(n6436), .A2(n9019), .ZN(n6437) );
  OR2_X1 U8216 ( .A1(n9110), .A2(n9005), .ZN(n6702) );
  NAND2_X1 U8217 ( .A1(n9110), .A2(n9005), .ZN(n6693) );
  NAND2_X1 U8218 ( .A1(n6702), .A2(n6693), .ZN(n9021) );
  AOI22_X1 U8219 ( .A1(n6451), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6450), .B2(
        n8863), .ZN(n6441) );
  NAND2_X1 U8220 ( .A1(n4502), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8221 ( .A1(n6507), .A2(n8855), .ZN(n6447) );
  NAND2_X1 U8222 ( .A1(n6443), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6444) );
  AND2_X1 U8223 ( .A1(n6454), .A2(n6444), .ZN(n9008) );
  OR2_X1 U8224 ( .A1(n6283), .A2(n9008), .ZN(n6446) );
  OR2_X1 U8225 ( .A1(n6436), .A2(n5205), .ZN(n6445) );
  NAND2_X1 U8226 ( .A1(n6813), .A2(n8993), .ZN(n6692) );
  NAND2_X1 U8227 ( .A1(n9009), .A2(n6708), .ZN(n8987) );
  NAND2_X1 U8228 ( .A1(n4533), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6449) );
  AOI22_X1 U8229 ( .A1(n6451), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7462), .B2(
        n6450), .ZN(n6452) );
  NAND2_X1 U8230 ( .A1(n4502), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6459) );
  INV_X1 U8231 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9102) );
  OR2_X1 U8232 ( .A1(n6507), .A2(n9102), .ZN(n6458) );
  NAND2_X1 U8233 ( .A1(n6454), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6455) );
  AND2_X1 U8234 ( .A1(n6503), .A2(n6455), .ZN(n8997) );
  OR2_X1 U8235 ( .A1(n6283), .A2(n8997), .ZN(n6457) );
  INV_X1 U8236 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8996) );
  OR2_X1 U8237 ( .A1(n6436), .A2(n8996), .ZN(n6456) );
  NAND2_X1 U8238 ( .A1(n9178), .A2(n9003), .ZN(n6711) );
  OR2_X1 U8239 ( .A1(n6558), .A2(n8138), .ZN(n6460) );
  INV_X1 U8240 ( .A(n9150), .ZN(n6818) );
  NAND2_X1 U8241 ( .A1(n6469), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8242 ( .A1(n6476), .A2(n6462), .ZN(n8942) );
  NAND2_X1 U8243 ( .A1(n8942), .A2(n6550), .ZN(n6465) );
  AOI22_X1 U8244 ( .A1(n6561), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n4502), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8245 ( .A1(n6267), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8246 ( .A1(n6818), .A2(n8921), .ZN(n6729) );
  OR2_X1 U8247 ( .A1(n6558), .A2(n8016), .ZN(n6466) );
  INV_X1 U8248 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U8249 ( .A1(n6496), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8250 ( .A1(n6469), .A2(n6468), .ZN(n8677) );
  NAND2_X1 U8251 ( .A1(n8677), .A2(n6550), .ZN(n6473) );
  NAND2_X1 U8252 ( .A1(n6561), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8253 ( .A1(n4502), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6470) );
  AND2_X1 U8254 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  OAI211_X1 U8255 ( .C1(n6436), .C2(n8605), .A(n6473), .B(n6472), .ZN(n8957)
         );
  NAND2_X1 U8256 ( .A1(n8681), .A2(n8940), .ZN(n8943) );
  AND2_X1 U8257 ( .A1(n6729), .A2(n8943), .ZN(n8929) );
  OR2_X1 U8258 ( .A1(n6558), .A2(n8224), .ZN(n6474) );
  NAND2_X1 U8259 ( .A1(n6476), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8260 ( .A1(n6524), .A2(n6477), .ZN(n8924) );
  NAND2_X1 U8261 ( .A1(n8924), .A2(n6550), .ZN(n6483) );
  INV_X1 U8262 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8263 ( .A1(n6561), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U8264 ( .A1(n4502), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6478) );
  OAI211_X1 U8265 ( .C1(n6480), .C2(n6436), .A(n6479), .B(n6478), .ZN(n6481)
         );
  INV_X1 U8266 ( .A(n6481), .ZN(n6482) );
  NAND2_X1 U8267 ( .A1(n8618), .A2(n8939), .ZN(n6573) );
  AND2_X1 U8268 ( .A1(n8929), .A2(n6573), .ZN(n6515) );
  INV_X1 U8269 ( .A(n6730), .ZN(n6514) );
  OR2_X1 U8270 ( .A1(n6558), .A2(n7868), .ZN(n6484) );
  NAND2_X1 U8271 ( .A1(n6505), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U8272 ( .A1(n6494), .A2(n6486), .ZN(n8966) );
  NAND2_X1 U8273 ( .A1(n6550), .A2(n8966), .ZN(n6491) );
  INV_X1 U8274 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9166) );
  OR2_X1 U8275 ( .A1(n6506), .A2(n9166), .ZN(n6490) );
  INV_X1 U8276 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9093) );
  OR2_X1 U8277 ( .A1(n6507), .A2(n9093), .ZN(n6489) );
  INV_X1 U8278 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6487) );
  OR2_X1 U8279 ( .A1(n6436), .A2(n6487), .ZN(n6488) );
  OR2_X1 U8280 ( .A1(n6558), .A2(n7999), .ZN(n6492) );
  NAND2_X1 U8281 ( .A1(n6494), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8282 ( .A1(n6496), .A2(n6495), .ZN(n8960) );
  NAND2_X1 U8283 ( .A1(n8960), .A2(n6550), .ZN(n6500) );
  NAND2_X1 U8284 ( .A1(n6561), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U8285 ( .A1(n4502), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8286 ( .A1(n6267), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8287 ( .A1(n9167), .A2(n8558), .ZN(n6575) );
  INV_X1 U8288 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7803) );
  OR2_X1 U8289 ( .A1(n6558), .A2(n7803), .ZN(n6501) );
  NAND2_X1 U8290 ( .A1(n6503), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8291 ( .A1(n6505), .A2(n6504), .ZN(n8982) );
  NAND2_X1 U8292 ( .A1(n6550), .A2(n8982), .ZN(n6512) );
  INV_X1 U8293 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9172) );
  OR2_X1 U8294 ( .A1(n6506), .A2(n9172), .ZN(n6511) );
  INV_X1 U8295 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9099) );
  OR2_X1 U8296 ( .A1(n6507), .A2(n9099), .ZN(n6510) );
  INV_X1 U8297 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6508) );
  OR2_X1 U8298 ( .A1(n6436), .A2(n6508), .ZN(n6509) );
  NAND2_X1 U8299 ( .A1(n8727), .A2(n8992), .ZN(n8963) );
  AND2_X1 U8300 ( .A1(n6575), .A2(n8963), .ZN(n8951) );
  OR2_X1 U8301 ( .A1(n5082), .A2(n8951), .ZN(n6513) );
  NAND2_X1 U8302 ( .A1(n9161), .A2(n8603), .ZN(n6722) );
  NAND2_X1 U8303 ( .A1(n6513), .A2(n6722), .ZN(n8597) );
  NAND2_X1 U8304 ( .A1(n6514), .A2(n8597), .ZN(n8927) );
  AND2_X1 U8305 ( .A1(n6515), .A2(n8927), .ZN(n6516) );
  AND2_X1 U8306 ( .A1(n8991), .A2(n6516), .ZN(n6518) );
  INV_X1 U8307 ( .A(n6516), .ZN(n6517) );
  INV_X1 U8308 ( .A(n6716), .ZN(n8950) );
  OR2_X1 U8309 ( .A1(n8950), .A2(n5082), .ZN(n8596) );
  AND2_X1 U8310 ( .A1(n5075), .A2(n8595), .ZN(n8925) );
  AOI21_X1 U8311 ( .B1(n8987), .B2(n6518), .A(n5067), .ZN(n6521) );
  INV_X1 U8312 ( .A(n6573), .ZN(n6736) );
  NAND2_X1 U8313 ( .A1(n9150), .A2(n8769), .ZN(n8930) );
  OR2_X1 U8314 ( .A1(n6736), .A2(n8930), .ZN(n6519) );
  OR2_X1 U8315 ( .A1(n6558), .A2(n8232), .ZN(n6522) );
  NAND2_X1 U8316 ( .A1(n6524), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8317 ( .A1(n6535), .A2(n6525), .ZN(n8912) );
  NAND2_X1 U8318 ( .A1(n8912), .A2(n6550), .ZN(n6531) );
  INV_X1 U8319 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8320 ( .A1(n4502), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8321 ( .A1(n6561), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6526) );
  OAI211_X1 U8322 ( .C1(n6528), .C2(n6436), .A(n6527), .B(n6526), .ZN(n6529)
         );
  INV_X1 U8323 ( .A(n6529), .ZN(n6530) );
  NOR2_X1 U8324 ( .A1(n6820), .A2(n8922), .ZN(n6740) );
  NAND2_X1 U8325 ( .A1(n6820), .A2(n8922), .ZN(n6572) );
  NAND2_X1 U8326 ( .A1(n6535), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8327 ( .A1(n6548), .A2(n6536), .ZN(n8901) );
  NAND2_X1 U8328 ( .A1(n8901), .A2(n6550), .ZN(n6542) );
  INV_X1 U8329 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8330 ( .A1(n6561), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U8331 ( .A1(n4502), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6537) );
  OAI211_X1 U8332 ( .C1(n6539), .C2(n6436), .A(n6538), .B(n6537), .ZN(n6540)
         );
  INV_X1 U8333 ( .A(n6540), .ZN(n6541) );
  NAND2_X2 U8334 ( .A1(n6542), .A2(n6541), .ZN(n8891) );
  INV_X1 U8335 ( .A(n6743), .ZN(n6543) );
  NAND2_X1 U8336 ( .A1(n6544), .A2(n6571), .ZN(n8887) );
  INV_X1 U8337 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6545) );
  OR2_X1 U8338 ( .A1(n6558), .A2(n6545), .ZN(n6546) );
  NAND2_X1 U8339 ( .A1(n6548), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8340 ( .A1(n8657), .A2(n6549), .ZN(n8897) );
  NAND2_X1 U8341 ( .A1(n8897), .A2(n6550), .ZN(n6555) );
  INV_X1 U8342 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U8343 ( .A1(n4502), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8344 ( .A1(n6561), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6551) );
  OAI211_X1 U8345 ( .C1(n8896), .C2(n6436), .A(n6552), .B(n6551), .ZN(n6553)
         );
  INV_X1 U8346 ( .A(n6553), .ZN(n6554) );
  NAND2_X1 U8347 ( .A1(n8887), .A2(n8888), .ZN(n6557) );
  OR2_X1 U8348 ( .A1(n9134), .A2(n6824), .ZN(n6556) );
  NAND2_X1 U8349 ( .A1(n6557), .A2(n6556), .ZN(n6830) );
  INV_X1 U8350 ( .A(n6830), .ZN(n6570) );
  OR2_X1 U8351 ( .A1(n6558), .A2(n9217), .ZN(n6559) );
  INV_X1 U8352 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U8353 ( .A1(n4502), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8354 ( .A1(n6561), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U8355 ( .C1(n6436), .C2(n8656), .A(n6563), .B(n6562), .ZN(n6564)
         );
  INV_X1 U8356 ( .A(n6564), .ZN(n6565) );
  INV_X1 U8357 ( .A(n9070), .ZN(n9127) );
  NAND2_X1 U8358 ( .A1(n8659), .A2(n8767), .ZN(n6749) );
  INV_X1 U8359 ( .A(n6749), .ZN(n6567) );
  AOI21_X1 U8360 ( .B1(n9127), .B2(n9128), .A(n6567), .ZN(n6568) );
  AOI21_X1 U8361 ( .B1(n6570), .B2(n6753), .A(n6569), .ZN(n6598) );
  INV_X1 U8362 ( .A(n6765), .ZN(n6596) );
  INV_X1 U8363 ( .A(n6829), .ZN(n6594) );
  INV_X1 U8364 ( .A(n6571), .ZN(n6744) );
  OR2_X2 U8365 ( .A1(n6744), .A2(n6743), .ZN(n8902) );
  INV_X1 U8366 ( .A(n6572), .ZN(n6741) );
  NAND2_X1 U8367 ( .A1(n8930), .A2(n6729), .ZN(n8945) );
  NAND2_X1 U8368 ( .A1(n6735), .A2(n6573), .ZN(n8933) );
  INV_X1 U8369 ( .A(n8943), .ZN(n6574) );
  NOR2_X1 U8370 ( .A1(n6730), .A2(n6574), .ZN(n8600) );
  NAND2_X1 U8371 ( .A1(n8952), .A2(n6575), .ZN(n8967) );
  INV_X1 U8372 ( .A(n8967), .ZN(n6590) );
  NAND2_X1 U8373 ( .A1(n6716), .A2(n8963), .ZN(n8980) );
  INV_X1 U8374 ( .A(n9021), .ZN(n9015) );
  NOR2_X1 U8375 ( .A1(n7556), .A2(n6776), .ZN(n6579) );
  XNOR2_X1 U8376 ( .A(n8776), .B(n6578), .ZN(n7694) );
  NAND4_X1 U8377 ( .A1(n6579), .A2(n6624), .A3(n7618), .A4(n7694), .ZN(n6581)
         );
  NAND2_X1 U8378 ( .A1(n8781), .A2(n7301), .ZN(n6601) );
  AND2_X1 U8379 ( .A1(n6601), .A2(n7461), .ZN(n7452) );
  NAND2_X1 U8380 ( .A1(n8775), .A2(n7710), .ZN(n6785) );
  NAND2_X1 U8381 ( .A1(n6789), .A2(n6785), .ZN(n7768) );
  NAND4_X1 U8382 ( .A1(n7452), .A2(n6336), .A3(n6604), .A4(n7768), .ZN(n6580)
         );
  NOR2_X1 U8383 ( .A1(n6581), .A2(n6580), .ZN(n6583) );
  INV_X1 U8384 ( .A(n6664), .ZN(n6582) );
  NOR2_X1 U8385 ( .A1(n6655), .A2(n6582), .ZN(n8085) );
  AND2_X1 U8386 ( .A1(n6651), .A2(n6645), .ZN(n7967) );
  NAND4_X1 U8387 ( .A1(n6583), .A2(n4752), .A3(n8085), .A4(n7967), .ZN(n6584)
         );
  NOR3_X1 U8388 ( .A1(n8171), .A2(n6584), .A3(n7982), .ZN(n6585) );
  NAND2_X1 U8389 ( .A1(n8227), .A2(n9056), .ZN(n6802) );
  NOR2_X1 U8390 ( .A1(n8227), .A2(n9056), .ZN(n6801) );
  OR2_X1 U8391 ( .A1(n4691), .A2(n6801), .ZN(n8209) );
  NAND4_X1 U8392 ( .A1(n9039), .A2(n9053), .A3(n6585), .A4(n8209), .ZN(n6586)
         );
  NAND2_X1 U8393 ( .A1(n6696), .A2(n6694), .ZN(n6808) );
  NOR2_X1 U8394 ( .A1(n6586), .A2(n6808), .ZN(n6587) );
  NAND4_X1 U8395 ( .A1(n8991), .A2(n9015), .A3(n9010), .A4(n6587), .ZN(n6588)
         );
  NOR2_X1 U8396 ( .A1(n8980), .A2(n6588), .ZN(n6589) );
  NAND4_X1 U8397 ( .A1(n8600), .A2(n8955), .A3(n6590), .A4(n6589), .ZN(n6591)
         );
  OR4_X1 U8398 ( .A1(n8609), .A2(n8945), .A3(n8933), .A4(n6591), .ZN(n6592) );
  NOR2_X1 U8399 ( .A1(n8902), .A2(n6592), .ZN(n6593) );
  NAND4_X1 U8400 ( .A1(n6594), .A2(n6593), .A3(n8888), .A4(n6754), .ZN(n6595)
         );
  OAI22_X1 U8401 ( .A1(n6598), .A2(n6597), .B1(n6596), .B2(n6595), .ZN(n6599)
         );
  NAND2_X1 U8402 ( .A1(n6601), .A2(n6865), .ZN(n6600) );
  NAND2_X1 U8403 ( .A1(n6600), .A2(n6881), .ZN(n6603) );
  NAND3_X1 U8404 ( .A1(n6601), .A2(n6613), .A3(n6831), .ZN(n6602) );
  NAND2_X1 U8405 ( .A1(n6603), .A2(n6602), .ZN(n6607) );
  NOR2_X1 U8406 ( .A1(n6613), .A2(n6837), .ZN(n6614) );
  NOR2_X1 U8407 ( .A1(n6614), .A2(n6779), .ZN(n6615) );
  NAND2_X1 U8408 ( .A1(n6616), .A2(n6615), .ZN(n6623) );
  NAND2_X1 U8409 ( .A1(n7629), .A2(n6617), .ZN(n6620) );
  NAND2_X1 U8410 ( .A1(n6632), .A2(n6618), .ZN(n6619) );
  MUX2_X1 U8411 ( .A(n6620), .B(n6619), .S(n6837), .Z(n6621) );
  INV_X1 U8412 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8413 ( .A1(n6623), .A2(n6622), .ZN(n6625) );
  NAND2_X1 U8414 ( .A1(n6625), .A2(n6624), .ZN(n6637) );
  INV_X1 U8415 ( .A(n7629), .ZN(n6627) );
  NAND2_X1 U8416 ( .A1(n8777), .A2(n6302), .ZN(n6626) );
  OAI211_X1 U8417 ( .C1(n6637), .C2(n6627), .A(n6626), .B(n6638), .ZN(n6630)
         );
  INV_X1 U8418 ( .A(n6628), .ZN(n6641) );
  NOR2_X1 U8419 ( .A1(n6633), .A2(n6641), .ZN(n6629) );
  AOI21_X1 U8420 ( .B1(n6630), .B2(n6629), .A(n6639), .ZN(n6631) );
  OR2_X1 U8421 ( .A1(n6631), .A2(n6881), .ZN(n6649) );
  INV_X1 U8422 ( .A(n6632), .ZN(n6636) );
  INV_X1 U8423 ( .A(n6633), .ZN(n6634) );
  OAI211_X1 U8424 ( .C1(n6637), .C2(n6636), .A(n6635), .B(n6634), .ZN(n6643)
         );
  INV_X1 U8425 ( .A(n6638), .ZN(n6640) );
  NOR2_X1 U8426 ( .A1(n6640), .A2(n6639), .ZN(n6642) );
  AOI21_X1 U8427 ( .B1(n6643), .B2(n6642), .A(n6641), .ZN(n6644) );
  OR2_X1 U8428 ( .A1(n6644), .A2(n6837), .ZN(n6648) );
  NAND2_X1 U8429 ( .A1(n6656), .A2(n6645), .ZN(n6646) );
  NOR2_X1 U8430 ( .A1(n6654), .A2(n7885), .ZN(n6647) );
  NAND3_X1 U8431 ( .A1(n6649), .A2(n6648), .A3(n6647), .ZN(n6663) );
  AND2_X1 U8432 ( .A1(n6651), .A2(n6650), .ZN(n6653) );
  OAI211_X1 U8433 ( .C1(n6654), .C2(n6653), .A(n6652), .B(n6664), .ZN(n6660)
         );
  INV_X1 U8434 ( .A(n6655), .ZN(n6667) );
  OAI211_X1 U8435 ( .C1(n6658), .C2(n6657), .A(n6667), .B(n6656), .ZN(n6659)
         );
  MUX2_X1 U8436 ( .A(n6660), .B(n6659), .S(n6881), .Z(n6661) );
  INV_X1 U8437 ( .A(n6661), .ZN(n6662) );
  NAND2_X1 U8438 ( .A1(n6663), .A2(n6662), .ZN(n6671) );
  AND2_X1 U8439 ( .A1(n8168), .A2(n6664), .ZN(n6666) );
  INV_X1 U8440 ( .A(n6668), .ZN(n6665) );
  AOI21_X1 U8441 ( .B1(n6671), .B2(n6666), .A(n6665), .ZN(n6673) );
  AND2_X1 U8442 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  AOI21_X1 U8443 ( .B1(n6671), .B2(n6670), .A(n6669), .ZN(n6672) );
  INV_X1 U8444 ( .A(n8171), .ZN(n6674) );
  MUX2_X1 U8445 ( .A(n6676), .B(n6675), .S(n6881), .Z(n6677) );
  MUX2_X1 U8446 ( .A(n9056), .B(n8227), .S(n6881), .Z(n6678) );
  NAND2_X1 U8447 ( .A1(n6679), .A2(n6801), .ZN(n6680) );
  NAND2_X1 U8448 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  NAND2_X1 U8449 ( .A1(n6682), .A2(n9053), .ZN(n6686) );
  MUX2_X1 U8450 ( .A(n6684), .B(n6683), .S(n6837), .Z(n6685) );
  NAND2_X1 U8451 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  NAND2_X1 U8452 ( .A1(n6687), .A2(n9039), .ZN(n6698) );
  INV_X1 U8453 ( .A(n6808), .ZN(n9027) );
  NAND2_X1 U8454 ( .A1(n6698), .A2(n5066), .ZN(n6690) );
  NAND2_X1 U8455 ( .A1(n6694), .A2(n6881), .ZN(n6689) );
  NAND2_X1 U8456 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NAND2_X1 U8457 ( .A1(n6691), .A2(n9015), .ZN(n6701) );
  OAI211_X1 U8458 ( .C1(n9021), .C2(n6694), .A(n6693), .B(n6692), .ZN(n6695)
         );
  NAND2_X1 U8459 ( .A1(n6695), .A2(n6837), .ZN(n6700) );
  NAND2_X1 U8460 ( .A1(n6696), .A2(n6881), .ZN(n6697) );
  AOI21_X1 U8461 ( .B1(n6698), .B2(n6419), .A(n6697), .ZN(n6699) );
  INV_X1 U8462 ( .A(n6702), .ZN(n6704) );
  NAND3_X1 U8463 ( .A1(n6813), .A2(n8993), .A3(n6881), .ZN(n6703) );
  OAI21_X1 U8464 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6709) );
  NAND3_X1 U8465 ( .A1(n6705), .A2(n8991), .A3(n6708), .ZN(n6707) );
  NAND2_X1 U8466 ( .A1(n6711), .A2(n6881), .ZN(n6706) );
  AOI22_X1 U8467 ( .A1(n6709), .A2(n6708), .B1(n6707), .B2(n6706), .ZN(n6715)
         );
  INV_X1 U8468 ( .A(n8980), .ZN(n6710) );
  NAND2_X1 U8469 ( .A1(n6710), .A2(n8595), .ZN(n6713) );
  NAND2_X1 U8470 ( .A1(n8963), .A2(n6711), .ZN(n6712) );
  MUX2_X1 U8471 ( .A(n6713), .B(n6712), .S(n6837), .Z(n6714) );
  OAI22_X1 U8472 ( .A1(n6715), .A2(n6714), .B1(n6837), .B2(n8951), .ZN(n6718)
         );
  AOI21_X1 U8473 ( .B1(n8952), .B2(n6716), .A(n6881), .ZN(n6717) );
  AOI21_X1 U8474 ( .B1(n6718), .B2(n8952), .A(n6717), .ZN(n6720) );
  INV_X1 U8475 ( .A(n9167), .ZN(n8699) );
  NAND2_X1 U8476 ( .A1(n8955), .A2(n5065), .ZN(n6719) );
  NOR2_X1 U8477 ( .A1(n6720), .A2(n6719), .ZN(n6728) );
  INV_X1 U8478 ( .A(n6721), .ZN(n6724) );
  NAND2_X1 U8479 ( .A1(n8943), .A2(n6722), .ZN(n6723) );
  MUX2_X1 U8480 ( .A(n6724), .B(n6723), .S(n6881), .Z(n6725) );
  INV_X1 U8481 ( .A(n8930), .ZN(n6731) );
  OAI21_X1 U8482 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6734) );
  INV_X1 U8483 ( .A(n8929), .ZN(n6732) );
  NAND2_X1 U8484 ( .A1(n6732), .A2(n8930), .ZN(n6733) );
  MUX2_X1 U8485 ( .A(n6734), .B(n6733), .S(n6837), .Z(n6739) );
  INV_X1 U8486 ( .A(n6735), .ZN(n6737) );
  MUX2_X1 U8487 ( .A(n6737), .B(n6736), .S(n6881), .Z(n6738) );
  MUX2_X1 U8488 ( .A(n6741), .B(n6740), .S(n6881), .Z(n6742) );
  MUX2_X1 U8489 ( .A(n6744), .B(n6743), .S(n6881), .Z(n6745) );
  MUX2_X1 U8490 ( .A(n6825), .B(n6824), .S(n6837), .Z(n6759) );
  NAND2_X1 U8491 ( .A1(n6760), .A2(n6759), .ZN(n6752) );
  NAND2_X1 U8492 ( .A1(n6752), .A2(n6748), .ZN(n6750) );
  NAND2_X1 U8493 ( .A1(n6752), .A2(n6825), .ZN(n6755) );
  OAI21_X1 U8494 ( .B1(n6755), .B2(n6829), .A(n5072), .ZN(n6756) );
  NAND2_X1 U8495 ( .A1(n6756), .A2(n6837), .ZN(n6757) );
  AOI21_X1 U8496 ( .B1(n6837), .B2(n6762), .A(n6761), .ZN(n6763) );
  OR2_X1 U8497 ( .A1(n6764), .A2(n6763), .ZN(n6768) );
  AOI21_X1 U8498 ( .B1(n6768), .B2(n6767), .A(n6766), .ZN(n6771) );
  NAND2_X1 U8499 ( .A1(n6769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6770) );
  OR2_X1 U8500 ( .A1(n6772), .A2(P2_U3151), .ZN(n8014) );
  NAND2_X1 U8501 ( .A1(n6831), .A2(n8869), .ZN(n6875) );
  INV_X1 U8502 ( .A(n6875), .ZN(n6773) );
  NAND2_X1 U8503 ( .A1(n6773), .A2(n7463), .ZN(n7255) );
  INV_X1 U8504 ( .A(n7255), .ZN(n7451) );
  NAND2_X1 U8505 ( .A1(n7258), .A2(n7451), .ZN(n7249) );
  NOR3_X1 U8506 ( .A1(n7249), .A2(n6834), .A3(n5208), .ZN(n6775) );
  OAI21_X1 U8507 ( .B1(n8014), .B2(n6831), .A(P2_B_REG_SCAN_IN), .ZN(n6774) );
  INV_X1 U8508 ( .A(n8992), .ZN(n8970) );
  INV_X1 U8509 ( .A(n9003), .ZN(n8977) );
  NAND2_X1 U8510 ( .A1(n8781), .A2(n7456), .ZN(n7464) );
  NAND2_X1 U8511 ( .A1(n6776), .A2(n7464), .ZN(n6778) );
  INV_X1 U8512 ( .A(n7953), .ZN(n7466) );
  OR2_X1 U8513 ( .A1(n7298), .A2(n7466), .ZN(n6777) );
  NAND2_X1 U8514 ( .A1(n6778), .A2(n6777), .ZN(n7619) );
  NAND2_X1 U8515 ( .A1(n7619), .A2(n6779), .ZN(n6782) );
  INV_X1 U8516 ( .A(n10024), .ZN(n6780) );
  OR2_X1 U8517 ( .A1(n8780), .A2(n6780), .ZN(n6781) );
  NAND2_X1 U8518 ( .A1(n6782), .A2(n6781), .ZN(n7557) );
  NAND2_X1 U8519 ( .A1(n7557), .A2(n7556), .ZN(n7634) );
  INV_X1 U8520 ( .A(n7958), .ZN(n7561) );
  OR2_X1 U8521 ( .A1(n8778), .A2(n7561), .ZN(n7633) );
  AND2_X1 U8522 ( .A1(n6783), .A2(n7633), .ZN(n6784) );
  NAND2_X1 U8523 ( .A1(n7634), .A2(n6784), .ZN(n7693) );
  NAND2_X1 U8524 ( .A1(n8776), .A2(n6578), .ZN(n7764) );
  AND2_X1 U8525 ( .A1(n7764), .A2(n6785), .ZN(n7880) );
  INV_X1 U8526 ( .A(n7948), .ZN(n10008) );
  NAND2_X1 U8527 ( .A1(n8774), .A2(n10008), .ZN(n6788) );
  NOR2_X1 U8528 ( .A1(n8776), .A2(n6578), .ZN(n7762) );
  OR2_X1 U8529 ( .A1(n8773), .A2(n8030), .ZN(n6790) );
  AND2_X1 U8530 ( .A1(n6790), .A2(n7965), .ZN(n6791) );
  NAND2_X1 U8531 ( .A1(n7966), .A2(n6791), .ZN(n6793) );
  NAND2_X1 U8532 ( .A1(n8773), .A2(n8030), .ZN(n6792) );
  NAND2_X1 U8533 ( .A1(n6793), .A2(n6792), .ZN(n8098) );
  OR2_X1 U8534 ( .A1(n8114), .A2(n8109), .ZN(n6794) );
  NAND2_X1 U8535 ( .A1(n8114), .A2(n8109), .ZN(n6795) );
  OR2_X1 U8536 ( .A1(n10039), .A2(n8772), .ZN(n6796) );
  NAND2_X1 U8537 ( .A1(n8158), .A2(n7982), .ZN(n6798) );
  INV_X1 U8538 ( .A(n8175), .ZN(n8771) );
  NAND2_X1 U8539 ( .A1(n10048), .A2(n8771), .ZN(n6797) );
  AND2_X1 U8540 ( .A1(n8179), .A2(n8770), .ZN(n6800) );
  NAND2_X1 U8541 ( .A1(n10055), .A2(n8210), .ZN(n6799) );
  NAND2_X1 U8542 ( .A1(n8206), .A2(n6802), .ZN(n9054) );
  OR2_X1 U8543 ( .A1(n9201), .A2(n9047), .ZN(n6803) );
  NAND2_X1 U8544 ( .A1(n9054), .A2(n6803), .ZN(n6805) );
  NAND2_X1 U8545 ( .A1(n9201), .A2(n9047), .ZN(n6804) );
  NAND2_X1 U8546 ( .A1(n6805), .A2(n6804), .ZN(n9041) );
  OR2_X1 U8547 ( .A1(n9194), .A2(n9058), .ZN(n6806) );
  NAND2_X1 U8548 ( .A1(n9194), .A2(n9058), .ZN(n9043) );
  NAND2_X1 U8549 ( .A1(n9188), .A2(n9016), .ZN(n6807) );
  AND2_X1 U8550 ( .A1(n9043), .A2(n6807), .ZN(n6810) );
  INV_X1 U8551 ( .A(n6807), .ZN(n6809) );
  INV_X1 U8552 ( .A(n9005), .ZN(n9029) );
  AND2_X1 U8553 ( .A1(n9110), .A2(n9029), .ZN(n6811) );
  AOI21_X1 U8554 ( .B1(n9014), .B2(n9021), .A(n6811), .ZN(n9002) );
  NAND2_X1 U8555 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8556 ( .A1(n9002), .A2(n6814), .ZN(n6816) );
  NAND2_X1 U8557 ( .A1(n8765), .A2(n8993), .ZN(n6815) );
  NAND2_X1 U8558 ( .A1(n6816), .A2(n6815), .ZN(n8990) );
  NOR2_X1 U8559 ( .A1(n8681), .A2(n8957), .ZN(n6817) );
  OAI22_X2 U8560 ( .A1(n8601), .A2(n6817), .B1(n9155), .B2(n8940), .ZN(n8937)
         );
  NOR2_X1 U8561 ( .A1(n9150), .A2(n8921), .ZN(n6819) );
  NAND2_X1 U8562 ( .A1(n8914), .A2(n8922), .ZN(n6821) );
  NAND2_X1 U8563 ( .A1(n9140), .A2(n8891), .ZN(n6823) );
  NOR2_X1 U8564 ( .A1(n9140), .A2(n8891), .ZN(n6822) );
  NAND2_X1 U8565 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  AOI22_X1 U8566 ( .A1(n8889), .A2(n6826), .B1(n8905), .B2(n9134), .ZN(n6827)
         );
  XNOR2_X1 U8567 ( .A(n6827), .B(n6829), .ZN(n6842) );
  NAND2_X1 U8568 ( .A1(n6831), .A2(n7462), .ZN(n6864) );
  OR2_X1 U8569 ( .A1(n6604), .A2(n7805), .ZN(n6828) );
  XNOR2_X1 U8570 ( .A(n6830), .B(n6829), .ZN(n8661) );
  INV_X1 U8571 ( .A(n7293), .ZN(n6832) );
  NAND2_X1 U8572 ( .A1(n6875), .A2(n6832), .ZN(n6833) );
  NAND2_X1 U8573 ( .A1(n8661), .A2(n8102), .ZN(n6840) );
  INV_X1 U8574 ( .A(n7288), .ZN(n6836) );
  NAND2_X1 U8575 ( .A1(n6261), .A2(P2_B_REG_SCAN_IN), .ZN(n6838) );
  AND2_X1 U8576 ( .A1(n9057), .A2(n6838), .ZN(n8878) );
  AOI22_X1 U8577 ( .A1(n9055), .A2(n8905), .B1(n8766), .B2(n8878), .ZN(n6839)
         );
  NAND2_X1 U8578 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  AND2_X1 U8579 ( .A1(n7805), .A2(n7462), .ZN(n6868) );
  INV_X1 U8580 ( .A(n10040), .ZN(n10034) );
  NAND2_X1 U8581 ( .A1(n8655), .A2(n6843), .ZN(n6887) );
  XNOR2_X1 U8582 ( .A(n6844), .B(P2_B_REG_SCAN_IN), .ZN(n6846) );
  NAND2_X1 U8583 ( .A1(n6846), .A2(n6845), .ZN(n6848) );
  NAND2_X1 U8584 ( .A1(n6845), .A2(n8233), .ZN(n6849) );
  NAND2_X1 U8585 ( .A1(n8233), .A2(n6844), .ZN(n7102) );
  INV_X2 U8586 ( .A(n6852), .ZN(n7292) );
  NOR2_X1 U8587 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6856) );
  NOR4_X1 U8588 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6855) );
  NOR4_X1 U8589 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6854) );
  NOR4_X1 U8590 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6853) );
  NAND4_X1 U8591 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6862)
         );
  NOR4_X1 U8592 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6860) );
  NOR4_X1 U8593 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6859) );
  NOR4_X1 U8594 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6858) );
  NOR4_X1 U8595 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6857) );
  NAND4_X1 U8596 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n6861)
         );
  NOR2_X1 U8597 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  NAND2_X1 U8598 ( .A1(n7449), .A2(n6882), .ZN(n7251) );
  INV_X1 U8599 ( .A(n7258), .ZN(n9206) );
  INV_X1 U8600 ( .A(n6864), .ZN(n6866) );
  NOR2_X1 U8601 ( .A1(n6865), .A2(n7805), .ZN(n7291) );
  NAND2_X1 U8602 ( .A1(n6866), .A2(n7291), .ZN(n7260) );
  AND2_X1 U8603 ( .A1(n6881), .A2(n10054), .ZN(n6867) );
  NAND2_X1 U8604 ( .A1(n7260), .A2(n6867), .ZN(n7262) );
  NAND2_X1 U8605 ( .A1(n9207), .A2(n7292), .ZN(n6883) );
  INV_X1 U8606 ( .A(n6882), .ZN(n6869) );
  NOR2_X1 U8607 ( .A1(n6883), .A2(n6869), .ZN(n7243) );
  NAND2_X1 U8608 ( .A1(n7260), .A2(n7255), .ZN(n6870) );
  NAND2_X1 U8609 ( .A1(n7264), .A2(n6870), .ZN(n6871) );
  OR2_X1 U8610 ( .A1(n10052), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6873) );
  OAI21_X1 U8611 ( .B1(n6887), .B2(n10061), .A(n6873), .ZN(n6874) );
  INV_X1 U8612 ( .A(n8659), .ZN(n6888) );
  NAND2_X1 U8613 ( .A1(n6874), .A2(n5063), .ZN(P2_U3456) );
  OR2_X1 U8614 ( .A1(n6875), .A2(n7805), .ZN(n6876) );
  NAND2_X1 U8615 ( .A1(n6876), .A2(n6881), .ZN(n6877) );
  NAND2_X1 U8616 ( .A1(n9207), .A2(n6877), .ZN(n6880) );
  INV_X1 U8617 ( .A(n6877), .ZN(n6878) );
  NAND2_X1 U8618 ( .A1(n7292), .A2(n6878), .ZN(n6879) );
  NAND2_X1 U8619 ( .A1(n6880), .A2(n6879), .ZN(n7450) );
  OR2_X1 U8620 ( .A1(n6881), .A2(n7293), .ZN(n7244) );
  NAND3_X1 U8621 ( .A1(n6882), .A2(n7258), .A3(n7244), .ZN(n7448) );
  NOR2_X1 U8622 ( .A1(n7448), .A2(n7257), .ZN(n6884) );
  INV_X2 U8623 ( .A(n10068), .ZN(n10065) );
  INV_X1 U8624 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U8625 ( .A1(n10068), .A2(n6885), .ZN(n6886) );
  OAI21_X1 U8626 ( .B1(n6887), .B2(n10068), .A(n6886), .ZN(n6889) );
  NAND2_X1 U8627 ( .A1(n6889), .A2(n5069), .ZN(P2_U3488) );
  OR2_X1 U8628 ( .A1(n9955), .A2(n6892), .ZN(n6894) );
  INV_X1 U8629 ( .A(n9993), .ZN(n9958) );
  AOI211_X1 U8630 ( .C1(n6895), .C2(n6894), .A(n9958), .B(n6893), .ZN(n6913)
         );
  NOR2_X1 U8631 ( .A1(n9983), .A2(n6935), .ZN(n6912) );
  INV_X1 U8632 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6896) );
  NOR2_X1 U8633 ( .A1(n9982), .A2(n6896), .ZN(n6911) );
  OAI21_X1 U8634 ( .B1(n6899), .B2(n6898), .A(n6897), .ZN(n6900) );
  NAND2_X1 U8635 ( .A1(n9994), .A2(n6900), .ZN(n6909) );
  INV_X1 U8636 ( .A(n6901), .ZN(n6903) );
  NAND3_X1 U8637 ( .A1(n9948), .A2(n6903), .A3(n6902), .ZN(n6904) );
  NAND2_X1 U8638 ( .A1(n6905), .A2(n6904), .ZN(n6906) );
  NAND2_X1 U8639 ( .A1(n9974), .A2(n6906), .ZN(n6908) );
  NOR2_X1 U8640 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10159), .ZN(n7550) );
  INV_X1 U8641 ( .A(n7550), .ZN(n6907) );
  NAND3_X1 U8642 ( .A1(n6909), .A2(n6908), .A3(n6907), .ZN(n6910) );
  OR4_X1 U8643 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(P2_U3186)
         );
  XNOR2_X1 U8644 ( .A(n6915), .B(n6914), .ZN(n6916) );
  NOR2_X1 U8645 ( .A1(n6916), .A2(n9958), .ZN(n6927) );
  NOR2_X1 U8646 ( .A1(n9983), .A2(n6945), .ZN(n6926) );
  XNOR2_X1 U8647 ( .A(n6918), .B(n6917), .ZN(n6919) );
  NOR2_X1 U8648 ( .A1(n8876), .A2(n6919), .ZN(n6925) );
  OAI21_X1 U8649 ( .B1(n6920), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7505), .ZN(
        n6921) );
  NAND2_X1 U8650 ( .A1(n9974), .A2(n6921), .ZN(n6923) );
  INV_X1 U8651 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10435) );
  NOR2_X1 U8652 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10435), .ZN(n7647) );
  INV_X1 U8653 ( .A(n7647), .ZN(n6922) );
  OAI211_X1 U8654 ( .C1(n9982), .C2(n10084), .A(n6923), .B(n6922), .ZN(n6924)
         );
  OR4_X1 U8655 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(P2_U3187)
         );
  AND2_X1 U8656 ( .A1(n6931), .A2(P1_U3086), .ZN(n8010) );
  INV_X2 U8657 ( .A(n8010), .ZN(n9826) );
  AOI22_X1 U8658 ( .A1(n9823), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n7098), .ZN(n6928) );
  OAI21_X1 U8659 ( .B1(n6937), .B2(n9826), .A(n6928), .ZN(P1_U3353) );
  AOI22_X1 U8660 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n9823), .B1(n9439), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6929) );
  OAI21_X1 U8661 ( .B1(n6932), .B2(n9826), .A(n6929), .ZN(P1_U3352) );
  AOI22_X1 U8662 ( .A1(n7077), .A2(P1_STATE_REG_SCAN_IN), .B1(n9823), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6930) );
  OAI21_X1 U8663 ( .B1(n6934), .B2(n9826), .A(n6930), .ZN(P1_U3351) );
  AND2_X1 U8664 ( .A1(n6931), .A2(P2_U3151), .ZN(n9219) );
  INV_X2 U8665 ( .A(n9219), .ZN(n9216) );
  NOR2_X1 U8666 ( .A1(n6931), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9213) );
  OAI222_X1 U8667 ( .A1(n9216), .A2(n6933), .B1(n9953), .B2(P2_U3151), .C1(
        n8665), .C2(n6932), .ZN(P2_U3292) );
  OAI222_X1 U8668 ( .A1(n9216), .A2(n6936), .B1(n6935), .B2(P2_U3151), .C1(
        n8665), .C2(n6934), .ZN(P2_U3291) );
  OAI222_X1 U8669 ( .A1(n9216), .A2(n5297), .B1(n9937), .B2(P2_U3151), .C1(
        n8665), .C2(n6937), .ZN(P2_U3293) );
  INV_X1 U8670 ( .A(n9428), .ZN(n6938) );
  INV_X1 U8671 ( .A(n9823), .ZN(n8653) );
  OAI222_X1 U8672 ( .A1(n6938), .A2(P1_U3086), .B1(n8653), .B2(n4713), .C1(
        n6943), .C2(n9826), .ZN(P1_U3354) );
  INV_X1 U8673 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6939) );
  OAI222_X1 U8674 ( .A1(P1_U3086), .A2(n9452), .B1(n9826), .B2(n6944), .C1(
        n6939), .C2(n8653), .ZN(P1_U3350) );
  OAI222_X1 U8675 ( .A1(P1_U3086), .A2(n7016), .B1(n9826), .B2(n6942), .C1(
        n4602), .C2(n8653), .ZN(P1_U3349) );
  OAI222_X1 U8676 ( .A1(n8665), .A2(n6942), .B1(n6941), .B2(P2_U3151), .C1(
        n6940), .C2(n9216), .ZN(P2_U3289) );
  OAI222_X1 U8677 ( .A1(n9216), .A2(n5293), .B1(n7150), .B2(P2_U3151), .C1(
        n8665), .C2(n6943), .ZN(P2_U3294) );
  OAI222_X1 U8678 ( .A1(n9216), .A2(n6946), .B1(n6945), .B2(P2_U3151), .C1(
        n8665), .C2(n6944), .ZN(P2_U3290) );
  OAI222_X1 U8679 ( .A1(n8665), .A2(n6949), .B1(n6948), .B2(P2_U3151), .C1(
        n6947), .C2(n9216), .ZN(P2_U3288) );
  INV_X1 U8680 ( .A(n7036), .ZN(n7032) );
  INV_X1 U8681 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10412) );
  OAI222_X1 U8682 ( .A1(P1_U3086), .A2(n7032), .B1(n9826), .B2(n6949), .C1(
        n10412), .C2(n8653), .ZN(P1_U3348) );
  INV_X1 U8683 ( .A(n6950), .ZN(n6953) );
  AOI22_X1 U8684 ( .A1(n7062), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9823), .ZN(n6951) );
  OAI21_X1 U8685 ( .B1(n6953), .B2(n9826), .A(n6951), .ZN(P1_U3347) );
  OAI222_X1 U8686 ( .A1(n9216), .A2(n6954), .B1(n8665), .B2(n6953), .C1(
        P2_U3151), .C2(n6952), .ZN(P2_U3287) );
  INV_X1 U8687 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6957) );
  AND2_X1 U8688 ( .A1(n6955), .A2(n9874), .ZN(n7328) );
  INV_X1 U8689 ( .A(n7328), .ZN(n6956) );
  OAI21_X1 U8690 ( .B1(n9874), .B2(n6957), .A(n6956), .ZN(P1_U3440) );
  INV_X1 U8691 ( .A(n6958), .ZN(n6960) );
  OAI222_X1 U8692 ( .A1(n8665), .A2(n6960), .B1(n9216), .B2(n5327), .C1(
        P2_U3151), .C2(n7782), .ZN(P2_U3286) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6959) );
  OAI222_X1 U8694 ( .A1(n8665), .A2(n6962), .B1(n7835), .B2(P2_U3151), .C1(
        n6959), .C2(n9216), .ZN(P2_U3285) );
  INV_X1 U8695 ( .A(n7120), .ZN(n7042) );
  OAI222_X1 U8696 ( .A1(n7042), .A2(P1_U3086), .B1(n8653), .B2(n5326), .C1(
        n6960), .C2(n9826), .ZN(P1_U3346) );
  INV_X1 U8697 ( .A(n7219), .ZN(n7211) );
  INV_X1 U8698 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6961) );
  OAI222_X1 U8699 ( .A1(P1_U3086), .A2(n7211), .B1(n9826), .B2(n6962), .C1(
        n6961), .C2(n8653), .ZN(P1_U3345) );
  NAND2_X1 U8700 ( .A1(n7862), .A2(P1_U3973), .ZN(n6963) );
  OAI21_X1 U8701 ( .B1(n5327), .B2(P1_U3973), .A(n6963), .ZN(P1_U3563) );
  AND2_X1 U8702 ( .A1(n7101), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8703 ( .A1(n7101), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8704 ( .A1(n7101), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8705 ( .A1(n7101), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8706 ( .A1(n7101), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8707 ( .A1(n7101), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8708 ( .A1(n7101), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8709 ( .A1(n7101), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8710 ( .A1(n7101), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8711 ( .A1(n7101), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8712 ( .A1(n7101), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8713 ( .A(n8011), .ZN(n6964) );
  OR2_X1 U8714 ( .A1(n5951), .A2(n6964), .ZN(n6965) );
  NAND2_X1 U8715 ( .A1(n6965), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8716 ( .A1(n8011), .A2(n8523), .ZN(n6967) );
  NAND2_X1 U8717 ( .A1(n6967), .A2(n6966), .ZN(n6969) );
  INV_X1 U8718 ( .A(n6969), .ZN(n6968) );
  INV_X1 U8719 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U8720 ( .A1(n6970), .A2(n6969), .ZN(n6988) );
  NAND3_X1 U8721 ( .A1(n9459), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5966), .ZN(
        n6974) );
  OAI21_X1 U8722 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n5926), .A(n7081), .ZN(
        n7082) );
  AOI21_X1 U8723 ( .B1(n5966), .B2(n5926), .A(n7082), .ZN(n6971) );
  MUX2_X1 U8724 ( .A(n7082), .B(n6971), .S(n4796), .Z(n6972) );
  AOI22_X1 U8725 ( .A1(n6988), .A2(n6972), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6973) );
  OAI211_X1 U8726 ( .C1(n9852), .C2(n6975), .A(n6974), .B(n6973), .ZN(P1_U3243) );
  INV_X1 U8727 ( .A(n7375), .ZN(n7379) );
  INV_X1 U8728 ( .A(n6976), .ZN(n6977) );
  INV_X1 U8729 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10437) );
  OAI222_X1 U8730 ( .A1(n7379), .A2(P1_U3086), .B1(n9826), .B2(n6977), .C1(
        n10437), .C2(n8653), .ZN(P1_U3344) );
  INV_X1 U8731 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U8732 ( .A1(n9216), .A2(n6978), .B1(n8665), .B2(n6977), .C1(
        P2_U3151), .C2(n7928), .ZN(P2_U3284) );
  NAND2_X1 U8733 ( .A1(n6988), .A2(n5922), .ZN(n9843) );
  INV_X1 U8734 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6979) );
  AND2_X1 U8735 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9433) );
  NAND2_X1 U8736 ( .A1(n9428), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6980) );
  INV_X1 U8737 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6981) );
  XNOR2_X1 U8738 ( .A(n7098), .B(n6981), .ZN(n7093) );
  NAND2_X1 U8739 ( .A1(n7092), .A2(n7093), .ZN(n7091) );
  NAND2_X1 U8740 ( .A1(n7098), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U8741 ( .A1(n7091), .A2(n6982), .ZN(n9442) );
  INV_X1 U8742 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6983) );
  XNOR2_X1 U8743 ( .A(n9439), .B(n6983), .ZN(n9443) );
  NAND2_X1 U8744 ( .A1(n9442), .A2(n9443), .ZN(n9441) );
  NAND2_X1 U8745 ( .A1(n9439), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U8746 ( .A1(n9441), .A2(n6984), .ZN(n7071) );
  INV_X1 U8747 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6985) );
  XNOR2_X1 U8748 ( .A(n7077), .B(n6985), .ZN(n7072) );
  NAND2_X1 U8749 ( .A1(n7071), .A2(n7072), .ZN(n7070) );
  NAND2_X1 U8750 ( .A1(n7077), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U8751 ( .A1(n7070), .A2(n6986), .ZN(n9456) );
  XNOR2_X1 U8752 ( .A(n9452), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9457) );
  XNOR2_X1 U8753 ( .A(n7020), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U8754 ( .A1(n7081), .A2(n6987), .ZN(n8535) );
  INV_X1 U8755 ( .A(n8535), .ZN(n7083) );
  AOI211_X1 U8756 ( .C1(n6990), .C2(n6989), .A(n7017), .B(n9471), .ZN(n7012)
         );
  INV_X1 U8757 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6991) );
  MUX2_X1 U8758 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6991), .S(n9428), .Z(n6993)
         );
  AND2_X1 U8759 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6992) );
  NAND2_X1 U8760 ( .A1(n6993), .A2(n6992), .ZN(n9431) );
  NAND2_X1 U8761 ( .A1(n9428), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8762 ( .A1(n9431), .A2(n6994), .ZN(n7089) );
  INV_X1 U8763 ( .A(n7089), .ZN(n6996) );
  INV_X1 U8764 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9914) );
  MUX2_X1 U8765 ( .A(n9914), .B(P1_REG1_REG_2__SCAN_IN), .S(n7098), .Z(n7090)
         );
  NAND2_X1 U8766 ( .A1(n7098), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U8767 ( .B1(n6996), .B2(n7090), .A(n6995), .ZN(n9445) );
  INV_X1 U8768 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6997) );
  MUX2_X1 U8769 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6997), .S(n9439), .Z(n9446)
         );
  NAND2_X1 U8770 ( .A1(n9445), .A2(n9446), .ZN(n9444) );
  NAND2_X1 U8771 ( .A1(n9439), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U8772 ( .A1(n9444), .A2(n6998), .ZN(n7069) );
  INV_X1 U8773 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6999) );
  MUX2_X1 U8774 ( .A(n6999), .B(P1_REG1_REG_4__SCAN_IN), .S(n7077), .Z(n7068)
         );
  INV_X1 U8775 ( .A(n7068), .ZN(n7000) );
  NAND2_X1 U8776 ( .A1(n7069), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U8777 ( .A1(n7077), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8778 ( .A1(n7002), .A2(n7001), .ZN(n9460) );
  INV_X1 U8779 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7003) );
  MUX2_X1 U8780 ( .A(n7003), .B(P1_REG1_REG_5__SCAN_IN), .S(n9452), .Z(n9461)
         );
  NAND2_X1 U8781 ( .A1(n9460), .A2(n9461), .ZN(n9458) );
  NAND2_X1 U8782 ( .A1(n7004), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U8783 ( .A1(n9458), .A2(n7008), .ZN(n7007) );
  INV_X1 U8784 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7005) );
  MUX2_X1 U8785 ( .A(n7005), .B(P1_REG1_REG_6__SCAN_IN), .S(n7016), .Z(n7006)
         );
  NAND2_X1 U8786 ( .A1(n7007), .A2(n7006), .ZN(n7026) );
  MUX2_X1 U8787 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7005), .S(n7016), .Z(n7009)
         );
  NAND3_X1 U8788 ( .A1(n7009), .A2(n9458), .A3(n7008), .ZN(n7010) );
  AND3_X1 U8789 ( .A1(n9459), .A2(n7026), .A3(n7010), .ZN(n7011) );
  NOR2_X1 U8790 ( .A1(n7012), .A2(n7011), .ZN(n7015) );
  INV_X1 U8791 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7013) );
  NOR2_X1 U8792 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7013), .ZN(n7536) );
  AOI21_X1 U8793 ( .B1(n9455), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7536), .ZN(
        n7014) );
  OAI211_X1 U8794 ( .C1(n7016), .C2(n9843), .A(n7015), .B(n7014), .ZN(P1_U3249) );
  XNOR2_X1 U8795 ( .A(n7036), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7018) );
  NOR2_X1 U8796 ( .A1(n7019), .A2(n7018), .ZN(n7033) );
  AOI211_X1 U8797 ( .C1(n7019), .C2(n7018), .A(n7033), .B(n9471), .ZN(n7029)
         );
  NAND2_X1 U8798 ( .A1(n7020), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8799 ( .A1(n7026), .A2(n7025), .ZN(n7023) );
  INV_X1 U8800 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7021) );
  MUX2_X1 U8801 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7021), .S(n7036), .Z(n7022)
         );
  NAND2_X1 U8802 ( .A1(n7023), .A2(n7022), .ZN(n7053) );
  MUX2_X1 U8803 ( .A(n7021), .B(P1_REG1_REG_7__SCAN_IN), .S(n7036), .Z(n7024)
         );
  NAND3_X1 U8804 ( .A1(n7026), .A2(n7025), .A3(n7024), .ZN(n7027) );
  AND3_X1 U8805 ( .A1(n9459), .A2(n7053), .A3(n7027), .ZN(n7028) );
  NOR2_X1 U8806 ( .A1(n7029), .A2(n7028), .ZN(n7031) );
  AND2_X1 U8807 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7574) );
  AOI21_X1 U8808 ( .B1(n9455), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7574), .ZN(
        n7030) );
  OAI211_X1 U8809 ( .C1(n7032), .C2(n9843), .A(n7031), .B(n7030), .ZN(P1_U3250) );
  XOR2_X1 U8810 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7120), .Z(n7035) );
  XNOR2_X1 U8811 ( .A(n7062), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7057) );
  OAI21_X1 U8812 ( .B1(n7035), .B2(n7034), .A(n7116), .ZN(n7044) );
  INV_X1 U8813 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U8814 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9919), .S(n7120), .Z(n7038)
         );
  NAND2_X1 U8815 ( .A1(n7036), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7052) );
  INV_X1 U8816 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9917) );
  MUX2_X1 U8817 ( .A(n9917), .B(P1_REG1_REG_8__SCAN_IN), .S(n7062), .Z(n7051)
         );
  AOI21_X1 U8818 ( .B1(n7053), .B2(n7052), .A(n7051), .ZN(n7065) );
  AOI21_X1 U8819 ( .B1(n7062), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7065), .ZN(
        n7037) );
  NAND2_X1 U8820 ( .A1(n7037), .A2(n7038), .ZN(n7119) );
  OAI21_X1 U8821 ( .B1(n7038), .B2(n7037), .A(n7119), .ZN(n7039) );
  NAND2_X1 U8822 ( .A1(n7039), .A2(n9459), .ZN(n7041) );
  AND2_X1 U8823 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7876) );
  AOI21_X1 U8824 ( .B1(n9455), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7876), .ZN(
        n7040) );
  OAI211_X1 U8825 ( .C1(n9843), .C2(n7042), .A(n7041), .B(n7040), .ZN(n7043)
         );
  AOI21_X1 U8826 ( .B1(n7044), .B2(n9849), .A(n7043), .ZN(n7045) );
  INV_X1 U8827 ( .A(n7045), .ZN(P1_U3252) );
  INV_X1 U8828 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7046) );
  OAI222_X1 U8829 ( .A1(n8665), .A2(n7048), .B1(n8047), .B2(P2_U3151), .C1(
        n7046), .C2(n9216), .ZN(P2_U3283) );
  INV_X1 U8830 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7047) );
  OAI222_X1 U8831 ( .A1(P1_U3086), .A2(n9844), .B1(n9826), .B2(n7048), .C1(
        n7047), .C2(n8653), .ZN(P1_U3343) );
  NOR2_X1 U8832 ( .A1(n7190), .A2(n9686), .ZN(n7333) );
  AND2_X1 U8833 ( .A1(n5964), .A2(n7337), .ZN(n8453) );
  NOR2_X1 U8834 ( .A1(n7109), .A2(n8453), .ZN(n8407) );
  AOI21_X1 U8835 ( .B1(n9786), .B2(n9681), .A(n8407), .ZN(n7049) );
  AOI211_X1 U8836 ( .C1(n7331), .C2(n7108), .A(n7333), .B(n7049), .ZN(n7128)
         );
  NAND2_X1 U8837 ( .A1(n9923), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7050) );
  OAI21_X1 U8838 ( .B1(n7128), .B2(n9923), .A(n7050), .ZN(P1_U3522) );
  NAND3_X1 U8839 ( .A1(n7053), .A2(n7052), .A3(n7051), .ZN(n7054) );
  NAND2_X1 U8840 ( .A1(n9459), .A2(n7054), .ZN(n7064) );
  INV_X1 U8841 ( .A(n9843), .ZN(n9440) );
  INV_X1 U8842 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7055) );
  NOR2_X1 U8843 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7055), .ZN(n7861) );
  AOI211_X1 U8844 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n9471), .ZN(n7059)
         );
  NOR2_X1 U8845 ( .A1(n7861), .A2(n7059), .ZN(n7060) );
  OAI21_X1 U8846 ( .B1(n9852), .B2(n10095), .A(n7060), .ZN(n7061) );
  AOI21_X1 U8847 ( .B1(n9440), .B2(n7062), .A(n7061), .ZN(n7063) );
  OAI21_X1 U8848 ( .B1(n7065), .B2(n7064), .A(n7063), .ZN(P1_U3251) );
  INV_X1 U8849 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7067) );
  AND2_X1 U8850 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7172) );
  INV_X1 U8851 ( .A(n7172), .ZN(n7066) );
  OAI21_X1 U8852 ( .B1(n9852), .B2(n7067), .A(n7066), .ZN(n7076) );
  XOR2_X1 U8853 ( .A(n7069), .B(n7068), .Z(n7074) );
  OAI211_X1 U8854 ( .C1(n7072), .C2(n7071), .A(n9849), .B(n7070), .ZN(n7073)
         );
  OAI21_X1 U8855 ( .B1(n9845), .B2(n7074), .A(n7073), .ZN(n7075) );
  AOI211_X1 U8856 ( .C1(n7077), .C2(n9440), .A(n7076), .B(n7075), .ZN(n7086)
         );
  OAI21_X1 U8857 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(n7193) );
  NAND3_X1 U8858 ( .A1(n7193), .A2(n7081), .A3(n5926), .ZN(n7085) );
  AOI22_X1 U8859 ( .A1(n7083), .A2(n9433), .B1(n7082), .B2(n4796), .ZN(n7084)
         );
  NAND3_X1 U8860 ( .A1(n7085), .A2(P1_U3973), .A3(n7084), .ZN(n7099) );
  NAND2_X1 U8861 ( .A1(n7086), .A2(n7099), .ZN(P1_U3247) );
  INV_X1 U8862 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7088) );
  INV_X1 U8863 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7087) );
  OAI22_X1 U8864 ( .A1(n9852), .A2(n7088), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7087), .ZN(n7097) );
  XOR2_X1 U8865 ( .A(n7090), .B(n7089), .Z(n7095) );
  OAI211_X1 U8866 ( .C1(n7093), .C2(n7092), .A(n9849), .B(n7091), .ZN(n7094)
         );
  OAI21_X1 U8867 ( .B1(n9845), .B2(n7095), .A(n7094), .ZN(n7096) );
  AOI211_X1 U8868 ( .C1(n7098), .C2(n9440), .A(n7097), .B(n7096), .ZN(n7100)
         );
  NAND2_X1 U8869 ( .A1(n7100), .A2(n7099), .ZN(P1_U3245) );
  INV_X1 U8870 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7104) );
  INV_X1 U8871 ( .A(n7102), .ZN(n7103) );
  AOI22_X1 U8872 ( .A1(n7101), .A2(n7104), .B1(n7254), .B2(n7103), .ZN(
        P2_U3376) );
  OAI21_X1 U8873 ( .B1(n7107), .B2(n7106), .A(n7105), .ZN(n8277) );
  AOI211_X1 U8874 ( .C1(n7108), .C2(n7185), .A(n9707), .B(n7351), .ZN(n8280)
         );
  INV_X1 U8875 ( .A(n8277), .ZN(n7113) );
  AOI22_X1 U8876 ( .A1(n5560), .A2(n9698), .B1(n9696), .B2(n5964), .ZN(n7112)
         );
  NAND2_X1 U8877 ( .A1(n7110), .A2(n9701), .ZN(n7111) );
  OAI211_X1 U8878 ( .C1(n7113), .C2(n7346), .A(n7112), .B(n7111), .ZN(n8276)
         );
  AOI211_X1 U8879 ( .C1(n7114), .C2(n8277), .A(n8280), .B(n8276), .ZN(n7136)
         );
  INV_X1 U8880 ( .A(n9780), .ZN(n7720) );
  AOI22_X1 U8881 ( .A1(n7720), .A2(n7185), .B1(n9923), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7115) );
  OAI21_X1 U8882 ( .B1(n7136), .B2(n9923), .A(n7115), .ZN(P1_U3523) );
  XNOR2_X1 U8883 ( .A(n7219), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7118) );
  OAI21_X1 U8884 ( .B1(n7120), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7116), .ZN(
        n7117) );
  NOR2_X1 U8885 ( .A1(n7117), .A2(n7118), .ZN(n7218) );
  AOI211_X1 U8886 ( .C1(n7118), .C2(n7117), .A(n9471), .B(n7218), .ZN(n7127)
         );
  OAI21_X1 U8887 ( .B1(n7120), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7119), .ZN(
        n7122) );
  INV_X1 U8888 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9921) );
  MUX2_X1 U8889 ( .A(n9921), .B(P1_REG1_REG_10__SCAN_IN), .S(n7219), .Z(n7121)
         );
  NOR2_X1 U8890 ( .A1(n7122), .A2(n7121), .ZN(n7217) );
  AOI211_X1 U8891 ( .C1(n7122), .C2(n7121), .A(n9845), .B(n7217), .ZN(n7126)
         );
  NOR2_X1 U8892 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7123), .ZN(n9268) );
  AOI21_X1 U8893 ( .B1(n9455), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9268), .ZN(
        n7124) );
  OAI21_X1 U8894 ( .B1(n9843), .B2(n7211), .A(n7124), .ZN(n7125) );
  OR3_X1 U8895 ( .A1(n7127), .A2(n7126), .A3(n7125), .ZN(P1_U3253) );
  INV_X1 U8896 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7130) );
  OR2_X1 U8897 ( .A1(n7128), .A2(n9911), .ZN(n7129) );
  OAI21_X1 U8898 ( .B1(n9913), .B2(n7130), .A(n7129), .ZN(P1_U3453) );
  NAND2_X1 U8899 ( .A1(n7298), .A2(P2_U3893), .ZN(n7131) );
  OAI21_X1 U8900 ( .B1(P2_U3893), .B2(n4713), .A(n7131), .ZN(P2_U3492) );
  NAND2_X1 U8901 ( .A1(n8114), .A2(P2_U3893), .ZN(n7132) );
  OAI21_X1 U8902 ( .B1(P2_U3893), .B2(n5326), .A(n7132), .ZN(P2_U3500) );
  AND2_X1 U8903 ( .A1(n7101), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8904 ( .A1(n7101), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8905 ( .A1(n7101), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8906 ( .A1(n7101), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8907 ( .A1(n7101), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8908 ( .A1(n7101), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8909 ( .A1(n7101), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8910 ( .A1(n7101), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8911 ( .A1(n7101), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8912 ( .A1(n7101), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8913 ( .A1(n7101), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8914 ( .A1(n7101), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8915 ( .A1(n7101), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8916 ( .A1(n7101), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8917 ( .A1(n7101), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8918 ( .A1(n7101), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8919 ( .A1(n7101), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8920 ( .A1(n7101), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8921 ( .A1(n7101), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  INV_X1 U8922 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7133) );
  OAI22_X1 U8923 ( .A1(n9814), .A2(n8454), .B1(n9913), .B2(n7133), .ZN(n7134)
         );
  INV_X1 U8924 ( .A(n7134), .ZN(n7135) );
  OAI21_X1 U8925 ( .B1(n7136), .B2(n9911), .A(n7135), .ZN(P1_U3456) );
  INV_X1 U8926 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7138) );
  INV_X1 U8927 ( .A(n7137), .ZN(n7140) );
  OAI222_X1 U8928 ( .A1(n9216), .A2(n7138), .B1(n8665), .B2(n7140), .C1(
        P2_U3151), .C2(n9963), .ZN(P2_U3282) );
  INV_X1 U8929 ( .A(n7731), .ZN(n7728) );
  INV_X1 U8930 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7139) );
  OAI222_X1 U8931 ( .A1(n7728), .A2(P1_U3086), .B1(n9826), .B2(n7140), .C1(
        n7139), .C2(n8653), .ZN(P1_U3342) );
  INV_X1 U8932 ( .A(n9982), .ZN(n8842) );
  OAI21_X1 U8933 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7141), .A(n7148), .ZN(n7142) );
  OAI21_X1 U8934 ( .B1(n9993), .B2(n7143), .A(n7142), .ZN(n7144) );
  OAI21_X1 U8935 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7269), .A(n7144), .ZN(n7145) );
  AOI21_X1 U8936 ( .B1(n8842), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7145), .ZN(
        n7146) );
  OAI21_X1 U8937 ( .B1(n7147), .B2(n9983), .A(n7146), .ZN(P2_U3182) );
  XNOR2_X1 U8938 ( .A(n7149), .B(n7148), .ZN(n7166) );
  NOR2_X1 U8939 ( .A1(n9983), .A2(n7150), .ZN(n7164) );
  NAND2_X1 U8940 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  NAND2_X1 U8941 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  NAND2_X1 U8942 ( .A1(n9994), .A2(n7155), .ZN(n7162) );
  NAND2_X1 U8943 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  NAND2_X1 U8944 ( .A1(n7159), .A2(n7158), .ZN(n7160) );
  NAND2_X1 U8945 ( .A1(n9974), .A2(n7160), .ZN(n7161) );
  OAI211_X1 U8946 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7319), .A(n7162), .B(n7161), .ZN(n7163) );
  AOI211_X1 U8947 ( .C1(n8842), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7164), .B(
        n7163), .ZN(n7165) );
  OAI21_X1 U8948 ( .B1(n9958), .B2(n7166), .A(n7165), .ZN(P2_U3183) );
  NAND2_X1 U8949 ( .A1(n7167), .A2(n9383), .ZN(n7176) );
  AOI21_X1 U8950 ( .B1(n7168), .B2(n7170), .A(n7169), .ZN(n7175) );
  AOI22_X1 U8951 ( .A1(n9386), .A2(n9427), .B1(n9391), .B2(n9425), .ZN(n7174)
         );
  NOR2_X1 U8952 ( .A1(n9299), .A2(n7443), .ZN(n7171) );
  AOI211_X1 U8953 ( .C1(n9393), .C2(n7440), .A(n7172), .B(n7171), .ZN(n7173)
         );
  OAI211_X1 U8954 ( .C1(n7176), .C2(n7175), .A(n7174), .B(n7173), .ZN(P1_U3230) );
  INV_X1 U8955 ( .A(n7177), .ZN(n7179) );
  OAI222_X1 U8956 ( .A1(n9216), .A2(n7178), .B1(n8665), .B2(n7179), .C1(
        P2_U3151), .C2(n9984), .ZN(P2_U3281) );
  INV_X1 U8957 ( .A(n7841), .ZN(n7180) );
  OAI222_X1 U8958 ( .A1(n7180), .A2(P1_U3086), .B1(n9826), .B2(n7179), .C1(
        n10206), .C2(n8653), .ZN(P1_U3341) );
  NAND2_X1 U8959 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  XNOR2_X1 U8960 ( .A(n7181), .B(n7184), .ZN(n7189) );
  AOI22_X1 U8961 ( .A1(n7185), .A2(n9407), .B1(n9391), .B2(n5560), .ZN(n7188)
         );
  NAND2_X1 U8962 ( .A1(n7186), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9367) );
  AOI22_X1 U8963 ( .A1(n9386), .A2(n5964), .B1(n9367), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7187) );
  OAI211_X1 U8964 ( .C1(n7189), .C2(n9402), .A(n7188), .B(n7187), .ZN(P1_U3222) );
  OAI22_X1 U8965 ( .A1(n9376), .A2(n7190), .B1(n9299), .B2(n7337), .ZN(n7191)
         );
  AOI21_X1 U8966 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9367), .A(n7191), .ZN(
        n7192) );
  OAI21_X1 U8967 ( .B1(n9402), .B2(n7193), .A(n7192), .ZN(P1_U3232) );
  OAI21_X1 U8968 ( .B1(n7195), .B2(n8405), .A(n7194), .ZN(n7445) );
  INV_X1 U8969 ( .A(n7275), .ZN(n7196) );
  AOI211_X1 U8970 ( .C1(n7198), .C2(n7230), .A(n9707), .B(n7196), .ZN(n7439)
         );
  XNOR2_X1 U8971 ( .A(n8295), .B(n8405), .ZN(n7197) );
  OAI222_X1 U8972 ( .A1(n9684), .A2(n7342), .B1(n9686), .B2(n7360), .C1(n7197), 
        .C2(n9681), .ZN(n7438) );
  AOI211_X1 U8973 ( .C1(n9909), .C2(n7445), .A(n7439), .B(n7438), .ZN(n7203)
         );
  AOI22_X1 U8974 ( .A1(n7720), .A2(n7198), .B1(n9923), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U8975 ( .B1(n7203), .B2(n9923), .A(n7199), .ZN(P1_U3526) );
  INV_X1 U8976 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7200) );
  OAI22_X1 U8977 ( .A1(n9814), .A2(n7443), .B1(n9913), .B2(n7200), .ZN(n7201)
         );
  INV_X1 U8978 ( .A(n7201), .ZN(n7202) );
  OAI21_X1 U8979 ( .B1(n7203), .B2(n9911), .A(n7202), .ZN(P1_U3465) );
  OAI21_X1 U8980 ( .B1(n7205), .B2(n7204), .A(n7168), .ZN(n7209) );
  AOI22_X1 U8981 ( .A1(n9386), .A2(n5560), .B1(n9391), .B2(n9426), .ZN(n7207)
         );
  AND2_X1 U8982 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9447) );
  AOI21_X1 U8983 ( .B1(n9407), .B2(n7235), .A(n9447), .ZN(n7206) );
  OAI211_X1 U8984 ( .C1(n9355), .C2(P1_REG3_REG_3__SCAN_IN), .A(n7207), .B(
        n7206), .ZN(n7208) );
  AOI21_X1 U8985 ( .B1(n7209), .B2(n9383), .A(n7208), .ZN(n7210) );
  INV_X1 U8986 ( .A(n7210), .ZN(P1_U3218) );
  NOR2_X1 U8987 ( .A1(n7211), .A2(n9921), .ZN(n7215) );
  INV_X1 U8988 ( .A(n7215), .ZN(n7213) );
  INV_X1 U8989 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7380) );
  MUX2_X1 U8990 ( .A(n7380), .B(P1_REG1_REG_11__SCAN_IN), .S(n7375), .Z(n7212)
         );
  NAND2_X1 U8991 ( .A1(n7213), .A2(n7212), .ZN(n7216) );
  MUX2_X1 U8992 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7380), .S(n7375), .Z(n7214)
         );
  OAI21_X1 U8993 ( .B1(n7217), .B2(n7215), .A(n7214), .ZN(n7378) );
  OAI211_X1 U8994 ( .C1(n7217), .C2(n7216), .A(n7378), .B(n9459), .ZN(n7224)
         );
  AND2_X1 U8995 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9357) );
  XNOR2_X1 U8996 ( .A(n7375), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7220) );
  AOI211_X1 U8997 ( .C1(n7221), .C2(n7220), .A(n7374), .B(n9471), .ZN(n7222)
         );
  AOI211_X1 U8998 ( .C1(n9455), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9357), .B(
        n7222), .ZN(n7223) );
  OAI211_X1 U8999 ( .C1(n9843), .C2(n7379), .A(n7224), .B(n7223), .ZN(P1_U3254) );
  NAND2_X1 U9000 ( .A1(n8957), .A2(P2_U3893), .ZN(n7225) );
  OAI21_X1 U9001 ( .B1(P2_U3893), .B2(n5368), .A(n7225), .ZN(P2_U3514) );
  INV_X1 U9002 ( .A(n7226), .ZN(n7270) );
  INV_X1 U9003 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7227) );
  OAI222_X1 U9004 ( .A1(n8665), .A2(n7270), .B1(n8811), .B2(P2_U3151), .C1(
        n7227), .C2(n9216), .ZN(P2_U3280) );
  OAI21_X1 U9005 ( .B1(n7228), .B2(n8404), .A(n7229), .ZN(n9862) );
  INV_X1 U9006 ( .A(n7352), .ZN(n7231) );
  AOI211_X1 U9007 ( .C1(n7235), .C2(n7231), .A(n9707), .B(n4874), .ZN(n9854)
         );
  XOR2_X1 U9008 ( .A(n8404), .B(n7232), .Z(n7233) );
  AOI222_X1 U9009 ( .A1(n9701), .A2(n7233), .B1(n5560), .B2(n9696), .C1(n9426), 
        .C2(n9698), .ZN(n9865) );
  INV_X1 U9010 ( .A(n9865), .ZN(n7234) );
  AOI211_X1 U9011 ( .C1(n9909), .C2(n9862), .A(n9854), .B(n7234), .ZN(n7240)
         );
  AOI22_X1 U9012 ( .A1(n7720), .A2(n7235), .B1(n9923), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7236) );
  OAI21_X1 U9013 ( .B1(n7240), .B2(n9923), .A(n7236), .ZN(P1_U3525) );
  INV_X1 U9014 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7237) );
  OAI22_X1 U9015 ( .A1(n9814), .A2(n9860), .B1(n9913), .B2(n7237), .ZN(n7238)
         );
  INV_X1 U9016 ( .A(n7238), .ZN(n7239) );
  OAI21_X1 U9017 ( .B1(n7240), .B2(n9911), .A(n7239), .ZN(P1_U3462) );
  INV_X1 U9018 ( .A(n7260), .ZN(n7241) );
  NAND2_X1 U9019 ( .A1(n7251), .A2(n7241), .ZN(n7247) );
  OR2_X1 U9020 ( .A1(n7243), .A2(n7242), .ZN(n7246) );
  NAND4_X1 U9021 ( .A1(n7247), .A2(n7246), .A3(n7245), .A4(n7244), .ZN(n7248)
         );
  NAND2_X1 U9022 ( .A1(n7248), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7253) );
  INV_X1 U9023 ( .A(n7249), .ZN(n7250) );
  NAND2_X1 U9024 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  AND2_X1 U9025 ( .A1(n7253), .A2(n7252), .ZN(n7390) );
  AND2_X1 U9026 ( .A1(n7390), .A2(n7254), .ZN(n7320) );
  OR2_X1 U9027 ( .A1(n7261), .A2(n7255), .ZN(n7289) );
  INV_X1 U9028 ( .A(n7289), .ZN(n7256) );
  NAND2_X1 U9029 ( .A1(n7264), .A2(n10047), .ZN(n7259) );
  INV_X1 U9030 ( .A(n8723), .ZN(n8764) );
  OR2_X1 U9031 ( .A1(n7261), .A2(n7260), .ZN(n7266) );
  INV_X1 U9032 ( .A(n7262), .ZN(n7263) );
  NAND2_X1 U9033 ( .A1(n7264), .A2(n7263), .ZN(n7265) );
  OAI22_X1 U9034 ( .A1(n8764), .A2(n7301), .B1(n8725), .B2(n7452), .ZN(n7267)
         );
  AOI21_X1 U9035 ( .B1(n8733), .B2(n7298), .A(n7267), .ZN(n7268) );
  OAI21_X1 U9036 ( .B1(n7320), .B2(n7269), .A(n7268), .ZN(P2_U3172) );
  INV_X1 U9037 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10396) );
  OAI222_X1 U9038 ( .A1(n8653), .A2(n10396), .B1(P1_U3086), .B2(n4678), .C1(
        n7270), .C2(n9826), .ZN(P1_U3340) );
  NOR2_X1 U9039 ( .A1(n7297), .A2(n9036), .ZN(n7453) );
  INV_X1 U9040 ( .A(n10045), .ZN(n10056) );
  AOI21_X1 U9041 ( .B1(n8989), .B2(n10056), .A(n7452), .ZN(n7271) );
  AOI211_X1 U9042 ( .C1(n10047), .C2(n7456), .A(n7453), .B(n7271), .ZN(n7652)
         );
  NAND2_X1 U9043 ( .A1(n10068), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7272) );
  OAI21_X1 U9044 ( .B1(n7652), .B2(n10068), .A(n7272), .ZN(P2_U3459) );
  OAI21_X1 U9045 ( .B1(n7274), .B2(n7276), .A(n7273), .ZN(n7435) );
  AOI211_X1 U9046 ( .C1(n7283), .C2(n7275), .A(n9707), .B(n7367), .ZN(n7429)
         );
  INV_X1 U9047 ( .A(n7276), .ZN(n8411) );
  XNOR2_X1 U9048 ( .A(n7277), .B(n8411), .ZN(n7278) );
  OAI222_X1 U9049 ( .A1(n9684), .A2(n7279), .B1(n9686), .B2(n7571), .C1(n9681), 
        .C2(n7278), .ZN(n7428) );
  AOI211_X1 U9050 ( .C1(n9909), .C2(n7435), .A(n7429), .B(n7428), .ZN(n7285)
         );
  INV_X1 U9051 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7280) );
  OAI22_X1 U9052 ( .A1(n9814), .A2(n7433), .B1(n9913), .B2(n7280), .ZN(n7281)
         );
  INV_X1 U9053 ( .A(n7281), .ZN(n7282) );
  OAI21_X1 U9054 ( .B1(n7285), .B2(n9911), .A(n7282), .ZN(P1_U3468) );
  AOI22_X1 U9055 ( .A1(n7720), .A2(n7283), .B1(n9923), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7284) );
  OAI21_X1 U9056 ( .B1(n7285), .B2(n9923), .A(n7284), .ZN(P1_U3527) );
  INV_X1 U9057 ( .A(n7286), .ZN(n7322) );
  OAI222_X1 U9058 ( .A1(n8665), .A2(n7322), .B1(n8832), .B2(P2_U3151), .C1(
        n7287), .C2(n9216), .ZN(P2_U3279) );
  INV_X1 U9059 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7309) );
  NOR2_X2 U9060 ( .A1(n7289), .A2(n7288), .ZN(n8761) );
  OAI22_X1 U9061 ( .A1(n8735), .A2(n7297), .B1(n10024), .B2(n8764), .ZN(n7290)
         );
  AOI21_X1 U9062 ( .B1(n8733), .B2(n8778), .A(n7290), .ZN(n7308) );
  NOR2_X1 U9063 ( .A1(n7463), .A2(n7293), .ZN(n7294) );
  XNOR2_X1 U9064 ( .A(n7678), .B(n10024), .ZN(n7393) );
  XNOR2_X1 U9065 ( .A(n7393), .B(n7391), .ZN(n7305) );
  XNOR2_X1 U9066 ( .A(n7678), .B(n7953), .ZN(n7299) );
  INV_X1 U9067 ( .A(n7299), .ZN(n7296) );
  NAND2_X1 U9068 ( .A1(n7297), .A2(n7296), .ZN(n7303) );
  NAND2_X1 U9069 ( .A1(n7299), .A2(n7298), .ZN(n7300) );
  AND2_X2 U9070 ( .A1(n7303), .A2(n7300), .ZN(n7312) );
  NAND2_X1 U9071 ( .A1(n8568), .A2(n7301), .ZN(n7302) );
  NAND2_X1 U9072 ( .A1(n7461), .A2(n7302), .ZN(n7313) );
  NAND2_X1 U9073 ( .A1(n7312), .A2(n7313), .ZN(n7314) );
  NAND2_X1 U9074 ( .A1(n7314), .A2(n7303), .ZN(n7304) );
  NAND2_X1 U9075 ( .A1(n7304), .A2(n7305), .ZN(n7395) );
  OAI21_X1 U9076 ( .B1(n7305), .B2(n7304), .A(n7395), .ZN(n7306) );
  NAND2_X1 U9077 ( .A1(n7306), .A2(n8754), .ZN(n7307) );
  OAI211_X1 U9078 ( .C1(n7320), .C2(n7309), .A(n7308), .B(n7307), .ZN(P2_U3177) );
  INV_X1 U9079 ( .A(n8781), .ZN(n7310) );
  OAI22_X1 U9080 ( .A1(n8735), .A2(n7310), .B1(n7953), .B2(n8764), .ZN(n7311)
         );
  AOI21_X1 U9081 ( .B1(n8733), .B2(n8780), .A(n7311), .ZN(n7318) );
  OAI21_X1 U9082 ( .B1(n7312), .B2(n7313), .A(n7315), .ZN(n7316) );
  NAND2_X1 U9083 ( .A1(n7316), .A2(n8754), .ZN(n7317) );
  OAI211_X1 U9084 ( .C1(n7320), .C2(n7319), .A(n7318), .B(n7317), .ZN(P2_U3162) );
  INV_X1 U9085 ( .A(n8076), .ZN(n8070) );
  OAI222_X1 U9086 ( .A1(P1_U3086), .A2(n8070), .B1(n9826), .B2(n7322), .C1(
        n7321), .C2(n8653), .ZN(P1_U3339) );
  NAND2_X1 U9087 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  NOR2_X1 U9088 ( .A1(n7326), .A2(n7325), .ZN(n7327) );
  NAND2_X1 U9089 ( .A1(n7328), .A2(n7327), .ZN(n7329) );
  INV_X4 U9090 ( .A(n9670), .ZN(n9866) );
  AOI21_X1 U9091 ( .B1(n9853), .B2(n7331), .A(n9492), .ZN(n7338) );
  AOI22_X1 U9092 ( .A1(n9866), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9856), .ZN(n7336) );
  NOR3_X1 U9093 ( .A1(n8407), .A2(n7332), .A3(n7331), .ZN(n7334) );
  OAI21_X1 U9094 ( .B1(n7334), .B2(n7333), .A(n9670), .ZN(n7335) );
  OAI211_X1 U9095 ( .C1(n7338), .C2(n7337), .A(n7336), .B(n7335), .ZN(P1_U3293) );
  INV_X1 U9096 ( .A(n8403), .ZN(n7339) );
  XNOR2_X1 U9097 ( .A(n7340), .B(n7339), .ZN(n7344) );
  NAND2_X1 U9098 ( .A1(n5545), .A2(n9696), .ZN(n7341) );
  OAI21_X1 U9099 ( .B1(n7342), .B2(n9686), .A(n7341), .ZN(n7343) );
  AOI21_X1 U9100 ( .B1(n7344), .B2(n9701), .A(n7343), .ZN(n9879) );
  NAND2_X1 U9101 ( .A1(n7345), .A2(n5457), .ZN(n8275) );
  AND2_X1 U9102 ( .A1(n7346), .A2(n8275), .ZN(n7347) );
  OR2_X1 U9103 ( .A1(n7348), .A2(n8403), .ZN(n7349) );
  NAND2_X1 U9104 ( .A1(n7350), .A2(n7349), .ZN(n9877) );
  INV_X1 U9105 ( .A(n9707), .ZN(n8200) );
  OAI21_X1 U9106 ( .B1(n7351), .B2(n5559), .A(n8200), .ZN(n7353) );
  OR2_X1 U9107 ( .A1(n7353), .A2(n7352), .ZN(n9875) );
  NAND2_X1 U9108 ( .A1(n9492), .A2(n9366), .ZN(n7355) );
  AOI22_X1 U9109 ( .A1(n9866), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9856), .ZN(n7354) );
  OAI211_X1 U9110 ( .C1(n9875), .C2(n9495), .A(n7355), .B(n7354), .ZN(n7356)
         );
  AOI21_X1 U9111 ( .B1(n9863), .B2(n9877), .A(n7356), .ZN(n7357) );
  OAI21_X1 U9112 ( .B1(n9866), .B2(n9879), .A(n7357), .ZN(P1_U3291) );
  XNOR2_X1 U9113 ( .A(n7358), .B(n8412), .ZN(n7359) );
  NAND2_X1 U9114 ( .A1(n7359), .A2(n9701), .ZN(n7363) );
  OAI22_X1 U9115 ( .A1(n7360), .A2(n9684), .B1(n7858), .B2(n9686), .ZN(n7361)
         );
  INV_X1 U9116 ( .A(n7361), .ZN(n7362) );
  NAND2_X1 U9117 ( .A1(n7363), .A2(n7362), .ZN(n9883) );
  INV_X1 U9118 ( .A(n9883), .ZN(n7372) );
  OAI21_X1 U9119 ( .B1(n7365), .B2(n8412), .A(n7364), .ZN(n9885) );
  INV_X1 U9120 ( .A(n7489), .ZN(n7366) );
  OAI211_X1 U9121 ( .C1(n9882), .C2(n7367), .A(n7366), .B(n8200), .ZN(n9881)
         );
  AOI22_X1 U9122 ( .A1(n9866), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7537), .B2(
        n9856), .ZN(n7369) );
  NAND2_X1 U9123 ( .A1(n9492), .A2(n7534), .ZN(n7368) );
  OAI211_X1 U9124 ( .C1(n9881), .C2(n9495), .A(n7369), .B(n7368), .ZN(n7370)
         );
  AOI21_X1 U9125 ( .B1(n9885), .B2(n9863), .A(n7370), .ZN(n7371) );
  OAI21_X1 U9126 ( .B1(n9866), .B2(n7372), .A(n7371), .ZN(P1_U3287) );
  NAND2_X1 U9127 ( .A1(n7731), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7373) );
  OAI21_X1 U9128 ( .B1(n7731), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7373), .ZN(
        n7377) );
  INV_X1 U9129 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7816) );
  AOI22_X1 U9130 ( .A1(n7381), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7816), .B2(
        n9844), .ZN(n9839) );
  OAI21_X1 U9131 ( .B1(n7381), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9837), .ZN(
        n7376) );
  NOR2_X1 U9132 ( .A1(n7377), .A2(n7376), .ZN(n7730) );
  AOI211_X1 U9133 ( .C1(n7377), .C2(n7376), .A(n7730), .B(n9471), .ZN(n7389)
         );
  INV_X1 U9134 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9924) );
  OAI21_X1 U9135 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n9842) );
  AOI22_X1 U9136 ( .A1(n7381), .A2(n9924), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n9844), .ZN(n9841) );
  NOR2_X1 U9137 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  AOI21_X1 U9138 ( .B1(n9844), .B2(n9924), .A(n9840), .ZN(n7384) );
  INV_X1 U9139 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7382) );
  MUX2_X1 U9140 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7382), .S(n7731), .Z(n7383)
         );
  NAND2_X1 U9141 ( .A1(n7383), .A2(n7384), .ZN(n7727) );
  OAI211_X1 U9142 ( .C1(n7384), .C2(n7383), .A(n9459), .B(n7727), .ZN(n7387)
         );
  NAND2_X1 U9143 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n8144) );
  INV_X1 U9144 ( .A(n8144), .ZN(n7385) );
  AOI21_X1 U9145 ( .B1(n9455), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7385), .ZN(
        n7386) );
  OAI211_X1 U9146 ( .C1(n9843), .C2(n7728), .A(n7387), .B(n7386), .ZN(n7388)
         );
  OR2_X1 U9147 ( .A1(n7389), .A2(n7388), .ZN(P1_U3256) );
  NOR2_X1 U9148 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7560), .ZN(n9946) );
  OAI22_X1 U9149 ( .A1(n8735), .A2(n7391), .B1(n6303), .B2(n8757), .ZN(n7392)
         );
  AOI211_X1 U9150 ( .C1(n7561), .C2(n8723), .A(n9946), .B(n7392), .ZN(n7402)
         );
  OR2_X1 U9151 ( .A1(n7393), .A2(n8780), .ZN(n7394) );
  NAND2_X1 U9152 ( .A1(n7395), .A2(n7394), .ZN(n7396) );
  XNOR2_X1 U9153 ( .A(n8639), .B(n7958), .ZN(n7541) );
  XNOR2_X1 U9154 ( .A(n7541), .B(n8778), .ZN(n7397) );
  AOI21_X1 U9155 ( .B1(n7396), .B2(n7397), .A(n8725), .ZN(n7400) );
  INV_X1 U9156 ( .A(n7396), .ZN(n7399) );
  NAND2_X1 U9157 ( .A1(n7399), .A2(n7398), .ZN(n7543) );
  NAND2_X1 U9158 ( .A1(n7400), .A2(n7543), .ZN(n7401) );
  OAI211_X1 U9159 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8758), .A(n7402), .B(
        n7401), .ZN(P2_U3158) );
  INV_X1 U9160 ( .A(n7404), .ZN(n7405) );
  AOI21_X1 U9161 ( .B1(n7406), .B2(n7403), .A(n7405), .ZN(n7410) );
  AOI22_X1 U9162 ( .A1(n9386), .A2(n9426), .B1(n9391), .B2(n9424), .ZN(n7409)
         );
  AND2_X1 U9163 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9454) );
  NOR2_X1 U9164 ( .A1(n9299), .A2(n7433), .ZN(n7407) );
  AOI211_X1 U9165 ( .C1(n9393), .C2(n7430), .A(n9454), .B(n7407), .ZN(n7408)
         );
  OAI211_X1 U9166 ( .C1(n7410), .C2(n9402), .A(n7409), .B(n7408), .ZN(P1_U3227) );
  INV_X1 U9167 ( .A(n7411), .ZN(n7412) );
  OAI222_X1 U9168 ( .A1(n8653), .A2(n10422), .B1(n9826), .B2(n7412), .C1(
        P1_U3086), .C2(n4666), .ZN(P1_U3338) );
  OAI222_X1 U9169 ( .A1(n9216), .A2(n7413), .B1(n8665), .B2(n7412), .C1(
        P2_U3151), .C2(n8845), .ZN(P2_U3278) );
  NAND2_X1 U9170 ( .A1(n7414), .A2(n8304), .ZN(n7485) );
  NOR2_X1 U9171 ( .A1(n7485), .A2(n8313), .ZN(n7484) );
  INV_X1 U9172 ( .A(n7484), .ZN(n7416) );
  NAND2_X1 U9173 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  XNOR2_X1 U9174 ( .A(n7417), .B(n7420), .ZN(n7418) );
  OAI222_X1 U9175 ( .A1(n9686), .A2(n9265), .B1(n9684), .B2(n7858), .C1(n7418), 
        .C2(n9681), .ZN(n9889) );
  INV_X1 U9176 ( .A(n9889), .ZN(n7427) );
  OAI21_X1 U9177 ( .B1(n7421), .B2(n7420), .A(n7419), .ZN(n9891) );
  INV_X1 U9178 ( .A(n7491), .ZN(n7422) );
  INV_X1 U9179 ( .A(n7863), .ZN(n9888) );
  OAI211_X1 U9180 ( .C1(n7422), .C2(n9888), .A(n8200), .B(n7474), .ZN(n9887)
         );
  AOI22_X1 U9181 ( .A1(n9866), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7857), .B2(
        n9856), .ZN(n7424) );
  NAND2_X1 U9182 ( .A1(n9492), .A2(n7863), .ZN(n7423) );
  OAI211_X1 U9183 ( .C1(n9887), .C2(n9495), .A(n7424), .B(n7423), .ZN(n7425)
         );
  AOI21_X1 U9184 ( .B1(n9891), .B2(n9863), .A(n7425), .ZN(n7426) );
  OAI21_X1 U9185 ( .B1(n7427), .B2(n9866), .A(n7426), .ZN(P1_U3285) );
  INV_X1 U9186 ( .A(n7428), .ZN(n7437) );
  NAND2_X1 U9187 ( .A1(n7429), .A2(n9853), .ZN(n7432) );
  AOI22_X1 U9188 ( .A1(n9866), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7430), .B2(
        n9856), .ZN(n7431) );
  OAI211_X1 U9189 ( .C1(n7433), .C2(n9859), .A(n7432), .B(n7431), .ZN(n7434)
         );
  AOI21_X1 U9190 ( .B1(n7435), .B2(n9863), .A(n7434), .ZN(n7436) );
  OAI21_X1 U9191 ( .B1(n7437), .B2(n9866), .A(n7436), .ZN(P1_U3288) );
  INV_X1 U9192 ( .A(n7438), .ZN(n7447) );
  NAND2_X1 U9193 ( .A1(n7439), .A2(n9853), .ZN(n7442) );
  AOI22_X1 U9194 ( .A1(n9866), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7440), .B2(
        n9856), .ZN(n7441) );
  OAI211_X1 U9195 ( .C1(n7443), .C2(n9859), .A(n7442), .B(n7441), .ZN(n7444)
         );
  AOI21_X1 U9196 ( .B1(n9863), .B2(n7445), .A(n7444), .ZN(n7446) );
  OAI21_X1 U9197 ( .B1(n7447), .B2(n9866), .A(n7446), .ZN(P1_U3289) );
  NOR3_X1 U9198 ( .A1(n7452), .A2(n7451), .A3(n10047), .ZN(n7454) );
  OAI21_X1 U9199 ( .B1(n7454), .B2(n7453), .A(n10023), .ZN(n7458) );
  AOI22_X1 U9200 ( .A1(n10017), .A2(n7456), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10019), .ZN(n7457) );
  OAI211_X1 U9201 ( .C1(n5214), .C2(n10023), .A(n7458), .B(n7457), .ZN(
        P2_U3233) );
  INV_X1 U9202 ( .A(n7459), .ZN(n7460) );
  AOI21_X1 U9203 ( .B1(n7461), .B2(n6776), .A(n7460), .ZN(n7516) );
  NAND2_X1 U9204 ( .A1(n7463), .A2(n7462), .ZN(n8091) );
  INV_X1 U9205 ( .A(n8091), .ZN(n7624) );
  XNOR2_X1 U9206 ( .A(n6776), .B(n7464), .ZN(n7465) );
  AOI222_X1 U9207 ( .A1(n9060), .A2(n7465), .B1(n8780), .B2(n9057), .C1(n8781), 
        .C2(n9055), .ZN(n7515) );
  MUX2_X1 U9208 ( .A(n7156), .B(n7515), .S(n10023), .Z(n7468) );
  AOI22_X1 U9209 ( .A1(n10017), .A2(n7466), .B1(n10019), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7467) );
  OAI211_X1 U9210 ( .C1(n7516), .C2(n9069), .A(n7468), .B(n7467), .ZN(P2_U3232) );
  OAI21_X1 U9211 ( .B1(n7484), .B2(n8310), .A(n8314), .ZN(n7469) );
  XNOR2_X1 U9212 ( .A(n7469), .B(n7472), .ZN(n7470) );
  AOI22_X1 U9213 ( .A1(n7470), .A2(n9701), .B1(n9696), .B2(n9422), .ZN(n9894)
         );
  OAI21_X1 U9214 ( .B1(n7473), .B2(n7472), .A(n7471), .ZN(n9897) );
  INV_X1 U9215 ( .A(n7480), .ZN(n9895) );
  XNOR2_X1 U9216 ( .A(n7474), .B(n9895), .ZN(n7476) );
  NOR2_X1 U9217 ( .A1(n9353), .A2(n9686), .ZN(n7475) );
  AOI21_X1 U9218 ( .B1(n7476), .B2(n8200), .A(n7475), .ZN(n9893) );
  INV_X1 U9219 ( .A(n7477), .ZN(n7874) );
  NAND2_X1 U9220 ( .A1(n9866), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7478) );
  OAI21_X1 U9221 ( .B1(n9490), .B2(n7874), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9222 ( .B1(n7480), .B2(n9492), .A(n7479), .ZN(n7481) );
  OAI21_X1 U9223 ( .B1(n9893), .B2(n9495), .A(n7481), .ZN(n7482) );
  AOI21_X1 U9224 ( .B1(n9897), .B2(n9863), .A(n7482), .ZN(n7483) );
  OAI21_X1 U9225 ( .B1(n9866), .B2(n9894), .A(n7483), .ZN(P1_U3284) );
  AOI21_X1 U9226 ( .B1(n8313), .B2(n7485), .A(n7484), .ZN(n7486) );
  OAI222_X1 U9227 ( .A1(n9686), .A2(n7873), .B1(n9684), .B2(n7571), .C1(n9681), 
        .C2(n7486), .ZN(n7519) );
  INV_X1 U9228 ( .A(n7519), .ZN(n7496) );
  OAI21_X1 U9229 ( .B1(n7488), .B2(n8313), .A(n7487), .ZN(n7521) );
  OR2_X1 U9230 ( .A1(n7489), .A2(n7577), .ZN(n7490) );
  AND3_X1 U9231 ( .A1(n7491), .A2(n7490), .A3(n8200), .ZN(n7520) );
  NAND2_X1 U9232 ( .A1(n7520), .A2(n9853), .ZN(n7493) );
  AOI22_X1 U9233 ( .A1(n9866), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7570), .B2(
        n9856), .ZN(n7492) );
  OAI211_X1 U9234 ( .C1(n7577), .C2(n9859), .A(n7493), .B(n7492), .ZN(n7494)
         );
  AOI21_X1 U9235 ( .B1(n7521), .B2(n9863), .A(n7494), .ZN(n7495) );
  OAI21_X1 U9236 ( .B1(n7496), .B2(n9866), .A(n7495), .ZN(P1_U3286) );
  AOI21_X1 U9237 ( .B1(n7498), .B2(n7497), .A(n7585), .ZN(n7514) );
  AOI21_X1 U9238 ( .B1(n7501), .B2(n7500), .A(n7499), .ZN(n7502) );
  NOR2_X1 U9239 ( .A1(n8876), .A2(n7502), .ZN(n7511) );
  INV_X1 U9240 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10087) );
  AND3_X1 U9241 ( .A1(n7505), .A2(n7504), .A3(n7503), .ZN(n7506) );
  OAI21_X1 U9242 ( .B1(n7507), .B2(n7506), .A(n9974), .ZN(n7509) );
  INV_X1 U9243 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10453) );
  NOR2_X1 U9244 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10453), .ZN(n7709) );
  INV_X1 U9245 ( .A(n7709), .ZN(n7508) );
  OAI211_X1 U9246 ( .C1(n10087), .C2(n9982), .A(n7509), .B(n7508), .ZN(n7510)
         );
  AOI211_X1 U9247 ( .C1(n8796), .C2(n7512), .A(n7511), .B(n7510), .ZN(n7513)
         );
  OAI21_X1 U9248 ( .B1(n7514), .B2(n9958), .A(n7513), .ZN(P2_U3188) );
  OAI21_X1 U9249 ( .B1(n10056), .B2(n7516), .A(n7515), .ZN(n7955) );
  OAI22_X1 U9250 ( .A1(n9101), .A2(n7953), .B1(n10065), .B2(n7151), .ZN(n7517)
         );
  AOI21_X1 U9251 ( .B1(n7955), .B2(n10065), .A(n7517), .ZN(n7518) );
  INV_X1 U9252 ( .A(n7518), .ZN(P2_U3460) );
  AOI211_X1 U9253 ( .C1(n9909), .C2(n7521), .A(n7520), .B(n7519), .ZN(n7527)
         );
  INV_X1 U9254 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7522) );
  OAI22_X1 U9255 ( .A1(n9814), .A2(n7577), .B1(n9913), .B2(n7522), .ZN(n7523)
         );
  INV_X1 U9256 ( .A(n7523), .ZN(n7524) );
  OAI21_X1 U9257 ( .B1(n7527), .B2(n9911), .A(n7524), .ZN(P1_U3474) );
  AOI22_X1 U9258 ( .A1(n7720), .A2(n7525), .B1(n9923), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7526) );
  OAI21_X1 U9259 ( .B1(n7527), .B2(n9923), .A(n7526), .ZN(P1_U3529) );
  INV_X1 U9260 ( .A(n7528), .ZN(n7530) );
  NOR2_X1 U9261 ( .A1(n7530), .A2(n7529), .ZN(n7533) );
  INV_X1 U9262 ( .A(n7531), .ZN(n7532) );
  AOI21_X1 U9263 ( .B1(n7533), .B2(n7404), .A(n7532), .ZN(n7540) );
  AOI22_X1 U9264 ( .A1(n7534), .A2(n9407), .B1(n9386), .B2(n9425), .ZN(n7539)
         );
  NOR2_X1 U9265 ( .A1(n9376), .A2(n7858), .ZN(n7535) );
  AOI211_X1 U9266 ( .C1(n9393), .C2(n7537), .A(n7536), .B(n7535), .ZN(n7538)
         );
  OAI211_X1 U9267 ( .C1(n7540), .C2(n9402), .A(n7539), .B(n7538), .ZN(P1_U3239) );
  NAND2_X1 U9268 ( .A1(n7541), .A2(n8778), .ZN(n7542) );
  XNOR2_X1 U9269 ( .A(n8639), .B(n10018), .ZN(n7544) );
  NAND2_X1 U9270 ( .A1(n6303), .A2(n7544), .ZN(n7672) );
  INV_X1 U9271 ( .A(n7544), .ZN(n7545) );
  NAND2_X1 U9272 ( .A1(n7545), .A2(n8777), .ZN(n7546) );
  AND2_X1 U9273 ( .A1(n7672), .A2(n7546), .ZN(n7668) );
  NAND2_X1 U9274 ( .A1(n7670), .A2(n7668), .ZN(n7642) );
  OAI21_X1 U9275 ( .B1(n7670), .B2(n7668), .A(n7642), .ZN(n7547) );
  NAND2_X1 U9276 ( .A1(n7547), .A2(n8754), .ZN(n7552) );
  INV_X1 U9277 ( .A(n8778), .ZN(n7548) );
  INV_X1 U9278 ( .A(n8776), .ZN(n7707) );
  OAI22_X1 U9279 ( .A1(n8735), .A2(n7548), .B1(n7707), .B2(n8757), .ZN(n7549)
         );
  AOI211_X1 U9280 ( .C1(n10018), .C2(n8723), .A(n7550), .B(n7549), .ZN(n7551)
         );
  OAI211_X1 U9281 ( .C1(n10016), .C2(n8758), .A(n7552), .B(n7551), .ZN(
        P2_U3170) );
  INV_X1 U9282 ( .A(n7553), .ZN(n7555) );
  INV_X1 U9283 ( .A(n7630), .ZN(n7554) );
  AOI21_X1 U9284 ( .B1(n7555), .B2(n7556), .A(n7554), .ZN(n7579) );
  XNOR2_X1 U9285 ( .A(n7557), .B(n7556), .ZN(n7558) );
  AOI222_X1 U9286 ( .A1(n9060), .A2(n7558), .B1(n8780), .B2(n9055), .C1(n8777), 
        .C2(n9057), .ZN(n7578) );
  MUX2_X1 U9287 ( .A(n7559), .B(n7578), .S(n10023), .Z(n7563) );
  AOI22_X1 U9288 ( .A1(n10017), .A2(n7561), .B1(n10019), .B2(n7560), .ZN(n7562) );
  OAI211_X1 U9289 ( .C1(n7579), .C2(n9069), .A(n7563), .B(n7562), .ZN(P2_U3230) );
  INV_X1 U9290 ( .A(n7564), .ZN(n7598) );
  OAI222_X1 U9291 ( .A1(n8665), .A2(n7598), .B1(n8858), .B2(P2_U3151), .C1(
        n7565), .C2(n9216), .ZN(P2_U3277) );
  OAI21_X1 U9292 ( .B1(n7568), .B2(n7566), .A(n7567), .ZN(n7569) );
  NAND2_X1 U9293 ( .A1(n7569), .A2(n9383), .ZN(n7576) );
  INV_X1 U9294 ( .A(n7570), .ZN(n7572) );
  OAI22_X1 U9295 ( .A1(n9355), .A2(n7572), .B1(n9396), .B2(n7571), .ZN(n7573)
         );
  AOI211_X1 U9296 ( .C1(n9391), .C2(n9422), .A(n7574), .B(n7573), .ZN(n7575)
         );
  OAI211_X1 U9297 ( .C1(n7577), .C2(n9299), .A(n7576), .B(n7575), .ZN(P1_U3213) );
  OAI21_X1 U9298 ( .B1(n7579), .B2(n10056), .A(n7578), .ZN(n7960) );
  OAI22_X1 U9299 ( .A1(n9101), .A2(n7958), .B1(n10065), .B2(n6284), .ZN(n7580)
         );
  AOI21_X1 U9300 ( .B1(n7960), .B2(n10065), .A(n7580), .ZN(n7581) );
  INV_X1 U9301 ( .A(n7581), .ZN(P2_U3462) );
  XNOR2_X1 U9302 ( .A(n7582), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7597) );
  INV_X1 U9303 ( .A(n8784), .ZN(n7587) );
  NOR3_X1 U9304 ( .A1(n7585), .A2(n7584), .A3(n7583), .ZN(n7586) );
  OAI21_X1 U9305 ( .B1(n7587), .B2(n7586), .A(n9993), .ZN(n7596) );
  INV_X1 U9306 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10090) );
  INV_X1 U9307 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10457) );
  NOR2_X1 U9308 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10457), .ZN(n7688) );
  INV_X1 U9309 ( .A(n7688), .ZN(n7588) );
  OAI21_X1 U9310 ( .B1(n9982), .B2(n10090), .A(n7588), .ZN(n7593) );
  AOI21_X1 U9311 ( .B1(n10012), .B2(n7589), .A(n7590), .ZN(n7591) );
  NOR2_X1 U9312 ( .A1(n7591), .A2(n9998), .ZN(n7592) );
  AOI211_X1 U9313 ( .C1(n8796), .C2(n7594), .A(n7593), .B(n7592), .ZN(n7595)
         );
  OAI211_X1 U9314 ( .C1(n7597), .C2(n8876), .A(n7596), .B(n7595), .ZN(P2_U3189) );
  INV_X1 U9315 ( .A(n8262), .ZN(n9480) );
  OAI222_X1 U9316 ( .A1(n8653), .A2(n10214), .B1(P1_U3086), .B2(n9480), .C1(
        n7598), .C2(n9826), .ZN(P1_U3337) );
  OAI21_X1 U9317 ( .B1(n7601), .B2(n7600), .A(n7599), .ZN(n7603) );
  OAI22_X1 U9318 ( .A1(n7809), .A2(n9686), .B1(n9265), .B2(n9684), .ZN(n7602)
         );
  AOI21_X1 U9319 ( .B1(n7603), .B2(n9701), .A(n7602), .ZN(n9900) );
  OAI21_X1 U9320 ( .B1(n7605), .B2(n8419), .A(n7604), .ZN(n9902) );
  NAND2_X1 U9321 ( .A1(n9902), .A2(n9863), .ZN(n7615) );
  INV_X1 U9322 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7607) );
  INV_X1 U9323 ( .A(n7606), .ZN(n9266) );
  OAI22_X1 U9324 ( .A1(n9670), .A2(n7607), .B1(n9266), .B2(n9490), .ZN(n7612)
         );
  INV_X1 U9325 ( .A(n7608), .ZN(n7610) );
  INV_X1 U9326 ( .A(n7609), .ZN(n7662) );
  OAI211_X1 U9327 ( .C1(n5670), .C2(n7610), .A(n7662), .B(n8200), .ZN(n9899)
         );
  NOR2_X1 U9328 ( .A1(n9899), .A2(n9495), .ZN(n7611) );
  AOI211_X1 U9329 ( .C1(n9492), .C2(n7613), .A(n7612), .B(n7611), .ZN(n7614)
         );
  OAI211_X1 U9330 ( .C1(n9866), .C2(n9900), .A(n7615), .B(n7614), .ZN(P1_U3283) );
  OAI21_X1 U9331 ( .B1(n7617), .B2(n7618), .A(n7616), .ZN(n10027) );
  OAI22_X1 U9332 ( .A1(n10024), .A2(n9063), .B1(n7309), .B2(n9061), .ZN(n7623)
         );
  XNOR2_X1 U9333 ( .A(n7619), .B(n7618), .ZN(n7622) );
  NAND2_X1 U9334 ( .A1(n10027), .A2(n8102), .ZN(n7621) );
  AOI22_X1 U9335 ( .A1(n9055), .A2(n7298), .B1(n8778), .B2(n9057), .ZN(n7620)
         );
  OAI211_X1 U9336 ( .C1(n8989), .C2(n7622), .A(n7621), .B(n7620), .ZN(n10025)
         );
  AOI211_X1 U9337 ( .C1(n7624), .C2(n10027), .A(n7623), .B(n10025), .ZN(n7625)
         );
  OR2_X1 U9338 ( .A1(n7625), .A2(n8033), .ZN(n7626) );
  OAI21_X1 U9339 ( .B1(n5152), .B2(n10023), .A(n7626), .ZN(P2_U3231) );
  INV_X1 U9340 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10192) );
  INV_X1 U9341 ( .A(n8880), .ZN(n7627) );
  NAND2_X1 U9342 ( .A1(n7627), .A2(P2_U3893), .ZN(n7628) );
  OAI21_X1 U9343 ( .B1(P2_U3893), .B2(n10192), .A(n7628), .ZN(P2_U3522) );
  NAND3_X1 U9344 ( .A1(n7630), .A2(n7636), .A3(n7629), .ZN(n7631) );
  AND2_X1 U9345 ( .A1(n7632), .A2(n7631), .ZN(n10014) );
  NAND2_X1 U9346 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  XNOR2_X1 U9347 ( .A(n7636), .B(n7635), .ZN(n7637) );
  AOI222_X1 U9348 ( .A1(n9060), .A2(n7637), .B1(n8778), .B2(n9055), .C1(n8776), 
        .C2(n9057), .ZN(n10013) );
  OAI21_X1 U9349 ( .B1(n10056), .B2(n10014), .A(n10013), .ZN(n7945) );
  OAI22_X1 U9350 ( .A1(n9101), .A2(n6302), .B1(n10065), .B2(n6295), .ZN(n7638)
         );
  AOI21_X1 U9351 ( .B1(n7945), .B2(n10065), .A(n7638), .ZN(n7639) );
  INV_X1 U9352 ( .A(n7639), .ZN(P2_U3463) );
  INV_X1 U9353 ( .A(n7642), .ZN(n7641) );
  INV_X1 U9354 ( .A(n7672), .ZN(n7640) );
  INV_X2 U9355 ( .A(n8568), .ZN(n8645) );
  XNOR2_X1 U9356 ( .A(n8645), .B(n6578), .ZN(n7674) );
  XNOR2_X1 U9357 ( .A(n7674), .B(n8776), .ZN(n7671) );
  NOR3_X1 U9358 ( .A1(n7641), .A2(n7640), .A3(n7671), .ZN(n7645) );
  NAND2_X1 U9359 ( .A1(n7642), .A2(n7672), .ZN(n7643) );
  NAND2_X1 U9360 ( .A1(n7643), .A2(n7671), .ZN(n7702) );
  INV_X1 U9361 ( .A(n7702), .ZN(n7644) );
  OAI21_X1 U9362 ( .B1(n7645), .B2(n7644), .A(n8754), .ZN(n7649) );
  INV_X1 U9363 ( .A(n8775), .ZN(n7686) );
  OAI22_X1 U9364 ( .A1(n8735), .A2(n6303), .B1(n7686), .B2(n8757), .ZN(n7646)
         );
  AOI211_X1 U9365 ( .C1(n6578), .C2(n8723), .A(n7647), .B(n7646), .ZN(n7648)
         );
  OAI211_X1 U9366 ( .C1(n7697), .C2(n8758), .A(n7649), .B(n7648), .ZN(P2_U3167) );
  INV_X1 U9367 ( .A(n7650), .ZN(n8654) );
  OAI222_X1 U9368 ( .A1(n9216), .A2(n7651), .B1(n8665), .B2(n8654), .C1(
        P2_U3151), .C2(n8869), .ZN(P2_U3276) );
  INV_X1 U9369 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7654) );
  OR2_X1 U9370 ( .A1(n7652), .A2(n10061), .ZN(n7653) );
  OAI21_X1 U9371 ( .B1(n7654), .B2(n10052), .A(n7653), .ZN(P2_U3390) );
  OAI21_X1 U9372 ( .B1(n7656), .B2(n7657), .A(n7655), .ZN(n7715) );
  INV_X1 U9373 ( .A(n7715), .ZN(n7667) );
  XNOR2_X1 U9374 ( .A(n7658), .B(n5917), .ZN(n7659) );
  NAND2_X1 U9375 ( .A1(n7659), .A2(n9701), .ZN(n7661) );
  AOI22_X1 U9376 ( .A1(n9421), .A2(n9696), .B1(n9698), .B2(n9419), .ZN(n7660)
         );
  NAND2_X1 U9377 ( .A1(n7661), .A2(n7660), .ZN(n7713) );
  AOI211_X1 U9378 ( .C1(n9358), .C2(n7662), .A(n9707), .B(n7818), .ZN(n7714)
         );
  NAND2_X1 U9379 ( .A1(n7714), .A2(n9853), .ZN(n7664) );
  AOI22_X1 U9380 ( .A1(n9866), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9352), .B2(
        n9856), .ZN(n7663) );
  OAI211_X1 U9381 ( .C1(n7717), .C2(n9859), .A(n7664), .B(n7663), .ZN(n7665)
         );
  AOI21_X1 U9382 ( .B1(n9670), .B2(n7713), .A(n7665), .ZN(n7666) );
  OAI21_X1 U9383 ( .B1(n7667), .B2(n9693), .A(n7666), .ZN(P1_U3282) );
  AND2_X1 U9384 ( .A1(n7668), .A2(n7671), .ZN(n7669) );
  NAND2_X1 U9385 ( .A1(n7670), .A2(n7669), .ZN(n7749) );
  INV_X1 U9386 ( .A(n7671), .ZN(n7673) );
  OR2_X1 U9387 ( .A1(n7673), .A2(n7672), .ZN(n7747) );
  AND2_X1 U9388 ( .A1(n7749), .A2(n7747), .ZN(n7676) );
  INV_X2 U9389 ( .A(n7678), .ZN(n8568) );
  INV_X2 U9390 ( .A(n8568), .ZN(n8623) );
  XNOR2_X1 U9391 ( .A(n10029), .B(n8623), .ZN(n7677) );
  XNOR2_X1 U9392 ( .A(n7677), .B(n8775), .ZN(n7703) );
  INV_X1 U9393 ( .A(n7703), .ZN(n7675) );
  NAND2_X1 U9394 ( .A1(n7707), .A2(n7674), .ZN(n7701) );
  AND2_X1 U9395 ( .A1(n7675), .A2(n7701), .ZN(n7745) );
  NAND2_X1 U9396 ( .A1(n7676), .A2(n7745), .ZN(n7682) );
  NAND2_X1 U9397 ( .A1(n7677), .A2(n8775), .ZN(n7681) );
  AND2_X1 U9398 ( .A1(n7682), .A2(n7681), .ZN(n7684) );
  XNOR2_X1 U9399 ( .A(n7678), .B(n7948), .ZN(n7679) );
  OR2_X1 U9400 ( .A1(n7679), .A2(n8774), .ZN(n7744) );
  NAND2_X1 U9401 ( .A1(n7679), .A2(n8774), .ZN(n7680) );
  AND2_X1 U9402 ( .A1(n7744), .A2(n7680), .ZN(n7683) );
  NAND2_X1 U9403 ( .A1(n7682), .A2(n7750), .ZN(n7742) );
  OAI21_X1 U9404 ( .B1(n7684), .B2(n7683), .A(n7742), .ZN(n7685) );
  NAND2_X1 U9405 ( .A1(n7685), .A2(n8754), .ZN(n7690) );
  OAI22_X1 U9406 ( .A1(n8735), .A2(n7686), .B1(n4688), .B2(n8757), .ZN(n7687)
         );
  AOI211_X1 U9407 ( .C1(n10008), .C2(n8723), .A(n7688), .B(n7687), .ZN(n7689)
         );
  OAI211_X1 U9408 ( .C1(n10007), .C2(n8758), .A(n7690), .B(n7689), .ZN(
        P2_U3153) );
  XOR2_X1 U9409 ( .A(n7694), .B(n7691), .Z(n7724) );
  AND2_X1 U9410 ( .A1(n7693), .A2(n7692), .ZN(n7763) );
  XOR2_X1 U9411 ( .A(n7763), .B(n7694), .Z(n7695) );
  AOI222_X1 U9412 ( .A1(n9060), .A2(n7695), .B1(n8775), .B2(n9057), .C1(n8777), 
        .C2(n9055), .ZN(n7723) );
  MUX2_X1 U9413 ( .A(n7696), .B(n7723), .S(n10023), .Z(n7700) );
  INV_X1 U9414 ( .A(n7697), .ZN(n7698) );
  AOI22_X1 U9415 ( .A1(n10017), .A2(n6578), .B1(n10019), .B2(n7698), .ZN(n7699) );
  OAI211_X1 U9416 ( .C1(n7724), .C2(n9069), .A(n7700), .B(n7699), .ZN(P2_U3228) );
  NAND2_X1 U9417 ( .A1(n7702), .A2(n7701), .ZN(n7704) );
  AOI21_X1 U9418 ( .B1(n7704), .B2(n7703), .A(n8725), .ZN(n7706) );
  OR2_X1 U9419 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  NAND2_X1 U9420 ( .A1(n7706), .A2(n7705), .ZN(n7712) );
  OAI22_X1 U9421 ( .A1(n8735), .A2(n7707), .B1(n4756), .B2(n8757), .ZN(n7708)
         );
  AOI211_X1 U9422 ( .C1(n7710), .C2(n8723), .A(n7709), .B(n7708), .ZN(n7711)
         );
  OAI211_X1 U9423 ( .C1(n7769), .C2(n8758), .A(n7712), .B(n7711), .ZN(P2_U3179) );
  AOI211_X1 U9424 ( .C1(n7715), .C2(n9909), .A(n7714), .B(n7713), .ZN(n7722)
         );
  INV_X1 U9425 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7716) );
  OAI22_X1 U9426 ( .A1(n7717), .A2(n9814), .B1(n9913), .B2(n7716), .ZN(n7718)
         );
  INV_X1 U9427 ( .A(n7718), .ZN(n7719) );
  OAI21_X1 U9428 ( .B1(n7722), .B2(n9911), .A(n7719), .ZN(P1_U3486) );
  AOI22_X1 U9429 ( .A1(n9358), .A2(n7720), .B1(n9923), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7721) );
  OAI21_X1 U9430 ( .B1(n7722), .B2(n9923), .A(n7721), .ZN(P1_U3533) );
  OAI21_X1 U9431 ( .B1(n10056), .B2(n7724), .A(n7723), .ZN(n7941) );
  OAI22_X1 U9432 ( .A1(n9101), .A2(n7939), .B1(n10065), .B2(n6917), .ZN(n7725)
         );
  AOI21_X1 U9433 ( .B1(n7941), .B2(n10065), .A(n7725), .ZN(n7726) );
  INV_X1 U9434 ( .A(n7726), .ZN(P2_U3464) );
  OAI21_X1 U9435 ( .B1(n7728), .B2(n7382), .A(n7727), .ZN(n7843) );
  XOR2_X1 U9436 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7841), .Z(n7842) );
  XNOR2_X1 U9437 ( .A(n7843), .B(n7842), .ZN(n7741) );
  INV_X1 U9438 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7738) );
  NOR2_X1 U9439 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7729), .ZN(n9245) );
  AOI21_X1 U9440 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7731), .A(n7730), .ZN(
        n7735) );
  NAND2_X1 U9441 ( .A1(n7841), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7845) );
  OR2_X1 U9442 ( .A1(n7841), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U9443 ( .A1(n7845), .A2(n7732), .ZN(n7734) );
  INV_X1 U9444 ( .A(n7846), .ZN(n7733) );
  AOI211_X1 U9445 ( .C1(n7735), .C2(n7734), .A(n7733), .B(n9471), .ZN(n7736)
         );
  NOR2_X1 U9446 ( .A1(n9245), .A2(n7736), .ZN(n7737) );
  OAI21_X1 U9447 ( .B1(n9852), .B2(n7738), .A(n7737), .ZN(n7739) );
  AOI21_X1 U9448 ( .B1(n9440), .B2(n7841), .A(n7739), .ZN(n7740) );
  OAI21_X1 U9449 ( .B1(n7741), .B2(n9845), .A(n7740), .ZN(P1_U3257) );
  INV_X1 U9450 ( .A(n7742), .ZN(n7743) );
  INV_X1 U9451 ( .A(n7744), .ZN(n7751) );
  XNOR2_X1 U9452 ( .A(n8030), .B(n8645), .ZN(n7788) );
  XNOR2_X1 U9453 ( .A(n7788), .B(n8773), .ZN(n7752) );
  NOR3_X1 U9454 ( .A1(n7743), .A2(n7751), .A3(n7752), .ZN(n7756) );
  AND2_X1 U9455 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  AND2_X1 U9456 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  NAND2_X1 U9457 ( .A1(n7749), .A2(n7748), .ZN(n7754) );
  AND2_X1 U9458 ( .A1(n4540), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U9459 ( .A1(n7754), .A2(n7753), .ZN(n7790) );
  INV_X1 U9460 ( .A(n7790), .ZN(n7755) );
  OAI21_X1 U9461 ( .B1(n7756), .B2(n7755), .A(n8754), .ZN(n7761) );
  INV_X1 U9462 ( .A(n8114), .ZN(n7758) );
  INV_X1 U9463 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U9464 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10201), .ZN(n8787) );
  AOI21_X1 U9465 ( .B1(n8761), .B2(n8774), .A(n8787), .ZN(n7757) );
  OAI21_X1 U9466 ( .B1(n7758), .B2(n8757), .A(n7757), .ZN(n7759) );
  AOI21_X1 U9467 ( .B1(n8030), .B2(n8723), .A(n7759), .ZN(n7760) );
  OAI211_X1 U9468 ( .C1(n8025), .C2(n8758), .A(n7761), .B(n7760), .ZN(P2_U3161) );
  OR2_X1 U9469 ( .A1(n7763), .A2(n7762), .ZN(n7881) );
  NAND2_X1 U9470 ( .A1(n7881), .A2(n7764), .ZN(n7765) );
  XNOR2_X1 U9471 ( .A(n7765), .B(n7768), .ZN(n7766) );
  AOI222_X1 U9472 ( .A1(n9060), .A2(n7766), .B1(n8774), .B2(n9057), .C1(n8776), 
        .C2(n9055), .ZN(n10028) );
  XOR2_X1 U9473 ( .A(n7768), .B(n7767), .Z(n10031) );
  NOR2_X1 U9474 ( .A1(n10023), .A2(n6314), .ZN(n7771) );
  OAI22_X1 U9475 ( .A1(n8984), .A2(n10029), .B1(n7769), .B2(n9061), .ZN(n7770)
         );
  AOI211_X1 U9476 ( .C1(n10031), .C2(n9023), .A(n7771), .B(n7770), .ZN(n7772)
         );
  OAI21_X1 U9477 ( .B1(n8033), .B2(n10028), .A(n7772), .ZN(P2_U3227) );
  AOI21_X1 U9478 ( .B1(n8107), .B2(n7774), .A(n7773), .ZN(n7787) );
  INV_X1 U9479 ( .A(n7828), .ZN(n7778) );
  NOR3_X1 U9480 ( .A1(n8786), .A2(n7776), .A3(n7775), .ZN(n7777) );
  OAI21_X1 U9481 ( .B1(n7778), .B2(n7777), .A(n9993), .ZN(n7786) );
  OAI21_X1 U9482 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7780), .A(n7779), .ZN(
        n7784) );
  NOR2_X1 U9483 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6215), .ZN(n7793) );
  AOI21_X1 U9484 ( .B1(n8842), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7793), .ZN(
        n7781) );
  OAI21_X1 U9485 ( .B1(n7782), .B2(n9983), .A(n7781), .ZN(n7783) );
  AOI21_X1 U9486 ( .B1(n7784), .B2(n9994), .A(n7783), .ZN(n7785) );
  OAI211_X1 U9487 ( .C1(n7787), .C2(n9998), .A(n7786), .B(n7785), .ZN(P2_U3191) );
  NAND2_X1 U9488 ( .A1(n7788), .A2(n4688), .ZN(n7789) );
  AND2_X2 U9489 ( .A1(n7790), .A2(n7789), .ZN(n7792) );
  XNOR2_X1 U9490 ( .A(n8109), .B(n8645), .ZN(n7977) );
  XNOR2_X1 U9491 ( .A(n7977), .B(n8114), .ZN(n7791) );
  OAI211_X1 U9492 ( .C1(n7792), .C2(n7791), .A(n7980), .B(n8754), .ZN(n7799)
         );
  AOI21_X1 U9493 ( .B1(n8761), .B2(n8773), .A(n7793), .ZN(n7796) );
  INV_X1 U9494 ( .A(n8106), .ZN(n7794) );
  NAND2_X1 U9495 ( .A1(n8747), .A2(n7794), .ZN(n7795) );
  OAI211_X1 U9496 ( .C1(n8100), .C2(n8757), .A(n7796), .B(n7795), .ZN(n7797)
         );
  INV_X1 U9497 ( .A(n7797), .ZN(n7798) );
  OAI211_X1 U9498 ( .C1(n10033), .C2(n8764), .A(n7799), .B(n7798), .ZN(
        P2_U3171) );
  INV_X1 U9499 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U9500 ( .A1(n7802), .A2(n8010), .ZN(n7801) );
  OAI211_X1 U9501 ( .C1(n10482), .C2(n8653), .A(n7801), .B(n7800), .ZN(
        P1_U3335) );
  INV_X1 U9502 ( .A(n7802), .ZN(n7806) );
  OAI222_X1 U9503 ( .A1(n8665), .A2(n7806), .B1(n7805), .B2(P2_U3151), .C1(
        n7803), .C2(n9216), .ZN(P2_U3275) );
  OAI21_X1 U9504 ( .B1(n8421), .B2(n7808), .A(n7807), .ZN(n7811) );
  OAI22_X1 U9505 ( .A1(n7809), .A2(n9684), .B1(n9242), .B2(n9686), .ZN(n7810)
         );
  AOI21_X1 U9506 ( .B1(n7811), .B2(n9701), .A(n7810), .ZN(n9905) );
  OAI21_X1 U9507 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n9910) );
  NAND2_X1 U9508 ( .A1(n9910), .A2(n9863), .ZN(n7822) );
  INV_X1 U9509 ( .A(n8055), .ZN(n7815) );
  OAI22_X1 U9510 ( .A1(n9670), .A2(n7816), .B1(n7815), .B2(n9490), .ZN(n7820)
         );
  INV_X1 U9511 ( .A(n7817), .ZN(n7900) );
  OAI211_X1 U9512 ( .C1(n9907), .C2(n7818), .A(n7900), .B(n8200), .ZN(n9904)
         );
  NOR2_X1 U9513 ( .A1(n9904), .A2(n9495), .ZN(n7819) );
  AOI211_X1 U9514 ( .C1(n9492), .C2(n8058), .A(n7820), .B(n7819), .ZN(n7821)
         );
  OAI211_X1 U9515 ( .C1(n9866), .C2(n9905), .A(n7822), .B(n7821), .ZN(P1_U3281) );
  AOI21_X1 U9516 ( .B1(n7825), .B2(n7824), .A(n7823), .ZN(n7840) );
  AND3_X1 U9517 ( .A1(n7828), .A2(n7827), .A3(n7826), .ZN(n7829) );
  OAI21_X1 U9518 ( .B1(n7830), .B2(n7829), .A(n9993), .ZN(n7839) );
  OAI21_X1 U9519 ( .B1(n7833), .B2(n7832), .A(n7831), .ZN(n7837) );
  AND2_X1 U9520 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8113) );
  AOI21_X1 U9521 ( .B1(n8842), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8113), .ZN(
        n7834) );
  OAI21_X1 U9522 ( .B1(n7835), .B2(n9983), .A(n7834), .ZN(n7836) );
  AOI21_X1 U9523 ( .B1(n7837), .B2(n9994), .A(n7836), .ZN(n7838) );
  OAI211_X1 U9524 ( .C1(n7840), .C2(n9998), .A(n7839), .B(n7838), .ZN(P2_U3192) );
  AOI22_X1 U9525 ( .A1(n7843), .A2(n7842), .B1(n7841), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n7906) );
  XOR2_X1 U9526 ( .A(n7848), .B(n7906), .Z(n7908) );
  XNOR2_X1 U9527 ( .A(n7908), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U9528 ( .A1(n9455), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9529 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9394) );
  OAI211_X1 U9530 ( .C1(n9843), .C2(n4678), .A(n7844), .B(n9394), .ZN(n7852)
         );
  INV_X1 U9531 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7850) );
  INV_X1 U9532 ( .A(n7912), .ZN(n7847) );
  NOR2_X1 U9533 ( .A1(n7850), .A2(n7849), .ZN(n7911) );
  AOI211_X1 U9534 ( .C1(n7850), .C2(n7849), .A(n7911), .B(n9471), .ZN(n7851)
         );
  AOI211_X1 U9535 ( .C1(n9459), .C2(n7853), .A(n7852), .B(n7851), .ZN(n7854)
         );
  INV_X1 U9536 ( .A(n7854), .ZN(P1_U3258) );
  AOI21_X1 U9537 ( .B1(n7855), .B2(n7856), .A(n4589), .ZN(n7866) );
  INV_X1 U9538 ( .A(n7857), .ZN(n7859) );
  OAI22_X1 U9539 ( .A1(n9355), .A2(n7859), .B1(n9396), .B2(n7858), .ZN(n7860)
         );
  AOI211_X1 U9540 ( .C1(n9391), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7865)
         );
  NAND2_X1 U9541 ( .A1(n9407), .A2(n7863), .ZN(n7864) );
  OAI211_X1 U9542 ( .C1(n7866), .C2(n9402), .A(n7865), .B(n7864), .ZN(P1_U3221) );
  INV_X1 U9543 ( .A(n7867), .ZN(n7892) );
  OAI222_X1 U9544 ( .A1(n8665), .A2(n7892), .B1(n6604), .B2(P2_U3151), .C1(
        n7868), .C2(n9216), .ZN(P2_U3274) );
  OAI21_X1 U9545 ( .B1(n7871), .B2(n7869), .A(n7870), .ZN(n7872) );
  NAND2_X1 U9546 ( .A1(n7872), .A2(n9383), .ZN(n7878) );
  OAI22_X1 U9547 ( .A1(n9355), .A2(n7874), .B1(n9396), .B2(n7873), .ZN(n7875)
         );
  AOI211_X1 U9548 ( .C1(n9391), .C2(n9421), .A(n7876), .B(n7875), .ZN(n7877)
         );
  OAI211_X1 U9549 ( .C1(n9895), .C2(n9299), .A(n7878), .B(n7877), .ZN(P1_U3231) );
  OAI21_X1 U9550 ( .B1(n7879), .B2(n6336), .A(n7963), .ZN(n10006) );
  NAND2_X1 U9551 ( .A1(n7881), .A2(n7880), .ZN(n7883) );
  AND2_X1 U9552 ( .A1(n7883), .A2(n6789), .ZN(n7886) );
  NAND2_X1 U9553 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  OAI211_X1 U9554 ( .C1(n7886), .C2(n7885), .A(n7884), .B(n9060), .ZN(n7888)
         );
  AOI22_X1 U9555 ( .A1(n9055), .A2(n8775), .B1(n8773), .B2(n9057), .ZN(n7887)
         );
  AND2_X1 U9556 ( .A1(n7888), .A2(n7887), .ZN(n10005) );
  OAI21_X1 U9557 ( .B1(n10006), .B2(n10056), .A(n10005), .ZN(n7950) );
  OAI22_X1 U9558 ( .A1(n9101), .A2(n7948), .B1(n10065), .B2(n6328), .ZN(n7889)
         );
  AOI21_X1 U9559 ( .B1(n7950), .B2(n10065), .A(n7889), .ZN(n7890) );
  INV_X1 U9560 ( .A(n7890), .ZN(P2_U3466) );
  OAI222_X1 U9561 ( .A1(P1_U3086), .A2(n8406), .B1(n9826), .B2(n7892), .C1(
        n7891), .C2(n8653), .ZN(P1_U3334) );
  OAI21_X1 U9562 ( .B1(n7894), .B2(n8423), .A(n7893), .ZN(n8019) );
  INV_X1 U9563 ( .A(n8019), .ZN(n7905) );
  XNOR2_X1 U9564 ( .A(n7895), .B(n5048), .ZN(n7896) );
  NAND2_X1 U9565 ( .A1(n7896), .A2(n9701), .ZN(n7898) );
  AOI22_X1 U9566 ( .A1(n9417), .A2(n9698), .B1(n9696), .B2(n9419), .ZN(n7897)
         );
  NAND2_X1 U9567 ( .A1(n7898), .A2(n7897), .ZN(n8017) );
  INV_X1 U9568 ( .A(n8005), .ZN(n7899) );
  AOI211_X1 U9569 ( .C1(n8147), .C2(n7900), .A(n9707), .B(n7899), .ZN(n8018)
         );
  NAND2_X1 U9570 ( .A1(n8018), .A2(n9853), .ZN(n7902) );
  AOI22_X1 U9571 ( .A1(n9866), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8143), .B2(
        n9856), .ZN(n7901) );
  OAI211_X1 U9572 ( .C1(n8024), .C2(n9859), .A(n7902), .B(n7901), .ZN(n7903)
         );
  AOI21_X1 U9573 ( .B1(n8017), .B2(n9670), .A(n7903), .ZN(n7904) );
  OAI21_X1 U9574 ( .B1(n7905), .B2(n9693), .A(n7904), .ZN(P1_U3280) );
  INV_X1 U9575 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7907) );
  OAI22_X1 U9576 ( .A1(n7908), .A2(n7907), .B1(n4678), .B2(n7906), .ZN(n7910)
         );
  XNOR2_X1 U9577 ( .A(n8076), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7909) );
  NOR2_X1 U9578 ( .A1(n7909), .A2(n7910), .ZN(n8069) );
  AOI21_X1 U9579 ( .B1(n7910), .B2(n7909), .A(n8069), .ZN(n7921) );
  NOR2_X1 U9580 ( .A1(n7912), .A2(n7911), .ZN(n7915) );
  NAND2_X1 U9581 ( .A1(n8076), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7913) );
  OAI21_X1 U9582 ( .B1(n8076), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7913), .ZN(
        n7914) );
  AOI211_X1 U9583 ( .C1(n7915), .C2(n7914), .A(n8075), .B(n9471), .ZN(n7916)
         );
  INV_X1 U9584 ( .A(n7916), .ZN(n7920) );
  INV_X1 U9585 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U9586 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9305) );
  OAI21_X1 U9587 ( .B1(n9852), .B2(n7917), .A(n9305), .ZN(n7918) );
  AOI21_X1 U9588 ( .B1(n9440), .B2(n8076), .A(n7918), .ZN(n7919) );
  OAI211_X1 U9589 ( .C1(n7921), .C2(n9845), .A(n7920), .B(n7919), .ZN(P1_U3259) );
  AOI21_X1 U9590 ( .B1(n7924), .B2(n7923), .A(n7922), .ZN(n7937) );
  OAI21_X1 U9591 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7926), .A(n7925), .ZN(
        n7935) );
  INV_X1 U9592 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U9593 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10438), .ZN(n8182) );
  AOI21_X1 U9594 ( .B1(n8842), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8182), .ZN(
        n7927) );
  OAI21_X1 U9595 ( .B1(n7928), .B2(n9983), .A(n7927), .ZN(n7934) );
  AOI21_X1 U9596 ( .B1(n7931), .B2(n7930), .A(n7929), .ZN(n7932) );
  NOR2_X1 U9597 ( .A1(n7932), .A2(n9998), .ZN(n7933) );
  AOI211_X1 U9598 ( .C1(n9994), .C2(n7935), .A(n7934), .B(n7933), .ZN(n7936)
         );
  OAI21_X1 U9599 ( .B1(n7937), .B2(n9958), .A(n7936), .ZN(P2_U3193) );
  INV_X1 U9600 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7938) );
  OAI22_X1 U9601 ( .A1(n9174), .A2(n7939), .B1(n7938), .B2(n10052), .ZN(n7940)
         );
  AOI21_X1 U9602 ( .B1(n7941), .B2(n10052), .A(n7940), .ZN(n7942) );
  INV_X1 U9603 ( .A(n7942), .ZN(P2_U3405) );
  INV_X1 U9604 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7943) );
  OAI22_X1 U9605 ( .A1(n9174), .A2(n6302), .B1(n7943), .B2(n10052), .ZN(n7944)
         );
  AOI21_X1 U9606 ( .B1(n7945), .B2(n10052), .A(n7944), .ZN(n7946) );
  INV_X1 U9607 ( .A(n7946), .ZN(P2_U3402) );
  INV_X1 U9608 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7947) );
  OAI22_X1 U9609 ( .A1(n9174), .A2(n7948), .B1(n7947), .B2(n10052), .ZN(n7949)
         );
  AOI21_X1 U9610 ( .B1(n7950), .B2(n10052), .A(n7949), .ZN(n7951) );
  INV_X1 U9611 ( .A(n7951), .ZN(P2_U3411) );
  INV_X1 U9612 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7952) );
  OAI22_X1 U9613 ( .A1(n9174), .A2(n7953), .B1(n7952), .B2(n10052), .ZN(n7954)
         );
  AOI21_X1 U9614 ( .B1(n7955), .B2(n10052), .A(n7954), .ZN(n7956) );
  INV_X1 U9615 ( .A(n7956), .ZN(P2_U3393) );
  INV_X1 U9616 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7957) );
  OAI22_X1 U9617 ( .A1(n9174), .A2(n7958), .B1(n7957), .B2(n10052), .ZN(n7959)
         );
  AOI21_X1 U9618 ( .B1(n7960), .B2(n10052), .A(n7959), .ZN(n7961) );
  INV_X1 U9619 ( .A(n7961), .ZN(P2_U3399) );
  NAND2_X1 U9620 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  XNOR2_X1 U9621 ( .A(n7964), .B(n7967), .ZN(n8027) );
  AND2_X1 U9622 ( .A1(n7966), .A2(n7965), .ZN(n7968) );
  XNOR2_X1 U9623 ( .A(n7968), .B(n7967), .ZN(n7969) );
  AOI222_X1 U9624 ( .A1(n9060), .A2(n7969), .B1(n8774), .B2(n9055), .C1(n8114), 
        .C2(n9057), .ZN(n8032) );
  OAI21_X1 U9625 ( .B1(n10056), .B2(n8027), .A(n8032), .ZN(n7975) );
  INV_X1 U9626 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7970) );
  OAI22_X1 U9627 ( .A1(n9174), .A2(n7973), .B1(n7970), .B2(n10052), .ZN(n7971)
         );
  AOI21_X1 U9628 ( .B1(n7975), .B2(n10052), .A(n7971), .ZN(n7972) );
  INV_X1 U9629 ( .A(n7972), .ZN(P2_U3414) );
  OAI22_X1 U9630 ( .A1(n9101), .A2(n7973), .B1(n10065), .B2(n6339), .ZN(n7974)
         );
  AOI21_X1 U9631 ( .B1(n7975), .B2(n10065), .A(n7974), .ZN(n7976) );
  INV_X1 U9632 ( .A(n7976), .ZN(P2_U3467) );
  XNOR2_X1 U9633 ( .A(n8094), .B(n8623), .ZN(n8120) );
  XNOR2_X1 U9634 ( .A(n7982), .B(n8623), .ZN(n8191) );
  INV_X1 U9635 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U9636 ( .A1(n7978), .A2(n8114), .ZN(n7979) );
  NOR3_X1 U9637 ( .A1(n10039), .A2(n8772), .A3(n8639), .ZN(n7981) );
  AOI211_X1 U9638 ( .C1(n8175), .C2(n8639), .A(n7981), .B(n8162), .ZN(n7985)
         );
  NOR3_X1 U9639 ( .A1(n8094), .A2(n8568), .A3(n8772), .ZN(n7983) );
  AOI211_X1 U9640 ( .C1(n8175), .C2(n8568), .A(n7983), .B(n7982), .ZN(n7984)
         );
  XNOR2_X1 U9641 ( .A(n8179), .B(n8645), .ZN(n7986) );
  XNOR2_X1 U9642 ( .A(n7986), .B(n8770), .ZN(n8151) );
  OAI21_X1 U9643 ( .B1(n7985), .B2(n7984), .A(n8151), .ZN(n7987) );
  XNOR2_X1 U9644 ( .A(n8227), .B(n8645), .ZN(n7988) );
  NOR2_X1 U9645 ( .A1(n7988), .A2(n8174), .ZN(n8061) );
  NAND2_X1 U9646 ( .A1(n7988), .A2(n8174), .ZN(n8062) );
  INV_X1 U9647 ( .A(n8062), .ZN(n7989) );
  NOR2_X1 U9648 ( .A1(n8061), .A2(n7989), .ZN(n7990) );
  XNOR2_X1 U9649 ( .A(n8063), .B(n7990), .ZN(n7996) );
  NAND2_X1 U9650 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9978) );
  INV_X1 U9651 ( .A(n9978), .ZN(n7992) );
  NOR2_X1 U9652 ( .A1(n8757), .A2(n8211), .ZN(n7991) );
  AOI211_X1 U9653 ( .C1(n8761), .C2(n8770), .A(n7992), .B(n7991), .ZN(n7993)
         );
  OAI21_X1 U9654 ( .B1(n8219), .B2(n8758), .A(n7993), .ZN(n7994) );
  AOI21_X1 U9655 ( .B1(n8227), .B2(n8723), .A(n7994), .ZN(n7995) );
  OAI21_X1 U9656 ( .B1(n7996), .B2(n8725), .A(n7995), .ZN(P2_U3174) );
  INV_X1 U9657 ( .A(n7997), .ZN(n8000) );
  OAI222_X1 U9658 ( .A1(n9216), .A2(n7999), .B1(n8665), .B2(n8000), .C1(
        P2_U3151), .C2(n7998), .ZN(P2_U3273) );
  OAI222_X1 U9659 ( .A1(n8001), .A2(P1_U3086), .B1(n9826), .B2(n8000), .C1(
        n10469), .C2(n8653), .ZN(P1_U3333) );
  INV_X1 U9660 ( .A(n8336), .ZN(n8424) );
  XNOR2_X1 U9661 ( .A(n8002), .B(n8424), .ZN(n9785) );
  AOI21_X1 U9662 ( .B1(n8336), .B2(n8003), .A(n4571), .ZN(n8004) );
  OAI222_X1 U9663 ( .A1(n9686), .A2(n9307), .B1(n9684), .B2(n9242), .C1(n9681), 
        .C2(n8004), .ZN(n9781) );
  AOI211_X1 U9664 ( .C1(n9783), .C2(n8005), .A(n9707), .B(n4565), .ZN(n9782)
         );
  NAND2_X1 U9665 ( .A1(n9782), .A2(n9853), .ZN(n8007) );
  AOI22_X1 U9666 ( .A1(n9866), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9241), .B2(
        n9856), .ZN(n8006) );
  OAI211_X1 U9667 ( .C1(n9248), .C2(n9859), .A(n8007), .B(n8006), .ZN(n8008)
         );
  AOI21_X1 U9668 ( .B1(n9781), .B2(n9670), .A(n8008), .ZN(n8009) );
  OAI21_X1 U9669 ( .B1(n9785), .B2(n9693), .A(n8009), .ZN(P1_U3279) );
  NAND2_X1 U9670 ( .A1(n8013), .A2(n8010), .ZN(n8012) );
  OR2_X1 U9671 ( .A1(n8011), .A2(P1_U3086), .ZN(n8540) );
  OAI211_X1 U9672 ( .C1(n5368), .C2(n8653), .A(n8012), .B(n8540), .ZN(P1_U3332) );
  NAND2_X1 U9673 ( .A1(n8013), .A2(n9213), .ZN(n8015) );
  OAI211_X1 U9674 ( .C1(n8016), .C2(n9216), .A(n8015), .B(n8014), .ZN(P2_U3272) );
  INV_X1 U9675 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8020) );
  AOI211_X1 U9676 ( .C1(n8019), .C2(n9909), .A(n8018), .B(n8017), .ZN(n8022)
         );
  MUX2_X1 U9677 ( .A(n8020), .B(n8022), .S(n9913), .Z(n8021) );
  OAI21_X1 U9678 ( .B1(n8024), .B2(n9814), .A(n8021), .ZN(P1_U3492) );
  MUX2_X1 U9679 ( .A(n7382), .B(n8022), .S(n9926), .Z(n8023) );
  OAI21_X1 U9680 ( .B1(n8024), .B2(n9780), .A(n8023), .ZN(P1_U3535) );
  OAI22_X1 U9681 ( .A1(n10023), .A2(n8026), .B1(n8025), .B2(n9061), .ZN(n8029)
         );
  NOR2_X1 U9682 ( .A1(n8027), .A2(n9069), .ZN(n8028) );
  AOI211_X1 U9683 ( .C1(n10017), .C2(n8030), .A(n8029), .B(n8028), .ZN(n8031)
         );
  OAI21_X1 U9684 ( .B1(n8033), .B2(n8032), .A(n8031), .ZN(P2_U3225) );
  AOI21_X1 U9685 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8052) );
  INV_X1 U9686 ( .A(n8037), .ZN(n8038) );
  NOR2_X1 U9687 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  NAND2_X1 U9688 ( .A1(n8042), .A2(n8041), .ZN(n8040) );
  OAI211_X1 U9689 ( .C1(n8042), .C2(n8041), .A(n9993), .B(n8040), .ZN(n8051)
         );
  OAI21_X1 U9690 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8049) );
  NOR2_X1 U9691 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10460), .ZN(n8153) );
  AOI21_X1 U9692 ( .B1(n8842), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8153), .ZN(
        n8046) );
  OAI21_X1 U9693 ( .B1(n8047), .B2(n9983), .A(n8046), .ZN(n8048) );
  AOI21_X1 U9694 ( .B1(n8049), .B2(n9994), .A(n8048), .ZN(n8050) );
  OAI211_X1 U9695 ( .C1(n8052), .C2(n9998), .A(n8051), .B(n8050), .ZN(P2_U3194) );
  XOR2_X1 U9696 ( .A(n8054), .B(n8053), .Z(n8060) );
  AOI22_X1 U9697 ( .A1(n9393), .A2(n8055), .B1(n9386), .B2(n9420), .ZN(n8056)
         );
  NAND2_X1 U9698 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9850) );
  OAI211_X1 U9699 ( .C1(n9242), .C2(n9376), .A(n8056), .B(n9850), .ZN(n8057)
         );
  AOI21_X1 U9700 ( .B1(n8058), .B2(n9407), .A(n8057), .ZN(n8059) );
  OAI21_X1 U9701 ( .B1(n8060), .B2(n9402), .A(n8059), .ZN(P1_U3224) );
  XNOR2_X1 U9702 ( .A(n9201), .B(n8645), .ZN(n8125) );
  XNOR2_X1 U9703 ( .A(n8125), .B(n9047), .ZN(n8127) );
  XOR2_X1 U9704 ( .A(n8128), .B(n8127), .Z(n8068) );
  INV_X1 U9705 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10480) );
  OAI22_X1 U9706 ( .A1(n8757), .A2(n8544), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10480), .ZN(n8064) );
  AOI21_X1 U9707 ( .B1(n8761), .B2(n9056), .A(n8064), .ZN(n8065) );
  OAI21_X1 U9708 ( .B1(n9062), .B2(n8758), .A(n8065), .ZN(n8066) );
  AOI21_X1 U9709 ( .B1(n9201), .B2(n8723), .A(n8066), .ZN(n8067) );
  OAI21_X1 U9710 ( .B1(n8068), .B2(n8725), .A(n8067), .ZN(P2_U3155) );
  INV_X1 U9711 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9778) );
  AOI21_X1 U9712 ( .B1(n8070), .B2(n9778), .A(n8069), .ZN(n8072) );
  XNOR2_X1 U9713 ( .A(n8261), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8071) );
  NOR2_X1 U9714 ( .A1(n8072), .A2(n8071), .ZN(n8259) );
  AOI21_X1 U9715 ( .B1(n8072), .B2(n8071), .A(n8259), .ZN(n8074) );
  NAND2_X1 U9716 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U9717 ( .A1(n9455), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n8073) );
  OAI211_X1 U9718 ( .C1(n9845), .C2(n8074), .A(n9312), .B(n8073), .ZN(n8081)
         );
  NOR2_X1 U9719 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n8261), .ZN(n8077) );
  AOI21_X1 U9720 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n8261), .A(n8077), .ZN(
        n8078) );
  AOI221_X1 U9721 ( .B1(n8079), .B2(n8252), .C1(n8078), .C2(n8252), .A(n9471), 
        .ZN(n8080) );
  AOI211_X1 U9722 ( .C1(n9440), .C2(n8261), .A(n8081), .B(n8080), .ZN(n8082)
         );
  INV_X1 U9723 ( .A(n8082), .ZN(P1_U3260) );
  INV_X1 U9724 ( .A(n8085), .ZN(n8083) );
  XNOR2_X1 U9725 ( .A(n8084), .B(n8083), .ZN(n10041) );
  XNOR2_X1 U9726 ( .A(n8086), .B(n8085), .ZN(n8087) );
  NAND2_X1 U9727 ( .A1(n8087), .A2(n9060), .ZN(n8089) );
  AOI22_X1 U9728 ( .A1(n8771), .A2(n9057), .B1(n9055), .B2(n8114), .ZN(n8088)
         );
  NAND2_X1 U9729 ( .A1(n8089), .A2(n8088), .ZN(n8090) );
  AOI21_X1 U9730 ( .B1(n10041), .B2(n8102), .A(n8090), .ZN(n10043) );
  NOR2_X1 U9731 ( .A1(n8033), .A2(n8091), .ZN(n8660) );
  INV_X1 U9732 ( .A(n8092), .ZN(n8115) );
  AOI22_X1 U9733 ( .A1(n8033), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10019), .B2(
        n8115), .ZN(n8093) );
  OAI21_X1 U9734 ( .B1(n8094), .B2(n8984), .A(n8093), .ZN(n8095) );
  AOI21_X1 U9735 ( .B1(n10041), .B2(n8660), .A(n8095), .ZN(n8096) );
  OAI21_X1 U9736 ( .B1(n10043), .B2(n8033), .A(n8096), .ZN(P2_U3223) );
  AOI21_X1 U9737 ( .B1(n8099), .B2(n8097), .A(n4591), .ZN(n8103) );
  INV_X1 U9738 ( .A(n8103), .ZN(n10035) );
  INV_X1 U9739 ( .A(n8660), .ZN(n8112) );
  XNOR2_X1 U9740 ( .A(n8098), .B(n8099), .ZN(n8105) );
  OAI22_X1 U9741 ( .A1(n8100), .A2(n9036), .B1(n4688), .B2(n9004), .ZN(n8101)
         );
  AOI21_X1 U9742 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8104) );
  OAI21_X1 U9743 ( .B1(n8989), .B2(n8105), .A(n8104), .ZN(n10037) );
  NAND2_X1 U9744 ( .A1(n10037), .A2(n10023), .ZN(n8111) );
  OAI22_X1 U9745 ( .A1(n10023), .A2(n8107), .B1(n8106), .B2(n9061), .ZN(n8108)
         );
  AOI21_X1 U9746 ( .B1(n10017), .B2(n8109), .A(n8108), .ZN(n8110) );
  OAI211_X1 U9747 ( .C1(n10035), .C2(n8112), .A(n8111), .B(n8110), .ZN(
        P2_U3224) );
  AOI21_X1 U9748 ( .B1(n8761), .B2(n8114), .A(n8113), .ZN(n8117) );
  NAND2_X1 U9749 ( .A1(n8747), .A2(n8115), .ZN(n8116) );
  OAI211_X1 U9750 ( .C1(n8175), .C2(n8757), .A(n8117), .B(n8116), .ZN(n8123)
         );
  XNOR2_X1 U9751 ( .A(n8118), .B(n8772), .ZN(n8119) );
  NOR2_X1 U9752 ( .A1(n8119), .A2(n8120), .ZN(n8188) );
  AOI21_X1 U9753 ( .B1(n8120), .B2(n8119), .A(n8188), .ZN(n8121) );
  NOR2_X1 U9754 ( .A1(n8121), .A2(n8725), .ZN(n8122) );
  AOI211_X1 U9755 ( .C1(n10039), .C2(n8723), .A(n8123), .B(n8122), .ZN(n8124)
         );
  INV_X1 U9756 ( .A(n8124), .ZN(P2_U3157) );
  INV_X1 U9757 ( .A(n9194), .ZN(n8136) );
  XNOR2_X1 U9758 ( .A(n9194), .B(n8623), .ZN(n8543) );
  XNOR2_X1 U9759 ( .A(n8543), .B(n9058), .ZN(n8129) );
  OAI211_X1 U9760 ( .C1(n8130), .C2(n8129), .A(n8542), .B(n8754), .ZN(n8135)
         );
  INV_X1 U9761 ( .A(n8131), .ZN(n9049) );
  NAND2_X1 U9762 ( .A1(n8761), .A2(n9047), .ZN(n8132) );
  NAND2_X1 U9763 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8809) );
  OAI211_X1 U9764 ( .C1(n8757), .C2(n9037), .A(n8132), .B(n8809), .ZN(n8133)
         );
  AOI21_X1 U9765 ( .B1(n9049), .B2(n8747), .A(n8133), .ZN(n8134) );
  OAI211_X1 U9766 ( .C1(n8136), .C2(n8764), .A(n8135), .B(n8134), .ZN(P2_U3181) );
  INV_X1 U9767 ( .A(n8137), .ZN(n8195) );
  OAI222_X1 U9768 ( .A1(n8665), .A2(n8195), .B1(P2_U3151), .B2(n6844), .C1(
        n8138), .C2(n9216), .ZN(P2_U3271) );
  NAND2_X1 U9769 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  XOR2_X1 U9770 ( .A(n8142), .B(n8141), .Z(n8149) );
  AOI22_X1 U9771 ( .A1(n9393), .A2(n8143), .B1(n9386), .B2(n9419), .ZN(n8145)
         );
  OAI211_X1 U9772 ( .C1(n9397), .C2(n9376), .A(n8145), .B(n8144), .ZN(n8146)
         );
  AOI21_X1 U9773 ( .B1(n8147), .B2(n9407), .A(n8146), .ZN(n8148) );
  OAI21_X1 U9774 ( .B1(n8149), .B2(n9402), .A(n8148), .ZN(P1_U3234) );
  NOR2_X1 U9775 ( .A1(n8118), .A2(n8772), .ZN(n8187) );
  NOR3_X1 U9776 ( .A1(n8188), .A2(n8187), .A3(n8191), .ZN(n8189) );
  AOI21_X1 U9777 ( .B1(n8771), .B2(n8191), .A(n8189), .ZN(n8150) );
  XOR2_X1 U9778 ( .A(n8151), .B(n8150), .Z(n8157) );
  NOR2_X1 U9779 ( .A1(n8757), .A2(n8174), .ZN(n8152) );
  AOI211_X1 U9780 ( .C1(n8761), .C2(n8771), .A(n8153), .B(n8152), .ZN(n8154)
         );
  OAI21_X1 U9781 ( .B1(n8176), .B2(n8758), .A(n8154), .ZN(n8155) );
  AOI21_X1 U9782 ( .B1(n8179), .B2(n8723), .A(n8155), .ZN(n8156) );
  OAI21_X1 U9783 ( .B1(n8157), .B2(n8725), .A(n8156), .ZN(P2_U3164) );
  XNOR2_X1 U9784 ( .A(n8158), .B(n8162), .ZN(n8159) );
  NAND2_X1 U9785 ( .A1(n8159), .A2(n9060), .ZN(n8161) );
  AOI22_X1 U9786 ( .A1(n9057), .A2(n8770), .B1(n8772), .B2(n9055), .ZN(n8160)
         );
  AND2_X1 U9787 ( .A1(n8161), .A2(n8160), .ZN(n10050) );
  OR2_X1 U9788 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  NAND2_X1 U9789 ( .A1(n8169), .A2(n8164), .ZN(n10046) );
  NAND2_X1 U9790 ( .A1(n10046), .A2(n9023), .ZN(n8167) );
  OAI22_X1 U9791 ( .A1(n10023), .A2(n7931), .B1(n8183), .B2(n9061), .ZN(n8165)
         );
  AOI21_X1 U9792 ( .B1(n10048), .B2(n10017), .A(n8165), .ZN(n8166) );
  OAI211_X1 U9793 ( .C1(n10050), .C2(n8033), .A(n8167), .B(n8166), .ZN(
        P2_U3222) );
  NAND2_X1 U9794 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  XNOR2_X1 U9795 ( .A(n8170), .B(n8171), .ZN(n10057) );
  XNOR2_X1 U9796 ( .A(n8172), .B(n8171), .ZN(n8173) );
  OAI222_X1 U9797 ( .A1(n9004), .A2(n8175), .B1(n9036), .B2(n8174), .C1(n8173), 
        .C2(n8989), .ZN(n10058) );
  NAND2_X1 U9798 ( .A1(n10058), .A2(n10023), .ZN(n8181) );
  OAI22_X1 U9799 ( .A1(n10023), .A2(n8177), .B1(n8176), .B2(n9061), .ZN(n8178)
         );
  AOI21_X1 U9800 ( .B1(n8179), .B2(n10017), .A(n8178), .ZN(n8180) );
  OAI211_X1 U9801 ( .C1(n10057), .C2(n9069), .A(n8181), .B(n8180), .ZN(
        P2_U3221) );
  AOI21_X1 U9802 ( .B1(n8761), .B2(n8772), .A(n8182), .ZN(n8186) );
  INV_X1 U9803 ( .A(n8183), .ZN(n8184) );
  NAND2_X1 U9804 ( .A1(n8747), .A2(n8184), .ZN(n8185) );
  OAI211_X1 U9805 ( .C1(n8210), .C2(n8757), .A(n8186), .B(n8185), .ZN(n8193)
         );
  OR2_X1 U9806 ( .A1(n8188), .A2(n8187), .ZN(n8190) );
  AOI211_X1 U9807 ( .C1(n8191), .C2(n8190), .A(n8725), .B(n8189), .ZN(n8192)
         );
  AOI211_X1 U9808 ( .C1(n10048), .C2(n8723), .A(n8193), .B(n8192), .ZN(n8194)
         );
  INV_X1 U9809 ( .A(n8194), .ZN(P2_U3176) );
  OAI222_X1 U9810 ( .A1(n5471), .A2(P1_U3086), .B1(n9826), .B2(n8195), .C1(
        n10414), .C2(n8653), .ZN(P1_U3331) );
  XNOR2_X1 U9811 ( .A(n8196), .B(n8426), .ZN(n8197) );
  AOI222_X1 U9812 ( .A1(n9701), .A2(n8197), .B1(n9416), .B2(n9698), .C1(n9417), 
        .C2(n9696), .ZN(n9831) );
  XOR2_X1 U9813 ( .A(n8198), .B(n8426), .Z(n9834) );
  NAND2_X1 U9814 ( .A1(n9834), .A2(n9863), .ZN(n8204) );
  OAI22_X1 U9815 ( .A1(n9670), .A2(n7850), .B1(n8199), .B2(n9490), .ZN(n8202)
         );
  OAI211_X1 U9816 ( .C1(n9832), .C2(n4565), .A(n8200), .B(n9708), .ZN(n9830)
         );
  NOR2_X1 U9817 ( .A1(n9830), .A2(n9495), .ZN(n8201) );
  AOI211_X1 U9818 ( .C1(n9492), .C2(n9408), .A(n8202), .B(n8201), .ZN(n8203)
         );
  OAI211_X1 U9819 ( .C1(n9866), .C2(n9831), .A(n8204), .B(n8203), .ZN(P1_U3278) );
  XNOR2_X1 U9820 ( .A(n8205), .B(n8209), .ZN(n8230) );
  INV_X1 U9821 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8214) );
  NOR2_X1 U9822 ( .A1(n8206), .A2(n4691), .ZN(n8207) );
  AOI211_X1 U9823 ( .C1(n8209), .C2(n8208), .A(n8989), .B(n8207), .ZN(n8213)
         );
  OAI22_X1 U9824 ( .A1(n8211), .A2(n9036), .B1(n8210), .B2(n9004), .ZN(n8212)
         );
  NOR2_X1 U9825 ( .A1(n8213), .A2(n8212), .ZN(n8225) );
  MUX2_X1 U9826 ( .A(n8214), .B(n8225), .S(n10052), .Z(n8216) );
  NAND2_X1 U9827 ( .A1(n8227), .A2(n9200), .ZN(n8215) );
  OAI211_X1 U9828 ( .C1(n8230), .C2(n9204), .A(n8216), .B(n8215), .ZN(P2_U3429) );
  INV_X1 U9829 ( .A(n8227), .ZN(n8217) );
  OAI21_X1 U9830 ( .B1(n8217), .B2(n9063), .A(n8225), .ZN(n8218) );
  NAND2_X1 U9831 ( .A1(n8218), .A2(n10023), .ZN(n8222) );
  INV_X1 U9832 ( .A(n8219), .ZN(n8220) );
  AOI22_X1 U9833 ( .A1(n8033), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10019), .B2(
        n8220), .ZN(n8221) );
  OAI211_X1 U9834 ( .C1(n8230), .C2(n9069), .A(n8222), .B(n8221), .ZN(P2_U3220) );
  INV_X1 U9835 ( .A(n8223), .ZN(n8541) );
  OAI222_X1 U9836 ( .A1(n8665), .A2(n8541), .B1(P2_U3151), .B2(n6845), .C1(
        n8224), .C2(n9216), .ZN(P2_U3270) );
  MUX2_X1 U9837 ( .A(n8226), .B(n8225), .S(n10065), .Z(n8229) );
  NAND2_X1 U9838 ( .A1(n8227), .A2(n9121), .ZN(n8228) );
  OAI211_X1 U9839 ( .C1(n9124), .C2(n8230), .A(n8229), .B(n8228), .ZN(P2_U3472) );
  INV_X1 U9840 ( .A(n8231), .ZN(n8234) );
  OAI222_X1 U9841 ( .A1(n8665), .A2(n8234), .B1(P2_U3151), .B2(n8233), .C1(
        n8232), .C2(n9216), .ZN(P2_U3269) );
  INV_X1 U9842 ( .A(n5473), .ZN(n8235) );
  OAI222_X1 U9843 ( .A1(n8235), .A2(P1_U3086), .B1(n9826), .B2(n8234), .C1(
        n10409), .C2(n8653), .ZN(P1_U3329) );
  INV_X1 U9844 ( .A(n8236), .ZN(n8240) );
  AOI21_X1 U9845 ( .B1(n9219), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8237), .ZN(
        n8238) );
  OAI21_X1 U9846 ( .B1(n8240), .B2(n8665), .A(n8238), .ZN(P2_U3268) );
  INV_X1 U9847 ( .A(P1_U3973), .ZN(n8239) );
  AND2_X1 U9848 ( .A1(n8239), .A2(n9852), .ZN(P1_U3085) );
  OAI222_X1 U9849 ( .A1(P1_U3086), .A2(n5926), .B1(n9826), .B2(n8240), .C1(
        n10182), .C2(n8653), .ZN(P1_U3328) );
  INV_X1 U9850 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8247) );
  XNOR2_X1 U9851 ( .A(n8241), .B(n8430), .ZN(n9585) );
  INV_X1 U9852 ( .A(n9578), .ZN(n8242) );
  AOI211_X1 U9853 ( .C1(n9256), .C2(n9596), .A(n9707), .B(n8242), .ZN(n9586)
         );
  OAI21_X1 U9854 ( .B1(n8430), .B2(n8243), .A(n9571), .ZN(n8244) );
  NAND2_X1 U9855 ( .A1(n8244), .A2(n9701), .ZN(n8246) );
  AOI22_X1 U9856 ( .A1(n9614), .A2(n9696), .B1(n9698), .B2(n9413), .ZN(n8245)
         );
  NAND2_X1 U9857 ( .A1(n8246), .A2(n8245), .ZN(n9592) );
  AOI211_X1 U9858 ( .C1(n9585), .C2(n9909), .A(n9586), .B(n9592), .ZN(n8249)
         );
  MUX2_X1 U9859 ( .A(n8247), .B(n8249), .S(n9913), .Z(n8248) );
  OAI21_X1 U9860 ( .B1(n9590), .B2(n9814), .A(n8248), .ZN(P1_U3513) );
  INV_X1 U9861 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8250) );
  MUX2_X1 U9862 ( .A(n8250), .B(n8249), .S(n9926), .Z(n8251) );
  OAI21_X1 U9863 ( .B1(n9590), .B2(n9780), .A(n8251), .ZN(P1_U3545) );
  NAND2_X1 U9864 ( .A1(n9480), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8255) );
  INV_X1 U9865 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U9866 ( .A1(n8262), .A2(n8253), .ZN(n8254) );
  AND2_X1 U9867 ( .A1(n8255), .A2(n8254), .ZN(n9473) );
  NOR2_X1 U9868 ( .A1(n9474), .A2(n9473), .ZN(n9472) );
  AND2_X1 U9869 ( .A1(n8262), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8256) );
  OR2_X1 U9870 ( .A1(n9472), .A2(n8256), .ZN(n8258) );
  INV_X1 U9871 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8257) );
  XNOR2_X1 U9872 ( .A(n8258), .B(n8257), .ZN(n8266) );
  XNOR2_X1 U9873 ( .A(n8262), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9468) );
  INV_X1 U9874 ( .A(n8259), .ZN(n8260) );
  OAI21_X1 U9875 ( .B1(n8261), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8260), .ZN(
        n9467) );
  OR2_X1 U9876 ( .A1(n9468), .A2(n9467), .ZN(n9465) );
  NAND2_X1 U9877 ( .A1(n8262), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U9878 ( .A1(n9465), .A2(n8263), .ZN(n8265) );
  INV_X1 U9879 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8264) );
  XNOR2_X1 U9880 ( .A(n8265), .B(n8264), .ZN(n8267) );
  AOI22_X1 U9881 ( .A1(n8266), .A2(n9849), .B1(n9459), .B2(n8267), .ZN(n8271)
         );
  INV_X1 U9882 ( .A(n8266), .ZN(n8269) );
  OAI21_X1 U9883 ( .B1(n9845), .B2(n8267), .A(n9843), .ZN(n8268) );
  AOI21_X1 U9884 ( .B1(n8269), .B2(n9849), .A(n8268), .ZN(n8270) );
  MUX2_X1 U9885 ( .A(n8271), .B(n8270), .S(n5457), .Z(n8274) );
  NOR2_X1 U9886 ( .A1(n8272), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9282) );
  INV_X1 U9887 ( .A(n9282), .ZN(n8273) );
  OAI211_X1 U9888 ( .C1(n4712), .C2(n9852), .A(n8274), .B(n8273), .ZN(P1_U3262) );
  INV_X1 U9889 ( .A(n8275), .ZN(n8278) );
  AOI21_X1 U9890 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8279) );
  MUX2_X1 U9891 ( .A(n6979), .B(n8279), .S(n9670), .Z(n8282) );
  AOI22_X1 U9892 ( .A1(n9853), .A2(n8280), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9856), .ZN(n8281) );
  OAI211_X1 U9893 ( .C1(n8454), .C2(n9859), .A(n8282), .B(n8281), .ZN(P1_U3292) );
  NAND2_X1 U9894 ( .A1(n9816), .A2(n5867), .ZN(n8284) );
  NAND2_X1 U9895 ( .A1(n8393), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U9896 ( .A1(n5870), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U9897 ( .A1(n5594), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9898 ( .A1(n8285), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8286) );
  NAND3_X1 U9899 ( .A1(n8288), .A2(n8287), .A3(n8286), .ZN(n9410) );
  NOR2_X1 U9900 ( .A1(n8592), .A2(n9410), .ZN(n8526) );
  INV_X1 U9901 ( .A(n8526), .ZN(n8504) );
  AOI21_X1 U9902 ( .B1(n9410), .B2(n4975), .A(n8402), .ZN(n8400) );
  INV_X1 U9903 ( .A(n8442), .ZN(n8365) );
  AOI21_X1 U9904 ( .B1(n9678), .B2(n9697), .A(n4976), .ZN(n8343) );
  INV_X1 U9905 ( .A(n8343), .ZN(n8346) );
  INV_X1 U9906 ( .A(n8341), .ZN(n8481) );
  OAI21_X1 U9907 ( .B1(n8481), .B2(n8339), .A(n9678), .ZN(n8345) );
  INV_X1 U9908 ( .A(n8304), .ZN(n8292) );
  INV_X1 U9909 ( .A(n8458), .ZN(n8291) );
  NOR3_X1 U9910 ( .A1(n8292), .A2(n8291), .A3(n8398), .ZN(n8309) );
  INV_X1 U9911 ( .A(n8459), .ZN(n8294) );
  INV_X1 U9912 ( .A(n8295), .ZN(n8297) );
  OAI211_X1 U9913 ( .C1(n8300), .C2(n8297), .A(n8302), .B(n8296), .ZN(n8308)
         );
  INV_X1 U9914 ( .A(n8301), .ZN(n8307) );
  INV_X1 U9915 ( .A(n8298), .ZN(n8299) );
  NAND3_X1 U9916 ( .A1(n8303), .A2(n8302), .A3(n8301), .ZN(n8305) );
  NAND2_X1 U9917 ( .A1(n8305), .A2(n8304), .ZN(n8306) );
  INV_X1 U9918 ( .A(n8310), .ZN(n8311) );
  MUX2_X1 U9919 ( .A(n8311), .B(n4530), .S(n8398), .Z(n8312) );
  INV_X1 U9920 ( .A(n8321), .ZN(n8316) );
  NAND2_X1 U9921 ( .A1(n8416), .A2(n8314), .ZN(n8315) );
  OAI21_X1 U9922 ( .B1(n8316), .B2(n8315), .A(n8320), .ZN(n8317) );
  NAND2_X1 U9923 ( .A1(n8325), .A2(n8322), .ZN(n8466) );
  AOI21_X1 U9924 ( .B1(n8317), .B2(n8463), .A(n8466), .ZN(n8318) );
  NAND2_X1 U9925 ( .A1(n8328), .A2(n8324), .ZN(n8467) );
  AOI21_X1 U9926 ( .B1(n8323), .B2(n8416), .A(n4912), .ZN(n8327) );
  NAND2_X1 U9927 ( .A1(n8324), .A2(n8463), .ZN(n8326) );
  OAI211_X1 U9928 ( .C1(n8327), .C2(n8326), .A(n8470), .B(n8325), .ZN(n8329)
         );
  NAND2_X1 U9929 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  INV_X1 U9930 ( .A(n8474), .ZN(n8332) );
  AOI211_X1 U9931 ( .C1(n8337), .C2(n8335), .A(n8332), .B(n8336), .ZN(n8334)
         );
  NAND2_X1 U9932 ( .A1(n9248), .A2(n9417), .ZN(n8333) );
  NAND2_X1 U9933 ( .A1(n8479), .A2(n8333), .ZN(n8473) );
  NOR3_X1 U9934 ( .A1(n8334), .A2(n8481), .A3(n8473), .ZN(n8344) );
  NAND2_X1 U9935 ( .A1(n8339), .A2(n8338), .ZN(n8478) );
  NAND2_X1 U9936 ( .A1(n8349), .A2(n8347), .ZN(n8484) );
  AND2_X1 U9937 ( .A1(n8354), .A2(n8348), .ZN(n8483) );
  OAI21_X1 U9938 ( .B1(n8351), .B2(n8484), .A(n8483), .ZN(n8353) );
  NAND2_X1 U9939 ( .A1(n8348), .A2(n8480), .ZN(n8350) );
  OAI211_X1 U9940 ( .C1(n8351), .C2(n8350), .A(n8492), .B(n8349), .ZN(n8352)
         );
  INV_X1 U9941 ( .A(n8360), .ZN(n8358) );
  AOI21_X1 U9942 ( .B1(n8360), .B2(n9653), .A(n8398), .ZN(n8356) );
  INV_X1 U9943 ( .A(n8354), .ZN(n8355) );
  OAI33_X1 U9944 ( .A1(n8398), .A2(n8358), .A3(n9663), .B1(n8357), .B2(n8356), 
        .B3(n8355), .ZN(n8362) );
  NAND2_X1 U9945 ( .A1(n8442), .A2(n8359), .ZN(n8487) );
  NAND2_X1 U9946 ( .A1(n8366), .A2(n8360), .ZN(n8443) );
  MUX2_X1 U9947 ( .A(n8487), .B(n8443), .S(n8398), .Z(n8361) );
  NAND2_X1 U9948 ( .A1(n9570), .A2(n8369), .ZN(n8445) );
  NAND2_X1 U9949 ( .A1(n8374), .A2(n8370), .ZN(n8371) );
  AND2_X1 U9950 ( .A1(n8371), .A2(n9570), .ZN(n8436) );
  MUX2_X1 U9951 ( .A(n8445), .B(n8436), .S(n8398), .Z(n8372) );
  OAI21_X1 U9952 ( .B1(n8398), .B2(n8374), .A(n8373), .ZN(n8376) );
  MUX2_X1 U9953 ( .A(n8447), .B(n8438), .S(n8398), .Z(n8375) );
  INV_X1 U9954 ( .A(n8448), .ZN(n8377) );
  NAND2_X1 U9955 ( .A1(n8509), .A2(n4976), .ZN(n8379) );
  AOI21_X1 U9956 ( .B1(n8398), .B2(n8389), .A(n8378), .ZN(n8388) );
  INV_X1 U9957 ( .A(n8389), .ZN(n8452) );
  INV_X1 U9958 ( .A(n8379), .ZN(n8381) );
  AND2_X1 U9959 ( .A1(n8490), .A2(n8441), .ZN(n8383) );
  INV_X1 U9960 ( .A(n8383), .ZN(n8380) );
  NAND3_X1 U9961 ( .A1(n8452), .A2(n8381), .A3(n8380), .ZN(n8387) );
  NAND2_X1 U9962 ( .A1(n8382), .A2(n8448), .ZN(n8384) );
  NAND4_X1 U9963 ( .A1(n8384), .A2(n8398), .A3(n8383), .A4(n8513), .ZN(n8386)
         );
  INV_X1 U9964 ( .A(n8509), .ZN(n8493) );
  NAND3_X1 U9965 ( .A1(n8513), .A2(n8398), .A3(n8493), .ZN(n8385) );
  OAI21_X1 U9966 ( .B1(n8389), .B2(n8513), .A(n8495), .ZN(n8390) );
  MUX2_X1 U9967 ( .A(n8496), .B(n8499), .S(n8398), .Z(n8391) );
  NAND2_X1 U9968 ( .A1(n8664), .A2(n5867), .ZN(n8395) );
  NAND2_X1 U9969 ( .A1(n8393), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8394) );
  INV_X1 U9970 ( .A(n8396), .ZN(n8397) );
  OAI21_X1 U9971 ( .B1(n8504), .B2(n5901), .A(n8401), .ZN(n8534) );
  AOI211_X1 U9972 ( .C1(n8402), .C2(n5457), .A(n8537), .B(n8505), .ZN(n8533)
         );
  INV_X1 U9973 ( .A(n8402), .ZN(n8520) );
  INV_X1 U9974 ( .A(n9642), .ZN(n9640) );
  INV_X1 U9975 ( .A(n9660), .ZN(n8429) );
  NOR2_X1 U9976 ( .A1(n8404), .A2(n8403), .ZN(n8409) );
  INV_X1 U9977 ( .A(n8405), .ZN(n8408) );
  NAND4_X1 U9978 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n8414)
         );
  NAND2_X1 U9979 ( .A1(n8411), .A2(n8410), .ZN(n8413) );
  NOR3_X1 U9980 ( .A1(n8414), .A2(n8413), .A3(n8412), .ZN(n8415) );
  NAND3_X1 U9981 ( .A1(n8416), .A2(n8415), .A3(n4530), .ZN(n8417) );
  NOR3_X1 U9982 ( .A1(n8419), .A2(n8418), .A3(n8417), .ZN(n8420) );
  NAND3_X1 U9983 ( .A1(n8421), .A2(n5917), .A3(n8420), .ZN(n8422) );
  NOR2_X1 U9984 ( .A1(n8423), .A2(n8422), .ZN(n8425) );
  NAND4_X1 U9985 ( .A1(n9704), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n8427)
         );
  NOR2_X1 U9986 ( .A1(n9683), .A2(n8427), .ZN(n8428) );
  AND3_X1 U9987 ( .A1(n9509), .A2(n9525), .A3(n8431), .ZN(n8433) );
  NAND2_X1 U9988 ( .A1(n9483), .A2(n8432), .ZN(n8500) );
  AND4_X1 U9989 ( .A1(n8434), .A2(n8516), .A3(n8433), .A4(n8500), .ZN(n8435)
         );
  INV_X1 U9990 ( .A(n8522), .ZN(n8507) );
  INV_X1 U9991 ( .A(n8436), .ZN(n8437) );
  NAND2_X1 U9992 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  NAND2_X1 U9993 ( .A1(n8439), .A2(n8447), .ZN(n8440) );
  NAND2_X1 U9994 ( .A1(n8441), .A2(n8440), .ZN(n8486) );
  AND2_X1 U9995 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  NOR2_X1 U9996 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  AND2_X1 U9997 ( .A1(n8447), .A2(n8446), .ZN(n8449) );
  OAI21_X1 U9998 ( .B1(n8486), .B2(n8449), .A(n8448), .ZN(n8450) );
  NAND3_X1 U9999 ( .A1(n8513), .A2(n8490), .A3(n8450), .ZN(n8451) );
  NAND2_X1 U10000 ( .A1(n8452), .A2(n8451), .ZN(n8511) );
  INV_X1 U10001 ( .A(n8511), .ZN(n8498) );
  INV_X1 U10002 ( .A(n8453), .ZN(n8456) );
  NAND2_X1 U10003 ( .A1(n5545), .A2(n8454), .ZN(n8455) );
  AND4_X1 U10004 ( .A1(n8457), .A2(n8456), .A3(n5944), .A4(n8455), .ZN(n8461)
         );
  AND4_X1 U10005 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n8464)
         );
  OAI211_X1 U10006 ( .C1(n8465), .C2(n8464), .A(n8463), .B(n8462), .ZN(n8469)
         );
  INV_X1 U10007 ( .A(n8466), .ZN(n8468) );
  AOI21_X1 U10008 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8472) );
  INV_X1 U10009 ( .A(n8470), .ZN(n8471) );
  NOR2_X1 U10010 ( .A1(n8472), .A2(n8471), .ZN(n8475) );
  AOI211_X1 U10011 ( .C1(n8475), .C2(n8474), .A(n4920), .B(n8473), .ZN(n8476)
         );
  AOI211_X1 U10012 ( .C1(n8479), .C2(n8478), .A(n8477), .B(n8476), .ZN(n8482)
         );
  NOR3_X1 U10013 ( .A1(n8482), .A2(n4907), .A3(n8481), .ZN(n8485) );
  OAI21_X1 U10014 ( .B1(n8485), .B2(n8484), .A(n8483), .ZN(n8491) );
  INV_X1 U10015 ( .A(n8486), .ZN(n8489) );
  INV_X1 U10016 ( .A(n8487), .ZN(n8488) );
  NAND3_X1 U10017 ( .A1(n8490), .A2(n8489), .A3(n8488), .ZN(n8510) );
  AOI21_X1 U10018 ( .B1(n8492), .B2(n8491), .A(n8510), .ZN(n8494) );
  OAI21_X1 U10019 ( .B1(n8494), .B2(n8493), .A(n8513), .ZN(n8497) );
  NAND2_X1 U10020 ( .A1(n8496), .A2(n8495), .ZN(n8514) );
  AOI21_X1 U10021 ( .B1(n8498), .B2(n8497), .A(n8514), .ZN(n8501) );
  NAND2_X1 U10022 ( .A1(n8500), .A2(n8499), .ZN(n8518) );
  OAI21_X1 U10023 ( .B1(n8501), .B2(n8518), .A(n8516), .ZN(n8502) );
  AOI21_X1 U10024 ( .B1(n8520), .B2(n8502), .A(n8526), .ZN(n8531) );
  NAND2_X1 U10025 ( .A1(n8504), .A2(n8503), .ZN(n8506) );
  OAI211_X1 U10026 ( .C1(n8507), .C2(n8506), .A(n5457), .B(n8505), .ZN(n8508)
         );
  AOI21_X1 U10027 ( .B1(n8531), .B2(n8525), .A(n8508), .ZN(n8529) );
  OAI21_X1 U10028 ( .B1(n8510), .B2(n9628), .A(n8509), .ZN(n8512) );
  AOI21_X1 U10029 ( .B1(n8513), .B2(n8512), .A(n8511), .ZN(n8515) );
  OAI22_X1 U10030 ( .A1(n8515), .A2(n8514), .B1(n9790), .B2(n9410), .ZN(n8519)
         );
  INV_X1 U10031 ( .A(n9410), .ZN(n8517) );
  OAI22_X1 U10032 ( .A1(n8519), .A2(n8518), .B1(n8517), .B2(n8516), .ZN(n8521)
         );
  NAND2_X1 U10033 ( .A1(n8521), .A2(n8520), .ZN(n8524) );
  AOI21_X1 U10034 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8527) );
  NOR4_X1 U10035 ( .A1(n8527), .A2(n5457), .A3(n8526), .A4(n8525), .ZN(n8528)
         );
  NOR2_X1 U10036 ( .A1(n8536), .A2(n8535), .ZN(n8539) );
  OAI21_X1 U10037 ( .B1(n8540), .B2(n8537), .A(P1_B_REG_SCAN_IN), .ZN(n8538)
         );
  OAI222_X1 U10038 ( .A1(n5472), .A2(P1_U3086), .B1(n9826), .B2(n8541), .C1(
        n10494), .C2(n8653), .ZN(P1_U3330) );
  XNOR2_X1 U10039 ( .A(n8765), .B(n8623), .ZN(n8550) );
  OAI21_X2 U10040 ( .B1(n8544), .B2(n8543), .A(n8542), .ZN(n8712) );
  INV_X1 U10041 ( .A(n8712), .ZN(n8547) );
  XOR2_X1 U10042 ( .A(n8623), .B(n9188), .Z(n8710) );
  INV_X1 U10043 ( .A(n8710), .ZN(n8546) );
  OAI21_X2 U10044 ( .B1(n8712), .B2(n8710), .A(n9016), .ZN(n8545) );
  XNOR2_X1 U10045 ( .A(n9110), .B(n8645), .ZN(n8548) );
  NAND2_X1 U10046 ( .A1(n8548), .A2(n9005), .ZN(n8549) );
  OAI21_X1 U10047 ( .B1(n8548), .B2(n9005), .A(n8549), .ZN(n8719) );
  INV_X1 U10048 ( .A(n8549), .ZN(n8752) );
  XNOR2_X1 U10049 ( .A(n8550), .B(n8993), .ZN(n8751) );
  INV_X1 U10050 ( .A(n8687), .ZN(n8552) );
  INV_X2 U10051 ( .A(n8568), .ZN(n8639) );
  XNOR2_X1 U10052 ( .A(n9178), .B(n8639), .ZN(n8554) );
  XNOR2_X1 U10053 ( .A(n8554), .B(n9003), .ZN(n8688) );
  INV_X1 U10054 ( .A(n8688), .ZN(n8551) );
  XNOR2_X1 U10055 ( .A(n8727), .B(n8639), .ZN(n8553) );
  NAND2_X1 U10056 ( .A1(n8553), .A2(n8992), .ZN(n8557) );
  OAI21_X1 U10057 ( .B1(n8553), .B2(n8992), .A(n8557), .ZN(n8728) );
  INV_X1 U10058 ( .A(n8554), .ZN(n8555) );
  AND2_X1 U10059 ( .A1(n8555), .A2(n8977), .ZN(n8729) );
  INV_X1 U10060 ( .A(n8557), .ZN(n8693) );
  XNOR2_X1 U10061 ( .A(n9167), .B(n8639), .ZN(n8559) );
  NAND2_X1 U10062 ( .A1(n8559), .A2(n8558), .ZN(n8739) );
  INV_X1 U10063 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U10064 ( .A1(n8560), .A2(n8978), .ZN(n8561) );
  AND2_X1 U10065 ( .A1(n8739), .A2(n8561), .ZN(n8692) );
  XNOR2_X1 U10066 ( .A(n9161), .B(n8639), .ZN(n8563) );
  XNOR2_X1 U10067 ( .A(n8563), .B(n8969), .ZN(n8740) );
  NAND2_X1 U10068 ( .A1(n8562), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U10069 ( .A1(n8563), .A2(n8603), .ZN(n8564) );
  NAND2_X1 U10070 ( .A1(n8742), .A2(n8564), .ZN(n8566) );
  XNOR2_X1 U10071 ( .A(n8681), .B(n8639), .ZN(n8565) );
  NAND2_X1 U10072 ( .A1(n8573), .A2(n8567), .ZN(n8676) );
  INV_X1 U10073 ( .A(n8573), .ZN(n8572) );
  XNOR2_X1 U10074 ( .A(n9150), .B(n8568), .ZN(n8569) );
  NAND2_X1 U10075 ( .A1(n8569), .A2(n8921), .ZN(n8700) );
  INV_X1 U10076 ( .A(n8569), .ZN(n8570) );
  NAND2_X1 U10077 ( .A1(n8570), .A2(n8769), .ZN(n8571) );
  NOR3_X1 U10078 ( .A1(n4508), .A2(n8572), .A3(n8574), .ZN(n8575) );
  INV_X1 U10079 ( .A(n8617), .ZN(n8703) );
  OAI21_X1 U10080 ( .B1(n8575), .B2(n8703), .A(n8754), .ZN(n8579) );
  INV_X1 U10081 ( .A(n8939), .ZN(n8768) );
  AOI22_X1 U10082 ( .A1(n8768), .A2(n8733), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8576) );
  OAI21_X1 U10083 ( .B1(n8940), .B2(n8735), .A(n8576), .ZN(n8577) );
  AOI21_X1 U10084 ( .B1(n8942), .B2(n8747), .A(n8577), .ZN(n8578) );
  OAI211_X1 U10085 ( .C1(n9150), .C2(n8764), .A(n8579), .B(n8578), .ZN(
        P2_U3169) );
  INV_X1 U10086 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8583) );
  XNOR2_X1 U10087 ( .A(n9481), .B(n8592), .ZN(n8580) );
  INV_X1 U10088 ( .A(n8581), .ZN(n8582) );
  NOR2_X1 U10089 ( .A1(n8588), .A2(n9715), .ZN(n8585) );
  MUX2_X1 U10090 ( .A(n8583), .B(n8585), .S(n9913), .Z(n8584) );
  OAI21_X1 U10091 ( .B1(n8592), .B2(n9814), .A(n8584), .ZN(P1_U3521) );
  INV_X1 U10092 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8586) );
  MUX2_X1 U10093 ( .A(n8586), .B(n8585), .S(n9926), .Z(n8587) );
  OAI21_X1 U10094 ( .B1(n8592), .B2(n9780), .A(n8587), .ZN(P1_U3553) );
  NAND2_X1 U10095 ( .A1(n8588), .A2(n9853), .ZN(n8591) );
  INV_X1 U10096 ( .A(n9715), .ZN(n8589) );
  NOR2_X1 U10097 ( .A1(n9866), .A2(n8589), .ZN(n9485) );
  AOI21_X1 U10098 ( .B1(n9866), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9485), .ZN(
        n8590) );
  OAI211_X1 U10099 ( .C1(n8592), .C2(n9859), .A(n8591), .B(n8590), .ZN(
        P1_U3263) );
  INV_X1 U10100 ( .A(n8593), .ZN(n9221) );
  INV_X1 U10101 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10456) );
  OAI222_X1 U10102 ( .A1(P1_U3086), .A2(n5922), .B1(n9826), .B2(n9221), .C1(
        n10456), .C2(n8653), .ZN(P1_U3327) );
  NAND2_X1 U10103 ( .A1(n8987), .A2(n8991), .ZN(n8926) );
  NAND2_X1 U10104 ( .A1(n8926), .A2(n8595), .ZN(n8981) );
  NOR2_X1 U10105 ( .A1(n8981), .A2(n8596), .ZN(n8598) );
  NOR2_X1 U10106 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  XNOR2_X1 U10107 ( .A(n8599), .B(n8600), .ZN(n9156) );
  XNOR2_X1 U10108 ( .A(n8601), .B(n8600), .ZN(n8602) );
  OAI222_X1 U10109 ( .A1(n9036), .A2(n8921), .B1(n9004), .B2(n8603), .C1(n8989), .C2(n8602), .ZN(n9154) );
  INV_X1 U10110 ( .A(n9154), .ZN(n8604) );
  MUX2_X1 U10111 ( .A(n8605), .B(n8604), .S(n10023), .Z(n8607) );
  AOI22_X1 U10112 ( .A1(n8681), .A2(n10017), .B1(n10019), .B2(n8677), .ZN(
        n8606) );
  OAI211_X1 U10113 ( .C1(n9156), .C2(n9069), .A(n8607), .B(n8606), .ZN(
        P2_U3210) );
  INV_X1 U10114 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8612) );
  XNOR2_X1 U10115 ( .A(n8608), .B(n8609), .ZN(n8916) );
  XNOR2_X1 U10116 ( .A(n8610), .B(n8609), .ZN(n8611) );
  OAI222_X1 U10117 ( .A1(n9004), .A2(n8939), .B1(n9036), .B2(n8640), .C1(n8989), .C2(n8611), .ZN(n8911) );
  AOI21_X1 U10118 ( .B1(n10045), .B2(n8916), .A(n8911), .ZN(n8614) );
  MUX2_X1 U10119 ( .A(n8612), .B(n8614), .S(n10052), .Z(n8613) );
  OAI21_X1 U10120 ( .B1(n8914), .B2(n9174), .A(n8613), .ZN(P2_U3453) );
  INV_X1 U10121 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8615) );
  MUX2_X1 U10122 ( .A(n8615), .B(n8614), .S(n10065), .Z(n8616) );
  OAI21_X1 U10123 ( .B1(n8914), .B2(n9101), .A(n8616), .ZN(P2_U3485) );
  NAND2_X1 U10124 ( .A1(n8617), .A2(n8700), .ZN(n8622) );
  XNOR2_X1 U10125 ( .A(n8618), .B(n8639), .ZN(n8619) );
  NAND2_X1 U10126 ( .A1(n8619), .A2(n8939), .ZN(n8625) );
  INV_X1 U10127 ( .A(n8619), .ZN(n8620) );
  NAND2_X1 U10128 ( .A1(n8620), .A2(n8768), .ZN(n8621) );
  NAND2_X1 U10129 ( .A1(n8622), .A2(n8701), .ZN(n8626) );
  INV_X1 U10130 ( .A(n8626), .ZN(n8704) );
  INV_X1 U10131 ( .A(n8625), .ZN(n8624) );
  XNOR2_X1 U10132 ( .A(n8914), .B(n8623), .ZN(n8635) );
  XNOR2_X1 U10133 ( .A(n8635), .B(n8922), .ZN(n8627) );
  NOR3_X1 U10134 ( .A1(n8704), .A2(n8624), .A3(n8627), .ZN(n8630) );
  NAND2_X1 U10135 ( .A1(n8626), .A2(n8625), .ZN(n8628) );
  INV_X1 U10136 ( .A(n8638), .ZN(n8629) );
  OAI21_X1 U10137 ( .B1(n8630), .B2(n8629), .A(n8754), .ZN(n8634) );
  AOI22_X1 U10138 ( .A1(n8768), .A2(n8761), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8631) );
  OAI21_X1 U10139 ( .B1(n8640), .B2(n8757), .A(n8631), .ZN(n8632) );
  AOI21_X1 U10140 ( .B1(n8912), .B2(n8747), .A(n8632), .ZN(n8633) );
  OAI211_X1 U10141 ( .C1(n8914), .C2(n8764), .A(n8634), .B(n8633), .ZN(
        P2_U3180) );
  INV_X1 U10142 ( .A(n8635), .ZN(n8636) );
  XNOR2_X1 U10143 ( .A(n9140), .B(n8639), .ZN(n8642) );
  XNOR2_X1 U10144 ( .A(n8642), .B(n8640), .ZN(n8668) );
  INV_X1 U10145 ( .A(n8642), .ZN(n8643) );
  NAND2_X1 U10146 ( .A1(n8643), .A2(n8891), .ZN(n8644) );
  NAND2_X1 U10147 ( .A1(n8669), .A2(n8644), .ZN(n8647) );
  XNOR2_X1 U10148 ( .A(n8888), .B(n8645), .ZN(n8646) );
  XNOR2_X1 U10149 ( .A(n8647), .B(n8646), .ZN(n8652) );
  AOI22_X1 U10150 ( .A1(n8891), .A2(n8761), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8649) );
  NAND2_X1 U10151 ( .A1(n8897), .A2(n8747), .ZN(n8648) );
  OAI211_X1 U10152 ( .C1(n8767), .C2(n8757), .A(n8649), .B(n8648), .ZN(n8650)
         );
  AOI21_X1 U10153 ( .B1(n9134), .B2(n8723), .A(n8650), .ZN(n8651) );
  OAI21_X1 U10154 ( .B1(n8652), .B2(n8725), .A(n8651), .ZN(P2_U3160) );
  OAI222_X1 U10155 ( .A1(n5901), .A2(P1_U3086), .B1(n9826), .B2(n8654), .C1(
        n10415), .C2(n8653), .ZN(P1_U3336) );
  NOR2_X1 U10156 ( .A1(n10023), .A2(n8656), .ZN(n8658) );
  NOR2_X1 U10157 ( .A1(n8657), .A2(n9061), .ZN(n8881) );
  AOI211_X1 U10158 ( .C1(n8659), .C2(n10017), .A(n8658), .B(n8881), .ZN(n8663)
         );
  NAND2_X1 U10159 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  OAI211_X1 U10160 ( .C1(n8655), .C2(n8033), .A(n8663), .B(n8662), .ZN(
        P2_U3204) );
  INV_X1 U10161 ( .A(n8664), .ZN(n9822) );
  OAI222_X1 U10162 ( .A1(n9216), .A2(n8666), .B1(n8665), .B2(n9822), .C1(
        P2_U3151), .C2(n6239), .ZN(P2_U3265) );
  INV_X1 U10163 ( .A(n9140), .ZN(n8675) );
  AOI21_X1 U10164 ( .B1(n8667), .B2(n8668), .A(n8725), .ZN(n8670) );
  NAND2_X1 U10165 ( .A1(n8670), .A2(n8669), .ZN(n8674) );
  AOI22_X1 U10166 ( .A1(n8905), .A2(n8733), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8671) );
  OAI21_X1 U10167 ( .B1(n8922), .B2(n8735), .A(n8671), .ZN(n8672) );
  AOI21_X1 U10168 ( .B1(n8901), .B2(n8747), .A(n8672), .ZN(n8673) );
  OAI211_X1 U10169 ( .C1(n8675), .C2(n8764), .A(n8674), .B(n8673), .ZN(
        P2_U3154) );
  AOI21_X1 U10170 ( .B1(n8957), .B2(n8676), .A(n4508), .ZN(n8683) );
  AOI22_X1 U10171 ( .A1(n8761), .A2(n8969), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8679) );
  NAND2_X1 U10172 ( .A1(n8747), .A2(n8677), .ZN(n8678) );
  OAI211_X1 U10173 ( .C1(n8921), .C2(n8757), .A(n8679), .B(n8678), .ZN(n8680)
         );
  AOI21_X1 U10174 ( .B1(n8681), .B2(n8723), .A(n8680), .ZN(n8682) );
  OAI21_X1 U10175 ( .B1(n8683), .B2(n8725), .A(n8682), .ZN(P2_U3156) );
  NAND2_X1 U10176 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8870) );
  OAI21_X1 U10177 ( .B1(n8757), .B2(n8992), .A(n8870), .ZN(n8684) );
  AOI21_X1 U10178 ( .B1(n8761), .B2(n6812), .A(n8684), .ZN(n8685) );
  OAI21_X1 U10179 ( .B1(n8997), .B2(n8758), .A(n8685), .ZN(n8690) );
  AOI211_X1 U10180 ( .C1(n8688), .C2(n8687), .A(n8725), .B(n8730), .ZN(n8689)
         );
  AOI211_X1 U10181 ( .C1(n9178), .C2(n8723), .A(n8690), .B(n8689), .ZN(n8691)
         );
  INV_X1 U10182 ( .A(n8691), .ZN(P2_U3159) );
  NOR3_X1 U10183 ( .A1(n4521), .A2(n8693), .A3(n8692), .ZN(n8694) );
  OAI21_X1 U10184 ( .B1(n4990), .B2(n8694), .A(n8754), .ZN(n8698) );
  AOI22_X1 U10185 ( .A1(n8733), .A2(n8969), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8695) );
  OAI21_X1 U10186 ( .B1(n8992), .B2(n8735), .A(n8695), .ZN(n8696) );
  AOI21_X1 U10187 ( .B1(n8966), .B2(n8747), .A(n8696), .ZN(n8697) );
  OAI211_X1 U10188 ( .C1(n8699), .C2(n8764), .A(n8698), .B(n8697), .ZN(
        P2_U3163) );
  INV_X1 U10189 ( .A(n8700), .ZN(n8702) );
  NOR3_X1 U10190 ( .A1(n8703), .A2(n8702), .A3(n8701), .ZN(n8705) );
  OAI21_X1 U10191 ( .B1(n8705), .B2(n8704), .A(n8754), .ZN(n8709) );
  AOI22_X1 U10192 ( .A1(n8904), .A2(n8733), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8706) );
  OAI21_X1 U10193 ( .B1(n8921), .B2(n8735), .A(n8706), .ZN(n8707) );
  AOI21_X1 U10194 ( .B1(n8924), .B2(n8747), .A(n8707), .ZN(n8708) );
  OAI211_X1 U10195 ( .C1(n9145), .C2(n8764), .A(n8709), .B(n8708), .ZN(
        P2_U3165) );
  XNOR2_X1 U10196 ( .A(n8710), .B(n9037), .ZN(n8711) );
  XNOR2_X1 U10197 ( .A(n8712), .B(n8711), .ZN(n8717) );
  INV_X1 U10198 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10470) );
  NOR2_X1 U10199 ( .A1(n10470), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8825) );
  NOR2_X1 U10200 ( .A1(n8757), .A2(n9005), .ZN(n8713) );
  AOI211_X1 U10201 ( .C1(n8761), .C2(n9058), .A(n8825), .B(n8713), .ZN(n8714)
         );
  OAI21_X1 U10202 ( .B1(n9031), .B2(n8758), .A(n8714), .ZN(n8715) );
  AOI21_X1 U10203 ( .B1(n9188), .B2(n8723), .A(n8715), .ZN(n8716) );
  OAI21_X1 U10204 ( .B1(n8717), .B2(n8725), .A(n8716), .ZN(P2_U3166) );
  AOI21_X1 U10205 ( .B1(n8719), .B2(n8718), .A(n8753), .ZN(n8726) );
  NOR2_X1 U10206 ( .A1(n8758), .A2(n9018), .ZN(n8722) );
  NAND2_X1 U10207 ( .A1(n8761), .A2(n9016), .ZN(n8720) );
  NAND2_X1 U10208 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8843) );
  OAI211_X1 U10209 ( .C1(n8757), .C2(n8993), .A(n8720), .B(n8843), .ZN(n8721)
         );
  AOI211_X1 U10210 ( .C1(n9110), .C2(n8723), .A(n8722), .B(n8721), .ZN(n8724)
         );
  OAI21_X1 U10211 ( .B1(n8726), .B2(n8725), .A(n8724), .ZN(P2_U3168) );
  OAI21_X1 U10212 ( .B1(n8730), .B2(n8729), .A(n8728), .ZN(n8731) );
  INV_X1 U10213 ( .A(n8731), .ZN(n8732) );
  OAI21_X1 U10214 ( .B1(n4521), .B2(n8732), .A(n8754), .ZN(n8738) );
  AOI22_X1 U10215 ( .A1(n8733), .A2(n8978), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8734) );
  OAI21_X1 U10216 ( .B1(n9003), .B2(n8735), .A(n8734), .ZN(n8736) );
  AOI21_X1 U10217 ( .B1(n8982), .B2(n8747), .A(n8736), .ZN(n8737) );
  OAI211_X1 U10218 ( .C1(n9175), .C2(n8764), .A(n8738), .B(n8737), .ZN(
        P2_U3173) );
  INV_X1 U10219 ( .A(n9161), .ZN(n8750) );
  INV_X1 U10220 ( .A(n8739), .ZN(n8741) );
  NOR3_X1 U10221 ( .A1(n4990), .A2(n8741), .A3(n8740), .ZN(n8744) );
  INV_X1 U10222 ( .A(n8742), .ZN(n8743) );
  OAI21_X1 U10223 ( .B1(n8744), .B2(n8743), .A(n8754), .ZN(n8749) );
  AOI22_X1 U10224 ( .A1(n8761), .A2(n8978), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8745) );
  OAI21_X1 U10225 ( .B1(n8940), .B2(n8757), .A(n8745), .ZN(n8746) );
  AOI21_X1 U10226 ( .B1(n8960), .B2(n8747), .A(n8746), .ZN(n8748) );
  OAI211_X1 U10227 ( .C1(n8750), .C2(n8764), .A(n8749), .B(n8748), .ZN(
        P2_U3175) );
  NOR3_X1 U10228 ( .A1(n8753), .A2(n8752), .A3(n8751), .ZN(n8755) );
  OAI21_X1 U10229 ( .B1(n4575), .B2(n8755), .A(n8754), .ZN(n8763) );
  OAI21_X1 U10230 ( .B1(n8757), .B2(n9003), .A(n8756), .ZN(n8760) );
  NOR2_X1 U10231 ( .A1(n8758), .A2(n9008), .ZN(n8759) );
  AOI211_X1 U10232 ( .C1(n8761), .C2(n9029), .A(n8760), .B(n8759), .ZN(n8762)
         );
  OAI211_X1 U10233 ( .C1(n8765), .C2(n8764), .A(n8763), .B(n8762), .ZN(
        P2_U3178) );
  MUX2_X1 U10234 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8766), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10235 ( .A(n8767), .ZN(n8890) );
  MUX2_X1 U10236 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8890), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10237 ( .A(n8905), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8779), .Z(
        P2_U3519) );
  MUX2_X1 U10238 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8891), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8904), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10241 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8769), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10242 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8969), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8978), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10244 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8970), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10245 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8977), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n6812), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10247 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9029), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10248 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9016), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10249 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9058), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10250 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9047), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10251 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9056), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10252 ( .A(n8770), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8779), .Z(
        P2_U3503) );
  MUX2_X1 U10253 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8771), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10254 ( .A(n8772), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8779), .Z(
        P2_U3501) );
  MUX2_X1 U10255 ( .A(n8773), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8779), .Z(
        P2_U3499) );
  MUX2_X1 U10256 ( .A(n8774), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8779), .Z(
        P2_U3498) );
  MUX2_X1 U10257 ( .A(n8775), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8779), .Z(
        P2_U3497) );
  MUX2_X1 U10258 ( .A(n8776), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8779), .Z(
        P2_U3496) );
  MUX2_X1 U10259 ( .A(n8777), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8779), .Z(
        P2_U3495) );
  MUX2_X1 U10260 ( .A(n8778), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8779), .Z(
        P2_U3494) );
  MUX2_X1 U10261 ( .A(n8780), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8779), .Z(
        P2_U3493) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8781), .S(P2_U3893), .Z(
        P2_U3491) );
  AND3_X1 U10263 ( .A1(n8784), .A2(n8783), .A3(n8782), .ZN(n8785) );
  OAI21_X1 U10264 ( .B1(n8786), .B2(n8785), .A(n9993), .ZN(n8803) );
  INV_X1 U10265 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10094) );
  INV_X1 U10266 ( .A(n8787), .ZN(n8788) );
  OAI21_X1 U10267 ( .B1(n9982), .B2(n10094), .A(n8788), .ZN(n8794) );
  AOI21_X1 U10268 ( .B1(n8791), .B2(n8790), .A(n8789), .ZN(n8792) );
  NOR2_X1 U10269 ( .A1(n8792), .A2(n9998), .ZN(n8793) );
  AOI211_X1 U10270 ( .C1(n8796), .C2(n8795), .A(n8794), .B(n8793), .ZN(n8802)
         );
  OAI21_X1 U10271 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8800) );
  NAND2_X1 U10272 ( .A1(n8800), .A2(n9994), .ZN(n8801) );
  NAND3_X1 U10273 ( .A1(n8803), .A2(n8802), .A3(n8801), .ZN(P2_U3190) );
  AOI21_X1 U10274 ( .B1(n9048), .B2(n8805), .A(n8804), .ZN(n8819) );
  OAI21_X1 U10275 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8813) );
  NAND2_X1 U10276 ( .A1(n8842), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8810) );
  OAI211_X1 U10277 ( .C1(n9983), .C2(n8811), .A(n8810), .B(n8809), .ZN(n8812)
         );
  AOI21_X1 U10278 ( .B1(n9993), .B2(n8813), .A(n8812), .ZN(n8818) );
  OAI21_X1 U10279 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8815), .A(n8814), .ZN(
        n8816) );
  NAND2_X1 U10280 ( .A1(n8816), .A2(n9994), .ZN(n8817) );
  OAI211_X1 U10281 ( .C1(n8819), .C2(n9998), .A(n8818), .B(n8817), .ZN(
        P2_U3197) );
  AOI21_X1 U10282 ( .B1(n4546), .B2(n8821), .A(n8820), .ZN(n8836) );
  OAI21_X1 U10283 ( .B1(n8824), .B2(n8823), .A(n8822), .ZN(n8834) );
  AOI21_X1 U10284 ( .B1(n8842), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8825), .ZN(
        n8831) );
  OAI21_X1 U10285 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8829) );
  NAND2_X1 U10286 ( .A1(n8829), .A2(n9993), .ZN(n8830) );
  OAI211_X1 U10287 ( .C1(n9983), .C2(n8832), .A(n8831), .B(n8830), .ZN(n8833)
         );
  AOI21_X1 U10288 ( .B1(n8834), .B2(n9994), .A(n8833), .ZN(n8835) );
  OAI21_X1 U10289 ( .B1(n8836), .B2(n9998), .A(n8835), .ZN(P2_U3198) );
  AOI21_X1 U10290 ( .B1(n9019), .B2(n8838), .A(n8837), .ZN(n8853) );
  OAI21_X1 U10291 ( .B1(n8841), .B2(n8840), .A(n8839), .ZN(n8847) );
  NAND2_X1 U10292 ( .A1(n8842), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8844) );
  OAI211_X1 U10293 ( .C1(n9983), .C2(n8845), .A(n8844), .B(n8843), .ZN(n8846)
         );
  AOI21_X1 U10294 ( .B1(n9993), .B2(n8847), .A(n8846), .ZN(n8852) );
  OAI21_X1 U10295 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8849), .A(n8848), .ZN(
        n8850) );
  NAND2_X1 U10296 ( .A1(n8850), .A2(n9994), .ZN(n8851) );
  OAI211_X1 U10297 ( .C1(n8853), .C2(n9998), .A(n8852), .B(n8851), .ZN(
        P2_U3199) );
  OAI21_X1 U10298 ( .B1(n8863), .B2(n8855), .A(n8854), .ZN(n8856) );
  XNOR2_X1 U10299 ( .A(n8869), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U10300 ( .A(n8856), .B(n8865), .ZN(n8877) );
  AOI21_X1 U10301 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8858), .A(n8857), .ZN(
        n8859) );
  XNOR2_X1 U10302 ( .A(n8869), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U10303 ( .A(n8859), .B(n8866), .ZN(n8860) );
  NAND2_X1 U10304 ( .A1(n8860), .A2(n9974), .ZN(n8875) );
  AOI21_X1 U10305 ( .B1(n8863), .B2(n8862), .A(n8861), .ZN(n8868) );
  MUX2_X1 U10306 ( .A(n8866), .B(n8865), .S(n8864), .Z(n8867) );
  XNOR2_X1 U10307 ( .A(n8868), .B(n8867), .ZN(n8873) );
  NOR2_X1 U10308 ( .A1(n9983), .A2(n8869), .ZN(n8872) );
  OAI21_X1 U10309 ( .B1(n9982), .B2(n4711), .A(n8870), .ZN(n8871) );
  AOI211_X1 U10310 ( .C1(n8873), .C2(n9993), .A(n8872), .B(n8871), .ZN(n8874)
         );
  OAI211_X1 U10311 ( .C1(n8877), .C2(n8876), .A(n8875), .B(n8874), .ZN(
        P2_U3201) );
  NAND2_X1 U10312 ( .A1(n9070), .A2(n10017), .ZN(n8882) );
  INV_X1 U10313 ( .A(n8878), .ZN(n8879) );
  NOR2_X1 U10314 ( .A1(n8880), .A2(n8879), .ZN(n9125) );
  AOI21_X1 U10315 ( .B1(n9125), .B2(n10023), .A(n8881), .ZN(n8884) );
  OAI211_X1 U10316 ( .C1(n10023), .C2(n8883), .A(n8882), .B(n8884), .ZN(
        P2_U3202) );
  NAND2_X1 U10317 ( .A1(n9128), .A2(n10017), .ZN(n8885) );
  OAI211_X1 U10318 ( .C1(n10023), .C2(n8886), .A(n8885), .B(n8884), .ZN(
        P2_U3203) );
  XNOR2_X1 U10319 ( .A(n8887), .B(n8888), .ZN(n9137) );
  XNOR2_X1 U10320 ( .A(n8889), .B(n8888), .ZN(n8895) );
  MUX2_X1 U10321 ( .A(n8896), .B(n9132), .S(n10023), .Z(n8899) );
  AOI22_X1 U10322 ( .A1(n9134), .A2(n10017), .B1(n10019), .B2(n8897), .ZN(
        n8898) );
  OAI211_X1 U10323 ( .C1(n9137), .C2(n9069), .A(n8899), .B(n8898), .ZN(
        P2_U3205) );
  XNOR2_X1 U10324 ( .A(n8900), .B(n8902), .ZN(n9143) );
  INV_X1 U10325 ( .A(n8901), .ZN(n8907) );
  XNOR2_X1 U10326 ( .A(n8903), .B(n8902), .ZN(n8906) );
  AOI222_X1 U10327 ( .A1(n9060), .A2(n8906), .B1(n8905), .B2(n9057), .C1(n8904), .C2(n9055), .ZN(n9138) );
  OAI21_X1 U10328 ( .B1(n8907), .B2(n9061), .A(n9138), .ZN(n8908) );
  NAND2_X1 U10329 ( .A1(n8908), .A2(n10023), .ZN(n8910) );
  AOI22_X1 U10330 ( .A1(n9140), .A2(n10017), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n8033), .ZN(n8909) );
  OAI211_X1 U10331 ( .C1(n9143), .C2(n9069), .A(n8910), .B(n8909), .ZN(
        P2_U3206) );
  INV_X1 U10332 ( .A(n8911), .ZN(n8918) );
  AOI22_X1 U10333 ( .A1(n8912), .A2(n10019), .B1(n8033), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8913) );
  OAI21_X1 U10334 ( .B1(n8914), .B2(n8984), .A(n8913), .ZN(n8915) );
  AOI21_X1 U10335 ( .B1(n8916), .B2(n9023), .A(n8915), .ZN(n8917) );
  OAI21_X1 U10336 ( .B1(n8918), .B2(n8033), .A(n8917), .ZN(P2_U3207) );
  NOR2_X1 U10337 ( .A1(n9145), .A2(n9063), .ZN(n8923) );
  XOR2_X1 U10338 ( .A(n8933), .B(n8919), .Z(n8920) );
  OAI222_X1 U10339 ( .A1(n9036), .A2(n8922), .B1(n9004), .B2(n8921), .C1(n8989), .C2(n8920), .ZN(n9144) );
  AOI211_X1 U10340 ( .C1(n10019), .C2(n8924), .A(n8923), .B(n9144), .ZN(n8936)
         );
  NAND2_X1 U10341 ( .A1(n8926), .A2(n8925), .ZN(n8928) );
  NAND2_X1 U10342 ( .A1(n8944), .A2(n8929), .ZN(n8931) );
  NAND2_X1 U10343 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  XOR2_X1 U10344 ( .A(n8933), .B(n8932), .Z(n9146) );
  INV_X1 U10345 ( .A(n9146), .ZN(n8934) );
  AOI22_X1 U10346 ( .A1(n8934), .A2(n9023), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8033), .ZN(n8935) );
  OAI21_X1 U10347 ( .B1(n8936), .B2(n8033), .A(n8935), .ZN(P2_U3208) );
  NOR2_X1 U10348 ( .A1(n9150), .A2(n9063), .ZN(n8941) );
  XNOR2_X1 U10349 ( .A(n8937), .B(n8945), .ZN(n8938) );
  OAI222_X1 U10350 ( .A1(n9004), .A2(n8940), .B1(n9036), .B2(n8939), .C1(n8938), .C2(n8989), .ZN(n9149) );
  AOI211_X1 U10351 ( .C1(n10019), .C2(n8942), .A(n8941), .B(n9149), .ZN(n8949)
         );
  NAND2_X1 U10352 ( .A1(n8944), .A2(n8943), .ZN(n8946) );
  XNOR2_X1 U10353 ( .A(n8946), .B(n8945), .ZN(n9151) );
  INV_X1 U10354 ( .A(n9151), .ZN(n8947) );
  AOI22_X1 U10355 ( .A1(n8947), .A2(n9023), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8033), .ZN(n8948) );
  OAI21_X1 U10356 ( .B1(n8949), .B2(n8033), .A(n8948), .ZN(P2_U3209) );
  NAND2_X1 U10357 ( .A1(n8964), .A2(n8951), .ZN(n8953) );
  NAND2_X1 U10358 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  XNOR2_X1 U10359 ( .A(n8954), .B(n8955), .ZN(n9164) );
  INV_X1 U10360 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U10361 ( .A(n8956), .B(n8955), .ZN(n8958) );
  AOI222_X1 U10362 ( .A1(n9060), .A2(n8958), .B1(n8957), .B2(n9057), .C1(n8978), .C2(n9055), .ZN(n9159) );
  MUX2_X1 U10363 ( .A(n8959), .B(n9159), .S(n10023), .Z(n8962) );
  AOI22_X1 U10364 ( .A1(n9161), .A2(n10017), .B1(n10019), .B2(n8960), .ZN(
        n8961) );
  OAI211_X1 U10365 ( .C1(n9164), .C2(n9069), .A(n8962), .B(n8961), .ZN(
        P2_U3211) );
  NAND2_X1 U10366 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  XNOR2_X1 U10367 ( .A(n8965), .B(n8967), .ZN(n9170) );
  INV_X1 U10368 ( .A(n8966), .ZN(n8972) );
  XNOR2_X1 U10369 ( .A(n8968), .B(n8967), .ZN(n8971) );
  AOI222_X1 U10370 ( .A1(n9060), .A2(n8971), .B1(n8970), .B2(n9055), .C1(n8969), .C2(n9057), .ZN(n9165) );
  OAI21_X1 U10371 ( .B1(n8972), .B2(n9061), .A(n9165), .ZN(n8973) );
  NAND2_X1 U10372 ( .A1(n8973), .A2(n10023), .ZN(n8975) );
  AOI22_X1 U10373 ( .A1(n9167), .A2(n10017), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n8033), .ZN(n8974) );
  OAI211_X1 U10374 ( .C1(n9170), .C2(n9069), .A(n8975), .B(n8974), .ZN(
        P2_U3212) );
  OAI21_X1 U10375 ( .B1(n4559), .B2(n8980), .A(n8976), .ZN(n8979) );
  AOI222_X1 U10376 ( .A1(n9060), .A2(n8979), .B1(n8978), .B2(n9057), .C1(n8977), .C2(n9055), .ZN(n9096) );
  XNOR2_X1 U10377 ( .A(n8981), .B(n8980), .ZN(n9098) );
  AOI22_X1 U10378 ( .A1(n8033), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n10019), 
        .B2(n8982), .ZN(n8983) );
  OAI21_X1 U10379 ( .B1(n9175), .B2(n8984), .A(n8983), .ZN(n8985) );
  AOI21_X1 U10380 ( .B1(n9098), .B2(n9023), .A(n8985), .ZN(n8986) );
  OAI21_X1 U10381 ( .B1(n9096), .B2(n8033), .A(n8986), .ZN(P2_U3213) );
  XNOR2_X1 U10382 ( .A(n8987), .B(n8991), .ZN(n9181) );
  AOI211_X1 U10383 ( .C1(n8991), .C2(n8990), .A(n8989), .B(n8988), .ZN(n8995)
         );
  OAI22_X1 U10384 ( .A1(n8993), .A2(n9004), .B1(n8992), .B2(n9036), .ZN(n8994)
         );
  NOR2_X1 U10385 ( .A1(n8995), .A2(n8994), .ZN(n9176) );
  MUX2_X1 U10386 ( .A(n8996), .B(n9176), .S(n10023), .Z(n9000) );
  INV_X1 U10387 ( .A(n8997), .ZN(n8998) );
  AOI22_X1 U10388 ( .A1(n9178), .A2(n10017), .B1(n10019), .B2(n8998), .ZN(
        n8999) );
  OAI211_X1 U10389 ( .C1(n9181), .C2(n9069), .A(n9000), .B(n8999), .ZN(
        P2_U3214) );
  INV_X1 U10390 ( .A(n9010), .ZN(n9001) );
  XNOR2_X1 U10391 ( .A(n9002), .B(n9001), .ZN(n9007) );
  OAI22_X1 U10392 ( .A1(n9005), .A2(n9004), .B1(n9003), .B2(n9036), .ZN(n9006)
         );
  AOI21_X1 U10393 ( .B1(n9007), .B2(n9060), .A(n9006), .ZN(n9106) );
  OAI22_X1 U10394 ( .A1(n10023), .A2(n5205), .B1(n9008), .B2(n9061), .ZN(n9012) );
  OAI21_X1 U10395 ( .B1(n4586), .B2(n9010), .A(n9009), .ZN(n9105) );
  NOR2_X1 U10396 ( .A1(n9105), .A2(n9069), .ZN(n9011) );
  AOI211_X1 U10397 ( .C1(n10017), .C2(n6813), .A(n9012), .B(n9011), .ZN(n9013)
         );
  OAI21_X1 U10398 ( .B1(n8033), .B2(n9106), .A(n9013), .ZN(P2_U3215) );
  XNOR2_X1 U10399 ( .A(n9014), .B(n9015), .ZN(n9017) );
  AOI222_X1 U10400 ( .A1(n9060), .A2(n9017), .B1(n6812), .B2(n9057), .C1(n9016), .C2(n9055), .ZN(n9113) );
  OAI22_X1 U10401 ( .A1(n10023), .A2(n9019), .B1(n9018), .B2(n9061), .ZN(n9020) );
  AOI21_X1 U10402 ( .B1(n9110), .B2(n10017), .A(n9020), .ZN(n9025) );
  XNOR2_X1 U10403 ( .A(n9022), .B(n9021), .ZN(n9111) );
  NAND2_X1 U10404 ( .A1(n9111), .A2(n9023), .ZN(n9024) );
  OAI211_X1 U10405 ( .C1(n9113), .C2(n8033), .A(n9025), .B(n9024), .ZN(
        P2_U3216) );
  XNOR2_X1 U10406 ( .A(n9026), .B(n9027), .ZN(n9191) );
  NAND2_X1 U10407 ( .A1(n9038), .A2(n9043), .ZN(n9028) );
  XNOR2_X1 U10408 ( .A(n9028), .B(n9027), .ZN(n9030) );
  AOI222_X1 U10409 ( .A1(n9060), .A2(n9030), .B1(n9029), .B2(n9057), .C1(n9058), .C2(n9055), .ZN(n9186) );
  MUX2_X1 U10410 ( .A(n5195), .B(n9186), .S(n10023), .Z(n9034) );
  INV_X1 U10411 ( .A(n9031), .ZN(n9032) );
  AOI22_X1 U10412 ( .A1(n9188), .A2(n10017), .B1(n10019), .B2(n9032), .ZN(
        n9033) );
  OAI211_X1 U10413 ( .C1(n9191), .C2(n9069), .A(n9034), .B(n9033), .ZN(
        P2_U3217) );
  XOR2_X1 U10414 ( .A(n9039), .B(n9035), .Z(n9197) );
  NOR2_X1 U10415 ( .A1(n9037), .A2(n9036), .ZN(n9046) );
  INV_X1 U10416 ( .A(n9038), .ZN(n9044) );
  INV_X1 U10417 ( .A(n9039), .ZN(n9040) );
  OAI21_X1 U10418 ( .B1(n9041), .B2(n9040), .A(n9060), .ZN(n9042) );
  AOI21_X1 U10419 ( .B1(n9044), .B2(n9043), .A(n9042), .ZN(n9045) );
  AOI211_X1 U10420 ( .C1(n9055), .C2(n9047), .A(n9046), .B(n9045), .ZN(n9192)
         );
  MUX2_X1 U10421 ( .A(n9048), .B(n9192), .S(n10023), .Z(n9051) );
  AOI22_X1 U10422 ( .A1(n9194), .A2(n10017), .B1(n10019), .B2(n9049), .ZN(
        n9050) );
  OAI211_X1 U10423 ( .C1(n9197), .C2(n9069), .A(n9051), .B(n9050), .ZN(
        P2_U3218) );
  XOR2_X1 U10424 ( .A(n9052), .B(n9053), .Z(n9205) );
  XNOR2_X1 U10425 ( .A(n9054), .B(n9053), .ZN(n9059) );
  AOI222_X1 U10426 ( .A1(n9060), .A2(n9059), .B1(n9058), .B2(n9057), .C1(n9056), .C2(n9055), .ZN(n9198) );
  INV_X1 U10427 ( .A(n9198), .ZN(n9066) );
  INV_X1 U10428 ( .A(n9201), .ZN(n9064) );
  OAI22_X1 U10429 ( .A1(n9064), .A2(n9063), .B1(n9062), .B2(n9061), .ZN(n9065)
         );
  OAI21_X1 U10430 ( .B1(n9066), .B2(n9065), .A(n10023), .ZN(n9068) );
  NAND2_X1 U10431 ( .A1(n8033), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9067) );
  OAI211_X1 U10432 ( .C1(n9205), .C2(n9069), .A(n9068), .B(n9067), .ZN(
        P2_U3219) );
  NAND2_X1 U10433 ( .A1(n9070), .A2(n9121), .ZN(n9071) );
  NAND2_X1 U10434 ( .A1(n9125), .A2(n10065), .ZN(n9073) );
  OAI211_X1 U10435 ( .C1(n10065), .C2(n9072), .A(n9071), .B(n9073), .ZN(
        P2_U3490) );
  INV_X1 U10436 ( .A(n9128), .ZN(n9075) );
  NAND2_X1 U10437 ( .A1(n10068), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U10438 ( .C1(n9075), .C2(n9101), .A(n9074), .B(n9073), .ZN(
        P2_U3489) );
  INV_X1 U10439 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U10440 ( .A1(n10068), .A2(n9076), .ZN(n9077) );
  NAND2_X1 U10441 ( .A1(n9134), .A2(n9121), .ZN(n9079) );
  OAI211_X1 U10442 ( .C1(n9137), .C2(n9124), .A(n9080), .B(n9079), .ZN(
        P2_U3487) );
  INV_X1 U10443 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9081) );
  MUX2_X1 U10444 ( .A(n9081), .B(n9138), .S(n10065), .Z(n9083) );
  NAND2_X1 U10445 ( .A1(n9140), .A2(n9121), .ZN(n9082) );
  OAI211_X1 U10446 ( .C1(n9124), .C2(n9143), .A(n9083), .B(n9082), .ZN(
        P2_U3486) );
  MUX2_X1 U10447 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9144), .S(n10065), .Z(
        n9085) );
  OAI22_X1 U10448 ( .A1(n9146), .A2(n9124), .B1(n9145), .B2(n9101), .ZN(n9084)
         );
  OR2_X1 U10449 ( .A1(n9085), .A2(n9084), .ZN(P2_U3484) );
  MUX2_X1 U10450 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9149), .S(n10065), .Z(
        n9087) );
  OAI22_X1 U10451 ( .A1(n9151), .A2(n9124), .B1(n9150), .B2(n9101), .ZN(n9086)
         );
  OR2_X1 U10452 ( .A1(n9087), .A2(n9086), .ZN(P2_U3483) );
  MUX2_X1 U10453 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9154), .S(n10065), .Z(
        n9089) );
  OAI22_X1 U10454 ( .A1(n9156), .A2(n9124), .B1(n9155), .B2(n9101), .ZN(n9088)
         );
  OR2_X1 U10455 ( .A1(n9089), .A2(n9088), .ZN(P2_U3482) );
  INV_X1 U10456 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9090) );
  MUX2_X1 U10457 ( .A(n9090), .B(n9159), .S(n10065), .Z(n9092) );
  NAND2_X1 U10458 ( .A1(n9161), .A2(n9121), .ZN(n9091) );
  OAI211_X1 U10459 ( .C1(n9164), .C2(n9124), .A(n9092), .B(n9091), .ZN(
        P2_U3481) );
  MUX2_X1 U10460 ( .A(n9093), .B(n9165), .S(n10065), .Z(n9095) );
  NAND2_X1 U10461 ( .A1(n9167), .A2(n9121), .ZN(n9094) );
  OAI211_X1 U10462 ( .C1(n9124), .C2(n9170), .A(n9095), .B(n9094), .ZN(
        P2_U3480) );
  INV_X1 U10463 ( .A(n9096), .ZN(n9097) );
  AOI21_X1 U10464 ( .B1(n10045), .B2(n9098), .A(n9097), .ZN(n9171) );
  MUX2_X1 U10465 ( .A(n9099), .B(n9171), .S(n10065), .Z(n9100) );
  OAI21_X1 U10466 ( .B1(n9175), .B2(n9101), .A(n9100), .ZN(P2_U3479) );
  MUX2_X1 U10467 ( .A(n9102), .B(n9176), .S(n10065), .Z(n9104) );
  NAND2_X1 U10468 ( .A1(n9178), .A2(n9121), .ZN(n9103) );
  OAI211_X1 U10469 ( .C1(n9181), .C2(n9124), .A(n9104), .B(n9103), .ZN(
        P2_U3478) );
  OR2_X1 U10470 ( .A1(n9105), .A2(n10056), .ZN(n9107) );
  NAND2_X1 U10471 ( .A1(n9107), .A2(n9106), .ZN(n9182) );
  MUX2_X1 U10472 ( .A(n9182), .B(P2_REG1_REG_18__SCAN_IN), .S(n10068), .Z(
        n9108) );
  AOI21_X1 U10473 ( .B1(n9121), .B2(n6813), .A(n9108), .ZN(n9109) );
  INV_X1 U10474 ( .A(n9109), .ZN(P2_U3477) );
  AOI22_X1 U10475 ( .A1(n9111), .A2(n10045), .B1(n10047), .B2(n9110), .ZN(
        n9112) );
  NAND2_X1 U10476 ( .A1(n9113), .A2(n9112), .ZN(n9185) );
  MUX2_X1 U10477 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9185), .S(n10065), .Z(
        P2_U3476) );
  MUX2_X1 U10478 ( .A(n9114), .B(n9186), .S(n10065), .Z(n9116) );
  NAND2_X1 U10479 ( .A1(n9188), .A2(n9121), .ZN(n9115) );
  OAI211_X1 U10480 ( .C1(n9191), .C2(n9124), .A(n9116), .B(n9115), .ZN(
        P2_U3475) );
  MUX2_X1 U10481 ( .A(n9117), .B(n9192), .S(n10065), .Z(n9119) );
  NAND2_X1 U10482 ( .A1(n9194), .A2(n9121), .ZN(n9118) );
  OAI211_X1 U10483 ( .C1(n9124), .C2(n9197), .A(n9119), .B(n9118), .ZN(
        P2_U3474) );
  MUX2_X1 U10484 ( .A(n9120), .B(n9198), .S(n10065), .Z(n9123) );
  NAND2_X1 U10485 ( .A1(n9201), .A2(n9121), .ZN(n9122) );
  OAI211_X1 U10486 ( .C1(n9124), .C2(n9205), .A(n9123), .B(n9122), .ZN(
        P2_U3473) );
  NAND2_X1 U10487 ( .A1(n9125), .A2(n10052), .ZN(n9129) );
  NAND2_X1 U10488 ( .A1(n10061), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9126) );
  OAI211_X1 U10489 ( .C1(n9127), .C2(n9174), .A(n9129), .B(n9126), .ZN(
        P2_U3458) );
  INV_X1 U10490 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U10491 ( .A1(n9128), .A2(n9200), .ZN(n9130) );
  OAI211_X1 U10492 ( .C1(n9131), .C2(n10052), .A(n9130), .B(n9129), .ZN(
        P2_U3457) );
  INV_X1 U10493 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9133) );
  MUX2_X1 U10494 ( .A(n9133), .B(n9132), .S(n10052), .Z(n9136) );
  NAND2_X1 U10495 ( .A1(n9134), .A2(n9200), .ZN(n9135) );
  OAI211_X1 U10496 ( .C1(n9137), .C2(n9204), .A(n9136), .B(n9135), .ZN(
        P2_U3455) );
  INV_X1 U10497 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9139) );
  MUX2_X1 U10498 ( .A(n9139), .B(n9138), .S(n10052), .Z(n9142) );
  NAND2_X1 U10499 ( .A1(n9140), .A2(n9200), .ZN(n9141) );
  OAI211_X1 U10500 ( .C1(n9143), .C2(n9204), .A(n9142), .B(n9141), .ZN(
        P2_U3454) );
  MUX2_X1 U10501 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9144), .S(n10052), .Z(
        n9148) );
  OAI22_X1 U10502 ( .A1(n9146), .A2(n9204), .B1(n9145), .B2(n9174), .ZN(n9147)
         );
  OR2_X1 U10503 ( .A1(n9148), .A2(n9147), .ZN(P2_U3452) );
  MUX2_X1 U10504 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9149), .S(n10052), .Z(
        n9153) );
  OAI22_X1 U10505 ( .A1(n9151), .A2(n9204), .B1(n9150), .B2(n9174), .ZN(n9152)
         );
  OR2_X1 U10506 ( .A1(n9153), .A2(n9152), .ZN(P2_U3451) );
  MUX2_X1 U10507 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9154), .S(n10052), .Z(
        n9158) );
  OAI22_X1 U10508 ( .A1(n9156), .A2(n9204), .B1(n9155), .B2(n9174), .ZN(n9157)
         );
  OR2_X1 U10509 ( .A1(n9158), .A2(n9157), .ZN(P2_U3450) );
  INV_X1 U10510 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9160) );
  MUX2_X1 U10511 ( .A(n9160), .B(n9159), .S(n10052), .Z(n9163) );
  NAND2_X1 U10512 ( .A1(n9161), .A2(n9200), .ZN(n9162) );
  OAI211_X1 U10513 ( .C1(n9164), .C2(n9204), .A(n9163), .B(n9162), .ZN(
        P2_U3449) );
  MUX2_X1 U10514 ( .A(n9166), .B(n9165), .S(n10052), .Z(n9169) );
  NAND2_X1 U10515 ( .A1(n9167), .A2(n9200), .ZN(n9168) );
  OAI211_X1 U10516 ( .C1(n9170), .C2(n9204), .A(n9169), .B(n9168), .ZN(
        P2_U3448) );
  MUX2_X1 U10517 ( .A(n9172), .B(n9171), .S(n10052), .Z(n9173) );
  OAI21_X1 U10518 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(P2_U3447) );
  INV_X1 U10519 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9177) );
  MUX2_X1 U10520 ( .A(n9177), .B(n9176), .S(n10052), .Z(n9180) );
  NAND2_X1 U10521 ( .A1(n9178), .A2(n9200), .ZN(n9179) );
  OAI211_X1 U10522 ( .C1(n9181), .C2(n9204), .A(n9180), .B(n9179), .ZN(
        P2_U3446) );
  MUX2_X1 U10523 ( .A(n9182), .B(P2_REG0_REG_18__SCAN_IN), .S(n10061), .Z(
        n9183) );
  AOI21_X1 U10524 ( .B1(n9200), .B2(n6813), .A(n9183), .ZN(n9184) );
  INV_X1 U10525 ( .A(n9184), .ZN(P2_U3444) );
  MUX2_X1 U10526 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9185), .S(n10052), .Z(
        P2_U3441) );
  INV_X1 U10527 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9187) );
  MUX2_X1 U10528 ( .A(n9187), .B(n9186), .S(n10052), .Z(n9190) );
  NAND2_X1 U10529 ( .A1(n9188), .A2(n9200), .ZN(n9189) );
  OAI211_X1 U10530 ( .C1(n9191), .C2(n9204), .A(n9190), .B(n9189), .ZN(
        P2_U3438) );
  INV_X1 U10531 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9193) );
  MUX2_X1 U10532 ( .A(n9193), .B(n9192), .S(n10052), .Z(n9196) );
  NAND2_X1 U10533 ( .A1(n9194), .A2(n9200), .ZN(n9195) );
  OAI211_X1 U10534 ( .C1(n9197), .C2(n9204), .A(n9196), .B(n9195), .ZN(
        P2_U3435) );
  INV_X1 U10535 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9199) );
  MUX2_X1 U10536 ( .A(n9199), .B(n9198), .S(n10052), .Z(n9203) );
  NAND2_X1 U10537 ( .A1(n9201), .A2(n9200), .ZN(n9202) );
  OAI211_X1 U10538 ( .C1(n9205), .C2(n9204), .A(n9203), .B(n9202), .ZN(
        P2_U3432) );
  MUX2_X1 U10539 ( .A(n9207), .B(P2_D_REG_1__SCAN_IN), .S(n9206), .Z(P2_U3377)
         );
  NAND3_X1 U10540 ( .A1(n9209), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9211) );
  OAI22_X1 U10541 ( .A1(n9208), .A2(n9211), .B1(n9210), .B2(n9216), .ZN(n9212)
         );
  AOI21_X1 U10542 ( .B1(n9816), .B2(n9213), .A(n9212), .ZN(n9214) );
  INV_X1 U10543 ( .A(n9214), .ZN(P2_U3264) );
  INV_X1 U10544 ( .A(n9215), .ZN(n9827) );
  OAI222_X1 U10545 ( .A1(n8665), .A2(n9827), .B1(n6240), .B2(P2_U3151), .C1(
        n9217), .C2(n9216), .ZN(P2_U3266) );
  AOI21_X1 U10546 ( .B1(n9219), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9218), .ZN(
        n9220) );
  OAI21_X1 U10547 ( .B1(n9221), .B2(n8665), .A(n9220), .ZN(P2_U3267) );
  MUX2_X1 U10548 ( .A(n9222), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10549 ( .A(n9223), .ZN(n9227) );
  AOI21_X1 U10550 ( .B1(n9382), .B2(n9225), .A(n9224), .ZN(n9226) );
  AOI22_X1 U10551 ( .A1(n9386), .A2(n9412), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9230) );
  AOI22_X1 U10552 ( .A1(n9393), .A2(n9530), .B1(n9391), .B2(n9411), .ZN(n9229)
         );
  NAND2_X1 U10553 ( .A1(n9529), .A2(n9407), .ZN(n9228) );
  INV_X1 U10554 ( .A(n9236), .ZN(n9240) );
  AND2_X1 U10555 ( .A1(n9233), .A2(n9232), .ZN(n9235) );
  AOI21_X1 U10556 ( .B1(n9236), .B2(n9235), .A(n9234), .ZN(n9237) );
  NOR2_X1 U10557 ( .A1(n9237), .A2(n9402), .ZN(n9238) );
  OAI21_X1 U10558 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9247) );
  INV_X1 U10559 ( .A(n9241), .ZN(n9243) );
  OAI22_X1 U10560 ( .A1(n9355), .A2(n9243), .B1(n9396), .B2(n9242), .ZN(n9244)
         );
  AOI211_X1 U10561 ( .C1(n9391), .C2(n9697), .A(n9245), .B(n9244), .ZN(n9246)
         );
  OAI211_X1 U10562 ( .C1(n9248), .C2(n9299), .A(n9247), .B(n9246), .ZN(
        P1_U3215) );
  AOI21_X1 U10563 ( .B1(n9251), .B2(n9250), .A(n9249), .ZN(n9258) );
  OAI22_X1 U10564 ( .A1(n9376), .A2(n9553), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9252), .ZN(n9255) );
  INV_X1 U10565 ( .A(n9587), .ZN(n9253) );
  OAI22_X1 U10566 ( .A1(n9355), .A2(n9253), .B1(n9396), .B2(n9290), .ZN(n9254)
         );
  OAI21_X1 U10567 ( .B1(n9258), .B2(n9402), .A(n9257), .ZN(P1_U3216) );
  INV_X1 U10568 ( .A(n9259), .ZN(n9261) );
  NOR2_X1 U10569 ( .A1(n9261), .A2(n9260), .ZN(n9345) );
  AOI21_X1 U10570 ( .B1(n9261), .B2(n9260), .A(n9345), .ZN(n9262) );
  NAND2_X1 U10571 ( .A1(n9262), .A2(n9263), .ZN(n9347) );
  OAI21_X1 U10572 ( .B1(n9263), .B2(n9262), .A(n9347), .ZN(n9264) );
  NAND2_X1 U10573 ( .A1(n9264), .A2(n9383), .ZN(n9270) );
  OAI22_X1 U10574 ( .A1(n9355), .A2(n9266), .B1(n9396), .B2(n9265), .ZN(n9267)
         );
  AOI211_X1 U10575 ( .C1(n9391), .C2(n9420), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI211_X1 U10576 ( .C1(n5670), .C2(n9299), .A(n9270), .B(n9269), .ZN(
        P1_U3217) );
  INV_X1 U10577 ( .A(n9271), .ZN(n9273) );
  NAND2_X1 U10578 ( .A1(n9273), .A2(n9272), .ZN(n9372) );
  NAND2_X1 U10579 ( .A1(n9372), .A2(n9373), .ZN(n9278) );
  NAND2_X1 U10580 ( .A1(n9271), .A2(n9274), .ZN(n9371) );
  AND2_X1 U10581 ( .A1(n9278), .A2(n9371), .ZN(n9280) );
  INV_X1 U10582 ( .A(n9275), .ZN(n9276) );
  XNOR2_X1 U10583 ( .A(n9277), .B(n9276), .ZN(n9279) );
  NAND3_X1 U10584 ( .A1(n9278), .A2(n9279), .A3(n9371), .ZN(n9325) );
  OAI211_X1 U10585 ( .C1(n9280), .C2(n9279), .A(n9383), .B(n9325), .ZN(n9284)
         );
  OAI22_X1 U10586 ( .A1(n9355), .A2(n9649), .B1(n9396), .B2(n9687), .ZN(n9281)
         );
  AOI211_X1 U10587 ( .C1(n9391), .C2(n9613), .A(n9282), .B(n9281), .ZN(n9283)
         );
  OAI211_X1 U10588 ( .C1(n9653), .C2(n9299), .A(n9284), .B(n9283), .ZN(
        P1_U3219) );
  XNOR2_X1 U10589 ( .A(n9286), .B(n9285), .ZN(n9287) );
  XNOR2_X1 U10590 ( .A(n9288), .B(n9287), .ZN(n9294) );
  INV_X1 U10591 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9289) );
  OAI22_X1 U10592 ( .A1(n9396), .A2(n9645), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9289), .ZN(n9292) );
  OAI22_X1 U10593 ( .A1(n9355), .A2(n9619), .B1(n9376), .B2(n9290), .ZN(n9291)
         );
  AOI211_X1 U10594 ( .C1(n9618), .C2(n9407), .A(n9292), .B(n9291), .ZN(n9293)
         );
  OAI21_X1 U10595 ( .B1(n9294), .B2(n9402), .A(n9293), .ZN(P1_U3223) );
  OAI21_X1 U10596 ( .B1(n9296), .B2(n9295), .A(n9381), .ZN(n9301) );
  AOI22_X1 U10597 ( .A1(n9391), .A2(n9412), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9298) );
  AOI22_X1 U10598 ( .A1(n9393), .A2(n9563), .B1(n9386), .B2(n9413), .ZN(n9297)
         );
  OAI211_X1 U10599 ( .C1(n9800), .C2(n9299), .A(n9298), .B(n9297), .ZN(n9300)
         );
  AOI21_X1 U10600 ( .B1(n9301), .B2(n9383), .A(n9300), .ZN(n9302) );
  INV_X1 U10601 ( .A(n9302), .ZN(P1_U3225) );
  XNOR2_X1 U10602 ( .A(n5080), .B(n9303), .ZN(n9304) );
  XNOR2_X1 U10603 ( .A(n4568), .B(n9304), .ZN(n9310) );
  AOI22_X1 U10604 ( .A1(n9393), .A2(n9710), .B1(n9391), .B2(n9699), .ZN(n9306)
         );
  OAI211_X1 U10605 ( .C1(n9307), .C2(n9396), .A(n9306), .B(n9305), .ZN(n9308)
         );
  AOI21_X1 U10606 ( .B1(n9709), .B2(n9407), .A(n9308), .ZN(n9309) );
  OAI21_X1 U10607 ( .B1(n9310), .B2(n9402), .A(n9309), .ZN(P1_U3226) );
  XOR2_X1 U10608 ( .A(n9311), .B(n4582), .Z(n9316) );
  AOI22_X1 U10609 ( .A1(n9393), .A2(n9675), .B1(n9386), .B2(n9416), .ZN(n9313)
         );
  OAI211_X1 U10610 ( .C1(n9687), .C2(n9376), .A(n9313), .B(n9312), .ZN(n9314)
         );
  AOI21_X1 U10611 ( .B1(n9770), .B2(n9407), .A(n9314), .ZN(n9315) );
  OAI21_X1 U10612 ( .B1(n9316), .B2(n9402), .A(n9315), .ZN(P1_U3228) );
  NOR3_X1 U10613 ( .A1(n9249), .A2(n9318), .A3(n9317), .ZN(n9319) );
  OAI21_X1 U10614 ( .B1(n4536), .B2(n9319), .A(n9383), .ZN(n9323) );
  AOI22_X1 U10615 ( .A1(n9391), .A2(n9544), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9322) );
  AOI22_X1 U10616 ( .A1(n9393), .A2(n9579), .B1(n9386), .B2(n4954), .ZN(n9321)
         );
  NAND2_X1 U10617 ( .A1(n9741), .A2(n9407), .ZN(n9320) );
  NAND4_X1 U10618 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(
        P1_U3229) );
  NAND2_X1 U10619 ( .A1(n9325), .A2(n9324), .ZN(n9329) );
  NOR2_X1 U10620 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  XNOR2_X1 U10621 ( .A(n9329), .B(n9328), .ZN(n9334) );
  INV_X1 U10622 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9330) );
  OAI22_X1 U10623 ( .A1(n9376), .A2(n9630), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9330), .ZN(n9332) );
  OAI22_X1 U10624 ( .A1(n9355), .A2(n9633), .B1(n9396), .B2(n9663), .ZN(n9331)
         );
  AOI211_X1 U10625 ( .C1(n9756), .C2(n9407), .A(n9332), .B(n9331), .ZN(n9333)
         );
  OAI21_X1 U10626 ( .B1(n9334), .B2(n9402), .A(n9333), .ZN(P1_U3233) );
  XNOR2_X1 U10627 ( .A(n9336), .B(n9335), .ZN(n9337) );
  XNOR2_X1 U10628 ( .A(n9338), .B(n9337), .ZN(n9344) );
  INV_X1 U10629 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9339) );
  OAI22_X1 U10630 ( .A1(n9396), .A2(n9630), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9339), .ZN(n9342) );
  INV_X1 U10631 ( .A(n9598), .ZN(n9340) );
  OAI22_X1 U10632 ( .A1(n9355), .A2(n9340), .B1(n9376), .B2(n9576), .ZN(n9341)
         );
  AOI211_X1 U10633 ( .C1(n9745), .C2(n9407), .A(n9342), .B(n9341), .ZN(n9343)
         );
  OAI21_X1 U10634 ( .B1(n9344), .B2(n9402), .A(n9343), .ZN(P1_U3235) );
  INV_X1 U10635 ( .A(n9345), .ZN(n9346) );
  NAND2_X1 U10636 ( .A1(n9347), .A2(n9346), .ZN(n9351) );
  NAND2_X1 U10637 ( .A1(n9349), .A2(n9348), .ZN(n9350) );
  XNOR2_X1 U10638 ( .A(n9351), .B(n9350), .ZN(n9361) );
  INV_X1 U10639 ( .A(n9352), .ZN(n9354) );
  OAI22_X1 U10640 ( .A1(n9355), .A2(n9354), .B1(n9396), .B2(n9353), .ZN(n9356)
         );
  AOI211_X1 U10641 ( .C1(n9391), .C2(n9419), .A(n9357), .B(n9356), .ZN(n9360)
         );
  NAND2_X1 U10642 ( .A1(n9358), .A2(n9407), .ZN(n9359) );
  OAI211_X1 U10643 ( .C1(n9361), .C2(n9402), .A(n9360), .B(n9359), .ZN(
        P1_U3236) );
  OAI21_X1 U10644 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9365) );
  NAND2_X1 U10645 ( .A1(n9365), .A2(n9383), .ZN(n9370) );
  AOI22_X1 U10646 ( .A1(n9366), .A2(n9407), .B1(n9391), .B2(n9427), .ZN(n9369)
         );
  AOI22_X1 U10647 ( .A1(n9386), .A2(n5545), .B1(n9367), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9368) );
  NAND3_X1 U10648 ( .A1(n9370), .A2(n9369), .A3(n9368), .ZN(P1_U3237) );
  NAND2_X1 U10649 ( .A1(n9372), .A2(n9371), .ZN(n9374) );
  XNOR2_X1 U10650 ( .A(n9374), .B(n9373), .ZN(n9379) );
  AOI22_X1 U10651 ( .A1(n9393), .A2(n9665), .B1(n9386), .B2(n9699), .ZN(n9375)
         );
  NAND2_X1 U10652 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9469) );
  OAI211_X1 U10653 ( .C1(n9663), .C2(n9376), .A(n9375), .B(n9469), .ZN(n9377)
         );
  AOI21_X1 U10654 ( .B1(n9766), .B2(n9407), .A(n9377), .ZN(n9378) );
  OAI21_X1 U10655 ( .B1(n9379), .B2(n9402), .A(n9378), .ZN(P1_U3238) );
  AND2_X1 U10656 ( .A1(n9381), .A2(n9380), .ZN(n9385) );
  OAI211_X1 U10657 ( .C1(n9385), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9390)
         );
  AOI22_X1 U10658 ( .A1(n9386), .A2(n9544), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9389) );
  AOI22_X1 U10659 ( .A1(n9393), .A2(n9538), .B1(n9391), .B2(n9545), .ZN(n9388)
         );
  NAND2_X1 U10660 ( .A1(n9730), .A2(n9407), .ZN(n9387) );
  NAND4_X1 U10661 ( .A1(n9390), .A2(n9389), .A3(n9388), .A4(n9387), .ZN(
        P1_U3240) );
  AOI22_X1 U10662 ( .A1(n9393), .A2(n9392), .B1(n9391), .B2(n9416), .ZN(n9395)
         );
  OAI211_X1 U10663 ( .C1(n9397), .C2(n9396), .A(n9395), .B(n9394), .ZN(n9406)
         );
  INV_X1 U10664 ( .A(n9398), .ZN(n9403) );
  AOI21_X1 U10665 ( .B1(n9403), .B2(n9400), .A(n9399), .ZN(n9401) );
  AOI211_X1 U10666 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9405)
         );
  AOI211_X1 U10667 ( .C1(n9408), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9409)
         );
  INV_X1 U10668 ( .A(n9409), .ZN(P1_U3241) );
  MUX2_X1 U10669 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9410), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10670 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n4975), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10671 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9511), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10672 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9411), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10673 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9545), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10674 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9412), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10675 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9544), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10676 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9413), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10677 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n4954), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10678 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9614), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10679 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9604), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10680 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9613), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10681 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9414), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10682 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9415), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10683 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9699), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10684 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9416), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9697), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9417), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10687 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9418), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10688 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9419), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9420), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9421), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9422), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9423), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9424), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9425), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9426), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9427), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5560), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5545), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10699 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n5964), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10700 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10071) );
  OR2_X1 U10701 ( .A1(n9852), .A2(n10071), .ZN(n9438) );
  AOI22_X1 U10702 ( .A1(n9440), .A2(n9428), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3086), .ZN(n9437) );
  MUX2_X1 U10703 ( .A(n6991), .B(P1_REG1_REG_1__SCAN_IN), .S(n9428), .Z(n9429)
         );
  OAI21_X1 U10704 ( .B1(n5966), .B2(n4796), .A(n9429), .ZN(n9430) );
  NAND3_X1 U10705 ( .A1(n9459), .A2(n9431), .A3(n9430), .ZN(n9436) );
  OAI211_X1 U10706 ( .C1(n9434), .C2(n9433), .A(n9849), .B(n9432), .ZN(n9435)
         );
  NAND4_X1 U10707 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(
        P1_U3244) );
  NAND2_X1 U10708 ( .A1(n9440), .A2(n9439), .ZN(n9451) );
  OAI211_X1 U10709 ( .C1(n9443), .C2(n9442), .A(n9849), .B(n9441), .ZN(n9450)
         );
  OAI211_X1 U10710 ( .C1(n9446), .C2(n9445), .A(n9459), .B(n9444), .ZN(n9449)
         );
  AOI21_X1 U10711 ( .B1(n9455), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9447), .ZN(
        n9448) );
  NAND4_X1 U10712 ( .A1(n9451), .A2(n9450), .A3(n9449), .A4(n9448), .ZN(
        P1_U3246) );
  NOR2_X1 U10713 ( .A1(n9843), .A2(n9452), .ZN(n9453) );
  AOI211_X1 U10714 ( .C1(n9455), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9454), .B(
        n9453), .ZN(n9464) );
  OAI211_X1 U10715 ( .C1(n9457), .C2(n9456), .A(n9849), .B(n4676), .ZN(n9463)
         );
  OAI211_X1 U10716 ( .C1(n9461), .C2(n9460), .A(n9459), .B(n9458), .ZN(n9462)
         );
  NAND3_X1 U10717 ( .A1(n9464), .A2(n9463), .A3(n9462), .ZN(P1_U3248) );
  INV_X1 U10718 ( .A(n9465), .ZN(n9466) );
  AOI211_X1 U10719 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9845), .ZN(n9478)
         );
  INV_X1 U10720 ( .A(n9469), .ZN(n9477) );
  INV_X1 U10721 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9470) );
  NOR2_X1 U10722 ( .A1(n9852), .A2(n9470), .ZN(n9476) );
  AOI211_X1 U10723 ( .C1(n9474), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9475)
         );
  NOR4_X1 U10724 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(n9479)
         );
  OAI21_X1 U10725 ( .B1(n9480), .B2(n9843), .A(n9479), .ZN(P1_U3261) );
  AOI211_X1 U10726 ( .C1(n9483), .C2(n9482), .A(n9707), .B(n9481), .ZN(n9716)
         );
  NAND2_X1 U10727 ( .A1(n9716), .A2(n9853), .ZN(n9487) );
  AND2_X1 U10728 ( .A1(n9866), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9484) );
  NOR2_X1 U10729 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  OAI211_X1 U10730 ( .C1(n9790), .C2(n9859), .A(n9487), .B(n9486), .ZN(
        P1_U3264) );
  NAND2_X1 U10731 ( .A1(n9866), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9488) );
  OAI21_X1 U10732 ( .B1(n9490), .B2(n9489), .A(n9488), .ZN(n9491) );
  AOI21_X1 U10733 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9494) );
  OAI21_X1 U10734 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  AOI21_X1 U10735 ( .B1(n9498), .B2(n9863), .A(n9497), .ZN(n9499) );
  OAI21_X1 U10736 ( .B1(n9500), .B2(n9866), .A(n9499), .ZN(P1_U3356) );
  OAI21_X1 U10737 ( .B1(n9502), .B2(n5893), .A(n9501), .ZN(n9723) );
  INV_X1 U10738 ( .A(n9503), .ZN(n9504) );
  AOI211_X1 U10739 ( .C1(n9720), .C2(n9527), .A(n9707), .B(n9504), .ZN(n9719)
         );
  AOI22_X1 U10740 ( .A1(n9866), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9505), .B2(
        n9856), .ZN(n9506) );
  OAI21_X1 U10741 ( .B1(n4875), .B2(n9859), .A(n9506), .ZN(n9515) );
  OAI21_X1 U10742 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9510) );
  AOI211_X1 U10743 ( .C1(n9719), .C2(n9853), .A(n9515), .B(n9514), .ZN(n9516)
         );
  OAI21_X1 U10744 ( .B1(n9723), .B2(n9693), .A(n9516), .ZN(P1_U3265) );
  OAI21_X1 U10745 ( .B1(n9525), .B2(n9518), .A(n9517), .ZN(n9519) );
  NAND2_X1 U10746 ( .A1(n9519), .A2(n9701), .ZN(n9523) );
  OAI22_X1 U10747 ( .A1(n9554), .A2(n9684), .B1(n9520), .B2(n9686), .ZN(n9521)
         );
  INV_X1 U10748 ( .A(n9521), .ZN(n9522) );
  NAND2_X1 U10749 ( .A1(n9523), .A2(n9522), .ZN(n9724) );
  INV_X1 U10750 ( .A(n9724), .ZN(n9535) );
  XNOR2_X1 U10751 ( .A(n9524), .B(n9525), .ZN(n9726) );
  NAND2_X1 U10752 ( .A1(n9726), .A2(n9863), .ZN(n9534) );
  INV_X1 U10753 ( .A(n9527), .ZN(n9528) );
  AOI211_X1 U10754 ( .C1(n9529), .C2(n4879), .A(n9707), .B(n9528), .ZN(n9725)
         );
  AOI22_X1 U10755 ( .A1(n9866), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9530), .B2(
        n9856), .ZN(n9531) );
  OAI21_X1 U10756 ( .B1(n9795), .B2(n9859), .A(n9531), .ZN(n9532) );
  AOI21_X1 U10757 ( .B1(n9725), .B2(n9853), .A(n9532), .ZN(n9533) );
  OAI211_X1 U10758 ( .C1(n9535), .C2(n9866), .A(n9534), .B(n9533), .ZN(
        P1_U3266) );
  XNOR2_X1 U10759 ( .A(n9537), .B(n9536), .ZN(n9733) );
  AOI211_X1 U10760 ( .C1(n9730), .C2(n9559), .A(n9707), .B(n9526), .ZN(n9729)
         );
  INV_X1 U10761 ( .A(n9730), .ZN(n9540) );
  AOI22_X1 U10762 ( .A1(n9866), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9538), .B2(
        n9856), .ZN(n9539) );
  OAI21_X1 U10763 ( .B1(n9540), .B2(n9859), .A(n9539), .ZN(n9548) );
  OAI21_X1 U10764 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9546) );
  AOI222_X1 U10765 ( .A1(n9701), .A2(n9546), .B1(n9545), .B2(n9698), .C1(n9544), .C2(n9696), .ZN(n9732) );
  NOR2_X1 U10766 ( .A1(n9732), .A2(n9866), .ZN(n9547) );
  AOI211_X1 U10767 ( .C1(n9729), .C2(n9853), .A(n9548), .B(n9547), .ZN(n9549)
         );
  OAI21_X1 U10768 ( .B1(n9733), .B2(n9693), .A(n9549), .ZN(P1_U3267) );
  NAND2_X1 U10769 ( .A1(n9550), .A2(n9558), .ZN(n9551) );
  AOI21_X1 U10770 ( .B1(n9552), .B2(n9551), .A(n9681), .ZN(n9556) );
  OAI22_X1 U10771 ( .A1(n9554), .A2(n9686), .B1(n9553), .B2(n9684), .ZN(n9555)
         );
  INV_X1 U10772 ( .A(n9734), .ZN(n9568) );
  XOR2_X1 U10773 ( .A(n9557), .B(n9558), .Z(n9736) );
  NAND2_X1 U10774 ( .A1(n9736), .A2(n9863), .ZN(n9567) );
  INV_X1 U10775 ( .A(n9577), .ZN(n9561) );
  INV_X1 U10776 ( .A(n9559), .ZN(n9560) );
  AOI211_X1 U10777 ( .C1(n9562), .C2(n9561), .A(n9707), .B(n9560), .ZN(n9735)
         );
  AOI22_X1 U10778 ( .A1(n9866), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9563), .B2(
        n9856), .ZN(n9564) );
  OAI21_X1 U10779 ( .B1(n9800), .B2(n9859), .A(n9564), .ZN(n9565) );
  AOI21_X1 U10780 ( .B1(n9735), .B2(n9853), .A(n9565), .ZN(n9566) );
  OAI211_X1 U10781 ( .C1(n9866), .C2(n9568), .A(n9567), .B(n9566), .ZN(
        P1_U3268) );
  OAI21_X1 U10782 ( .B1(n4538), .B2(n9572), .A(n9569), .ZN(n9743) );
  NAND2_X1 U10783 ( .A1(n9571), .A2(n9570), .ZN(n9573) );
  XNOR2_X1 U10784 ( .A(n9573), .B(n9572), .ZN(n9574) );
  OAI222_X1 U10785 ( .A1(n9684), .A2(n9576), .B1(n9686), .B2(n9575), .C1(n9574), .C2(n9681), .ZN(n9739) );
  INV_X1 U10786 ( .A(n9741), .ZN(n9582) );
  AOI211_X1 U10787 ( .C1(n9741), .C2(n9578), .A(n9707), .B(n9577), .ZN(n9740)
         );
  NAND2_X1 U10788 ( .A1(n9740), .A2(n9853), .ZN(n9581) );
  AOI22_X1 U10789 ( .A1(n9866), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9579), .B2(
        n9856), .ZN(n9580) );
  OAI211_X1 U10790 ( .C1(n9582), .C2(n9859), .A(n9581), .B(n9580), .ZN(n9583)
         );
  AOI21_X1 U10791 ( .B1(n9739), .B2(n9670), .A(n9583), .ZN(n9584) );
  OAI21_X1 U10792 ( .B1(n9743), .B2(n9693), .A(n9584), .ZN(P1_U3269) );
  INV_X1 U10793 ( .A(n9585), .ZN(n9594) );
  NAND2_X1 U10794 ( .A1(n9586), .A2(n9853), .ZN(n9589) );
  AOI22_X1 U10795 ( .A1(n9866), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9587), .B2(
        n9856), .ZN(n9588) );
  OAI211_X1 U10796 ( .C1(n9590), .C2(n9859), .A(n9589), .B(n9588), .ZN(n9591)
         );
  AOI21_X1 U10797 ( .B1(n9670), .B2(n9592), .A(n9591), .ZN(n9593) );
  OAI21_X1 U10798 ( .B1(n9594), .B2(n9693), .A(n9593), .ZN(P1_U3270) );
  XOR2_X1 U10799 ( .A(n9595), .B(n9603), .Z(n9748) );
  INV_X1 U10800 ( .A(n9596), .ZN(n9597) );
  AOI211_X1 U10801 ( .C1(n9745), .C2(n4883), .A(n9707), .B(n9597), .ZN(n9744)
         );
  AOI22_X1 U10802 ( .A1(n9866), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9598), .B2(
        n9856), .ZN(n9599) );
  OAI21_X1 U10803 ( .B1(n9600), .B2(n9859), .A(n9599), .ZN(n9607) );
  OAI21_X1 U10804 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9605) );
  AOI222_X1 U10805 ( .A1(n9701), .A2(n9605), .B1(n4954), .B2(n9698), .C1(n9604), .C2(n9696), .ZN(n9747) );
  NOR2_X1 U10806 ( .A1(n9747), .A2(n9866), .ZN(n9606) );
  AOI211_X1 U10807 ( .C1(n9744), .C2(n9853), .A(n9607), .B(n9606), .ZN(n9608)
         );
  OAI21_X1 U10808 ( .B1(n9748), .B2(n9693), .A(n9608), .ZN(P1_U3271) );
  XOR2_X1 U10809 ( .A(n9609), .B(n9611), .Z(n9751) );
  INV_X1 U10810 ( .A(n9751), .ZN(n9625) );
  OAI21_X1 U10811 ( .B1(n9611), .B2(n4563), .A(n9610), .ZN(n9612) );
  NAND2_X1 U10812 ( .A1(n9612), .A2(n9701), .ZN(n9616) );
  AOI22_X1 U10813 ( .A1(n9614), .A2(n9698), .B1(n9696), .B2(n9613), .ZN(n9615)
         );
  NAND2_X1 U10814 ( .A1(n9616), .A2(n9615), .ZN(n9749) );
  AOI211_X1 U10815 ( .C1(n9618), .C2(n9631), .A(n9707), .B(n9617), .ZN(n9750)
         );
  NAND2_X1 U10816 ( .A1(n9750), .A2(n9853), .ZN(n9622) );
  INV_X1 U10817 ( .A(n9619), .ZN(n9620) );
  AOI22_X1 U10818 ( .A1(n9866), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9620), .B2(
        n9856), .ZN(n9621) );
  OAI211_X1 U10819 ( .C1(n9806), .C2(n9859), .A(n9622), .B(n9621), .ZN(n9623)
         );
  AOI21_X1 U10820 ( .B1(n9670), .B2(n9749), .A(n9623), .ZN(n9624) );
  OAI21_X1 U10821 ( .B1(n9625), .B2(n9693), .A(n9624), .ZN(P1_U3272) );
  XOR2_X1 U10822 ( .A(n9626), .B(n9627), .Z(n9758) );
  XNOR2_X1 U10823 ( .A(n9628), .B(n9627), .ZN(n9629) );
  OAI222_X1 U10824 ( .A1(n9686), .A2(n9630), .B1(n9684), .B2(n9663), .C1(n9681), .C2(n9629), .ZN(n9754) );
  INV_X1 U10825 ( .A(n9631), .ZN(n9632) );
  AOI211_X1 U10826 ( .C1(n9756), .C2(n9646), .A(n9707), .B(n9632), .ZN(n9755)
         );
  NAND2_X1 U10827 ( .A1(n9755), .A2(n9853), .ZN(n9636) );
  INV_X1 U10828 ( .A(n9633), .ZN(n9634) );
  AOI22_X1 U10829 ( .A1(n9866), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9634), .B2(
        n9856), .ZN(n9635) );
  OAI211_X1 U10830 ( .C1(n9637), .C2(n9859), .A(n9636), .B(n9635), .ZN(n9638)
         );
  AOI21_X1 U10831 ( .B1(n9754), .B2(n9670), .A(n9638), .ZN(n9639) );
  OAI21_X1 U10832 ( .B1(n9758), .B2(n9693), .A(n9639), .ZN(P1_U3273) );
  XNOR2_X1 U10833 ( .A(n9641), .B(n9640), .ZN(n9763) );
  XNOR2_X1 U10834 ( .A(n9643), .B(n9642), .ZN(n9644) );
  OAI222_X1 U10835 ( .A1(n9686), .A2(n9645), .B1(n9684), .B2(n9687), .C1(n9644), .C2(n9681), .ZN(n9759) );
  INV_X1 U10836 ( .A(n9664), .ZN(n9648) );
  INV_X1 U10837 ( .A(n9646), .ZN(n9647) );
  AOI211_X1 U10838 ( .C1(n9761), .C2(n9648), .A(n9707), .B(n9647), .ZN(n9760)
         );
  NAND2_X1 U10839 ( .A1(n9760), .A2(n9853), .ZN(n9652) );
  INV_X1 U10840 ( .A(n9649), .ZN(n9650) );
  AOI22_X1 U10841 ( .A1(n9866), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9650), .B2(
        n9856), .ZN(n9651) );
  OAI211_X1 U10842 ( .C1(n9653), .C2(n9859), .A(n9652), .B(n9651), .ZN(n9654)
         );
  AOI21_X1 U10843 ( .B1(n9759), .B2(n9670), .A(n9654), .ZN(n9655) );
  OAI21_X1 U10844 ( .B1(n9763), .B2(n9693), .A(n9655), .ZN(P1_U3274) );
  XNOR2_X1 U10845 ( .A(n9656), .B(n9660), .ZN(n9768) );
  INV_X1 U10846 ( .A(n9657), .ZN(n9658) );
  AOI21_X1 U10847 ( .B1(n9660), .B2(n9659), .A(n9658), .ZN(n9661) );
  OAI222_X1 U10848 ( .A1(n9686), .A2(n9663), .B1(n9684), .B2(n9662), .C1(n9681), .C2(n9661), .ZN(n9764) );
  AOI211_X1 U10849 ( .C1(n9766), .C2(n9673), .A(n9707), .B(n9664), .ZN(n9765)
         );
  NAND2_X1 U10850 ( .A1(n9765), .A2(n9853), .ZN(n9667) );
  AOI22_X1 U10851 ( .A1(n9866), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9665), .B2(
        n9856), .ZN(n9666) );
  OAI211_X1 U10852 ( .C1(n9668), .C2(n9859), .A(n9667), .B(n9666), .ZN(n9669)
         );
  AOI21_X1 U10853 ( .B1(n9764), .B2(n9670), .A(n9669), .ZN(n9671) );
  OAI21_X1 U10854 ( .B1(n9768), .B2(n9693), .A(n9671), .ZN(P1_U3275) );
  XOR2_X1 U10855 ( .A(n9683), .B(n9672), .Z(n9773) );
  INV_X1 U10856 ( .A(n9673), .ZN(n9674) );
  AOI211_X1 U10857 ( .C1(n9770), .C2(n9705), .A(n9707), .B(n9674), .ZN(n9769)
         );
  AOI22_X1 U10858 ( .A1(n9866), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9675), .B2(
        n9856), .ZN(n9676) );
  OAI21_X1 U10859 ( .B1(n9677), .B2(n9859), .A(n9676), .ZN(n9691) );
  NAND2_X1 U10860 ( .A1(n9694), .A2(n9678), .ZN(n9682) );
  INV_X1 U10861 ( .A(n9679), .ZN(n9680) );
  AOI211_X1 U10862 ( .C1(n9683), .C2(n9682), .A(n9681), .B(n9680), .ZN(n9689)
         );
  OAI22_X1 U10863 ( .A1(n9687), .A2(n9686), .B1(n9685), .B2(n9684), .ZN(n9688)
         );
  NOR2_X1 U10864 ( .A1(n9689), .A2(n9688), .ZN(n9772) );
  NOR2_X1 U10865 ( .A1(n9772), .A2(n9866), .ZN(n9690) );
  AOI211_X1 U10866 ( .C1(n9769), .C2(n9853), .A(n9691), .B(n9690), .ZN(n9692)
         );
  OAI21_X1 U10867 ( .B1(n9773), .B2(n9693), .A(n9692), .ZN(P1_U3276) );
  OAI21_X1 U10868 ( .B1(n9704), .B2(n9695), .A(n9694), .ZN(n9700) );
  AOI222_X1 U10869 ( .A1(n9701), .A2(n9700), .B1(n9699), .B2(n9698), .C1(n9697), .C2(n9696), .ZN(n9774) );
  AOI21_X1 U10870 ( .B1(n9704), .B2(n9703), .A(n9702), .ZN(n9777) );
  NAND2_X1 U10871 ( .A1(n9777), .A2(n9863), .ZN(n9714) );
  INV_X1 U10872 ( .A(n9705), .ZN(n9706) );
  AOI211_X1 U10873 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9776)
         );
  AOI22_X1 U10874 ( .A1(n9866), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9710), .B2(
        n9856), .ZN(n9711) );
  OAI21_X1 U10875 ( .B1(n4884), .B2(n9859), .A(n9711), .ZN(n9712) );
  AOI21_X1 U10876 ( .B1(n9776), .B2(n9853), .A(n9712), .ZN(n9713) );
  OAI211_X1 U10877 ( .C1(n9866), .C2(n9774), .A(n9714), .B(n9713), .ZN(
        P1_U3277) );
  INV_X1 U10878 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9717) );
  NOR2_X1 U10879 ( .A1(n9716), .A2(n9715), .ZN(n9787) );
  MUX2_X1 U10880 ( .A(n9717), .B(n9787), .S(n9926), .Z(n9718) );
  OAI21_X1 U10881 ( .B1(n9790), .B2(n9780), .A(n9718), .ZN(P1_U3552) );
  AOI21_X1 U10882 ( .B1(n9829), .B2(n9720), .A(n9719), .ZN(n9721) );
  OAI211_X1 U10883 ( .C1(n9723), .C2(n9786), .A(n9722), .B(n9721), .ZN(n9791)
         );
  MUX2_X1 U10884 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9791), .S(n9926), .Z(
        P1_U3550) );
  INV_X1 U10885 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9727) );
  AOI211_X1 U10886 ( .C1(n9726), .C2(n9909), .A(n9725), .B(n9724), .ZN(n9792)
         );
  MUX2_X1 U10887 ( .A(n9727), .B(n9792), .S(n9926), .Z(n9728) );
  OAI21_X1 U10888 ( .B1(n9795), .B2(n9780), .A(n9728), .ZN(P1_U3549) );
  AOI21_X1 U10889 ( .B1(n9829), .B2(n9730), .A(n9729), .ZN(n9731) );
  OAI211_X1 U10890 ( .C1(n9733), .C2(n9786), .A(n9732), .B(n9731), .ZN(n9796)
         );
  MUX2_X1 U10891 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9796), .S(n9926), .Z(
        P1_U3548) );
  INV_X1 U10892 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9737) );
  AOI211_X1 U10893 ( .C1(n9736), .C2(n9909), .A(n9735), .B(n9734), .ZN(n9797)
         );
  MUX2_X1 U10894 ( .A(n9737), .B(n9797), .S(n9926), .Z(n9738) );
  OAI21_X1 U10895 ( .B1(n9800), .B2(n9780), .A(n9738), .ZN(P1_U3547) );
  AOI211_X1 U10896 ( .C1(n9829), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9742)
         );
  OAI21_X1 U10897 ( .B1(n9743), .B2(n9786), .A(n9742), .ZN(n9801) );
  MUX2_X1 U10898 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9801), .S(n9926), .Z(
        P1_U3546) );
  AOI21_X1 U10899 ( .B1(n9829), .B2(n9745), .A(n9744), .ZN(n9746) );
  OAI211_X1 U10900 ( .C1(n9748), .C2(n9786), .A(n9747), .B(n9746), .ZN(n9802)
         );
  MUX2_X1 U10901 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9802), .S(n9926), .Z(
        P1_U3544) );
  AOI211_X1 U10902 ( .C1(n9751), .C2(n9909), .A(n9750), .B(n9749), .ZN(n9803)
         );
  MUX2_X1 U10903 ( .A(n9752), .B(n9803), .S(n9926), .Z(n9753) );
  OAI21_X1 U10904 ( .B1(n9806), .B2(n9780), .A(n9753), .ZN(P1_U3543) );
  AOI211_X1 U10905 ( .C1(n9829), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9757)
         );
  OAI21_X1 U10906 ( .B1(n9758), .B2(n9786), .A(n9757), .ZN(n9807) );
  MUX2_X1 U10907 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9807), .S(n9926), .Z(
        P1_U3542) );
  AOI211_X1 U10908 ( .C1(n9829), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9762)
         );
  OAI21_X1 U10909 ( .B1(n9763), .B2(n9786), .A(n9762), .ZN(n9808) );
  MUX2_X1 U10910 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9808), .S(n9926), .Z(
        P1_U3541) );
  AOI211_X1 U10911 ( .C1(n9829), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9767)
         );
  OAI21_X1 U10912 ( .B1(n9768), .B2(n9786), .A(n9767), .ZN(n9809) );
  MUX2_X1 U10913 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9809), .S(n9926), .Z(
        P1_U3540) );
  AOI21_X1 U10914 ( .B1(n9829), .B2(n9770), .A(n9769), .ZN(n9771) );
  OAI211_X1 U10915 ( .C1(n9773), .C2(n9786), .A(n9772), .B(n9771), .ZN(n9810)
         );
  MUX2_X1 U10916 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9810), .S(n9926), .Z(
        P1_U3539) );
  INV_X1 U10917 ( .A(n9774), .ZN(n9775) );
  AOI211_X1 U10918 ( .C1(n9777), .C2(n9909), .A(n9776), .B(n9775), .ZN(n9811)
         );
  MUX2_X1 U10919 ( .A(n9778), .B(n9811), .S(n9926), .Z(n9779) );
  OAI21_X1 U10920 ( .B1(n4884), .B2(n9780), .A(n9779), .ZN(P1_U3538) );
  AOI211_X1 U10921 ( .C1(n9829), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9784)
         );
  OAI21_X1 U10922 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9815) );
  MUX2_X1 U10923 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9815), .S(n9926), .Z(
        P1_U3536) );
  INV_X1 U10924 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9788) );
  MUX2_X1 U10925 ( .A(n9788), .B(n9787), .S(n9913), .Z(n9789) );
  OAI21_X1 U10926 ( .B1(n9790), .B2(n9814), .A(n9789), .ZN(P1_U3520) );
  MUX2_X1 U10927 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9791), .S(n9913), .Z(
        P1_U3518) );
  INV_X1 U10928 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U10929 ( .A(n9793), .B(n9792), .S(n9913), .Z(n9794) );
  OAI21_X1 U10930 ( .B1(n9795), .B2(n9814), .A(n9794), .ZN(P1_U3517) );
  MUX2_X1 U10931 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9796), .S(n9913), .Z(
        P1_U3516) );
  INV_X1 U10932 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U10933 ( .A(n9798), .B(n9797), .S(n9913), .Z(n9799) );
  OAI21_X1 U10934 ( .B1(n9800), .B2(n9814), .A(n9799), .ZN(P1_U3515) );
  MUX2_X1 U10935 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9801), .S(n9913), .Z(
        P1_U3514) );
  MUX2_X1 U10936 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9802), .S(n9913), .Z(
        P1_U3512) );
  INV_X1 U10937 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9804) );
  MUX2_X1 U10938 ( .A(n9804), .B(n9803), .S(n9913), .Z(n9805) );
  OAI21_X1 U10939 ( .B1(n9806), .B2(n9814), .A(n9805), .ZN(P1_U3511) );
  MUX2_X1 U10940 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9807), .S(n9913), .Z(
        P1_U3510) );
  MUX2_X1 U10941 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9808), .S(n9913), .Z(
        P1_U3509) );
  MUX2_X1 U10942 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9809), .S(n9913), .Z(
        P1_U3507) );
  MUX2_X1 U10943 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9810), .S(n9913), .Z(
        P1_U3504) );
  INV_X1 U10944 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9812) );
  MUX2_X1 U10945 ( .A(n9812), .B(n9811), .S(n9913), .Z(n9813) );
  OAI21_X1 U10946 ( .B1(n4884), .B2(n9814), .A(n9813), .ZN(P1_U3501) );
  MUX2_X1 U10947 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9815), .S(n9913), .Z(
        P1_U3495) );
  INV_X1 U10948 ( .A(n9816), .ZN(n9820) );
  NOR4_X1 U10949 ( .A1(n9817), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5625), .ZN(n9818) );
  AOI21_X1 U10950 ( .B1(n9823), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9818), .ZN(
        n9819) );
  OAI21_X1 U10951 ( .B1(n9820), .B2(n9826), .A(n9819), .ZN(P1_U3324) );
  AOI22_X1 U10952 ( .A1(n5497), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9823), .ZN(n9821) );
  OAI21_X1 U10953 ( .B1(n9822), .B2(n9826), .A(n9821), .ZN(P1_U3325) );
  AOI22_X1 U10954 ( .A1(n9824), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9823), .ZN(n9825) );
  OAI21_X1 U10955 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(P1_U3326) );
  MUX2_X1 U10956 ( .A(n9828), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10957 ( .A(n9829), .ZN(n9906) );
  OAI211_X1 U10958 ( .C1(n9832), .C2(n9906), .A(n9831), .B(n9830), .ZN(n9833)
         );
  AOI21_X1 U10959 ( .B1(n9834), .B2(n9909), .A(n9833), .ZN(n9836) );
  AOI22_X1 U10960 ( .A1(n9926), .A2(n9836), .B1(n7907), .B2(n9923), .ZN(
        P1_U3537) );
  INV_X1 U10961 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10962 ( .A1(n9913), .A2(n9836), .B1(n9835), .B2(n9911), .ZN(
        P1_U3498) );
  XNOR2_X1 U10963 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10964 ( .A(P1_RD_REG_SCAN_IN), .B(n4788), .Z(U126) );
  INV_X1 U10965 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10111) );
  OAI21_X1 U10966 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(n9848) );
  AOI21_X1 U10967 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9846) );
  OAI22_X1 U10968 ( .A1(n9846), .A2(n9845), .B1(n9844), .B2(n9843), .ZN(n9847)
         );
  AOI21_X1 U10969 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9851) );
  OAI211_X1 U10970 ( .C1(n9852), .C2(n10111), .A(n9851), .B(n9850), .ZN(
        P1_U3255) );
  NAND2_X1 U10971 ( .A1(n9854), .A2(n9853), .ZN(n9858) );
  AOI22_X1 U10972 ( .A1(n9866), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9856), .B2(
        n9855), .ZN(n9857) );
  OAI211_X1 U10973 ( .C1(n9860), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9861)
         );
  AOI21_X1 U10974 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9864) );
  OAI21_X1 U10975 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(P1_U3290) );
  AND2_X1 U10976 ( .A1(n9874), .A2(n9867), .ZN(n9871) );
  AND2_X1 U10977 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9868), .ZN(P1_U3294) );
  AND2_X1 U10978 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9868), .ZN(P1_U3295) );
  AND2_X1 U10979 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9868), .ZN(P1_U3296) );
  AND2_X1 U10980 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9868), .ZN(P1_U3297) );
  AND2_X1 U10981 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9868), .ZN(P1_U3298) );
  AND2_X1 U10982 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9868), .ZN(P1_U3299) );
  AND2_X1 U10983 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9868), .ZN(P1_U3300) );
  AND2_X1 U10984 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9868), .ZN(P1_U3301) );
  AND2_X1 U10985 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9868), .ZN(P1_U3302) );
  AND2_X1 U10986 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9868), .ZN(P1_U3303) );
  AND2_X1 U10987 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9868), .ZN(P1_U3304) );
  AND2_X1 U10988 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9868), .ZN(P1_U3305) );
  AND2_X1 U10989 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9868), .ZN(P1_U3306) );
  AND2_X1 U10990 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9868), .ZN(P1_U3307) );
  AND2_X1 U10991 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9868), .ZN(P1_U3308) );
  AND2_X1 U10992 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9868), .ZN(P1_U3309) );
  AND2_X1 U10993 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9868), .ZN(P1_U3310) );
  AND2_X1 U10994 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9868), .ZN(P1_U3311) );
  AND2_X1 U10995 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9868), .ZN(P1_U3312) );
  AND2_X1 U10996 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9868), .ZN(P1_U3313) );
  AND2_X1 U10997 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9868), .ZN(P1_U3314) );
  AND2_X1 U10998 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9868), .ZN(P1_U3315) );
  AND2_X1 U10999 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9868), .ZN(P1_U3316) );
  AND2_X1 U11000 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9868), .ZN(P1_U3317) );
  AND2_X1 U11001 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9868), .ZN(P1_U3318) );
  AND2_X1 U11002 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9868), .ZN(P1_U3319) );
  NOR2_X1 U11003 ( .A1(n9871), .A2(n9869), .ZN(P1_U3320) );
  NOR2_X1 U11004 ( .A1(n9871), .A2(n9870), .ZN(P1_U3321) );
  NOR2_X1 U11005 ( .A1(n9871), .A2(n10392), .ZN(P1_U3322) );
  NOR2_X1 U11006 ( .A1(n9871), .A2(n10428), .ZN(P1_U3323) );
  INV_X1 U11007 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9873) );
  OAI21_X1 U11008 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(P1_U3439) );
  OAI21_X1 U11009 ( .B1(n5559), .B2(n9906), .A(n9875), .ZN(n9876) );
  AOI21_X1 U11010 ( .B1(n9877), .B2(n9909), .A(n9876), .ZN(n9878) );
  AND2_X1 U11011 ( .A1(n9879), .A2(n9878), .ZN(n9915) );
  INV_X1 U11012 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U11013 ( .A1(n9913), .A2(n9915), .B1(n9880), .B2(n9911), .ZN(
        P1_U3459) );
  OAI21_X1 U11014 ( .B1(n9882), .B2(n9906), .A(n9881), .ZN(n9884) );
  AOI211_X1 U11015 ( .C1(n9909), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9916)
         );
  INV_X1 U11016 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9886) );
  AOI22_X1 U11017 ( .A1(n9913), .A2(n9916), .B1(n9886), .B2(n9911), .ZN(
        P1_U3471) );
  OAI21_X1 U11018 ( .B1(n9888), .B2(n9906), .A(n9887), .ZN(n9890) );
  AOI211_X1 U11019 ( .C1(n9909), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9918)
         );
  INV_X1 U11020 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U11021 ( .A1(n9913), .A2(n9918), .B1(n9892), .B2(n9911), .ZN(
        P1_U3477) );
  OAI211_X1 U11022 ( .C1(n9895), .C2(n9906), .A(n9894), .B(n9893), .ZN(n9896)
         );
  AOI21_X1 U11023 ( .B1(n9909), .B2(n9897), .A(n9896), .ZN(n9920) );
  INV_X1 U11024 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U11025 ( .A1(n9913), .A2(n9920), .B1(n9898), .B2(n9911), .ZN(
        P1_U3480) );
  OAI211_X1 U11026 ( .C1(n5670), .C2(n9906), .A(n9900), .B(n9899), .ZN(n9901)
         );
  AOI21_X1 U11027 ( .B1(n9902), .B2(n9909), .A(n9901), .ZN(n9922) );
  INV_X1 U11028 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U11029 ( .A1(n9913), .A2(n9922), .B1(n9903), .B2(n9911), .ZN(
        P1_U3483) );
  OAI211_X1 U11030 ( .C1(n9907), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9908)
         );
  AOI21_X1 U11031 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9925) );
  INV_X1 U11032 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U11033 ( .A1(n9913), .A2(n9925), .B1(n9912), .B2(n9911), .ZN(
        P1_U3489) );
  AOI22_X1 U11034 ( .A1(n9926), .A2(n9915), .B1(n9914), .B2(n9923), .ZN(
        P1_U3524) );
  AOI22_X1 U11035 ( .A1(n9926), .A2(n9916), .B1(n7005), .B2(n9923), .ZN(
        P1_U3528) );
  AOI22_X1 U11036 ( .A1(n9926), .A2(n9918), .B1(n9917), .B2(n9923), .ZN(
        P1_U3530) );
  AOI22_X1 U11037 ( .A1(n9926), .A2(n9920), .B1(n9919), .B2(n9923), .ZN(
        P1_U3531) );
  AOI22_X1 U11038 ( .A1(n9926), .A2(n9922), .B1(n9921), .B2(n9923), .ZN(
        P1_U3532) );
  AOI22_X1 U11039 ( .A1(n9926), .A2(n9925), .B1(n9924), .B2(n9923), .ZN(
        P1_U3534) );
  INV_X1 U11040 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10077) );
  OAI21_X1 U11041 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  NAND2_X1 U11042 ( .A1(n9994), .A2(n9930), .ZN(n9936) );
  OAI21_X1 U11043 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9934) );
  NAND2_X1 U11044 ( .A1(n9974), .A2(n9934), .ZN(n9935) );
  OAI211_X1 U11045 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7309), .A(n9936), .B(
        n9935), .ZN(n9939) );
  NOR2_X1 U11046 ( .A1(n9983), .A2(n9937), .ZN(n9938) );
  NOR2_X1 U11047 ( .A1(n9939), .A2(n9938), .ZN(n9944) );
  XOR2_X1 U11048 ( .A(n9941), .B(n9940), .Z(n9942) );
  NAND2_X1 U11049 ( .A1(n9942), .A2(n9993), .ZN(n9943) );
  OAI211_X1 U11050 ( .C1(n10077), .C2(n9982), .A(n9944), .B(n9943), .ZN(
        P2_U3184) );
  INV_X1 U11051 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10073) );
  XNOR2_X1 U11052 ( .A(n9945), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9947) );
  AOI21_X1 U11053 ( .B1(n9994), .B2(n9947), .A(n9946), .ZN(n9952) );
  OAI21_X1 U11054 ( .B1(n9949), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9948), .ZN(
        n9950) );
  NAND2_X1 U11055 ( .A1(n9974), .A2(n9950), .ZN(n9951) );
  OAI211_X1 U11056 ( .C1(n9983), .C2(n9953), .A(n9952), .B(n9951), .ZN(n9954)
         );
  INV_X1 U11057 ( .A(n9954), .ZN(n9961) );
  AOI21_X1 U11058 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(n9959) );
  OR2_X1 U11059 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  OAI211_X1 U11060 ( .C1(n10073), .C2(n9982), .A(n9961), .B(n9960), .ZN(
        P2_U3185) );
  INV_X1 U11061 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9962) );
  OAI22_X1 U11062 ( .A1(n9963), .A2(n9983), .B1(n9982), .B2(n9962), .ZN(n9964)
         );
  INV_X1 U11063 ( .A(n9964), .ZN(n9980) );
  OAI21_X1 U11064 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9966), .A(n9965), .ZN(
        n9971) );
  OAI21_X1 U11065 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9970) );
  AOI22_X1 U11066 ( .A1(n9971), .A2(n9994), .B1(n9993), .B2(n9970), .ZN(n9979)
         );
  INV_X1 U11067 ( .A(n9972), .ZN(n9973) );
  NOR2_X1 U11068 ( .A1(n9973), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9976) );
  OAI21_X1 U11069 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9977) );
  NAND4_X1 U11070 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(
        P2_U3195) );
  INV_X1 U11071 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9981) );
  OAI22_X1 U11072 ( .A1(n9984), .A2(n9983), .B1(n9982), .B2(n9981), .ZN(n9985)
         );
  INV_X1 U11073 ( .A(n9985), .ZN(n10003) );
  OAI21_X1 U11074 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9995) );
  OAI21_X1 U11075 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9992) );
  AOI22_X1 U11076 ( .A1(n9995), .A2(n9994), .B1(n9993), .B2(n9992), .ZN(n10002) );
  NAND2_X1 U11077 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10001)
         );
  AOI21_X1 U11078 ( .B1(n4570), .B2(n9997), .A(n9996), .ZN(n9999) );
  OR2_X1 U11079 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND4_X1 U11080 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        P2_U3196) );
  INV_X1 U11081 ( .A(n10004), .ZN(n10015) );
  OAI21_X1 U11082 ( .B1(n10006), .B2(n10015), .A(n10005), .ZN(n10010) );
  INV_X1 U11083 ( .A(n10007), .ZN(n10009) );
  AOI222_X1 U11084 ( .A1(n10023), .A2(n10010), .B1(n10009), .B2(n10019), .C1(
        n10008), .C2(n10017), .ZN(n10011) );
  OAI21_X1 U11085 ( .B1(n10023), .B2(n10012), .A(n10011), .ZN(P2_U3226) );
  OAI21_X1 U11086 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10021) );
  INV_X1 U11087 ( .A(n10016), .ZN(n10020) );
  AOI222_X1 U11088 ( .A1(n10023), .A2(n10021), .B1(n10020), .B2(n10019), .C1(
        n10018), .C2(n10017), .ZN(n10022) );
  OAI21_X1 U11089 ( .B1(n10023), .B2(n6293), .A(n10022), .ZN(P2_U3229) );
  NOR2_X1 U11090 ( .A1(n10024), .A2(n10054), .ZN(n10026) );
  AOI211_X1 U11091 ( .C1(n10040), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10062) );
  AOI22_X1 U11092 ( .A1(n10061), .A2(n6274), .B1(n10062), .B2(n10052), .ZN(
        P2_U3396) );
  INV_X1 U11093 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10032) );
  OAI21_X1 U11094 ( .B1(n10029), .B2(n10054), .A(n10028), .ZN(n10030) );
  AOI21_X1 U11095 ( .B1(n10031), .B2(n10045), .A(n10030), .ZN(n10063) );
  AOI22_X1 U11096 ( .A1(n10061), .A2(n10032), .B1(n10063), .B2(n10052), .ZN(
        P2_U3408) );
  INV_X1 U11097 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10038) );
  OAI22_X1 U11098 ( .A1(n10035), .A2(n10034), .B1(n10033), .B2(n10054), .ZN(
        n10036) );
  NOR2_X1 U11099 ( .A1(n10037), .A2(n10036), .ZN(n10064) );
  AOI22_X1 U11100 ( .A1(n10061), .A2(n10038), .B1(n10064), .B2(n10052), .ZN(
        P2_U3417) );
  INV_X1 U11101 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11102 ( .A1(n10041), .A2(n10040), .B1(n10047), .B2(n10039), .ZN(
        n10042) );
  AND2_X1 U11103 ( .A1(n10043), .A2(n10042), .ZN(n10066) );
  AOI22_X1 U11104 ( .A1(n10061), .A2(n10044), .B1(n10066), .B2(n10052), .ZN(
        P2_U3420) );
  INV_X1 U11105 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U11106 ( .A1(n10046), .A2(n10045), .ZN(n10051) );
  NAND2_X1 U11107 ( .A1(n10048), .A2(n10047), .ZN(n10049) );
  AOI22_X1 U11108 ( .A1(n10061), .A2(n10053), .B1(n10067), .B2(n10052), .ZN(
        P2_U3423) );
  INV_X1 U11109 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10060) );
  OAI22_X1 U11110 ( .A1(n10057), .A2(n10056), .B1(n10055), .B2(n10054), .ZN(
        n10059) );
  NOR2_X1 U11111 ( .A1(n10059), .A2(n10058), .ZN(n10069) );
  AOI22_X1 U11112 ( .A1(n10061), .A2(n10060), .B1(n10069), .B2(n10052), .ZN(
        P2_U3426) );
  AOI22_X1 U11113 ( .A1(n10065), .A2(n10062), .B1(n6275), .B2(n10068), .ZN(
        P2_U3461) );
  AOI22_X1 U11114 ( .A1(n10065), .A2(n10063), .B1(n6317), .B2(n10068), .ZN(
        P2_U3465) );
  AOI22_X1 U11115 ( .A1(n10065), .A2(n10064), .B1(n6346), .B2(n10068), .ZN(
        P2_U3468) );
  AOI22_X1 U11116 ( .A1(n10065), .A2(n10066), .B1(n6359), .B2(n10068), .ZN(
        P2_U3469) );
  AOI22_X1 U11117 ( .A1(n10065), .A2(n10067), .B1(n6370), .B2(n10068), .ZN(
        P2_U3470) );
  AOI22_X1 U11118 ( .A1(n10065), .A2(n10069), .B1(n6380), .B2(n10068), .ZN(
        P2_U3471) );
  AOI21_X1 U11119 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U11120 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10070) );
  NOR2_X1 U11121 ( .A1(n10071), .A2(n10070), .ZN(n10074) );
  NOR2_X1 U11122 ( .A1(n10076), .A2(n10074), .ZN(n10072) );
  XOR2_X1 U11123 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10072), .Z(ADD_1068_U5) );
  XOR2_X1 U11124 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11125 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10123) );
  NOR2_X1 U11126 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10121) );
  NOR2_X1 U11127 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10119) );
  NOR2_X1 U11128 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10117) );
  NOR2_X1 U11129 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10115) );
  NOR2_X1 U11130 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10113) );
  NOR2_X1 U11131 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10109) );
  NOR2_X1 U11132 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10105) );
  NOR2_X1 U11133 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10101) );
  NOR2_X1 U11134 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10097) );
  NOR2_X1 U11135 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10093) );
  NOR2_X1 U11136 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10089) );
  NOR2_X1 U11137 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10086) );
  NOR2_X1 U11138 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10083) );
  NAND2_X1 U11139 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10081) );
  XNOR2_X1 U11140 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n10073), .ZN(n10535) );
  NAND2_X1 U11141 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10079) );
  NOR2_X1 U11142 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10074), .ZN(n10075) );
  NOR2_X1 U11143 ( .A1(n10076), .A2(n10075), .ZN(n10525) );
  XNOR2_X1 U11144 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n10077), .ZN(n10524) );
  NAND2_X1 U11145 ( .A1(n10525), .A2(n10524), .ZN(n10078) );
  NAND2_X1 U11146 ( .A1(n10079), .A2(n10078), .ZN(n10534) );
  NAND2_X1 U11147 ( .A1(n10535), .A2(n10534), .ZN(n10080) );
  NAND2_X1 U11148 ( .A1(n10081), .A2(n10080), .ZN(n10537) );
  XNOR2_X1 U11149 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10536) );
  NOR2_X1 U11150 ( .A1(n10537), .A2(n10536), .ZN(n10082) );
  NOR2_X1 U11151 ( .A1(n10083), .A2(n10082), .ZN(n10527) );
  XOR2_X1 U11152 ( .A(n10084), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10526) );
  NOR2_X1 U11153 ( .A1(n10527), .A2(n10526), .ZN(n10085) );
  NOR2_X1 U11154 ( .A1(n10086), .A2(n10085), .ZN(n10533) );
  XOR2_X1 U11155 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10087), .Z(n10532) );
  NOR2_X1 U11156 ( .A1(n10533), .A2(n10532), .ZN(n10088) );
  NOR2_X1 U11157 ( .A1(n10089), .A2(n10088), .ZN(n10529) );
  INV_X1 U11158 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11159 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10091), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n10090), .ZN(n10528) );
  NOR2_X1 U11160 ( .A1(n10529), .A2(n10528), .ZN(n10092) );
  NOR2_X1 U11161 ( .A1(n10093), .A2(n10092), .ZN(n10531) );
  INV_X1 U11162 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11163 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10095), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10094), .ZN(n10530) );
  NOR2_X1 U11164 ( .A1(n10531), .A2(n10530), .ZN(n10096) );
  NOR2_X1 U11165 ( .A1(n10097), .A2(n10096), .ZN(n10523) );
  INV_X1 U11166 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10099) );
  INV_X1 U11167 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U11168 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10099), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10098), .ZN(n10522) );
  NOR2_X1 U11169 ( .A1(n10523), .A2(n10522), .ZN(n10100) );
  NOR2_X1 U11170 ( .A1(n10101), .A2(n10100), .ZN(n10140) );
  INV_X1 U11171 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10103) );
  INV_X1 U11172 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U11173 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10103), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10102), .ZN(n10139) );
  NOR2_X1 U11174 ( .A1(n10140), .A2(n10139), .ZN(n10104) );
  NOR2_X1 U11175 ( .A1(n10105), .A2(n10104), .ZN(n10138) );
  INV_X1 U11176 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10107) );
  INV_X1 U11177 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11178 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10107), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10106), .ZN(n10137) );
  NOR2_X1 U11179 ( .A1(n10138), .A2(n10137), .ZN(n10108) );
  NOR2_X1 U11180 ( .A1(n10109), .A2(n10108), .ZN(n10136) );
  INV_X1 U11181 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11182 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10111), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10110), .ZN(n10135) );
  NOR2_X1 U11183 ( .A1(n10136), .A2(n10135), .ZN(n10112) );
  NOR2_X1 U11184 ( .A1(n10113), .A2(n10112), .ZN(n10134) );
  XNOR2_X1 U11185 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10133) );
  NOR2_X1 U11186 ( .A1(n10134), .A2(n10133), .ZN(n10114) );
  NOR2_X1 U11187 ( .A1(n10115), .A2(n10114), .ZN(n10132) );
  XNOR2_X1 U11188 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10131) );
  NOR2_X1 U11189 ( .A1(n10132), .A2(n10131), .ZN(n10116) );
  NOR2_X1 U11190 ( .A1(n10117), .A2(n10116), .ZN(n10130) );
  XNOR2_X1 U11191 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10129) );
  NOR2_X1 U11192 ( .A1(n10130), .A2(n10129), .ZN(n10118) );
  NOR2_X1 U11193 ( .A1(n10119), .A2(n10118), .ZN(n10128) );
  XNOR2_X1 U11194 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10127) );
  NOR2_X1 U11195 ( .A1(n10128), .A2(n10127), .ZN(n10120) );
  NOR2_X1 U11196 ( .A1(n10121), .A2(n10120), .ZN(n10126) );
  XNOR2_X1 U11197 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10125) );
  NOR2_X1 U11198 ( .A1(n10126), .A2(n10125), .ZN(n10122) );
  NOR2_X1 U11199 ( .A1(n10123), .A2(n10122), .ZN(n10141) );
  NAND2_X1 U11200 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10141), .ZN(n10142) );
  OAI21_X1 U11201 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10141), .A(n10142), 
        .ZN(n10124) );
  XOR2_X1 U11202 ( .A(n10124), .B(n10144), .Z(ADD_1068_U55) );
  XNOR2_X1 U11203 ( .A(n10126), .B(n10125), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11204 ( .A(n10128), .B(n10127), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11205 ( .A(n10130), .B(n10129), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11206 ( .A(n10132), .B(n10131), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11207 ( .A(n10134), .B(n10133), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11208 ( .A(n10136), .B(n10135), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11209 ( .A(n10138), .B(n10137), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11210 ( .A(n10140), .B(n10139), .ZN(ADD_1068_U63) );
  NOR2_X1 U11211 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10141), .ZN(n10143) );
  OAI21_X1 U11212 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10521) );
  OAI22_X1 U11213 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .ZN(n10145) );
  AOI221_X1 U11214 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        keyinput_g77), .C2(P2_DATAO_REG_19__SCAN_IN), .A(n10145), .ZN(n10152)
         );
  OAI22_X1 U11215 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_g116), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .ZN(n10146) );
  AOI221_X1 U11216 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g83), .C2(P2_DATAO_REG_13__SCAN_IN), .A(n10146), .ZN(n10151)
         );
  OAI22_X1 U11217 ( .A1(SI_21_), .A2(keyinput_g11), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n10147) );
  AOI221_X1 U11218 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g17), .C2(
        SI_15_), .A(n10147), .ZN(n10150) );
  OAI22_X1 U11219 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g104), .B1(
        keyinput_g8), .B2(SI_24_), .ZN(n10148) );
  AOI221_X1 U11220 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_24_), .C2(keyinput_g8), .A(n10148), .ZN(n10149) );
  NAND4_X1 U11221 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10281) );
  OAI22_X1 U11222 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g112), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_g114), .ZN(n10153) );
  AOI221_X1 U11223 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g114), .C2(P1_IR_REG_24__SCAN_IN), .A(n10153), .ZN(n10179) );
  OAI22_X1 U11224 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g40), .B2(P2_REG3_REG_3__SCAN_IN), .ZN(n10154) );
  AOI221_X1 U11225 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n10154), .ZN(n10157) );
  OAI22_X1 U11226 ( .A1(SI_27_), .A2(keyinput_g5), .B1(SI_30_), .B2(
        keyinput_g2), .ZN(n10155) );
  AOI221_X1 U11227 ( .B1(SI_27_), .B2(keyinput_g5), .C1(keyinput_g2), .C2(
        SI_30_), .A(n10155), .ZN(n10156) );
  OAI211_X1 U11228 ( .C1(n10159), .C2(keyinput_g52), .A(n10157), .B(n10156), 
        .ZN(n10158) );
  AOI21_X1 U11229 ( .B1(n10159), .B2(keyinput_g52), .A(n10158), .ZN(n10178) );
  AOI22_X1 U11230 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(SI_2_), .B2(
        keyinput_g30), .ZN(n10160) );
  OAI221_X1 U11231 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(SI_2_), 
        .C2(keyinput_g30), .A(n10160), .ZN(n10167) );
  AOI22_X1 U11232 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(SI_3_), .B2(keyinput_g29), .ZN(n10161) );
  OAI221_X1 U11233 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        SI_3_), .C2(keyinput_g29), .A(n10161), .ZN(n10166) );
  AOI22_X1 U11234 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_g119), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_g90), .ZN(n10162) );
  OAI221_X1 U11235 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_g119), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_g90), .A(n10162), .ZN(n10165) );
  AOI22_X1 U11236 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10163) );
  OAI221_X1 U11237 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n10163), .ZN(n10164)
         );
  NOR4_X1 U11238 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10177) );
  AOI22_X1 U11239 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput_g127), .ZN(n10168) );
  OAI221_X1 U11240 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput_g127), .A(n10168), .ZN(n10175) );
  AOI22_X1 U11241 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        SI_26_), .B2(keyinput_g6), .ZN(n10169) );
  OAI221_X1 U11242 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        SI_26_), .C2(keyinput_g6), .A(n10169), .ZN(n10174) );
  AOI22_X1 U11243 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .ZN(n10170) );
  OAI221_X1 U11244 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g94), .A(n10170), .ZN(n10173) );
  AOI22_X1 U11245 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_g123), .ZN(n10171) );
  OAI221_X1 U11246 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_g123), .A(n10171), .ZN(n10172) );
  NOR4_X1 U11247 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10176) );
  NAND4_X1 U11248 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10280) );
  AOI22_X1 U11249 ( .A1(n10414), .A2(keyinput_g72), .B1(keyinput_g58), .B2(
        n10438), .ZN(n10180) );
  OAI221_X1 U11250 ( .B1(n10414), .B2(keyinput_g72), .C1(n10438), .C2(
        keyinput_g58), .A(n10180), .ZN(n10189) );
  AOI22_X1 U11251 ( .A1(n10482), .A2(keyinput_g76), .B1(n10182), .B2(
        keyinput_g69), .ZN(n10181) );
  OAI221_X1 U11252 ( .B1(n10482), .B2(keyinput_g76), .C1(n10182), .C2(
        keyinput_g69), .A(n10181), .ZN(n10188) );
  AOI22_X1 U11253 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_g95), .ZN(n10183) );
  OAI221_X1 U11254 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_g95), .A(n10183), .ZN(n10187) );
  XOR2_X1 U11255 ( .A(n7309), .B(keyinput_g59), .Z(n10185) );
  XNOR2_X1 U11256 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g111), .ZN(n10184)
         );
  NAND2_X1 U11257 ( .A1(n10185), .A2(n10184), .ZN(n10186) );
  NOR4_X1 U11258 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10227) );
  INV_X1 U11259 ( .A(SI_16_), .ZN(n10421) );
  AOI22_X1 U11260 ( .A1(n10469), .A2(keyinput_g74), .B1(keyinput_g16), .B2(
        n10421), .ZN(n10190) );
  OAI221_X1 U11261 ( .B1(n10469), .B2(keyinput_g74), .C1(n10421), .C2(
        keyinput_g16), .A(n10190), .ZN(n10199) );
  AOI22_X1 U11262 ( .A1(n10192), .A2(keyinput_g65), .B1(n10408), .B2(
        keyinput_g106), .ZN(n10191) );
  OAI221_X1 U11263 ( .B1(n10192), .B2(keyinput_g65), .C1(n10408), .C2(
        keyinput_g106), .A(n10191), .ZN(n10198) );
  XOR2_X1 U11264 ( .A(n5368), .B(keyinput_g73), .Z(n10196) );
  XNOR2_X1 U11265 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n10195) );
  XNOR2_X1 U11266 ( .A(SI_6_), .B(keyinput_g26), .ZN(n10194) );
  XNOR2_X1 U11267 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g101), .ZN(n10193)
         );
  NAND4_X1 U11268 ( .A1(n10196), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10197) );
  NOR3_X1 U11269 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10226) );
  INV_X1 U11270 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U11271 ( .A1(n10484), .A2(keyinput_g42), .B1(keyinput_g43), .B2(
        n10201), .ZN(n10200) );
  OAI221_X1 U11272 ( .B1(n10484), .B2(keyinput_g42), .C1(n10201), .C2(
        keyinput_g43), .A(n10200), .ZN(n10212) );
  INV_X1 U11273 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11274 ( .A1(n10204), .A2(keyinput_g41), .B1(n10203), .B2(
        keyinput_g38), .ZN(n10202) );
  OAI221_X1 U11275 ( .B1(n10204), .B2(keyinput_g41), .C1(n10203), .C2(
        keyinput_g38), .A(n10202), .ZN(n10211) );
  AOI22_X1 U11276 ( .A1(n10206), .A2(keyinput_g82), .B1(keyinput_g46), .B2(
        n10460), .ZN(n10205) );
  OAI221_X1 U11277 ( .B1(n10206), .B2(keyinput_g82), .C1(n10460), .C2(
        keyinput_g46), .A(n10205), .ZN(n10210) );
  XNOR2_X1 U11278 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g92), .ZN(n10208) );
  XNOR2_X1 U11279 ( .A(SI_5_), .B(keyinput_g27), .ZN(n10207) );
  NAND2_X1 U11280 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  NOR4_X1 U11281 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10225) );
  AOI22_X1 U11282 ( .A1(n10428), .A2(keyinput_g124), .B1(keyinput_g78), .B2(
        n10214), .ZN(n10213) );
  OAI221_X1 U11283 ( .B1(n10428), .B2(keyinput_g124), .C1(n10214), .C2(
        keyinput_g78), .A(n10213), .ZN(n10223) );
  INV_X1 U11284 ( .A(SI_13_), .ZN(n10479) );
  AOI22_X1 U11285 ( .A1(n10479), .A2(keyinput_g19), .B1(n10318), .B2(
        keyinput_g107), .ZN(n10215) );
  OAI221_X1 U11286 ( .B1(n10479), .B2(keyinput_g19), .C1(n10318), .C2(
        keyinput_g107), .A(n10215), .ZN(n10222) );
  AOI22_X1 U11287 ( .A1(n10409), .A2(keyinput_g70), .B1(keyinput_g25), .B2(
        n10217), .ZN(n10216) );
  OAI221_X1 U11288 ( .B1(n10409), .B2(keyinput_g70), .C1(n10217), .C2(
        keyinput_g25), .A(n10216), .ZN(n10221) );
  XNOR2_X1 U11289 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g117), .ZN(n10219)
         );
  XNOR2_X1 U11290 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n10218) );
  NAND2_X1 U11291 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  NOR4_X1 U11292 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10224) );
  NAND4_X1 U11293 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10279) );
  AOI22_X1 U11294 ( .A1(n5326), .A2(keyinput_g87), .B1(keyinput_g1), .B2(
        n10229), .ZN(n10228) );
  OAI221_X1 U11295 ( .B1(n5326), .B2(keyinput_g87), .C1(n10229), .C2(
        keyinput_g1), .A(n10228), .ZN(n10239) );
  XNOR2_X1 U11296 ( .A(n10230), .B(keyinput_g100), .ZN(n10238) );
  XNOR2_X1 U11297 ( .A(n10231), .B(keyinput_g47), .ZN(n10237) );
  XNOR2_X1 U11298 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g110), .ZN(n10235)
         );
  XNOR2_X1 U11299 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g105), .ZN(n10234)
         );
  XNOR2_X1 U11300 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g91), .ZN(n10233) );
  XNOR2_X1 U11301 ( .A(SI_14_), .B(keyinput_g18), .ZN(n10232) );
  NAND4_X1 U11302 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10236) );
  NOR4_X1 U11303 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10277) );
  AOI22_X1 U11304 ( .A1(n10457), .A2(keyinput_g35), .B1(n10241), .B2(
        keyinput_g10), .ZN(n10240) );
  OAI221_X1 U11305 ( .B1(n10457), .B2(keyinput_g35), .C1(n10241), .C2(
        keyinput_g10), .A(n10240), .ZN(n10251) );
  INV_X1 U11306 ( .A(SI_12_), .ZN(n10243) );
  AOI22_X1 U11307 ( .A1(n10243), .A2(keyinput_g20), .B1(keyinput_g23), .B2(
        n10454), .ZN(n10242) );
  OAI221_X1 U11308 ( .B1(n10243), .B2(keyinput_g20), .C1(n10454), .C2(
        keyinput_g23), .A(n10242), .ZN(n10250) );
  AOI22_X1 U11309 ( .A1(n10245), .A2(keyinput_g24), .B1(n10494), .B2(
        keyinput_g71), .ZN(n10244) );
  OAI221_X1 U11310 ( .B1(n10245), .B2(keyinput_g24), .C1(n10494), .C2(
        keyinput_g71), .A(n10244), .ZN(n10249) );
  XNOR2_X1 U11311 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g120), .ZN(n10247)
         );
  XNOR2_X1 U11312 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n10246)
         );
  NAND2_X1 U11313 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  NOR4_X1 U11314 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10276) );
  AOI22_X1 U11315 ( .A1(n6215), .A2(keyinput_g53), .B1(keyinput_g61), .B2(
        n10453), .ZN(n10252) );
  OAI221_X1 U11316 ( .B1(n6215), .B2(keyinput_g53), .C1(n10453), .C2(
        keyinput_g61), .A(n10252), .ZN(n10261) );
  AOI22_X1 U11317 ( .A1(n10382), .A2(keyinput_g98), .B1(keyinput_g51), .B2(
        n10254), .ZN(n10253) );
  OAI221_X1 U11318 ( .B1(n10382), .B2(keyinput_g98), .C1(n10254), .C2(
        keyinput_g51), .A(n10253), .ZN(n10260) );
  XNOR2_X1 U11319 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_g80), .ZN(n10258) );
  XNOR2_X1 U11320 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n10257)
         );
  XNOR2_X1 U11321 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g93), .ZN(n10256) );
  XNOR2_X1 U11322 ( .A(SI_4_), .B(keyinput_g28), .ZN(n10255) );
  NAND4_X1 U11323 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10259) );
  NOR3_X1 U11324 ( .A1(n10261), .A2(n10260), .A3(n10259), .ZN(n10275) );
  AOI22_X1 U11325 ( .A1(n10456), .A2(keyinput_g68), .B1(n10263), .B2(
        keyinput_g21), .ZN(n10262) );
  OAI221_X1 U11326 ( .B1(n10456), .B2(keyinput_g68), .C1(n10263), .C2(
        keyinput_g21), .A(n10262), .ZN(n10273) );
  INV_X1 U11327 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U11328 ( .A1(n10440), .A2(keyinput_g99), .B1(keyinput_g9), .B2(
        n10265), .ZN(n10264) );
  OAI221_X1 U11329 ( .B1(n10440), .B2(keyinput_g99), .C1(n10265), .C2(
        keyinput_g9), .A(n10264), .ZN(n10272) );
  INV_X1 U11330 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10267) );
  INV_X1 U11331 ( .A(SI_18_), .ZN(n10424) );
  AOI22_X1 U11332 ( .A1(n10267), .A2(keyinput_g57), .B1(n10424), .B2(
        keyinput_g14), .ZN(n10266) );
  OAI221_X1 U11333 ( .B1(n10267), .B2(keyinput_g57), .C1(n10424), .C2(
        keyinput_g14), .A(n10266), .ZN(n10271) );
  XOR2_X1 U11334 ( .A(n10435), .B(keyinput_g49), .Z(n10269) );
  XNOR2_X1 U11335 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g96), .ZN(n10268) );
  NAND2_X1 U11336 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  NOR4_X1 U11337 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10274) );
  NAND4_X1 U11338 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NOR4_X1 U11339 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10517) );
  OAI22_X1 U11340 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g86), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10282) );
  AOI221_X1 U11341 ( .B1(SI_25_), .B2(keyinput_g7), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n10282), .ZN(n10289)
         );
  OAI22_X1 U11342 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_g108), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .ZN(n10283) );
  AOI221_X1 U11343 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_g108), .C1(
        keyinput_g44), .C2(P2_REG3_REG_1__SCAN_IN), .A(n10283), .ZN(n10288) );
  OAI22_X1 U11344 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10284) );
  AOI221_X1 U11345 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        keyinput_g48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n10284), .ZN(n10287)
         );
  OAI22_X1 U11346 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_g125), .B1(
        keyinput_g67), .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10285) );
  AOI221_X1 U11347 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_g125), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_g67), .A(n10285), .ZN(n10286)
         );
  NAND4_X1 U11348 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10317) );
  OAI22_X1 U11349 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g113), .B1(SI_1_), 
        .B2(keyinput_g31), .ZN(n10290) );
  AOI221_X1 U11350 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g31), .C2(SI_1_), .A(n10290), .ZN(n10297) );
  OAI22_X1 U11351 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g102), .B1(
        keyinput_g32), .B2(SI_0_), .ZN(n10291) );
  AOI221_X1 U11352 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g102), .C1(SI_0_), .C2(keyinput_g32), .A(n10291), .ZN(n10296) );
  OAI22_X1 U11353 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_g121), .B1(
        keyinput_g79), .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n10292) );
  AOI221_X1 U11354 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_g121), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n10292), .ZN(n10295)
         );
  OAI22_X1 U11355 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g45), .B2(P2_REG3_REG_21__SCAN_IN), .ZN(n10293) );
  AOI221_X1 U11356 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n10293), .ZN(n10294)
         );
  NAND4_X1 U11357 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10316) );
  OAI22_X1 U11358 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g126), .B1(SI_28_), 
        .B2(keyinput_g4), .ZN(n10298) );
  AOI221_X1 U11359 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g4), .C2(SI_28_), .A(n10298), .ZN(n10305) );
  OAI22_X1 U11360 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_g122), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput_g118), .ZN(n10299) );
  AOI221_X1 U11361 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g118), .C2(P1_IR_REG_28__SCAN_IN), .A(n10299), .ZN(n10304) );
  OAI22_X1 U11362 ( .A1(SI_29_), .A2(keyinput_g3), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .ZN(n10300) );
  AOI221_X1 U11363 ( .B1(SI_29_), .B2(keyinput_g3), .C1(keyinput_g66), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n10300), .ZN(n10303) );
  OAI22_X1 U11364 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g37), .B2(
        P2_REG3_REG_14__SCAN_IN), .ZN(n10301) );
  AOI221_X1 U11365 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10301), .ZN(n10302)
         );
  NAND4_X1 U11366 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10315) );
  OAI22_X1 U11367 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g109), .B1(
        keyinput_g103), .B2(P1_IR_REG_13__SCAN_IN), .ZN(n10306) );
  AOI221_X1 U11368 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g109), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g103), .A(n10306), .ZN(n10313) );
  OAI22_X1 U11369 ( .A1(SI_17_), .A2(keyinput_g15), .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n10307) );
  AOI221_X1 U11370 ( .B1(SI_17_), .B2(keyinput_g15), .C1(keyinput_g54), .C2(
        P2_REG3_REG_0__SCAN_IN), .A(n10307), .ZN(n10312) );
  OAI22_X1 U11371 ( .A1(SI_20_), .A2(keyinput_g12), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n10308) );
  AOI221_X1 U11372 ( .B1(SI_20_), .B2(keyinput_g12), .C1(keyinput_g88), .C2(
        P2_DATAO_REG_8__SCAN_IN), .A(n10308), .ZN(n10311) );
  OAI22_X1 U11373 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n10309) );
  AOI221_X1 U11374 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g63), .C2(P2_REG3_REG_15__SCAN_IN), .A(n10309), .ZN(n10310)
         );
  NAND4_X1 U11375 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10314) );
  NOR4_X1 U11376 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10516) );
  XNOR2_X1 U11377 ( .A(n10318), .B(keyinput_f107), .ZN(n10325) );
  AOI22_X1 U11378 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .ZN(n10319) );
  OAI221_X1 U11379 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_f114), .A(n10319), .ZN(n10324) );
  AOI22_X1 U11380 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P1_IR_REG_18__SCAN_IN), 
        .B2(keyinput_f108), .ZN(n10320) );
  OAI221_X1 U11381 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P1_IR_REG_18__SCAN_IN), 
        .C2(keyinput_f108), .A(n10320), .ZN(n10323) );
  AOI22_X1 U11382 ( .A1(SI_8_), .A2(keyinput_f24), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .ZN(n10321) );
  OAI221_X1 U11383 ( .B1(SI_8_), .B2(keyinput_f24), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_f82), .A(n10321), .ZN(n10322)
         );
  NOR4_X1 U11384 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10353) );
  AOI22_X1 U11385 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_f104), .ZN(n10326) );
  OAI221_X1 U11386 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_f104), .A(n10326), .ZN(n10333) );
  AOI22_X1 U11387 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_f94), .ZN(n10327) );
  OAI221_X1 U11388 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f94), .A(n10327), .ZN(n10332) );
  AOI22_X1 U11389 ( .A1(SI_11_), .A2(keyinput_f21), .B1(P1_IR_REG_26__SCAN_IN), 
        .B2(keyinput_f116), .ZN(n10328) );
  OAI221_X1 U11390 ( .B1(SI_11_), .B2(keyinput_f21), .C1(P1_IR_REG_26__SCAN_IN), .C2(keyinput_f116), .A(n10328), .ZN(n10331) );
  AOI22_X1 U11391 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n10329) );
  OAI221_X1 U11392 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n10329), .ZN(n10330)
         );
  NOR4_X1 U11393 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10352) );
  AOI22_X1 U11394 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_f69), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .ZN(n10334) );
  OAI221_X1 U11395 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_f103), .A(n10334), .ZN(n10341) );
  AOI22_X1 U11396 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .ZN(n10335) );
  OAI221_X1 U11397 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_f117), .A(n10335), .ZN(n10340) );
  AOI22_X1 U11398 ( .A1(SI_31_), .A2(keyinput_f1), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10336) );
  OAI221_X1 U11399 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10336), .ZN(n10339)
         );
  AOI22_X1 U11400 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10337) );
  OAI221_X1 U11401 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10337), .ZN(n10338) );
  NOR4_X1 U11402 ( .A1(n10341), .A2(n10340), .A3(n10339), .A4(n10338), .ZN(
        n10351) );
  AOI22_X1 U11403 ( .A1(SI_4_), .A2(keyinput_f28), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n10342) );
  OAI221_X1 U11404 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_25_), .C2(
        keyinput_f7), .A(n10342), .ZN(n10349) );
  AOI22_X1 U11405 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .ZN(n10343) );
  OAI221_X1 U11406 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f102), .A(n10343), .ZN(n10348) );
  AOI22_X1 U11407 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n10344) );
  OAI221_X1 U11408 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10344), .ZN(n10347)
         );
  AOI22_X1 U11409 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput_f119), .ZN(n10345) );
  OAI221_X1 U11410 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput_f119), .A(n10345), .ZN(n10346) );
  NOR4_X1 U11411 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NAND4_X1 U11412 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10510) );
  AOI22_X1 U11413 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .ZN(n10354) );
  OAI221_X1 U11414 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f101), .A(n10354), .ZN(n10361) );
  AOI22_X1 U11415 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n10355) );
  OAI221_X1 U11416 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n10355), .ZN(n10360)
         );
  AOI22_X1 U11417 ( .A1(SI_1_), .A2(keyinput_f31), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_f109), .ZN(n10356) );
  OAI221_X1 U11418 ( .B1(SI_1_), .B2(keyinput_f31), .C1(P1_IR_REG_19__SCAN_IN), 
        .C2(keyinput_f109), .A(n10356), .ZN(n10359) );
  AOI22_X1 U11419 ( .A1(SI_5_), .A2(keyinput_f27), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n10357) );
  OAI221_X1 U11420 ( .B1(SI_5_), .B2(keyinput_f27), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n10357), .ZN(n10358)
         );
  NOR4_X1 U11421 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10390) );
  AOI22_X1 U11422 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n10362) );
  OAI221_X1 U11423 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n10362), .ZN(n10369) );
  AOI22_X1 U11424 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10363) );
  OAI221_X1 U11425 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10363), .ZN(n10368)
         );
  AOI22_X1 U11426 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        SI_26_), .B2(keyinput_f6), .ZN(n10364) );
  OAI221_X1 U11427 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        SI_26_), .C2(keyinput_f6), .A(n10364), .ZN(n10367) );
  AOI22_X1 U11428 ( .A1(SI_14_), .A2(keyinput_f18), .B1(SI_19_), .B2(
        keyinput_f13), .ZN(n10365) );
  OAI221_X1 U11429 ( .B1(SI_14_), .B2(keyinput_f18), .C1(SI_19_), .C2(
        keyinput_f13), .A(n10365), .ZN(n10366) );
  NOR4_X1 U11430 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10389) );
  AOI22_X1 U11431 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_f122), .ZN(n10370) );
  OAI221_X1 U11432 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f122), .A(n10370), .ZN(n10377) );
  AOI22_X1 U11433 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput_f127), .ZN(n10371) );
  OAI221_X1 U11434 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput_f127), .A(n10371), .ZN(n10376) );
  AOI22_X1 U11435 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_f115), .ZN(n10372) );
  OAI221_X1 U11436 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput_f115), .A(n10372), .ZN(n10375) );
  AOI22_X1 U11437 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P1_IR_REG_5__SCAN_IN), 
        .B2(keyinput_f95), .ZN(n10373) );
  OAI221_X1 U11438 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P1_IR_REG_5__SCAN_IN), 
        .C2(keyinput_f95), .A(n10373), .ZN(n10374) );
  NOR4_X1 U11439 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10388) );
  AOI22_X1 U11440 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_f93), .ZN(n10378) );
  OAI221_X1 U11441 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_f93), .A(n10378), .ZN(n10386) );
  AOI22_X1 U11442 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10379) );
  OAI221_X1 U11443 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n10379), .ZN(n10385)
         );
  AOI22_X1 U11444 ( .A1(SI_15_), .A2(keyinput_f17), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_f126), .ZN(n10380) );
  OAI221_X1 U11445 ( .B1(SI_15_), .B2(keyinput_f17), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_f126), .A(n10380), .ZN(n10384) );
  AOI22_X1 U11446 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        n10382), .B2(keyinput_f98), .ZN(n10381) );
  OAI221_X1 U11447 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        n10382), .C2(keyinput_f98), .A(n10381), .ZN(n10383) );
  NOR4_X1 U11448 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  NAND4_X1 U11449 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10509) );
  AOI22_X1 U11450 ( .A1(n10392), .A2(keyinput_f125), .B1(keyinput_f4), .B2(
        n5393), .ZN(n10391) );
  OAI221_X1 U11451 ( .B1(n10392), .B2(keyinput_f125), .C1(n5393), .C2(
        keyinput_f4), .A(n10391), .ZN(n10403) );
  INV_X1 U11452 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U11453 ( .A1(n5368), .A2(keyinput_f73), .B1(keyinput_f55), .B2(
        n10394), .ZN(n10393) );
  OAI221_X1 U11454 ( .B1(n5368), .B2(keyinput_f73), .C1(n10394), .C2(
        keyinput_f55), .A(n10393), .ZN(n10402) );
  AOI22_X1 U11455 ( .A1(n10397), .A2(keyinput_f8), .B1(keyinput_f81), .B2(
        n10396), .ZN(n10395) );
  OAI221_X1 U11456 ( .B1(n10397), .B2(keyinput_f8), .C1(n10396), .C2(
        keyinput_f81), .A(n10395), .ZN(n10401) );
  XNOR2_X1 U11457 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .ZN(n10399)
         );
  XNOR2_X1 U11458 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f92), .ZN(n10398) );
  NAND2_X1 U11459 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  NOR4_X1 U11460 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10451) );
  INV_X1 U11461 ( .A(SI_21_), .ZN(n10405) );
  AOI22_X1 U11462 ( .A1(n10406), .A2(keyinput_f5), .B1(keyinput_f11), .B2(
        n10405), .ZN(n10404) );
  OAI221_X1 U11463 ( .B1(n10406), .B2(keyinput_f5), .C1(n10405), .C2(
        keyinput_f11), .A(n10404), .ZN(n10419) );
  AOI22_X1 U11464 ( .A1(n10409), .A2(keyinput_f70), .B1(n10408), .B2(
        keyinput_f106), .ZN(n10407) );
  OAI221_X1 U11465 ( .B1(n10409), .B2(keyinput_f70), .C1(n10408), .C2(
        keyinput_f106), .A(n10407), .ZN(n10418) );
  AOI22_X1 U11466 ( .A1(n10412), .A2(keyinput_f89), .B1(n10411), .B2(
        keyinput_f15), .ZN(n10410) );
  OAI221_X1 U11467 ( .B1(n10412), .B2(keyinput_f89), .C1(n10411), .C2(
        keyinput_f15), .A(n10410), .ZN(n10417) );
  AOI22_X1 U11468 ( .A1(n10415), .A2(keyinput_f77), .B1(n10414), .B2(
        keyinput_f72), .ZN(n10413) );
  OAI221_X1 U11469 ( .B1(n10415), .B2(keyinput_f77), .C1(n10414), .C2(
        keyinput_f72), .A(n10413), .ZN(n10416) );
  NOR4_X1 U11470 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10450) );
  AOI22_X1 U11471 ( .A1(n10422), .A2(keyinput_f79), .B1(keyinput_f16), .B2(
        n10421), .ZN(n10420) );
  OAI221_X1 U11472 ( .B1(n10422), .B2(keyinput_f79), .C1(n10421), .C2(
        keyinput_f16), .A(n10420), .ZN(n10432) );
  AOI22_X1 U11473 ( .A1(n7319), .A2(keyinput_f44), .B1(n10424), .B2(
        keyinput_f14), .ZN(n10423) );
  OAI221_X1 U11474 ( .B1(n7319), .B2(keyinput_f44), .C1(n10424), .C2(
        keyinput_f14), .A(n10423), .ZN(n10431) );
  XNOR2_X1 U11475 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10427) );
  XNOR2_X1 U11476 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f100), .ZN(n10426)
         );
  XNOR2_X1 U11477 ( .A(SI_23_), .B(keyinput_f9), .ZN(n10425) );
  NAND3_X1 U11478 ( .A1(n10427), .A2(n10426), .A3(n10425), .ZN(n10430) );
  XNOR2_X1 U11479 ( .A(n10428), .B(keyinput_f124), .ZN(n10429) );
  NOR4_X1 U11480 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .ZN(
        n10449) );
  AOI22_X1 U11481 ( .A1(n10435), .A2(keyinput_f49), .B1(n10434), .B2(
        keyinput_f26), .ZN(n10433) );
  OAI221_X1 U11482 ( .B1(n10435), .B2(keyinput_f49), .C1(n10434), .C2(
        keyinput_f26), .A(n10433), .ZN(n10447) );
  AOI22_X1 U11483 ( .A1(n10438), .A2(keyinput_f58), .B1(n10437), .B2(
        keyinput_f85), .ZN(n10436) );
  OAI221_X1 U11484 ( .B1(n10438), .B2(keyinput_f58), .C1(n10437), .C2(
        keyinput_f85), .A(n10436), .ZN(n10446) );
  AOI22_X1 U11485 ( .A1(n10441), .A2(keyinput_f3), .B1(n10440), .B2(
        keyinput_f99), .ZN(n10439) );
  OAI221_X1 U11486 ( .B1(n10441), .B2(keyinput_f3), .C1(n10440), .C2(
        keyinput_f99), .A(n10439), .ZN(n10445) );
  XNOR2_X1 U11487 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_f113), .ZN(n10443)
         );
  XNOR2_X1 U11488 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f105), .ZN(n10442)
         );
  NAND2_X1 U11489 ( .A1(n10443), .A2(n10442), .ZN(n10444) );
  NOR4_X1 U11490 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  NAND4_X1 U11491 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10508) );
  AOI22_X1 U11492 ( .A1(n10454), .A2(keyinput_f23), .B1(keyinput_f61), .B2(
        n10453), .ZN(n10452) );
  OAI221_X1 U11493 ( .B1(n10454), .B2(keyinput_f23), .C1(n10453), .C2(
        keyinput_f61), .A(n10452), .ZN(n10466) );
  AOI22_X1 U11494 ( .A1(n10457), .A2(keyinput_f35), .B1(n10456), .B2(
        keyinput_f68), .ZN(n10455) );
  OAI221_X1 U11495 ( .B1(n10457), .B2(keyinput_f35), .C1(n10456), .C2(
        keyinput_f68), .A(n10455), .ZN(n10465) );
  AOI22_X1 U11496 ( .A1(n10460), .A2(keyinput_f46), .B1(n10459), .B2(
        keyinput_f63), .ZN(n10458) );
  OAI221_X1 U11497 ( .B1(n10460), .B2(keyinput_f46), .C1(n10459), .C2(
        keyinput_f63), .A(n10458), .ZN(n10464) );
  XNOR2_X1 U11498 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f97), .ZN(n10462) );
  XNOR2_X1 U11499 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_f86), .ZN(n10461) );
  NAND2_X1 U11500 ( .A1(n10462), .A2(n10461), .ZN(n10463) );
  NOR4_X1 U11501 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10506) );
  AOI22_X1 U11502 ( .A1(n4788), .A2(keyinput_f33), .B1(keyinput_f59), .B2(
        n7309), .ZN(n10467) );
  OAI221_X1 U11503 ( .B1(n4788), .B2(keyinput_f33), .C1(n7309), .C2(
        keyinput_f59), .A(n10467), .ZN(n10477) );
  AOI22_X1 U11504 ( .A1(n10470), .A2(keyinput_f48), .B1(n10469), .B2(
        keyinput_f74), .ZN(n10468) );
  OAI221_X1 U11505 ( .B1(n10470), .B2(keyinput_f48), .C1(n10469), .C2(
        keyinput_f74), .A(n10468), .ZN(n10476) );
  XNOR2_X1 U11506 ( .A(SI_22_), .B(keyinput_f10), .ZN(n10474) );
  XNOR2_X1 U11507 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f96), .ZN(n10473) );
  XNOR2_X1 U11508 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f110), .ZN(n10472)
         );
  XNOR2_X1 U11509 ( .A(SI_12_), .B(keyinput_f20), .ZN(n10471) );
  NAND4_X1 U11510 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  NOR3_X1 U11511 ( .A1(n10477), .A2(n10476), .A3(n10475), .ZN(n10505) );
  AOI22_X1 U11512 ( .A1(n10480), .A2(keyinput_f37), .B1(n10479), .B2(
        keyinput_f19), .ZN(n10478) );
  OAI221_X1 U11513 ( .B1(n10480), .B2(keyinput_f37), .C1(n10479), .C2(
        keyinput_f19), .A(n10478), .ZN(n10492) );
  AOI22_X1 U11514 ( .A1(n10483), .A2(keyinput_f12), .B1(keyinput_f76), .B2(
        n10482), .ZN(n10481) );
  OAI221_X1 U11515 ( .B1(n10483), .B2(keyinput_f12), .C1(n10482), .C2(
        keyinput_f76), .A(n10481), .ZN(n10491) );
  XOR2_X1 U11516 ( .A(n10484), .B(keyinput_f42), .Z(n10489) );
  INV_X1 U11517 ( .A(SI_0_), .ZN(n10485) );
  XOR2_X1 U11518 ( .A(n10485), .B(keyinput_f32), .Z(n10488) );
  XNOR2_X1 U11519 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10487) );
  XNOR2_X1 U11520 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f90), .ZN(n10486) );
  NAND4_X1 U11521 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10490) );
  NOR3_X1 U11522 ( .A1(n10492), .A2(n10491), .A3(n10490), .ZN(n10504) );
  AOI22_X1 U11523 ( .A1(P2_U3151), .A2(keyinput_f34), .B1(n10494), .B2(
        keyinput_f71), .ZN(n10493) );
  OAI221_X1 U11524 ( .B1(P2_U3151), .B2(keyinput_f34), .C1(n10494), .C2(
        keyinput_f71), .A(n10493), .ZN(n10502) );
  XOR2_X1 U11525 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f91), .Z(n10501) );
  XNOR2_X1 U11526 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_f112), .ZN(n10498)
         );
  XNOR2_X1 U11527 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_f57), .ZN(n10497)
         );
  XNOR2_X1 U11528 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_f50), .ZN(n10496)
         );
  XNOR2_X1 U11529 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_f111), .ZN(n10495)
         );
  NAND4_X1 U11530 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10500) );
  XNOR2_X1 U11531 ( .A(keyinput_f56), .B(n6218), .ZN(n10499) );
  NOR4_X1 U11532 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  NAND4_X1 U11533 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10507) );
  OR4_X1 U11534 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10512) );
  AOI21_X1 U11535 ( .B1(keyinput_f22), .B2(n10512), .A(SI_10_), .ZN(n10514) );
  INV_X1 U11536 ( .A(keyinput_f22), .ZN(n10511) );
  AOI21_X1 U11537 ( .B1(n10512), .B2(n10511), .A(keyinput_g22), .ZN(n10513) );
  AOI22_X1 U11538 ( .A1(keyinput_g22), .A2(n10514), .B1(SI_10_), .B2(n10513), 
        .ZN(n10515) );
  AOI21_X1 U11539 ( .B1(n10517), .B2(n10516), .A(n10515), .ZN(n10519) );
  XNOR2_X1 U11540 ( .A(n4711), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10518) );
  XNOR2_X1 U11541 ( .A(n10519), .B(n10518), .ZN(n10520) );
  XNOR2_X1 U11542 ( .A(n10521), .B(n10520), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11543 ( .A(n10523), .B(n10522), .ZN(ADD_1068_U47) );
  XOR2_X1 U11544 ( .A(n10525), .B(n10524), .Z(ADD_1068_U54) );
  XNOR2_X1 U11545 ( .A(n10527), .B(n10526), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11546 ( .A(n10529), .B(n10528), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11547 ( .A(n10531), .B(n10530), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11548 ( .A(n10533), .B(n10532), .ZN(ADD_1068_U50) );
  XOR2_X1 U11549 ( .A(n10535), .B(n10534), .Z(ADD_1068_U53) );
  XNOR2_X1 U11550 ( .A(n10537), .B(n10536), .ZN(ADD_1068_U52) );
  AOI22_X1 U6462 ( .A1(n9626), .A2(n5791), .B1(n9613), .B2(n9756), .ZN(n9609)
         );
endmodule

