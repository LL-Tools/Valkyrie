

module b22_C_AntiSAT_k_128_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15250, n15253;

  INV_X4 U7228 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  XNOR2_X1 U7229 ( .A(n14093), .B(n11776), .ZN(n14085) );
  NAND2_X1 U7230 ( .A1(n8158), .A2(n8157), .ZN(n13532) );
  AND2_X2 U7231 ( .A1(n12325), .A2(n12324), .ZN(n12758) );
  XNOR2_X1 U7232 ( .A(n8901), .B(n8508), .ZN(n11564) );
  INV_X2 U7233 ( .A(n14246), .ZN(n14340) );
  INV_X1 U7234 ( .A(n12153), .ZN(n12194) );
  INV_X2 U7236 ( .A(n13798), .ZN(n13752) );
  CLKBUF_X1 U7237 ( .A(n12026), .Z(n11998) );
  BUF_X1 U7238 ( .A(n8143), .Z(n6486) );
  OR2_X1 U7239 ( .A1(n8928), .A2(n8542), .ZN(n8547) );
  NAND2_X1 U7240 ( .A1(n7668), .A2(n10922), .ZN(n10183) );
  XNOR2_X1 U7241 ( .A(n8514), .B(n8513), .ZN(n13050) );
  CLKBUF_X2 U7242 ( .A(n11152), .Z(n6491) );
  INV_X2 U7243 ( .A(n6686), .ZN(n12025) );
  INV_X2 U7244 ( .A(n7529), .ZN(n12006) );
  CLKBUF_X2 U7245 ( .A(n12023), .Z(n12013) );
  AND2_X1 U7246 ( .A1(n7425), .A2(n7424), .ZN(n7613) );
  NOR2_X2 U7247 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7712) );
  NOR2_X1 U7248 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9048) );
  CLKBUF_X1 U7249 ( .A(n15250), .Z(P1_U4016) );
  NOR2_X1 U7250 ( .A1(n9822), .A2(n9118), .ZN(n15250) );
  INV_X1 U7251 ( .A(n12026), .ZN(n11953) );
  NOR2_X1 U7252 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7424) );
  INV_X1 U7253 ( .A(n10386), .ZN(n9012) );
  NAND2_X1 U7254 ( .A1(n8559), .A2(n10826), .ZN(n8979) );
  OR2_X1 U7255 ( .A1(n12023), .A2(n9518), .ZN(n9521) );
  AND3_X1 U7256 ( .A1(n7120), .A2(n9147), .A3(n7416), .ZN(n9175) );
  NAND2_X1 U7257 ( .A1(n9978), .A2(n13042), .ZN(n9981) );
  INV_X1 U7258 ( .A(n12108), .ZN(n8460) );
  NOR2_X1 U7259 ( .A1(n8845), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8856) );
  INV_X2 U7260 ( .A(n13690), .ZN(n6487) );
  AOI22_X1 U7261 ( .A1(n6652), .A2(n14085), .B1(n7404), .B2(n6504), .ZN(n14087) );
  AOI21_X1 U7262 ( .B1(n11512), .B2(n7422), .A(n6547), .ZN(n14240) );
  INV_X1 U7263 ( .A(n11685), .ZN(n11645) );
  OR2_X1 U7264 ( .A1(n12571), .A2(n12570), .ZN(n12573) );
  NAND2_X1 U7265 ( .A1(n7028), .A2(n7034), .ZN(n8901) );
  OAI22_X1 U7266 ( .A1(n12012), .A2(n8255), .B1(n6653), .B2(n7022), .ZN(n8307)
         );
  INV_X1 U7267 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7709) );
  AND4_X1 U7268 ( .A1(n8627), .A2(n8626), .A3(n8625), .A4(n8624), .ZN(n10779)
         );
  NAND2_X1 U7269 ( .A1(n12820), .A2(n12433), .ZN(n12807) );
  XNOR2_X1 U7270 ( .A(n8889), .B(n8888), .ZN(n13053) );
  INV_X1 U7271 ( .A(n9005), .ZN(n12544) );
  INV_X1 U7272 ( .A(n10911), .ZN(n10055) );
  NAND2_X2 U7273 ( .A1(n13909), .A2(n13910), .ZN(n13908) );
  NAND2_X1 U7274 ( .A1(n13789), .A2(n13706), .ZN(n13866) );
  INV_X2 U7275 ( .A(n9188), .ZN(n11656) );
  AND2_X1 U7276 ( .A1(n6640), .A2(n6695), .ZN(n12548) );
  INV_X1 U7277 ( .A(n10959), .ZN(n12558) );
  INV_X2 U7278 ( .A(n9671), .ZN(n12623) );
  INV_X1 U7279 ( .A(n11835), .ZN(n14044) );
  XOR2_X1 U7280 ( .A(n10685), .B(n13206), .Z(n6481) );
  AOI21_X2 U7281 ( .B1(n6503), .B2(n6866), .A(n11110), .ZN(n6864) );
  NOR2_X4 U7282 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9959) );
  AND2_X2 U7283 ( .A1(n14006), .A2(n14007), .ZN(n14004) );
  NOR2_X2 U7284 ( .A1(n14898), .A2(n8692), .ZN(n14897) );
  NAND4_X4 U7285 ( .A1(n8546), .A2(n8547), .A3(n8545), .A4(n8544), .ZN(n12564)
         );
  NAND4_X2 U7286 ( .A1(n9192), .A2(n9191), .A3(n9190), .A4(n9189), .ZN(n11844)
         );
  NOR2_X2 U7287 ( .A1(n8941), .A2(n8940), .ZN(n13052) );
  NAND2_X2 U7288 ( .A1(n9822), .A2(n9510), .ZN(n13682) );
  XNOR2_X2 U7289 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n8370) );
  NAND2_X2 U7290 ( .A1(n8475), .A2(n8474), .ZN(n8601) );
  OAI222_X1 U7291 ( .A1(P3_U3151), .A2(n8459), .B1(n13054), .B2(n12114), .C1(
        n13057), .C2(n12113), .ZN(P3_U3265) );
  INV_X2 U7292 ( .A(n8459), .ZN(n8461) );
  OAI21_X2 U7293 ( .B1(n11812), .B2(n11811), .A(n11810), .ZN(n13501) );
  XNOR2_X1 U7294 ( .A(n8392), .B(n8393), .ZN(n14417) );
  NAND2_X1 U7295 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  OAI21_X2 U7296 ( .B1(n8156), .B2(n7314), .A(n7313), .ZN(n8175) );
  INV_X1 U7297 ( .A(n6686), .ZN(n6482) );
  BUF_X4 U7298 ( .A(n12478), .Z(n6483) );
  INV_X1 U7299 ( .A(n8515), .ZN(n12478) );
  OAI222_X1 U7300 ( .A1(n13057), .A2(n11565), .B1(P3_U3151), .B2(n12542), .C1(
        n15044), .C2(n13054), .ZN(P3_U3267) );
  OAI21_X2 U7301 ( .B1(n11093), .B2(n11092), .A(n11094), .ZN(n11199) );
  NAND2_X2 U7302 ( .A1(n11059), .A2(n11058), .ZN(n11093) );
  XNOR2_X2 U7303 ( .A(n12617), .B(n14411), .ZN(n12612) );
  XNOR2_X2 U7304 ( .A(n7631), .B(n7626), .ZN(n10922) );
  OR2_X1 U7305 ( .A1(n14848), .A2(n10072), .ZN(n10911) );
  AND2_X2 U7307 ( .A1(n12313), .A2(n8998), .ZN(n12530) );
  OR2_X2 U7308 ( .A1(n12200), .A2(n8926), .ZN(n12313) );
  OR2_X2 U7309 ( .A1(n7649), .A2(n7709), .ZN(n7652) );
  NAND2_X2 U7310 ( .A1(n13045), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8454) );
  OAI21_X2 U7311 ( .B1(n11024), .B2(n7075), .A(n7071), .ZN(n11298) );
  OAI21_X2 U7312 ( .B1(n10983), .B2(n8987), .A(n8988), .ZN(n11024) );
  NAND2_X2 U7313 ( .A1(n7793), .A2(n7792), .ZN(n14878) );
  OAI21_X2 U7314 ( .B1(n14205), .B2(n7131), .A(n7129), .ZN(n14168) );
  AND2_X2 U7315 ( .A1(n7654), .A2(n13630), .ZN(n7683) );
  AOI21_X2 U7316 ( .B1(n6810), .B2(n6807), .A(n6806), .ZN(n6805) );
  XNOR2_X2 U7317 ( .A(n10490), .B(n10491), .ZN(n10323) );
  NOR2_X2 U7318 ( .A1(n11172), .A2(n7079), .ZN(n11173) );
  NAND2_X1 U7319 ( .A1(n8459), .A2(n8460), .ZN(n8928) );
  BUF_X4 U7320 ( .A(n8143), .Z(n6485) );
  XNOR2_X2 U7321 ( .A(n10472), .B(n10491), .ZN(n10326) );
  OAI21_X2 U7322 ( .B1(n14925), .B2(n7086), .A(n7085), .ZN(n12596) );
  NOR2_X4 U7323 ( .A1(n7701), .A2(n7700), .ZN(n9383) );
  NAND3_X2 U7324 ( .A1(n7686), .A2(n6716), .A3(n7684), .ZN(n13213) );
  AOI21_X2 U7325 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10709), .A(n9604), .ZN(
        n9609) );
  XNOR2_X2 U7326 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8539) );
  NAND4_X2 U7327 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n13211)
         );
  NOR2_X2 U7328 ( .A1(n8379), .A2(n8380), .ZN(n8383) );
  NOR2_X2 U7329 ( .A1(n14529), .A2(n14530), .ZN(n14528) );
  NAND2_X2 U7330 ( .A1(n14419), .A2(n6651), .ZN(n14529) );
  XNOR2_X2 U7331 ( .A(n6669), .B(n9757), .ZN(n9750) );
  NAND2_X2 U7332 ( .A1(n9850), .A2(n9731), .ZN(n6669) );
  XNOR2_X2 U7333 ( .A(n8496), .B(n10923), .ZN(n8829) );
  NAND2_X2 U7334 ( .A1(n6941), .A2(n8495), .ZN(n8496) );
  XNOR2_X2 U7335 ( .A(n8396), .B(n7097), .ZN(n14418) );
  INV_X2 U7336 ( .A(n6885), .ZN(n8396) );
  AOI21_X2 U7337 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n13999), .A(n14004), .ZN(
        n9309) );
  OAI22_X2 U7338 ( .A1(n14388), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(n8433), .B2(
        n8434), .ZN(n6878) );
  XNOR2_X2 U7339 ( .A(n6880), .B(n6879), .ZN(n14388) );
  XNOR2_X2 U7340 ( .A(n12627), .B(n12628), .ZN(n12597) );
  NOR2_X2 U7341 ( .A1(n12600), .A2(n12596), .ZN(n12627) );
  OR2_X1 U7342 ( .A1(n14128), .A2(n14127), .ZN(n14130) );
  NAND2_X1 U7343 ( .A1(n8023), .A2(n8022), .ZN(n13571) );
  OR2_X1 U7344 ( .A1(n11429), .A2(n11428), .ZN(n11430) );
  NAND2_X1 U7345 ( .A1(n10522), .A2(n10521), .ZN(n10520) );
  NAND2_X1 U7346 ( .A1(n12561), .A2(n14965), .ZN(n12347) );
  INV_X2 U7347 ( .A(n14945), .ZN(n12561) );
  AND4_X2 U7348 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n10844)
         );
  INV_X1 U7349 ( .A(n13207), .ZN(n10597) );
  NAND2_X2 U7350 ( .A1(n12544), .A2(n12329), .ZN(n12463) );
  BUF_X2 U7351 ( .A(n8564), .Z(n6498) );
  NAND2_X1 U7352 ( .A1(n9909), .A2(n9908), .ZN(n11862) );
  NAND4_X1 U7353 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n13950)
         );
  INV_X4 U7354 ( .A(n7820), .ZN(n8214) );
  NAND2_X2 U7355 ( .A1(n11685), .A2(n9517), .ZN(n12023) );
  AND2_X1 U7356 ( .A1(n9181), .A2(n14373), .ZN(n11152) );
  NAND2_X4 U7357 ( .A1(n9158), .A2(n14378), .ZN(n11685) );
  NAND2_X2 U7358 ( .A1(n8336), .A2(n11800), .ZN(n7678) );
  INV_X2 U7359 ( .A(n9517), .ZN(n9515) );
  XNOR2_X1 U7360 ( .A(n8570), .B(n8569), .ZN(n9076) );
  AND2_X2 U7361 ( .A1(n6825), .A2(n7410), .ZN(n6814) );
  AOI21_X1 U7362 ( .B1(n12487), .B2(n12531), .A(n12534), .ZN(n12489) );
  MUX2_X1 U7363 ( .A(n12465), .B(n12464), .S(n12463), .Z(n12487) );
  NOR2_X1 U7364 ( .A1(n7525), .A2(n12539), .ZN(n6641) );
  NAND2_X1 U7365 ( .A1(n12729), .A2(n6535), .ZN(n12913) );
  AND2_X1 U7366 ( .A1(n7352), .A2(n7350), .ZN(n12730) );
  NAND2_X1 U7367 ( .A1(n6902), .A2(n6900), .ZN(n12214) );
  INV_X1 U7368 ( .A(n6898), .ZN(n6900) );
  NAND2_X1 U7369 ( .A1(n6923), .A2(n6921), .ZN(n6916) );
  NAND2_X1 U7370 ( .A1(n6896), .A2(n12158), .ZN(n6898) );
  AND2_X1 U7371 ( .A1(n14140), .A2(n11713), .ZN(n14111) );
  NAND3_X1 U7372 ( .A1(n12771), .A2(n6509), .A3(n7052), .ZN(n7049) );
  NAND3_X1 U7373 ( .A1(n8193), .A2(n8192), .A3(n8191), .ZN(n13625) );
  NAND2_X1 U7374 ( .A1(n7002), .A2(n11797), .ZN(n13309) );
  XNOR2_X1 U7375 ( .A(n8253), .B(n8252), .ZN(n12012) );
  AND2_X1 U7376 ( .A1(n11823), .A2(n8288), .ZN(n13304) );
  NAND2_X1 U7377 ( .A1(n11631), .A2(n11630), .ZN(n14270) );
  NAND2_X1 U7378 ( .A1(n12182), .A2(n6909), .ZN(n12253) );
  XNOR2_X1 U7379 ( .A(n8200), .B(n8199), .ZN(n13631) );
  INV_X1 U7380 ( .A(n14085), .ZN(n6488) );
  NAND2_X1 U7381 ( .A1(n8517), .A2(n8516), .ZN(n12200) );
  NOR2_X1 U7382 ( .A1(n7259), .A2(n13873), .ZN(n7258) );
  NAND2_X1 U7383 ( .A1(n12283), .A2(n12282), .ZN(n12281) );
  NAND2_X2 U7384 ( .A1(n8139), .A2(n8138), .ZN(n13526) );
  OAI21_X1 U7385 ( .B1(n7033), .B2(n7032), .A(n7042), .ZN(n8519) );
  INV_X1 U7386 ( .A(n13352), .ZN(n13537) );
  CLKBUF_X1 U7387 ( .A(n13412), .Z(n6649) );
  NAND2_X1 U7388 ( .A1(n8107), .A2(n8106), .ZN(n13369) );
  NAND2_X1 U7389 ( .A1(n11706), .A2(n11705), .ZN(n14295) );
  NAND2_X1 U7390 ( .A1(n12846), .A2(n7343), .ZN(n8828) );
  AND2_X1 U7391 ( .A1(n8123), .A2(n8122), .ZN(n13352) );
  XNOR2_X1 U7392 ( .A(n8175), .B(n8137), .ZN(n11737) );
  NAND2_X1 U7393 ( .A1(n11717), .A2(n11716), .ZN(n14290) );
  AND2_X1 U7394 ( .A1(n8879), .A2(n8878), .ZN(n12152) );
  NAND2_X1 U7395 ( .A1(n14195), .A2(n11764), .ZN(n14180) );
  NAND2_X1 U7396 ( .A1(n8505), .A2(n8504), .ZN(n8536) );
  OAI21_X2 U7397 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8156) );
  NAND2_X1 U7398 ( .A1(n6967), .A2(n6972), .ZN(n8136) );
  CLKBUF_X1 U7399 ( .A(n11526), .Z(n6742) );
  XNOR2_X1 U7400 ( .A(n6925), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8877) );
  INV_X1 U7401 ( .A(n13549), .ZN(n13388) );
  INV_X1 U7402 ( .A(n13427), .ZN(n6489) );
  NAND2_X2 U7403 ( .A1(n7625), .A2(n7624), .ZN(n13561) );
  NAND2_X2 U7404 ( .A1(n11674), .A2(n11673), .ZN(n14314) );
  AND2_X1 U7405 ( .A1(n8084), .A2(n8083), .ZN(n13549) );
  CLKBUF_X1 U7406 ( .A(n11568), .Z(n6753) );
  NAND2_X1 U7407 ( .A1(n8066), .A2(n8065), .ZN(n13557) );
  NOR2_X1 U7408 ( .A1(n8853), .A2(n8852), .ZN(n8501) );
  OR2_X1 U7409 ( .A1(n11402), .A2(n11403), .ZN(n11536) );
  NAND2_X1 U7410 ( .A1(n14473), .A2(n11464), .ZN(n14499) );
  OR2_X1 U7411 ( .A1(n14232), .A2(n13849), .ZN(n11949) );
  NOR2_X1 U7412 ( .A1(n6620), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U7413 ( .A1(n8004), .A2(n8003), .ZN(n13576) );
  OR4_X1 U7414 ( .A1(n11497), .A2(n11483), .A3(n11312), .A4(n8299), .ZN(n8300)
         );
  OR2_X1 U7415 ( .A1(n14533), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6890) );
  AND2_X1 U7416 ( .A1(n11636), .A2(n11635), .ZN(n14246) );
  OAI211_X1 U7417 ( .C1(n12573), .C2(n12575), .A(n6715), .B(n7184), .ZN(n14914) );
  XNOR2_X1 U7418 ( .A(n8018), .B(n8000), .ZN(n11638) );
  NAND2_X1 U7419 ( .A1(n10985), .A2(n12368), .ZN(n10984) );
  NAND2_X1 U7420 ( .A1(n11121), .A2(n11120), .ZN(n11142) );
  NAND2_X1 U7421 ( .A1(n8016), .A2(n7999), .ZN(n8018) );
  OR2_X1 U7422 ( .A1(n7998), .A2(n9641), .ZN(n8016) );
  NAND2_X1 U7423 ( .A1(n10778), .A2(n10777), .ZN(n10776) );
  OR2_X1 U7424 ( .A1(n14554), .A2(n14553), .ZN(n6729) );
  NAND2_X1 U7425 ( .A1(n7874), .A2(n7873), .ZN(n11291) );
  NAND2_X1 U7426 ( .A1(n10843), .A2(n10842), .ZN(n10841) );
  NAND2_X1 U7427 ( .A1(n11147), .A2(n11146), .ZN(n14492) );
  NAND2_X1 U7428 ( .A1(n8985), .A2(n12356), .ZN(n10837) );
  NAND2_X1 U7429 ( .A1(n11036), .A2(n11035), .ZN(n14503) );
  NAND2_X1 U7430 ( .A1(n6650), .A2(n6555), .ZN(n7081) );
  NAND2_X1 U7431 ( .A1(n10367), .A2(n10366), .ZN(n10444) );
  AOI21_X1 U7432 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n14778), .A(n14779), .ZN(
        n14793) );
  NAND2_X1 U7433 ( .A1(n6944), .A2(n7026), .ZN(n8771) );
  NAND4_X1 U7434 ( .A1(n8528), .A2(n8527), .A3(n8526), .A4(n8525), .ZN(n12746)
         );
  NAND2_X1 U7435 ( .A1(n10520), .A2(n10422), .ZN(n10423) );
  OAI21_X1 U7436 ( .B1(n7868), .B2(n7297), .A(n7294), .ZN(n7907) );
  BUF_X1 U7437 ( .A(n10685), .Z(n6727) );
  NAND2_X1 U7438 ( .A1(n6740), .A2(n8492), .ZN(n8756) );
  NAND2_X1 U7439 ( .A1(n7835), .A2(n7834), .ZN(n10927) );
  CLKBUF_X1 U7440 ( .A(n13173), .Z(n13185) );
  NOR2_X1 U7441 ( .A1(n10076), .A2(n10075), .ZN(n13181) );
  OR2_X1 U7442 ( .A1(n8882), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8892) );
  NAND2_X2 U7443 ( .A1(n10189), .A2(n13473), .ZN(n13476) );
  XNOR2_X1 U7444 ( .A(n6767), .B(n9791), .ZN(n9777) );
  NAND2_X1 U7445 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  NAND2_X1 U7446 ( .A1(n9776), .A2(n9775), .ZN(n6767) );
  INV_X2 U7447 ( .A(n14671), .ZN(n14646) );
  NAND2_X2 U7448 ( .A1(n11757), .A2(n14662), .ZN(n14671) );
  NAND2_X1 U7449 ( .A1(n7186), .A2(n7185), .ZN(n9776) );
  OAI21_X2 U7450 ( .B1(n9992), .B2(n9991), .A(n14940), .ZN(n9993) );
  OR2_X1 U7451 ( .A1(n9735), .A2(n9734), .ZN(n9790) );
  OR2_X1 U7452 ( .A1(n9754), .A2(n9697), .ZN(n7186) );
  INV_X2 U7453 ( .A(n8908), .ZN(n8847) );
  NAND2_X1 U7454 ( .A1(n7552), .A2(n7551), .ZN(n7768) );
  INV_X2 U7455 ( .A(n12463), .ZN(n12446) );
  BUF_X2 U7456 ( .A(n8564), .Z(n6497) );
  XNOR2_X1 U7457 ( .A(n9696), .B(n7084), .ZN(n9755) );
  BUF_X2 U7458 ( .A(n12481), .Z(n6490) );
  NAND4_X2 U7459 ( .A1(n9586), .A2(n9585), .A3(n9584), .A4(n9583), .ZN(n13947)
         );
  AND2_X1 U7460 ( .A1(n9846), .A2(n9695), .ZN(n9696) );
  BUF_X1 U7461 ( .A(n8292), .Z(n6667) );
  NAND4_X1 U7462 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n13946)
         );
  NAND4_X1 U7463 ( .A1(n7759), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n13209)
         );
  XNOR2_X1 U7464 ( .A(n11555), .B(n13950), .ZN(n12063) );
  INV_X1 U7465 ( .A(n11544), .ZN(n11555) );
  OR2_X1 U7466 ( .A1(n9848), .A2(n9847), .ZN(n9850) );
  CLKBUF_X2 U7467 ( .A(n6517), .Z(n7820) );
  INV_X4 U7468 ( .A(n11656), .ZN(n11039) );
  NOR2_X1 U7469 ( .A1(n10016), .A2(n9703), .ZN(n10015) );
  XNOR2_X1 U7470 ( .A(n8457), .B(n8456), .ZN(n12108) );
  CLKBUF_X2 U7471 ( .A(n12011), .Z(n6686) );
  AND2_X2 U7472 ( .A1(n9181), .A2(n9182), .ZN(n11743) );
  XNOR2_X1 U7473 ( .A(n7082), .B(n9726), .ZN(n10016) );
  NAND2_X1 U7474 ( .A1(n9060), .A2(n9059), .ZN(n11322) );
  INV_X1 U7475 ( .A(n12031), .ZN(n14385) );
  AND2_X1 U7476 ( .A1(n7653), .A2(n11566), .ZN(n7682) );
  CLKBUF_X1 U7477 ( .A(n8254), .Z(n6653) );
  AND2_X2 U7478 ( .A1(n7654), .A2(n7653), .ZN(n8143) );
  CLKBUF_X1 U7479 ( .A(n13472), .Z(n6754) );
  CLKBUF_X1 U7480 ( .A(n9491), .Z(n6682) );
  INV_X1 U7481 ( .A(n9491), .ZN(n8263) );
  INV_X1 U7482 ( .A(n11566), .ZN(n7654) );
  OR2_X1 U7483 ( .A1(n9725), .A2(n7083), .ZN(n7082) );
  NAND2_X2 U7484 ( .A1(n9515), .A2(P1_U3086), .ZN(n14382) );
  XNOR2_X1 U7485 ( .A(n6875), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9491) );
  NAND2_X2 U7486 ( .A1(n9515), .A2(P3_U3151), .ZN(n13057) );
  XNOR2_X1 U7487 ( .A(n7554), .B(SI_6_), .ZN(n7767) );
  NAND2_X2 U7488 ( .A1(n9517), .A2(P3_U3151), .ZN(n13054) );
  XNOR2_X1 U7489 ( .A(n8342), .B(n7090), .ZN(n8375) );
  NAND2_X1 U7490 ( .A1(n14367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9177) );
  NAND2_X2 U7491 ( .A1(n9517), .A2(P2_U3088), .ZN(n13637) );
  CLKBUF_X1 U7492 ( .A(n8336), .Z(n9494) );
  NAND2_X1 U7493 ( .A1(n9517), .A2(P1_U3086), .ZN(n14379) );
  NAND2_X1 U7494 ( .A1(n6644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U7495 ( .A1(n7093), .A2(n7091), .ZN(n8342) );
  NOR2_X2 U7496 ( .A1(n7627), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7629) );
  AND4_X1 U7497 ( .A1(n7077), .A2(n8447), .A3(n7078), .A4(n8442), .ZN(n8937)
         );
  NAND2_X1 U7498 ( .A1(n9095), .A2(n9107), .ZN(n13968) );
  OR2_X1 U7499 ( .A1(n8945), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n8814) );
  BUF_X2 U7500 ( .A(n9147), .Z(n9287) );
  INV_X1 U7501 ( .A(n7001), .ZN(n7620) );
  NAND2_X2 U7502 ( .A1(n6978), .A2(n6977), .ZN(n11682) );
  AND3_X1 U7503 ( .A1(n6999), .A2(n6599), .A3(n7889), .ZN(n6846) );
  BUF_X2 U7504 ( .A(n9076), .Z(n6500) );
  AND2_X2 U7505 ( .A1(n8713), .A2(n8446), .ZN(n8447) );
  INV_X2 U7506 ( .A(n7734), .ZN(n6492) );
  NAND2_X1 U7507 ( .A1(n9138), .A2(n9137), .ZN(n9519) );
  NAND2_X1 U7508 ( .A1(n6668), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6978) );
  INV_X1 U7509 ( .A(n8597), .ZN(n8442) );
  AND4_X1 U7510 ( .A1(n8725), .A2(n8741), .A3(n8715), .A4(n8443), .ZN(n8446)
         );
  AND2_X1 U7511 ( .A1(n7089), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8371) );
  AND4_X1 U7512 ( .A1(n8444), .A2(n8445), .A3(n8642), .A4(n15098), .ZN(n8713)
         );
  OR2_X1 U7513 ( .A1(n9666), .A2(n6496), .ZN(n8570) );
  INV_X1 U7514 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8441) );
  NOR2_X1 U7515 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8440) );
  NOR2_X2 U7516 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9666) );
  INV_X1 U7517 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8912) );
  INV_X1 U7518 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8642) );
  NOR2_X1 U7519 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8444) );
  NOR2_X1 U7520 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8445) );
  INV_X1 U7521 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8715) );
  INV_X4 U7522 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7523 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8741) );
  INV_X1 U7524 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8725) );
  INV_X1 U7525 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7532) );
  INV_X1 U7526 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14048) );
  INV_X1 U7527 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7533) );
  NOR2_X1 U7528 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8448) );
  NOR2_X1 U7529 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8449) );
  NOR2_X1 U7530 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n8450) );
  INV_X1 U7531 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n15098) );
  NOR2_X2 U7532 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7713) );
  INV_X4 U7533 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U7534 ( .A1(n12076), .A2(n11113), .ZN(n7172) );
  INV_X1 U7535 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6493) );
  AOI21_X2 U7536 ( .B1(n13168), .B2(n13167), .A(n11583), .ZN(n13076) );
  NOR2_X2 U7537 ( .A1(n13114), .A2(n11579), .ZN(n13168) );
  NAND2_X1 U7538 ( .A1(n8459), .A2(n8460), .ZN(n6494) );
  INV_X1 U7539 ( .A(n6494), .ZN(n6495) );
  NOR2_X2 U7540 ( .A1(n14546), .A2(n8422), .ZN(n14433) );
  INV_X1 U7541 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n6496) );
  INV_X2 U7542 ( .A(n12564), .ZN(n8559) );
  INV_X2 U7543 ( .A(n10147), .ZN(n6914) );
  AND2_X1 U7544 ( .A1(n8459), .A2(n12108), .ZN(n8564) );
  NAND2_X1 U7545 ( .A1(n8461), .A2(n8460), .ZN(n6499) );
  MUX2_X1 U7546 ( .A(n9211), .B(P1_REG2_REG_2__SCAN_IN), .S(n13968), .Z(n13974) );
  NOR2_X2 U7547 ( .A1(n8634), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U7548 ( .A(n14015), .B(n14583), .ZN(n14578) );
  NOR2_X2 U7549 ( .A1(n14567), .A2(n6730), .ZN(n14015) );
  NAND2_X1 U7550 ( .A1(n8461), .A2(n12108), .ZN(n12481) );
  INV_X1 U7551 ( .A(n8768), .ZN(n7328) );
  XNOR2_X1 U7552 ( .A(n8247), .B(n13292), .ZN(n8304) );
  NOR2_X1 U7553 ( .A1(n13349), .A2(n13532), .ZN(n7003) );
  INV_X1 U7554 ( .A(n6497), .ZN(n8908) );
  BUF_X1 U7555 ( .A(n12481), .Z(n6694) );
  NAND2_X1 U7556 ( .A1(n9005), .A2(n12332), .ZN(n15004) );
  AOI21_X1 U7557 ( .B1(n6504), .B2(n11775), .A(n6569), .ZN(n7402) );
  AOI22_X1 U7558 ( .A1(n6517), .A2(n13081), .B1(n6748), .B2(n8093), .ZN(n7688)
         );
  OAI22_X1 U7559 ( .A1(n11861), .A2(n11860), .B1(n7239), .B2(n11863), .ZN(
        n7237) );
  NOR2_X1 U7560 ( .A1(n7530), .A2(n11935), .ZN(n11936) );
  NOR2_X1 U7561 ( .A1(n11934), .A2(n11998), .ZN(n11935) );
  INV_X1 U7562 ( .A(n7938), .ZN(n6855) );
  NAND2_X1 U7563 ( .A1(n7978), .A2(n6550), .ZN(n7520) );
  NOR2_X1 U7564 ( .A1(n13304), .A2(n13320), .ZN(n6665) );
  INV_X1 U7565 ( .A(n7867), .ZN(n7572) );
  NAND2_X1 U7566 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7092), .ZN(n7091) );
  INV_X1 U7567 ( .A(n12332), .ZN(n12329) );
  INV_X1 U7568 ( .A(n7046), .ZN(n12535) );
  AND2_X1 U7569 ( .A1(n6500), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7083) );
  INV_X1 U7570 ( .A(n7334), .ZN(n7333) );
  OAI21_X1 U7571 ( .B1(n12511), .B2(n7335), .A(n8706), .ZN(n7334) );
  OR2_X1 U7572 ( .A1(n9036), .A2(n12720), .ZN(n12491) );
  INV_X1 U7573 ( .A(n12863), .ZN(n7330) );
  AND2_X1 U7574 ( .A1(n6590), .A2(n7385), .ZN(n7078) );
  OAI21_X1 U7575 ( .B1(n8866), .B2(n8865), .A(n6637), .ZN(n6925) );
  NOR2_X1 U7576 ( .A1(n8814), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8913) );
  AOI21_X1 U7577 ( .B1(n8640), .B2(n8480), .A(n6613), .ZN(n6939) );
  NOR2_X1 U7578 ( .A1(n13304), .A2(n7147), .ZN(n7141) );
  NOR2_X1 U7579 ( .A1(n13449), .A2(n6672), .ZN(n6516) );
  INV_X1 U7580 ( .A(n11791), .ZN(n6672) );
  NOR2_X1 U7581 ( .A1(n8292), .A2(n14847), .ZN(n9496) );
  OAI21_X2 U7582 ( .B1(n9493), .B2(n9492), .A(n13472), .ZN(n10043) );
  AND2_X1 U7583 ( .A1(n10183), .A2(n9491), .ZN(n9492) );
  AND2_X1 U7584 ( .A1(n6808), .A2(n13749), .ZN(n6807) );
  NOR2_X1 U7585 ( .A1(n7258), .A2(n13781), .ZN(n7255) );
  NAND2_X1 U7586 ( .A1(n7252), .A2(n6811), .ZN(n6810) );
  NAND2_X1 U7587 ( .A1(n7124), .A2(n7126), .ZN(n7122) );
  NAND2_X1 U7588 ( .A1(n11685), .A2(n9515), .ZN(n12011) );
  AND2_X1 U7589 ( .A1(n7526), .A2(n7273), .ZN(n7119) );
  NOR3_X1 U7590 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U7591 ( .A1(n7942), .A2(n7587), .ZN(n7961) );
  AND2_X1 U7592 ( .A1(n7592), .A2(n7591), .ZN(n7960) );
  NAND2_X1 U7593 ( .A1(n7907), .A2(n7527), .ZN(n7582) );
  XNOR2_X1 U7594 ( .A(n7566), .B(SI_10_), .ZN(n7852) );
  XNOR2_X1 U7595 ( .A(n7560), .B(SI_8_), .ZN(n7811) );
  XNOR2_X1 U7596 ( .A(n8345), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n8366) );
  OAI21_X1 U7597 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9324), .A(n8355), .ZN(
        n8395) );
  NOR2_X1 U7598 ( .A1(n9981), .A2(n10826), .ZN(n6684) );
  AND2_X1 U7599 ( .A1(n9646), .A2(n9068), .ZN(n8574) );
  OR2_X1 U7600 ( .A1(n12333), .A2(n12153), .ZN(n9984) );
  NAND2_X1 U7601 ( .A1(n12253), .A2(n7384), .ZN(n12204) );
  AND2_X1 U7602 ( .A1(n12205), .A2(n12145), .ZN(n7384) );
  NAND2_X1 U7603 ( .A1(n12281), .A2(n6617), .ZN(n12182) );
  INV_X1 U7604 ( .A(n12185), .ZN(n6911) );
  AND2_X1 U7605 ( .A1(n7046), .A2(n7045), .ZN(n12494) );
  OR2_X1 U7606 ( .A1(n10014), .A2(n9704), .ZN(n6768) );
  NOR2_X1 U7607 ( .A1(n12629), .A2(n12630), .ZN(n12632) );
  NAND2_X1 U7608 ( .A1(n7352), .A2(n7353), .ZN(n12731) );
  INV_X1 U7609 ( .A(n8575), .ZN(n8515) );
  INV_X1 U7610 ( .A(n12758), .ZN(n12327) );
  NAND2_X1 U7611 ( .A1(n8677), .A2(n8676), .ZN(n8707) );
  AOI21_X1 U7612 ( .B1(n7064), .B2(n7066), .A(n7062), .ZN(n7061) );
  INV_X1 U7613 ( .A(n12364), .ZN(n7062) );
  NAND2_X1 U7614 ( .A1(n12491), .A2(n12461), .ZN(n12533) );
  OR2_X1 U7615 ( .A1(n12944), .A2(n12858), .ZN(n12830) );
  INV_X1 U7616 ( .A(n14944), .ZN(n12896) );
  AND3_X1 U7617 ( .A1(n9664), .A2(n12446), .A3(n9646), .ZN(n12898) );
  OR2_X1 U7618 ( .A1(n9015), .A2(n9014), .ZN(n9996) );
  AND2_X1 U7619 ( .A1(n13041), .A2(n9967), .ZN(n9995) );
  AND2_X1 U7620 ( .A1(n7037), .A2(n7035), .ZN(n7034) );
  NAND2_X1 U7621 ( .A1(n8536), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U7622 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7036), .ZN(n7035) );
  NAND2_X1 U7623 ( .A1(n8536), .A2(n8506), .ZN(n7031) );
  XNOR2_X1 U7624 ( .A(n8916), .B(n8915), .ZN(n9005) );
  NAND2_X1 U7625 ( .A1(n8447), .A2(n8612), .ZN(n8786) );
  NAND2_X1 U7626 ( .A1(n7637), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7877) );
  INV_X1 U7627 ( .A(n7837), .ZN(n7637) );
  NAND2_X1 U7628 ( .A1(n7678), .A2(n9515), .ZN(n8254) );
  NOR2_X1 U7629 ( .A1(n10389), .A2(n7480), .ZN(n7479) );
  INV_X1 U7630 ( .A(n10248), .ZN(n7480) );
  NOR2_X1 U7631 ( .A1(n8312), .A2(n6688), .ZN(n6687) );
  INV_X1 U7632 ( .A(n6689), .ZN(n6688) );
  INV_X1 U7633 ( .A(n13515), .ZN(n11809) );
  INV_X1 U7634 ( .A(n13322), .ZN(n7002) );
  XNOR2_X1 U7635 ( .A(n13515), .B(n13305), .ZN(n11824) );
  XOR2_X1 U7636 ( .A(n13191), .B(n13526), .Z(n13320) );
  AOI21_X1 U7637 ( .B1(n7435), .B2(n13413), .A(n6561), .ZN(n7434) );
  NAND2_X1 U7638 ( .A1(n13434), .A2(n11794), .ZN(n13414) );
  OAI211_X1 U7639 ( .C1(n10599), .C2(n7116), .A(n10688), .B(n7115), .ZN(n10815) );
  OR2_X1 U7640 ( .A1(n7117), .A2(n7116), .ZN(n7115) );
  INV_X1 U7641 ( .A(n10686), .ZN(n7116) );
  NAND2_X1 U7642 ( .A1(n10599), .A2(n7117), .ZN(n10687) );
  NAND2_X1 U7643 ( .A1(n10524), .A2(n10428), .ZN(n10596) );
  INV_X2 U7644 ( .A(n8255), .ZN(n8236) );
  INV_X2 U7645 ( .A(n8254), .ZN(n8021) );
  NAND2_X1 U7646 ( .A1(n13866), .A2(n7255), .ZN(n7254) );
  AOI22_X1 U7647 ( .A1(n12005), .A2(n12004), .B1(n12003), .B2(n12002), .ZN(
        n12045) );
  AND4_X1 U7648 ( .A1(n11157), .A2(n11156), .A3(n11155), .A4(n11154), .ZN(
        n13661) );
  XNOR2_X1 U7649 ( .A(n14266), .B(n11625), .ZN(n12089) );
  NAND2_X1 U7650 ( .A1(n11739), .A2(n11738), .ZN(n14093) );
  AND2_X1 U7651 ( .A1(n14127), .A2(n11702), .ZN(n7160) );
  OR2_X1 U7652 ( .A1(n14345), .A2(n13674), .ZN(n11934) );
  NAND2_X1 U7653 ( .A1(n11118), .A2(n11117), .ZN(n11121) );
  NOR2_X1 U7654 ( .A1(n14385), .A2(n12019), .ZN(n14658) );
  NAND2_X1 U7655 ( .A1(n11648), .A2(n11647), .ZN(n14327) );
  OAI21_X1 U7656 ( .B1(n14417), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6539), .ZN(
        n6885) );
  AND4_X1 U7657 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(n12850)
         );
  OAI21_X1 U7658 ( .B1(n10076), .B2(n10187), .A(n13473), .ZN(n13173) );
  NOR2_X1 U7659 ( .A1(n7453), .A2(n7734), .ZN(n7632) );
  INV_X1 U7660 ( .A(n7451), .ZN(n7453) );
  NAND2_X1 U7661 ( .A1(n13631), .A2(n12025), .ZN(n11631) );
  NAND2_X1 U7662 ( .A1(n7209), .A2(n11839), .ZN(n7208) );
  AND2_X1 U7663 ( .A1(n7238), .A2(n11867), .ZN(n7236) );
  NAND2_X1 U7664 ( .A1(n7806), .A2(n7805), .ZN(n6859) );
  NAND2_X1 U7665 ( .A1(n7810), .A2(n7809), .ZN(n6858) );
  INV_X1 U7666 ( .A(n7830), .ZN(n6861) );
  NOR2_X1 U7667 ( .A1(n11905), .A2(n11902), .ZN(n6831) );
  OAI21_X1 U7668 ( .B1(n11903), .B2(n6831), .A(n6661), .ZN(n11909) );
  NOR2_X1 U7669 ( .A1(n11908), .A2(n6662), .ZN(n6661) );
  INV_X1 U7670 ( .A(n6830), .ZN(n6662) );
  INV_X1 U7671 ( .A(n11911), .ZN(n7228) );
  AND2_X1 U7672 ( .A1(n7517), .A2(n7846), .ZN(n7514) );
  AND2_X1 U7673 ( .A1(n7517), .A2(n7850), .ZN(n7512) );
  NAND2_X1 U7674 ( .A1(n7866), .A2(n7516), .ZN(n7515) );
  INV_X1 U7675 ( .A(n6549), .ZN(n7516) );
  INV_X1 U7676 ( .A(n11936), .ZN(n7216) );
  AOI21_X1 U7677 ( .B1(n11936), .B2(n6544), .A(n6508), .ZN(n7215) );
  AND2_X1 U7678 ( .A1(n6849), .A2(n6852), .ZN(n7958) );
  OAI21_X1 U7679 ( .B1(n6854), .B2(n6574), .A(n6853), .ZN(n6852) );
  INV_X1 U7680 ( .A(n7996), .ZN(n6873) );
  INV_X1 U7681 ( .A(n7997), .ZN(n6874) );
  NOR2_X1 U7682 ( .A1(n7503), .A2(n6572), .ZN(n7501) );
  NAND2_X1 U7683 ( .A1(n8015), .A2(n8012), .ZN(n7510) );
  NOR2_X1 U7684 ( .A1(n6519), .A2(n6870), .ZN(n6869) );
  NAND2_X1 U7685 ( .A1(n7224), .A2(n11980), .ZN(n7223) );
  NAND2_X1 U7686 ( .A1(n6660), .A2(n6659), .ZN(n11978) );
  NAND2_X1 U7687 ( .A1(n11979), .A2(n7221), .ZN(n7220) );
  INV_X1 U7688 ( .A(n11980), .ZN(n7221) );
  NAND2_X1 U7689 ( .A1(n6862), .A2(n7504), .ZN(n8096) );
  NAND2_X1 U7690 ( .A1(n8075), .A2(n8076), .ZN(n7504) );
  OR2_X1 U7691 ( .A1(n8059), .A2(n6863), .ZN(n6862) );
  INV_X1 U7692 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8486) );
  OR4_X1 U7693 ( .A1(n8301), .A2(n13393), .A3(n13411), .A4(n13432), .ZN(n8302)
         );
  NAND3_X1 U7694 ( .A1(n7713), .A2(n7615), .A3(n7000), .ZN(n7001) );
  AND4_X1 U7695 ( .A1(n7616), .A2(n7619), .A3(n7618), .A4(n7617), .ZN(n7000)
         );
  NOR2_X1 U7696 ( .A1(n6681), .A2(n7709), .ZN(n6673) );
  INV_X1 U7697 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6681) );
  INV_X1 U7698 ( .A(n13857), .ZN(n6811) );
  INV_X1 U7699 ( .A(n7396), .ZN(n7395) );
  OAI21_X1 U7700 ( .B1(n11141), .B2(n7397), .A(n12077), .ZN(n7396) );
  INV_X1 U7701 ( .A(n11144), .ZN(n7397) );
  INV_X1 U7702 ( .A(n7592), .ZN(n6955) );
  INV_X1 U7703 ( .A(n6954), .ZN(n6953) );
  OAI21_X1 U7704 ( .B1(n7960), .B2(n6955), .A(n9549), .ZN(n6954) );
  AOI21_X1 U7705 ( .B1(n6952), .B2(n6956), .A(n6951), .ZN(n6950) );
  INV_X1 U7706 ( .A(n7979), .ZN(n6951) );
  INV_X1 U7707 ( .A(n7960), .ZN(n6952) );
  AND2_X1 U7708 ( .A1(n7103), .A2(n7102), .ZN(n7526) );
  NOR2_X1 U7709 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n7103) );
  NOR2_X1 U7710 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7102) );
  OAI22_X1 U7711 ( .A1(n6502), .A2(n7924), .B1(n7581), .B2(SI_14_), .ZN(n7301)
         );
  NAND2_X1 U7712 ( .A1(n7578), .A2(n14403), .ZN(n7581) );
  AOI21_X1 U7713 ( .B1(n7788), .B2(n7559), .A(n7811), .ZN(n6962) );
  OAI21_X1 U7714 ( .B1(n9517), .B2(n6691), .A(n6690), .ZN(n7558) );
  NAND2_X1 U7715 ( .A1(n9517), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6690) );
  AND2_X1 U7716 ( .A1(n9980), .A2(n10826), .ZN(n7379) );
  INV_X1 U7717 ( .A(n11326), .ZN(n7377) );
  NAND2_X1 U7718 ( .A1(n6908), .A2(n10943), .ZN(n6906) );
  INV_X1 U7719 ( .A(n12159), .ZN(n6901) );
  AOI21_X1 U7720 ( .B1(n14438), .B2(n12493), .A(n12492), .ZN(n7045) );
  AND2_X1 U7721 ( .A1(n6500), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U7722 ( .A1(n12634), .A2(n12875), .ZN(n6765) );
  NAND2_X1 U7723 ( .A1(n8620), .A2(n8604), .ZN(n7347) );
  AND2_X1 U7724 ( .A1(n12355), .A2(n12356), .ZN(n12506) );
  NAND2_X1 U7725 ( .A1(n8979), .A2(n8980), .ZN(n14936) );
  AOI21_X1 U7726 ( .B1(n7339), .B2(n12784), .A(n6570), .ZN(n7338) );
  NOR2_X1 U7727 ( .A1(n7059), .A2(n6553), .ZN(n7057) );
  INV_X1 U7728 ( .A(n12438), .ZN(n7059) );
  INV_X1 U7729 ( .A(n8996), .ZN(n7058) );
  INV_X1 U7730 ( .A(n12439), .ZN(n7055) );
  OR2_X1 U7731 ( .A1(n12991), .A2(n12812), .ZN(n12439) );
  INV_X1 U7732 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8452) );
  INV_X1 U7733 ( .A(n8944), .ZN(n7077) );
  INV_X1 U7734 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n6703) );
  INV_X1 U7735 ( .A(n8670), .ZN(n6935) );
  AOI21_X1 U7736 ( .B1(n6931), .B2(n8476), .A(n6612), .ZN(n6930) );
  INV_X1 U7737 ( .A(n8476), .ZN(n6932) );
  INV_X1 U7738 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7386) );
  INV_X1 U7739 ( .A(n13061), .ZN(n7466) );
  INV_X1 U7740 ( .A(n11607), .ZN(n7464) );
  INV_X1 U7741 ( .A(n11597), .ZN(n7473) );
  NOR2_X1 U7742 ( .A1(n13178), .A2(n7468), .ZN(n7467) );
  INV_X1 U7743 ( .A(n7470), .ZN(n7468) );
  INV_X1 U7744 ( .A(n11612), .ZN(n11604) );
  AND2_X1 U7745 ( .A1(n13292), .A2(n8215), .ZN(n7499) );
  AOI21_X1 U7746 ( .B1(n7495), .B2(n7496), .A(n6877), .ZN(n6876) );
  AND2_X1 U7747 ( .A1(n8173), .A2(n7497), .ZN(n7496) );
  INV_X1 U7748 ( .A(n6528), .ZN(n7138) );
  NOR2_X1 U7749 ( .A1(n7140), .A2(n7137), .ZN(n7136) );
  NOR2_X1 U7750 ( .A1(n13334), .A2(n7138), .ZN(n7137) );
  NAND2_X1 U7751 ( .A1(n7143), .A2(n7145), .ZN(n7140) );
  INV_X1 U7752 ( .A(n7141), .ZN(n7139) );
  NAND2_X1 U7753 ( .A1(n11797), .A2(n13190), .ZN(n7145) );
  INV_X1 U7754 ( .A(n13320), .ZN(n7143) );
  INV_X1 U7755 ( .A(n13385), .ZN(n6723) );
  AND2_X1 U7756 ( .A1(n7712), .A2(n7614), .ZN(n7615) );
  INV_X1 U7757 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7614) );
  NOR2_X1 U7758 ( .A1(n6538), .A2(n7107), .ZN(n7106) );
  NOR2_X1 U7759 ( .A1(n11205), .A2(n7108), .ZN(n7107) );
  INV_X1 U7760 ( .A(n11310), .ZN(n7108) );
  NAND2_X1 U7761 ( .A1(n7157), .A2(n11056), .ZN(n7155) );
  OR2_X1 U7762 ( .A1(n11255), .A2(n8290), .ZN(n11203) );
  NOR2_X1 U7763 ( .A1(n11066), .A2(n7158), .ZN(n7157) );
  INV_X1 U7764 ( .A(n11063), .ZN(n7158) );
  AND2_X1 U7765 ( .A1(n7118), .A2(n10598), .ZN(n7117) );
  NAND2_X1 U7766 ( .A1(n7439), .A2(n13137), .ZN(n7438) );
  NAND2_X1 U7767 ( .A1(n13503), .A2(n7440), .ZN(n13477) );
  NOR2_X1 U7768 ( .A1(n13480), .A2(n7441), .ZN(n7440) );
  INV_X1 U7769 ( .A(n11813), .ZN(n7441) );
  AND2_X1 U7770 ( .A1(n10922), .A2(n11500), .ZN(n8305) );
  INV_X1 U7771 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U7772 ( .A1(n6811), .A2(n6809), .ZN(n6808) );
  INV_X1 U7773 ( .A(n13858), .ZN(n6809) );
  AOI21_X1 U7774 ( .B1(n7255), .B2(n6526), .A(n7253), .ZN(n7252) );
  INV_X1 U7775 ( .A(n13780), .ZN(n7253) );
  AND2_X1 U7776 ( .A1(n13812), .A2(n6540), .ZN(n7262) );
  AND2_X1 U7777 ( .A1(n12042), .A2(n12041), .ZN(n12048) );
  OR2_X1 U7778 ( .A1(n14283), .A2(n11774), .ZN(n7403) );
  NOR2_X1 U7779 ( .A1(n14145), .A2(n7407), .ZN(n7406) );
  INV_X1 U7780 ( .A(n11766), .ZN(n7407) );
  NOR2_X1 U7781 ( .A1(n11637), .A2(n7128), .ZN(n7127) );
  INV_X1 U7782 ( .A(n11632), .ZN(n7128) );
  INV_X1 U7783 ( .A(n12072), .ZN(n7420) );
  OR2_X1 U7784 ( .A1(n10750), .A2(n10756), .ZN(n7421) );
  OR2_X1 U7785 ( .A1(n7402), .A2(n7400), .ZN(n7399) );
  INV_X1 U7786 ( .A(n11779), .ZN(n7400) );
  NOR2_X1 U7787 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9055) );
  AND3_X1 U7788 ( .A1(n9054), .A2(n9099), .A3(n9053), .ZN(n6825) );
  OR2_X1 U7789 ( .A1(n9175), .A2(n14366), .ZN(n9154) );
  OAI21_X1 U7790 ( .B1(n8175), .B2(n8174), .A(n6965), .ZN(n8200) );
  AOI21_X1 U7791 ( .B1(n7314), .B2(n7313), .A(n7312), .ZN(n7311) );
  AND2_X1 U7792 ( .A1(n9092), .A2(n9055), .ZN(n6815) );
  NAND2_X1 U7793 ( .A1(n6969), .A2(n6968), .ZN(n6967) );
  INV_X1 U7794 ( .A(n8103), .ZN(n6968) );
  NAND2_X1 U7795 ( .A1(n7582), .A2(n7581), .ZN(n7299) );
  AOI21_X1 U7796 ( .B1(n7296), .B2(n7298), .A(n7295), .ZN(n7294) );
  INV_X1 U7797 ( .A(n7577), .ZN(n7295) );
  INV_X1 U7798 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U7799 ( .A(n7558), .B(SI_7_), .ZN(n7788) );
  NAND2_X1 U7800 ( .A1(n7556), .A2(n7555), .ZN(n7789) );
  INV_X1 U7801 ( .A(n7767), .ZN(n7553) );
  INV_X1 U7802 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9099) );
  INV_X1 U7803 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7090) );
  OAI21_X1 U7804 ( .B1(n8366), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n8346), .ZN(
        n8347) );
  XOR2_X1 U7805 ( .A(n8347), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n8381) );
  AOI22_X1 U7806 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9249), .B1(n8386), .B2(
        n8350), .ZN(n8352) );
  AOI21_X1 U7807 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n10352), .A(n8359), .ZN(
        n8403) );
  NOR2_X1 U7808 ( .A1(n8400), .A2(n8399), .ZN(n8359) );
  AND2_X1 U7809 ( .A1(n7364), .A2(n12215), .ZN(n7363) );
  INV_X1 U7810 ( .A(n12290), .ZN(n7364) );
  NAND2_X1 U7811 ( .A1(n12161), .A2(n12218), .ZN(n7367) );
  OR2_X1 U7812 ( .A1(n12290), .A2(n7368), .ZN(n7365) );
  AND2_X1 U7813 ( .A1(n11082), .A2(n11080), .ZN(n6908) );
  AND2_X1 U7814 ( .A1(n9646), .A2(n9517), .ZN(n8575) );
  NOR2_X1 U7815 ( .A1(n12128), .A2(n7383), .ZN(n7382) );
  INV_X1 U7816 ( .A(n12126), .ZN(n7383) );
  INV_X1 U7817 ( .A(n12155), .ZN(n12240) );
  AND2_X1 U7818 ( .A1(n9983), .A2(n10828), .ZN(n6676) );
  NOR2_X1 U7819 ( .A1(n12159), .A2(n12551), .ZN(n6903) );
  NOR2_X1 U7820 ( .A1(n12489), .A2(n12535), .ZN(n12541) );
  NAND4_X1 U7821 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n12563)
         );
  OR2_X1 U7822 ( .A1(n6490), .A2(n9652), .ZN(n8568) );
  OR2_X1 U7823 ( .A1(n6494), .A2(n9651), .ZN(n8566) );
  OR2_X1 U7824 ( .A1(n8905), .A2(n8549), .ZN(n8553) );
  INV_X1 U7825 ( .A(n9843), .ZN(n7178) );
  INV_X1 U7826 ( .A(n7082), .ZN(n9727) );
  INV_X1 U7827 ( .A(n9700), .ZN(n7185) );
  NOR2_X1 U7828 ( .A1(n10491), .A2(n10490), .ZN(n10493) );
  NOR2_X1 U7829 ( .A1(n10489), .A2(n10478), .ZN(n7079) );
  AND2_X1 U7830 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  OAI21_X1 U7831 ( .B1(n12652), .B2(n12651), .A(n12650), .ZN(n12653) );
  NOR2_X1 U7832 ( .A1(n12634), .A2(n12949), .ZN(n7088) );
  INV_X1 U7833 ( .A(n13050), .ZN(n9671) );
  AOI21_X1 U7834 ( .B1(n7350), .B2(n8897), .A(n6568), .ZN(n7349) );
  INV_X1 U7835 ( .A(n6945), .ZN(n7052) );
  INV_X1 U7836 ( .A(n12528), .ZN(n12744) );
  NAND2_X1 U7837 ( .A1(n12822), .A2(n12821), .ZN(n7322) );
  AND4_X1 U7838 ( .A1(n8826), .A2(n8825), .A3(n8824), .A4(n8823), .ZN(n12851)
         );
  AOI21_X1 U7839 ( .B1(n7074), .B2(n7073), .A(n7072), .ZN(n7071) );
  INV_X1 U7840 ( .A(n12376), .ZN(n7072) );
  AOI21_X1 U7841 ( .B1(n7333), .B2(n7335), .A(n6621), .ZN(n7332) );
  AND4_X1 U7842 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n12264)
         );
  NAND2_X1 U7843 ( .A1(n11021), .A2(n12511), .ZN(n11020) );
  INV_X1 U7844 ( .A(n14399), .ZN(n10491) );
  AND4_X1 U7845 ( .A1(n8682), .A2(n8681), .A3(n8680), .A4(n8679), .ZN(n11274)
         );
  AND4_X1 U7846 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n11085)
         );
  AND2_X1 U7847 ( .A1(n12369), .A2(n12370), .ZN(n12505) );
  NAND2_X1 U7848 ( .A1(n10837), .A2(n12503), .ZN(n10839) );
  INV_X1 U7849 ( .A(n7347), .ZN(n7346) );
  INV_X1 U7850 ( .A(n12506), .ZN(n8620) );
  NAND2_X1 U7851 ( .A1(n10112), .A2(n10113), .ZN(n10111) );
  INV_X1 U7852 ( .A(n12898), .ZN(n14943) );
  NAND2_X1 U7853 ( .A1(n7047), .A2(n12479), .ZN(n12488) );
  NAND2_X1 U7854 ( .A1(n13043), .A2(n12477), .ZN(n7047) );
  NAND2_X1 U7855 ( .A1(n8864), .A2(n8863), .ZN(n12789) );
  AND2_X1 U7856 ( .A1(n12319), .A2(n12321), .ZN(n12775) );
  INV_X1 U7857 ( .A(n7320), .ZN(n7319) );
  AOI21_X1 U7858 ( .B1(n7320), .B2(n7318), .A(n7317), .ZN(n7316) );
  NOR2_X1 U7859 ( .A1(n8839), .A2(n7321), .ZN(n7320) );
  AND2_X1 U7860 ( .A1(n12439), .A2(n12438), .ZN(n12799) );
  INV_X1 U7861 ( .A(n12525), .ZN(n12808) );
  NAND2_X1 U7862 ( .A1(n8819), .A2(n8818), .ZN(n12522) );
  NAND2_X1 U7863 ( .A1(n8995), .A2(n6506), .ZN(n12845) );
  AND4_X1 U7864 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n12858)
         );
  AOI21_X1 U7865 ( .B1(n6501), .B2(n7327), .A(n6622), .ZN(n7326) );
  CLKBUF_X1 U7866 ( .A(n12881), .Z(n12882) );
  INV_X1 U7867 ( .A(n12861), .ZN(n14947) );
  NAND2_X1 U7868 ( .A1(n7370), .A2(n13052), .ZN(n9170) );
  NAND2_X1 U7869 ( .A1(n8950), .A2(n11388), .ZN(n7370) );
  NAND2_X1 U7870 ( .A1(n12471), .A2(n12470), .ZN(n7023) );
  AOI21_X1 U7871 ( .B1(n7025), .B2(n12112), .A(n7024), .ZN(n12471) );
  AND2_X1 U7872 ( .A1(n11622), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7024) );
  INV_X1 U7873 ( .A(n12111), .ZN(n7025) );
  INV_X1 U7874 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U7875 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n7043), .ZN(n7042) );
  NOR2_X1 U7876 ( .A1(n7040), .A2(n7041), .ZN(n7039) );
  INV_X1 U7877 ( .A(n8888), .ZN(n7040) );
  NAND2_X1 U7878 ( .A1(n8877), .A2(n11704), .ZN(n8505) );
  INV_X1 U7879 ( .A(n6925), .ZN(n8503) );
  NOR2_X1 U7880 ( .A1(n8945), .A2(n8942), .ZN(n8943) );
  NAND2_X1 U7881 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7388) );
  NAND2_X1 U7882 ( .A1(n8499), .A2(n6639), .ZN(n8853) );
  NAND2_X1 U7883 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n15204), .ZN(n6639) );
  NAND2_X1 U7884 ( .A1(n8917), .A2(n8918), .ZN(n8955) );
  INV_X1 U7885 ( .A(n8924), .ZN(n8917) );
  NAND2_X1 U7886 ( .A1(n6942), .A2(n7012), .ZN(n8813) );
  NAND2_X1 U7887 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7013), .ZN(n7012) );
  XNOR2_X1 U7888 ( .A(n8816), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12690) );
  NAND3_X1 U7889 ( .A1(n8447), .A2(n6912), .A3(n7385), .ZN(n8945) );
  NOR2_X1 U7890 ( .A1(n8597), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U7891 ( .A1(n6943), .A2(n8493), .ZN(n8785) );
  NAND2_X1 U7892 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10126), .ZN(n8493) );
  NAND2_X1 U7893 ( .A1(n8490), .A2(n8489), .ZN(n8739) );
  INV_X1 U7894 ( .A(n8487), .ZN(n7019) );
  XNOR2_X1 U7895 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8670) );
  AOI21_X1 U7896 ( .B1(n6939), .B2(n6937), .A(n6577), .ZN(n6936) );
  INV_X1 U7897 ( .A(n8480), .ZN(n6937) );
  INV_X1 U7898 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8481) );
  INV_X1 U7899 ( .A(n6939), .ZN(n6938) );
  CLKBUF_X1 U7900 ( .A(n8641), .Z(n6751) );
  NAND2_X1 U7901 ( .A1(n15157), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8476) );
  XNOR2_X1 U7902 ( .A(n7183), .B(P3_IR_REG_1__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U7903 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7183) );
  AND2_X1 U7904 ( .A1(n8470), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8555) );
  INV_X1 U7905 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U7906 ( .A1(n6735), .A2(n7819), .ZN(n10685) );
  NAND2_X1 U7907 ( .A1(n10708), .A2(n8236), .ZN(n6735) );
  AND2_X1 U7908 ( .A1(n10046), .A2(n10045), .ZN(n13084) );
  OR2_X1 U7909 ( .A1(n7877), .A2(n7638), .ZN(n7895) );
  AND2_X1 U7910 ( .A1(n11569), .A2(n11570), .ZN(n7488) );
  AND2_X1 U7911 ( .A1(n7487), .A2(n7486), .ZN(n7485) );
  INV_X1 U7912 ( .A(n13108), .ZN(n7486) );
  OR2_X1 U7913 ( .A1(n7488), .A2(n7489), .ZN(n7487) );
  AND2_X1 U7914 ( .A1(n11239), .A2(n11236), .ZN(n7482) );
  INV_X1 U7915 ( .A(n7682), .ZN(n7969) );
  INV_X1 U7916 ( .A(n7683), .ZN(n7775) );
  INV_X1 U7917 ( .A(n7969), .ZN(n7794) );
  AND2_X1 U7918 ( .A1(n7685), .A2(n7447), .ZN(n6716) );
  NAND3_X1 U7919 ( .A1(n7664), .A2(n7665), .A3(n7666), .ZN(n8292) );
  AND2_X1 U7920 ( .A1(n7663), .A2(n7662), .ZN(n7665) );
  NAND2_X1 U7921 ( .A1(n8027), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7666) );
  AND2_X1 U7922 ( .A1(n9339), .A2(n9382), .ZN(n9384) );
  AND2_X1 U7923 ( .A1(n8245), .A2(n8244), .ZN(n13305) );
  NAND2_X1 U7924 ( .A1(n7144), .A2(n7143), .ZN(n7142) );
  OR2_X1 U7925 ( .A1(n13520), .A2(n13190), .ZN(n8288) );
  XNOR2_X1 U7926 ( .A(n13532), .B(n13192), .ZN(n13334) );
  OR2_X1 U7927 ( .A1(n6649), .A2(n13413), .ZN(n7437) );
  NAND2_X1 U7928 ( .A1(n11793), .A2(n11792), .ZN(n13434) );
  AOI21_X1 U7929 ( .B1(n6516), .B2(n11790), .A(n7175), .ZN(n7174) );
  NAND2_X1 U7930 ( .A1(n11789), .A2(n11788), .ZN(n13468) );
  NAND2_X1 U7931 ( .A1(n6720), .A2(n6545), .ZN(n11789) );
  NAND2_X1 U7932 ( .A1(n13501), .A2(n13500), .ZN(n13503) );
  NAND2_X1 U7933 ( .A1(n7615), .A2(n7713), .ZN(n7734) );
  OR3_X1 U7934 ( .A1(n7930), .A2(n7929), .A3(n11404), .ZN(n7947) );
  NAND2_X1 U7935 ( .A1(n11206), .A2(n11205), .ZN(n11311) );
  NAND2_X1 U7936 ( .A1(n10817), .A2(n10816), .ZN(n11064) );
  NAND2_X1 U7937 ( .A1(n10596), .A2(n10595), .ZN(n10599) );
  INV_X1 U7938 ( .A(n6481), .ZN(n7118) );
  NAND2_X1 U7939 ( .A1(n10423), .A2(n10429), .ZN(n10590) );
  NOR2_X1 U7940 ( .A1(n7430), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U7941 ( .A1(n9945), .A2(n9944), .ZN(n10266) );
  NAND2_X1 U7942 ( .A1(n9942), .A2(n9941), .ZN(n10405) );
  XNOR2_X1 U7943 ( .A(n8293), .B(n13158), .ZN(n9625) );
  NAND2_X1 U7944 ( .A1(n9626), .A2(n9625), .ZN(n9942) );
  INV_X1 U7945 ( .A(n13445), .ZN(n13435) );
  AND2_X1 U7946 ( .A1(n10063), .A2(n9494), .ZN(n13437) );
  NAND2_X1 U7947 ( .A1(n7315), .A2(n8238), .ZN(n13515) );
  NAND2_X1 U7948 ( .A1(n13629), .A2(n8236), .ZN(n7315) );
  AND2_X1 U7949 ( .A1(n13310), .A2(n13309), .ZN(n13519) );
  OR2_X1 U7950 ( .A1(n10952), .A2(n8255), .ZN(n8066) );
  NAND2_X1 U7951 ( .A1(n7859), .A2(n7858), .ZN(n11062) );
  NAND2_X1 U7952 ( .A1(n7774), .A2(n7773), .ZN(n10567) );
  INV_X1 U7953 ( .A(n10336), .ZN(n10093) );
  INV_X1 U7954 ( .A(n14859), .ZN(n14877) );
  NOR2_X1 U7955 ( .A1(n7648), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7649) );
  NAND3_X1 U7956 ( .A1(n7451), .A2(n7446), .A3(n7620), .ZN(n7648) );
  AND2_X1 U7957 ( .A1(n7622), .A2(n7646), .ZN(n7446) );
  INV_X1 U7958 ( .A(n8063), .ZN(n6983) );
  INV_X1 U7959 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6848) );
  AOI21_X1 U7960 ( .B1(n13772), .B2(n13769), .A(n13796), .ZN(n6787) );
  AOI21_X1 U7961 ( .B1(n14270), .B2(n9526), .A(n7276), .ZN(n13799) );
  NAND2_X1 U7962 ( .A1(n13866), .A2(n13865), .ZN(n7263) );
  NAND2_X1 U7963 ( .A1(n14499), .A2(n11468), .ZN(n11474) );
  NAND2_X1 U7964 ( .A1(n7263), .A2(n7262), .ZN(n13875) );
  NAND2_X1 U7965 ( .A1(n6507), .A2(n7269), .ZN(n7268) );
  INV_X1 U7966 ( .A(n13834), .ZN(n7269) );
  NAND2_X1 U7967 ( .A1(n6582), .A2(n6507), .ZN(n7267) );
  NAND2_X1 U7968 ( .A1(n6779), .A2(n7265), .ZN(n13885) );
  AND2_X1 U7969 ( .A1(n13887), .A2(n7266), .ZN(n7265) );
  NAND2_X1 U7970 ( .A1(n13908), .A2(n7267), .ZN(n6779) );
  NAND2_X1 U7971 ( .A1(n7267), .A2(n7268), .ZN(n7266) );
  NAND2_X1 U7972 ( .A1(n10441), .A2(n10440), .ZN(n10446) );
  INV_X1 U7973 ( .A(n6812), .ZN(n7250) );
  OAI21_X1 U7974 ( .B1(n10445), .B2(n7251), .A(n10660), .ZN(n6812) );
  OAI21_X1 U7975 ( .B1(n6800), .B2(n6799), .A(n6798), .ZN(n13895) );
  AOI21_X1 U7976 ( .B1(n6805), .B2(n6803), .A(n6802), .ZN(n6798) );
  INV_X1 U7977 ( .A(n6805), .ZN(n6799) );
  OR2_X1 U7978 ( .A1(n13677), .A2(n13676), .ZN(n13910) );
  NAND2_X1 U7979 ( .A1(n11743), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U7980 ( .A1(n11152), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U7981 ( .A1(n11653), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9295) );
  INV_X1 U7982 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13983) );
  OR2_X1 U7983 ( .A1(n14090), .A2(n14270), .ZN(n14072) );
  OR2_X1 U7984 ( .A1(n14089), .A2(n14093), .ZN(n14090) );
  NAND2_X1 U7985 ( .A1(n14130), .A2(n11771), .ZN(n14112) );
  NAND2_X1 U7986 ( .A1(n6757), .A2(n14145), .ZN(n14147) );
  NAND2_X1 U7987 ( .A1(n14179), .A2(n11766), .ZN(n14161) );
  NAND2_X1 U7988 ( .A1(n14180), .A2(n14181), .ZN(n14179) );
  NAND2_X1 U7989 ( .A1(n14205), .A2(n14204), .ZN(n14203) );
  NOR2_X1 U7990 ( .A1(n14204), .A2(n7412), .ZN(n7411) );
  INV_X1 U7991 ( .A(n11763), .ZN(n7412) );
  NAND2_X1 U7992 ( .A1(n14222), .A2(n7413), .ZN(n14215) );
  NOR2_X1 U7993 ( .A1(n11657), .A2(n7414), .ZN(n7413) );
  INV_X1 U7994 ( .A(n11949), .ZN(n7414) );
  AND2_X1 U7995 ( .A1(n11641), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U7996 ( .A1(n14239), .A2(n11761), .ZN(n14223) );
  NAND2_X1 U7997 ( .A1(n14223), .A2(n6836), .ZN(n14222) );
  NAND2_X1 U7998 ( .A1(n6742), .A2(n12083), .ZN(n11633) );
  NAND2_X1 U7999 ( .A1(n11430), .A2(n6511), .ZN(n11512) );
  NAND2_X1 U8000 ( .A1(n6756), .A2(n6755), .ZN(n7159) );
  NAND2_X1 U8001 ( .A1(n6743), .A2(n6534), .ZN(n7173) );
  NAND2_X1 U8002 ( .A1(n11032), .A2(n11031), .ZN(n11118) );
  AND2_X1 U8003 ( .A1(n10450), .A2(n10449), .ZN(n11865) );
  AOI21_X1 U8004 ( .B1(n13625), .B2(n12025), .A(n12024), .ZN(n14258) );
  NAND2_X1 U8005 ( .A1(n11624), .A2(n11623), .ZN(n14266) );
  AND2_X1 U8006 ( .A1(n14384), .A2(n11685), .ZN(n14308) );
  NAND2_X1 U8007 ( .A1(n11116), .A2(n11115), .ZN(n14424) );
  AND2_X1 U8008 ( .A1(n7417), .A2(n9061), .ZN(n7416) );
  NOR2_X1 U8009 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7417) );
  NAND2_X1 U8010 ( .A1(n8234), .A2(n8233), .ZN(n8250) );
  AND2_X1 U8011 ( .A1(n9287), .A2(n7274), .ZN(n7271) );
  INV_X1 U8012 ( .A(n6967), .ZN(n6966) );
  NAND2_X1 U8013 ( .A1(n8102), .A2(SI_24_), .ZN(n6972) );
  XNOR2_X1 U8014 ( .A(n9151), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U8015 ( .A1(n6648), .A2(SI_20_), .ZN(n7600) );
  NAND2_X1 U8016 ( .A1(n7241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9289) );
  NOR2_X1 U8017 ( .A1(n7244), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U8018 ( .A1(n6958), .A2(n7592), .ZN(n7981) );
  NAND2_X1 U8019 ( .A1(n7961), .A2(n7960), .ZN(n6958) );
  XNOR2_X1 U8020 ( .A(n7961), .B(n7960), .ZN(n11509) );
  XNOR2_X1 U8021 ( .A(n7888), .B(n7528), .ZN(n11114) );
  NAND2_X1 U8022 ( .A1(n7870), .A2(n7573), .ZN(n7888) );
  XNOR2_X1 U8023 ( .A(n8370), .B(n8371), .ZN(n8372) );
  NAND2_X1 U8024 ( .A1(n6894), .A2(n6893), .ZN(n6892) );
  NAND2_X1 U8025 ( .A1(n8374), .A2(n14394), .ZN(n6893) );
  INV_X1 U8026 ( .A(n14391), .ZN(n6894) );
  XNOR2_X1 U8027 ( .A(n9306), .B(n8381), .ZN(n8382) );
  NAND2_X1 U8028 ( .A1(n14408), .A2(n14407), .ZN(n7099) );
  AOI21_X1 U8029 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9603), .A(n8356), .ZN(
        n8362) );
  NOR2_X1 U8030 ( .A1(n8395), .A2(n8394), .ZN(n8356) );
  AOI21_X1 U8031 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n15069), .A(n8360), .ZN(
        n8407) );
  NOR2_X1 U8032 ( .A1(n8403), .A2(n8402), .ZN(n8360) );
  OR2_X1 U8033 ( .A1(n14535), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6889) );
  AND3_X1 U8034 ( .A1(n8690), .A2(n8689), .A3(n8688), .ZN(n11089) );
  AND4_X1 U8035 ( .A1(n8639), .A2(n8638), .A3(n8637), .A4(n8636), .ZN(n10959)
         );
  AND2_X1 U8036 ( .A1(n12253), .A2(n12145), .ZN(n12206) );
  NAND2_X1 U8037 ( .A1(n12231), .A2(n12136), .ZN(n12283) );
  INV_X1 U8038 ( .A(n12303), .ZN(n12294) );
  OAI211_X1 U8039 ( .C1(n6902), .C2(n6899), .A(n7368), .B(n6897), .ZN(n6904)
         );
  INV_X1 U8040 ( .A(n12215), .ZN(n6899) );
  NAND2_X1 U8041 ( .A1(n6898), .A2(n12215), .ZN(n6897) );
  NAND2_X1 U8042 ( .A1(n9988), .A2(n9995), .ZN(n12311) );
  INV_X1 U8043 ( .A(n12257), .ZN(n12307) );
  INV_X1 U8044 ( .A(n12858), .ZN(n12834) );
  INV_X1 U8045 ( .A(n12299), .ZN(n12897) );
  AND2_X1 U8046 ( .A1(n12665), .A2(n12666), .ZN(n6771) );
  OAI21_X1 U8047 ( .B1(n12681), .B2(n14928), .A(n6774), .ZN(n6773) );
  AOI21_X1 U8048 ( .B1(n12669), .B2(n12688), .A(n6775), .ZN(n6774) );
  NAND2_X1 U8049 ( .A1(n12667), .A2(n12668), .ZN(n6775) );
  OR2_X1 U8050 ( .A1(n9672), .A2(n9671), .ZN(n14926) );
  NAND2_X1 U8051 ( .A1(n12913), .A2(n14993), .ZN(n12733) );
  INV_X1 U8052 ( .A(n12154), .ZN(n12926) );
  NAND2_X1 U8053 ( .A1(n8844), .A2(n8843), .ZN(n12933) );
  NAND2_X1 U8054 ( .A1(n8803), .A2(n8802), .ZN(n12944) );
  AND3_X1 U8055 ( .A1(n8619), .A2(n8618), .A3(n8617), .ZN(n14976) );
  NAND2_X1 U8056 ( .A1(n6579), .A2(n6916), .ZN(n12495) );
  NAND2_X1 U8057 ( .A1(n8774), .A2(n8773), .ZN(n13021) );
  OR2_X1 U8058 ( .A1(n15012), .A2(n15004), .ZN(n13039) );
  AOI21_X1 U8059 ( .B1(n7479), .B2(n7477), .A(n7476), .ZN(n7475) );
  INV_X1 U8060 ( .A(n10253), .ZN(n7476) );
  NAND2_X1 U8061 ( .A1(n11737), .A2(n8236), .ZN(n8139) );
  NAND2_X1 U8062 ( .A1(n13156), .A2(n6667), .ZN(n7456) );
  NAND2_X1 U8063 ( .A1(n13155), .A2(n13212), .ZN(n7457) );
  NAND2_X1 U8064 ( .A1(n9332), .A2(n9466), .ZN(n7165) );
  NAND2_X1 U8065 ( .A1(n7164), .A2(n9515), .ZN(n7162) );
  NAND2_X1 U8066 ( .A1(n10067), .A2(n10066), .ZN(n10087) );
  INV_X1 U8067 ( .A(n10069), .ZN(n10066) );
  OR2_X1 U8068 ( .A1(n11659), .A2(n8255), .ZN(n8043) );
  AND2_X1 U8069 ( .A1(n10071), .A2(n10065), .ZN(n13162) );
  INV_X1 U8070 ( .A(n8316), .ZN(n6866) );
  NAND2_X1 U8071 ( .A1(n6503), .A2(n8287), .ZN(n6867) );
  XNOR2_X1 U8072 ( .A(n7450), .B(n11824), .ZN(n13518) );
  NAND2_X1 U8073 ( .A1(n13301), .A2(n11823), .ZN(n7450) );
  OR2_X1 U8074 ( .A1(n11703), .A2(n8255), .ZN(n8107) );
  AND2_X1 U8075 ( .A1(n10190), .A2(n6754), .ZN(n13507) );
  NAND2_X1 U8076 ( .A1(n14843), .A2(n10074), .ZN(n13473) );
  CLKBUF_X1 U8077 ( .A(n13392), .Z(n13509) );
  NAND2_X1 U8078 ( .A1(n10792), .A2(n10791), .ZN(n10797) );
  NAND2_X1 U8079 ( .A1(n11348), .A2(n11347), .ZN(n14518) );
  NAND2_X1 U8080 ( .A1(n9821), .A2(n9820), .ZN(n10367) );
  INV_X1 U8081 ( .A(n14475), .ZN(n14504) );
  NAND2_X1 U8082 ( .A1(n6581), .A2(n6647), .ZN(n14275) );
  NAND2_X1 U8083 ( .A1(n7398), .A2(n7402), .ZN(n14066) );
  INV_X1 U8084 ( .A(n14088), .ZN(n6645) );
  NAND2_X1 U8085 ( .A1(n14276), .A2(n14723), .ZN(n6646) );
  NAND2_X1 U8086 ( .A1(n11696), .A2(n11695), .ZN(n14156) );
  OR2_X1 U8087 ( .A1(n11659), .A2(n6686), .ZN(n11662) );
  XNOR2_X1 U8088 ( .A(n8372), .B(n6887), .ZN(n15245) );
  INV_X1 U8089 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6887) );
  XNOR2_X1 U8090 ( .A(n6892), .B(n8376), .ZN(n15243) );
  INV_X1 U8091 ( .A(n8397), .ZN(n7097) );
  XNOR2_X1 U8092 ( .A(n8404), .B(n8405), .ZN(n14533) );
  NAND2_X1 U8093 ( .A1(n8093), .A2(n14847), .ZN(n7669) );
  NAND2_X1 U8094 ( .A1(n6832), .A2(n11843), .ZN(n11856) );
  OAI211_X1 U8095 ( .C1(n11852), .C2(n12026), .A(n7208), .B(n11841), .ZN(n6832) );
  NAND2_X1 U8096 ( .A1(n11863), .A2(n7239), .ZN(n7238) );
  OAI21_X1 U8097 ( .B1(n7493), .B2(n7492), .A(n7491), .ZN(n7724) );
  NAND2_X1 U8098 ( .A1(n6573), .A2(n7707), .ZN(n7491) );
  NOR2_X1 U8099 ( .A1(n6573), .A2(n7707), .ZN(n7493) );
  NAND2_X1 U8100 ( .A1(n11874), .A2(n7213), .ZN(n7212) );
  OR2_X1 U8101 ( .A1(n7745), .A2(n7747), .ZN(n7522) );
  NAND2_X1 U8102 ( .A1(n6831), .A2(n6830), .ZN(n6828) );
  NAND2_X1 U8103 ( .A1(n11905), .A2(n11902), .ZN(n6830) );
  NAND2_X1 U8104 ( .A1(n6589), .A2(n6861), .ZN(n6860) );
  NAND2_X1 U8105 ( .A1(n7518), .A2(n6549), .ZN(n7517) );
  NAND2_X1 U8106 ( .A1(n6658), .A2(n6657), .ZN(n11939) );
  OR2_X1 U8107 ( .A1(n13933), .A2(n11998), .ZN(n6657) );
  NAND2_X1 U8108 ( .A1(n11944), .A2(n11937), .ZN(n6658) );
  NAND2_X1 U8109 ( .A1(n7227), .A2(n11911), .ZN(n7226) );
  INV_X1 U8110 ( .A(n11912), .ZN(n7227) );
  OAI22_X1 U8111 ( .A1(n6523), .A2(n7505), .B1(n7887), .B2(n7506), .ZN(n7905)
         );
  AND2_X1 U8112 ( .A1(n7506), .A2(n7887), .ZN(n7505) );
  INV_X1 U8113 ( .A(n7921), .ZN(n7494) );
  AND2_X1 U8114 ( .A1(n6853), .A2(n6556), .ZN(n6850) );
  NAND2_X1 U8115 ( .A1(n6522), .A2(n6855), .ZN(n6853) );
  NOR2_X1 U8116 ( .A1(n6522), .A2(n6855), .ZN(n6854) );
  NOR2_X1 U8117 ( .A1(n7216), .A2(n11922), .ZN(n7214) );
  INV_X1 U8118 ( .A(n11963), .ZN(n7230) );
  AND2_X1 U8119 ( .A1(n7235), .A2(n11959), .ZN(n7234) );
  INV_X1 U8120 ( .A(n11958), .ZN(n7235) );
  NAND2_X1 U8121 ( .A1(n7233), .A2(n11958), .ZN(n7232) );
  INV_X1 U8122 ( .A(n11959), .ZN(n7233) );
  OAI21_X1 U8123 ( .B1(n11960), .B2(n7234), .A(n6841), .ZN(n11969) );
  NOR2_X1 U8124 ( .A1(n6842), .A2(n11963), .ZN(n6841) );
  INV_X1 U8125 ( .A(n7232), .ZN(n6842) );
  NOR2_X1 U8126 ( .A1(n7997), .A2(n7996), .ZN(n6870) );
  NAND2_X1 U8127 ( .A1(n6580), .A2(n6872), .ZN(n6871) );
  NAND2_X1 U8128 ( .A1(n6873), .A2(n7520), .ZN(n6872) );
  INV_X1 U8129 ( .A(n11977), .ZN(n6659) );
  OAI21_X1 U8130 ( .B1(n7500), .B2(n8034), .A(n7502), .ZN(n8058) );
  NAND2_X1 U8131 ( .A1(n6572), .A2(n7503), .ZN(n7502) );
  OR2_X1 U8132 ( .A1(n8037), .A2(n7501), .ZN(n7500) );
  NOR2_X1 U8133 ( .A1(n11984), .A2(n11981), .ZN(n6845) );
  INV_X1 U8134 ( .A(n11981), .ZN(n6844) );
  NAND2_X1 U8135 ( .A1(n12530), .A2(n6924), .ZN(n12317) );
  INV_X1 U8136 ( .A(n8876), .ZN(n7341) );
  OR4_X1 U8137 ( .A1(n11202), .A2(n11056), .A3(n11198), .A4(n8298), .ZN(n8299)
         );
  NAND2_X1 U8138 ( .A1(n12315), .A2(n12446), .ZN(n6642) );
  NOR2_X1 U8139 ( .A1(n7340), .A2(n7337), .ZN(n7336) );
  INV_X1 U8140 ( .A(n8863), .ZN(n7337) );
  NAND2_X1 U8141 ( .A1(n7042), .A2(n6636), .ZN(n7038) );
  AOI21_X1 U8142 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8097) );
  OR2_X1 U8143 ( .A1(n8118), .A2(n8119), .ZN(n7498) );
  NAND2_X1 U8144 ( .A1(n8118), .A2(n8119), .ZN(n7497) );
  NOR2_X1 U8145 ( .A1(n8246), .A2(n7308), .ZN(n7307) );
  AND2_X1 U8146 ( .A1(n8269), .A2(n8270), .ZN(n7308) );
  AND2_X1 U8147 ( .A1(n10410), .A2(n10093), .ZN(n6995) );
  NAND2_X1 U8148 ( .A1(n14044), .A2(n12031), .ZN(n11836) );
  NOR2_X1 U8149 ( .A1(n8153), .A2(SI_26_), .ZN(n7314) );
  NAND2_X1 U8150 ( .A1(n8153), .A2(SI_26_), .ZN(n7313) );
  INV_X1 U8151 ( .A(n7573), .ZN(n7298) );
  NAND2_X1 U8152 ( .A1(n7574), .A2(n9124), .ZN(n7577) );
  OAI21_X1 U8153 ( .B1(n9517), .B2(n6738), .A(n6737), .ZN(n7550) );
  NAND2_X1 U8154 ( .A1(n9517), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6737) );
  OAI21_X1 U8155 ( .B1(n11682), .B2(n7545), .A(n7544), .ZN(n7547) );
  NAND2_X1 U8156 ( .A1(n11682), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7544) );
  OAI21_X1 U8157 ( .B1(n11682), .B2(n6734), .A(n6733), .ZN(n7541) );
  NAND2_X1 U8158 ( .A1(n11682), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6733) );
  OAI21_X1 U8159 ( .B1(n11682), .B2(n6726), .A(n6725), .ZN(n7538) );
  NAND2_X1 U8160 ( .A1(n11682), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6725) );
  INV_X1 U8161 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U8162 ( .A1(n8343), .A2(n8344), .ZN(n8345) );
  OR2_X1 U8163 ( .A1(n10146), .A2(n7375), .ZN(n7372) );
  INV_X1 U8164 ( .A(n10143), .ZN(n7375) );
  OR2_X1 U8165 ( .A1(n12488), .A2(n12709), .ZN(n7046) );
  NAND2_X1 U8166 ( .A1(n6920), .A2(n6918), .ZN(n6917) );
  NOR2_X1 U8167 ( .A1(n12496), .A2(n6919), .ZN(n6918) );
  INV_X1 U8168 ( .A(n12313), .ZN(n6919) );
  OR2_X1 U8169 ( .A1(n8905), .A2(n8563), .ZN(n8567) );
  NOR2_X1 U8170 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9674), .ZN(n9677) );
  NAND2_X1 U8171 ( .A1(n12753), .A2(n12763), .ZN(n7353) );
  NOR2_X1 U8172 ( .A1(n6924), .A2(n7351), .ZN(n7350) );
  INV_X1 U8173 ( .A(n7353), .ZN(n7351) );
  INV_X1 U8174 ( .A(n8811), .ZN(n7344) );
  NAND2_X1 U8175 ( .A1(n8776), .A2(n8775), .ZN(n8792) );
  INV_X1 U8176 ( .A(n8691), .ZN(n7335) );
  INV_X1 U8177 ( .A(n7065), .ZN(n7064) );
  INV_X1 U8178 ( .A(n12360), .ZN(n7066) );
  INV_X1 U8179 ( .A(n10112), .ZN(n12514) );
  NAND2_X1 U8180 ( .A1(n7049), .A2(n6924), .ZN(n6923) );
  OR2_X1 U8181 ( .A1(n12975), .A2(n12292), .ZN(n12325) );
  INV_X1 U8182 ( .A(n12434), .ZN(n7321) );
  INV_X1 U8183 ( .A(n12435), .ZN(n7317) );
  INV_X1 U8184 ( .A(n12538), .ZN(n9978) );
  NOR2_X1 U8185 ( .A1(n7038), .A2(n7030), .ZN(n7029) );
  INV_X1 U8186 ( .A(n8506), .ZN(n7030) );
  OR2_X1 U8187 ( .A1(n7039), .A2(n7038), .ZN(n7037) );
  NAND2_X1 U8188 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10950), .ZN(n8495) );
  NAND2_X1 U8189 ( .A1(n6940), .A2(n7015), .ZN(n8488) );
  AOI21_X1 U8190 ( .B1(n7018), .B2(n7019), .A(n7016), .ZN(n7015) );
  NOR2_X1 U8191 ( .A1(n9314), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7016) );
  XNOR2_X1 U8192 ( .A(n11612), .B(n13081), .ZN(n10047) );
  AOI21_X1 U8193 ( .B1(n8307), .B2(n8306), .A(n6754), .ZN(n6689) );
  NAND2_X1 U8194 ( .A1(n8304), .A2(n6663), .ZN(n8312) );
  NOR2_X1 U8195 ( .A1(n11824), .A2(n6664), .ZN(n6663) );
  OAI211_X1 U8196 ( .C1(n8306), .C2(n8307), .A(n6524), .B(n6665), .ZN(n6664)
         );
  INV_X1 U8197 ( .A(n13630), .ZN(n7653) );
  INV_X1 U8198 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n15187) );
  INV_X1 U8199 ( .A(n11796), .ZN(n7152) );
  INV_X1 U8200 ( .A(n11795), .ZN(n7149) );
  INV_X1 U8201 ( .A(n13431), .ZN(n7175) );
  OR2_X1 U8202 ( .A1(n13468), .A2(n11790), .ZN(n7177) );
  INV_X1 U8203 ( .A(n13486), .ZN(n6720) );
  OR2_X1 U8204 ( .A1(n7822), .A2(n7821), .ZN(n7837) );
  NAND2_X1 U8205 ( .A1(n6994), .A2(n6995), .ZN(n6996) );
  NOR2_X1 U8206 ( .A1(n14868), .A2(n10567), .ZN(n6994) );
  INV_X1 U8207 ( .A(n10265), .ZN(n7430) );
  INV_X1 U8208 ( .A(n9943), .ZN(n7428) );
  NAND2_X1 U8209 ( .A1(n8292), .A2(n10377), .ZN(n9488) );
  NOR2_X1 U8210 ( .A1(n13421), .A2(n13557), .ZN(n13399) );
  NAND2_X1 U8211 ( .A1(n6489), .A2(n7439), .ZN(n13421) );
  NAND2_X1 U8212 ( .A1(n7011), .A2(n7008), .ZN(n11417) );
  NAND2_X1 U8213 ( .A1(n10403), .A2(n9943), .ZN(n9945) );
  INV_X1 U8214 ( .A(n6993), .ZN(n10280) );
  NOR2_X2 U8215 ( .A1(n10407), .A2(n10406), .ZN(n10410) );
  XNOR2_X1 U8216 ( .A(n7621), .B(n7646), .ZN(n8336) );
  OAI21_X1 U8217 ( .B1(n6998), .B2(n7001), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7621) );
  AND2_X1 U8218 ( .A1(n7629), .A2(n8318), .ZN(n8322) );
  NOR2_X1 U8219 ( .A1(n7628), .A2(n7629), .ZN(n7668) );
  NAND2_X1 U8220 ( .A1(n6680), .A2(n6679), .ZN(n7628) );
  NAND2_X1 U8221 ( .A1(n6681), .A2(n7709), .ZN(n6679) );
  AND2_X1 U8222 ( .A1(n13923), .A2(n10452), .ZN(n7276) );
  AND2_X1 U8223 ( .A1(n11350), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11431) );
  INV_X1 U8224 ( .A(n11845), .ZN(n9510) );
  NOR2_X1 U8225 ( .A1(n7279), .A2(n6793), .ZN(n6792) );
  INV_X1 U8226 ( .A(n10791), .ZN(n6793) );
  INV_X1 U8227 ( .A(n7280), .ZN(n7279) );
  INV_X1 U8228 ( .A(n10796), .ZN(n7278) );
  NAND2_X1 U8229 ( .A1(n6792), .A2(n6795), .ZN(n6790) );
  INV_X1 U8230 ( .A(n13760), .ZN(n6802) );
  NAND2_X1 U8231 ( .A1(n7219), .A2(n11997), .ZN(n7217) );
  OR2_X1 U8232 ( .A1(n11656), .A2(n14744), .ZN(n9293) );
  INV_X1 U8233 ( .A(n11671), .ZN(n7133) );
  AND2_X1 U8234 ( .A1(n11663), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11675) );
  OR2_X1 U8235 ( .A1(n14340), .A2(n13681), .ZN(n11761) );
  INV_X1 U8236 ( .A(n6837), .ZN(n6836) );
  NOR2_X1 U8237 ( .A1(n11352), .A2(n11351), .ZN(n11350) );
  OR2_X1 U8238 ( .A1(n14424), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U8239 ( .A1(n11913), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U8240 ( .A1(n10513), .A2(n11865), .ZN(n10649) );
  AND2_X1 U8241 ( .A1(n12019), .A2(n12030), .ZN(n11845) );
  NAND2_X1 U8242 ( .A1(n7392), .A2(n7393), .ZN(n11429) );
  AOI21_X1 U8243 ( .B1(n7395), .B2(n7397), .A(n6566), .ZN(n7393) );
  AND3_X2 U8244 ( .A1(n9522), .A2(n9521), .A3(n9520), .ZN(n11544) );
  NAND2_X1 U8245 ( .A1(n7272), .A2(n9287), .ZN(n9149) );
  INV_X1 U8246 ( .A(SI_22_), .ZN(n6982) );
  INV_X1 U8247 ( .A(n9149), .ZN(n6818) );
  INV_X1 U8248 ( .A(n7290), .ZN(n7289) );
  OAI21_X1 U8249 ( .B1(n7594), .B2(n6610), .A(n7602), .ZN(n7290) );
  OR2_X1 U8250 ( .A1(n7595), .A2(n6610), .ZN(n7291) );
  NAND2_X1 U8251 ( .A1(n6948), .A2(n6947), .ZN(n7998) );
  AOI22_X1 U8252 ( .A1(n6950), .A2(n6957), .B1(n6953), .B2(n6955), .ZN(n6947)
         );
  OR2_X1 U8253 ( .A1(n6950), .A2(n6953), .ZN(n6949) );
  AND2_X1 U8254 ( .A1(n6815), .A2(n7526), .ZN(n6813) );
  NAND2_X1 U8255 ( .A1(n7288), .A2(n7287), .ZN(n7603) );
  AOI21_X1 U8256 ( .B1(n7594), .B2(n7595), .A(n6610), .ZN(n7287) );
  NAND2_X1 U8257 ( .A1(n7998), .A2(n7594), .ZN(n7288) );
  NAND2_X1 U8258 ( .A1(n15253), .A2(n7240), .ZN(n7244) );
  AND2_X1 U8259 ( .A1(n9288), .A2(n7245), .ZN(n7240) );
  INV_X1 U8260 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7245) );
  INV_X1 U8261 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9288) );
  NOR2_X1 U8262 ( .A1(n7303), .A2(n15172), .ZN(n7302) );
  INV_X1 U8263 ( .A(n7301), .ZN(n7300) );
  AND2_X1 U8264 ( .A1(n7587), .A2(n7586), .ZN(n7939) );
  NAND2_X1 U8265 ( .A1(n7573), .A2(n7571), .ZN(n7867) );
  INV_X1 U8266 ( .A(n7852), .ZN(n7565) );
  OR2_X1 U8267 ( .A1(n7868), .A2(n7867), .ZN(n7870) );
  XNOR2_X1 U8268 ( .A(n7562), .B(SI_9_), .ZN(n7831) );
  INV_X1 U8269 ( .A(n7559), .ZN(n6963) );
  AND2_X1 U8270 ( .A1(n9051), .A2(n9052), .ZN(n7410) );
  INV_X1 U8271 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U8272 ( .A1(n11682), .A2(n9069), .ZN(n6739) );
  NAND2_X1 U8273 ( .A1(n8354), .A2(n8353), .ZN(n8365) );
  OR2_X1 U8274 ( .A1(n8388), .A2(n9237), .ZN(n8353) );
  AND2_X1 U8275 ( .A1(n12192), .A2(n7363), .ZN(n7362) );
  NOR2_X1 U8276 ( .A1(n7360), .A2(n6542), .ZN(n7358) );
  NOR2_X1 U8277 ( .A1(n6518), .A2(n7361), .ZN(n7360) );
  INV_X1 U8278 ( .A(n12192), .ZN(n7361) );
  NOR2_X1 U8279 ( .A1(n8892), .A2(n8463), .ZN(n8523) );
  INV_X1 U8280 ( .A(n12746), .ZN(n12197) );
  XNOR2_X1 U8281 ( .A(n12153), .B(n6914), .ZN(n10163) );
  NAND2_X1 U8282 ( .A1(n10155), .A2(n7374), .ZN(n10166) );
  INV_X1 U8283 ( .A(n7372), .ZN(n7374) );
  NAND2_X1 U8284 ( .A1(n6907), .A2(n6905), .ZN(n11368) );
  AND2_X1 U8285 ( .A1(n6626), .A2(n6906), .ZN(n6905) );
  INV_X1 U8286 ( .A(n10165), .ZN(n7373) );
  NAND2_X1 U8287 ( .A1(n12151), .A2(n6901), .ZN(n6896) );
  AND4_X1 U8288 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .ZN(n8926)
         );
  NOR2_X1 U8289 ( .A1(n9749), .A2(n9733), .ZN(n9735) );
  INV_X1 U8290 ( .A(n6669), .ZN(n9732) );
  NOR2_X1 U8291 ( .A1(n9878), .A2(n9879), .ZN(n9882) );
  NAND2_X1 U8292 ( .A1(n7189), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7188) );
  INV_X1 U8293 ( .A(n10495), .ZN(n7189) );
  NOR2_X1 U8294 ( .A1(n10323), .A2(n10309), .ZN(n10492) );
  NOR2_X1 U8295 ( .A1(n14903), .A2(n14902), .ZN(n14901) );
  INV_X1 U8296 ( .A(n14900), .ZN(n11188) );
  NOR3_X1 U8297 ( .A1(n14920), .A2(n14919), .A3(n14923), .ZN(n14921) );
  NOR2_X1 U8298 ( .A1(n12632), .A2(n12631), .ZN(n12643) );
  AND2_X1 U8299 ( .A1(n8523), .A2(n12196), .ZN(n12706) );
  INV_X1 U8300 ( .A(n12530), .ZN(n12723) );
  NAND2_X1 U8301 ( .A1(n7051), .A2(n6509), .ZN(n7050) );
  NAND2_X1 U8302 ( .A1(n6946), .A2(n12453), .ZN(n7051) );
  AND2_X1 U8303 ( .A1(n12975), .A2(n12778), .ZN(n6638) );
  OR2_X1 U8304 ( .A1(n8880), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U8305 ( .A1(n8869), .A2(n15199), .ZN(n8880) );
  INV_X1 U8306 ( .A(n12764), .ZN(n12791) );
  AND2_X1 U8307 ( .A1(n8868), .A2(n8867), .ZN(n12154) );
  AND2_X1 U8308 ( .A1(n8856), .A2(n12273), .ZN(n8869) );
  OR2_X1 U8309 ( .A1(n8833), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8845) );
  NOR2_X1 U8310 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(n8805), .ZN(n8821) );
  AND2_X1 U8311 ( .A1(n8746), .A2(n12169), .ZN(n8762) );
  NOR2_X1 U8312 ( .A1(n8729), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8746) );
  OR3_X1 U8313 ( .A1(n8707), .A2(P3_REG3_REG_12__SCAN_IN), .A3(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8729) );
  AND2_X1 U8314 ( .A1(n8663), .A2(n8462), .ZN(n8677) );
  INV_X1 U8315 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n8676) );
  AND2_X1 U8316 ( .A1(n8675), .A2(n12388), .ZN(n12368) );
  AND4_X1 U8317 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n10986)
         );
  NAND2_X1 U8318 ( .A1(n7345), .A2(n6693), .ZN(n10843) );
  NAND2_X1 U8319 ( .A1(n7347), .A2(n8621), .ZN(n6693) );
  NOR2_X1 U8320 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8605) );
  AND3_X1 U8321 ( .A1(n8590), .A2(n8589), .A3(n8588), .ZN(n10216) );
  AOI21_X1 U8322 ( .B1(n14941), .B2(n14942), .A(n6530), .ZN(n7523) );
  NAND2_X1 U8323 ( .A1(n12468), .A2(n12467), .ZN(n14438) );
  OR2_X1 U8324 ( .A1(n7050), .A2(n12314), .ZN(n6920) );
  NAND2_X1 U8325 ( .A1(n8903), .A2(n8902), .ZN(n9036) );
  AOI21_X1 U8326 ( .B1(n7057), .B2(n7060), .A(n7055), .ZN(n7054) );
  INV_X1 U8327 ( .A(n8997), .ZN(n7060) );
  INV_X1 U8328 ( .A(n7068), .ZN(n7067) );
  OAI21_X1 U8329 ( .B1(n6506), .B2(n7069), .A(n12429), .ZN(n7068) );
  INV_X1 U8330 ( .A(n12420), .ZN(n7069) );
  INV_X1 U8331 ( .A(n15004), .ZN(n15001) );
  AOI21_X1 U8332 ( .B1(n8901), .B2(n8900), .A(n8899), .ZN(n12111) );
  AND2_X1 U8333 ( .A1(n14374), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8899) );
  AND2_X1 U8334 ( .A1(n7078), .A2(n8452), .ZN(n6760) );
  NAND2_X1 U8335 ( .A1(n8949), .A2(n6702), .ZN(n6701) );
  NAND2_X1 U8336 ( .A1(n13044), .A2(n6703), .ZN(n6702) );
  AND2_X1 U8337 ( .A1(n10953), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6926) );
  INV_X1 U8338 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U8339 ( .A1(n8494), .A2(n7014), .ZN(n8800) );
  NAND2_X1 U8340 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n10304), .ZN(n7014) );
  NAND2_X1 U8341 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U8342 ( .A1(n8483), .A2(n8482), .ZN(n8684) );
  AOI21_X1 U8343 ( .B1(n6936), .B2(n6938), .A(n6935), .ZN(n6934) );
  XNOR2_X1 U8344 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8683) );
  OR2_X1 U8345 ( .A1(n8653), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8654) );
  NOR2_X1 U8346 ( .A1(n8654), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8686) );
  AOI21_X1 U8347 ( .B1(n6930), .B2(n6932), .A(n6575), .ZN(n6928) );
  NAND2_X1 U8348 ( .A1(n8442), .A2(n8441), .ZN(n8613) );
  NAND2_X1 U8349 ( .A1(n9132), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8473) );
  XNOR2_X1 U8350 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8582) );
  XNOR2_X1 U8351 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8571) );
  INV_X1 U8352 ( .A(n10103), .ZN(n7477) );
  OR2_X1 U8353 ( .A1(n7465), .A2(n13097), .ZN(n7460) );
  NAND2_X1 U8354 ( .A1(n7466), .A2(n11607), .ZN(n7465) );
  AOI21_X1 U8355 ( .B1(n7466), .B2(n7463), .A(n7462), .ZN(n7461) );
  NOR2_X1 U8356 ( .A1(n11610), .A2(n11609), .ZN(n7462) );
  NOR2_X1 U8357 ( .A1(n7467), .A2(n7464), .ZN(n7463) );
  NAND2_X1 U8358 ( .A1(n9515), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U8359 ( .A1(n9516), .A2(n7164), .ZN(n7163) );
  INV_X1 U8360 ( .A(n7947), .ZN(n7640) );
  OR2_X1 U8361 ( .A1(n11569), .A2(n11570), .ZN(n7489) );
  NAND2_X1 U8362 ( .A1(n7641), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7990) );
  INV_X1 U8363 ( .A(n7971), .ZN(n7641) );
  INV_X1 U8364 ( .A(n8086), .ZN(n8085) );
  AOI21_X1 U8365 ( .B1(n11596), .B2(n7471), .A(n6614), .ZN(n13123) );
  NAND2_X1 U8366 ( .A1(n7473), .A2(n7472), .ZN(n7471) );
  INV_X1 U8367 ( .A(n13066), .ZN(n7472) );
  NAND2_X1 U8368 ( .A1(n13492), .A2(n6667), .ZN(n10376) );
  NAND2_X1 U8369 ( .A1(n7643), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8046) );
  INV_X1 U8370 ( .A(n8044), .ZN(n7643) );
  OR2_X1 U8371 ( .A1(n7990), .A2(n13118), .ZN(n8006) );
  NAND2_X1 U8372 ( .A1(n11602), .A2(n11603), .ZN(n7470) );
  NOR2_X1 U8373 ( .A1(n8248), .A2(n7499), .ZN(n7309) );
  INV_X1 U8374 ( .A(n8274), .ZN(n8277) );
  NOR2_X1 U8375 ( .A1(n9384), .A2(n6677), .ZN(n14765) );
  NOR2_X1 U8376 ( .A1(n14765), .A2(n14764), .ZN(n14763) );
  AOI21_X1 U8377 ( .B1(n9352), .B2(P2_REG1_REG_4__SCAN_IN), .A(n9551), .ZN(
        n9369) );
  OAI21_X1 U8378 ( .B1(n9403), .B2(n9343), .A(n9342), .ZN(n9414) );
  AOI21_X1 U8379 ( .B1(n9444), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9439), .ZN(
        n9441) );
  NAND2_X1 U8380 ( .A1(n7139), .A2(n7145), .ZN(n6675) );
  NAND2_X1 U8381 ( .A1(n7136), .A2(n7138), .ZN(n6674) );
  INV_X1 U8382 ( .A(n11824), .ZN(n11798) );
  NAND2_X1 U8383 ( .A1(n13524), .A2(n11822), .ZN(n13302) );
  NAND2_X1 U8384 ( .A1(n13526), .A2(n13191), .ZN(n11822) );
  NAND2_X1 U8385 ( .A1(n7003), .A2(n11821), .ZN(n13322) );
  INV_X1 U8386 ( .A(n7003), .ZN(n13338) );
  AND2_X1 U8387 ( .A1(n8204), .A2(n8142), .ZN(n13324) );
  OAI22_X1 U8388 ( .A1(n13345), .A2(n13344), .B1(n13352), .B2(n13193), .ZN(
        n13330) );
  AND2_X1 U8389 ( .A1(n13369), .A2(n13377), .ZN(n6685) );
  AOI22_X1 U8390 ( .A1(n13358), .A2(n13363), .B1(n13099), .B2(n13369), .ZN(
        n13345) );
  NAND2_X1 U8391 ( .A1(n13381), .A2(n6722), .ZN(n13358) );
  NAND2_X1 U8392 ( .A1(n13388), .A2(n13126), .ZN(n6722) );
  OAI21_X1 U8393 ( .B1(n13414), .B2(n7150), .A(n7148), .ZN(n13379) );
  INV_X1 U8394 ( .A(n7151), .ZN(n7150) );
  AOI21_X1 U8395 ( .B1(n7151), .B2(n7149), .A(n6564), .ZN(n7148) );
  NOR2_X1 U8396 ( .A1(n13393), .A2(n7152), .ZN(n7151) );
  NAND2_X1 U8397 ( .A1(n6724), .A2(n6723), .ZN(n13381) );
  INV_X1 U8398 ( .A(n13379), .ZN(n6724) );
  NOR2_X1 U8399 ( .A1(n6723), .A2(n7432), .ZN(n7431) );
  INV_X1 U8400 ( .A(n7434), .ZN(n7432) );
  NOR2_X1 U8401 ( .A1(n13405), .A2(n7436), .ZN(n7435) );
  INV_X1 U8402 ( .A(n7438), .ZN(n7436) );
  NAND2_X1 U8403 ( .A1(n7005), .A2(n7004), .ZN(n13427) );
  NAND2_X1 U8404 ( .A1(n8289), .A2(n13431), .ZN(n13449) );
  NAND2_X1 U8405 ( .A1(n7177), .A2(n11791), .ZN(n13450) );
  NAND2_X1 U8406 ( .A1(n7177), .A2(n6516), .ZN(n13453) );
  INV_X1 U8407 ( .A(n7007), .ZN(n13466) );
  INV_X1 U8408 ( .A(n11497), .ZN(n11811) );
  AOI21_X1 U8409 ( .B1(n7106), .B2(n7108), .A(n6563), .ZN(n7104) );
  INV_X1 U8410 ( .A(n11483), .ZN(n11492) );
  NAND2_X1 U8411 ( .A1(n7639), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7930) );
  INV_X1 U8412 ( .A(n7010), .ZN(n11210) );
  OAI21_X1 U8413 ( .B1(n10817), .B2(n7156), .A(n7154), .ZN(n11204) );
  INV_X1 U8414 ( .A(n7157), .ZN(n7156) );
  AND2_X1 U8415 ( .A1(n11097), .A2(n7155), .ZN(n7154) );
  OR2_X1 U8416 ( .A1(n10694), .A2(n10927), .ZN(n10821) );
  NOR2_X2 U8417 ( .A1(n10821), .A2(n11062), .ZN(n11070) );
  NAND2_X1 U8418 ( .A1(n10812), .A2(n10811), .ZN(n11057) );
  NOR2_X2 U8419 ( .A1(n6996), .A2(n14878), .ZN(n10592) );
  NAND2_X1 U8420 ( .A1(n6993), .A2(n6997), .ZN(n10532) );
  INV_X1 U8421 ( .A(n9488), .ZN(n10044) );
  NAND2_X1 U8422 ( .A1(n7437), .A2(n7438), .ZN(n13406) );
  NAND2_X1 U8423 ( .A1(n13503), .A2(n11813), .ZN(n13479) );
  AOI22_X1 U8424 ( .A1(n13435), .A2(n6667), .B1(n13212), .B2(n13437), .ZN(
        n9502) );
  AND2_X1 U8425 ( .A1(n8305), .A2(n8263), .ZN(n14855) );
  AND2_X1 U8426 ( .A1(n9472), .A2(n9471), .ZN(n14838) );
  XNOR2_X1 U8427 ( .A(n7623), .B(n7622), .ZN(n11800) );
  NAND2_X1 U8428 ( .A1(n8324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7623) );
  OR2_X1 U8429 ( .A1(n8326), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8328) );
  OR2_X1 U8430 ( .A1(n7629), .A2(n7709), .ZN(n6875) );
  BUF_X1 U8431 ( .A(n7668), .Z(n9497) );
  INV_X1 U8432 ( .A(n11500), .ZN(n13472) );
  INV_X1 U8433 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7984) );
  OR3_X1 U8434 ( .A1(n7813), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_6__SCAN_IN), .ZN(n7815) );
  AND2_X1 U8435 ( .A1(n7714), .A2(n7732), .ZN(n9351) );
  NOR2_X1 U8436 ( .A1(n10975), .A2(n7281), .ZN(n7280) );
  INV_X1 U8437 ( .A(n10972), .ZN(n7281) );
  NAND2_X1 U8438 ( .A1(n9514), .A2(n9513), .ZN(n7283) );
  INV_X1 U8439 ( .A(n13826), .ZN(n6806) );
  INV_X1 U8440 ( .A(n6807), .ZN(n6803) );
  NAND2_X1 U8441 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  OR2_X1 U8442 ( .A1(n13908), .A2(n13834), .ZN(n7270) );
  NAND2_X1 U8443 ( .A1(n6804), .A2(n6808), .ZN(n13825) );
  INV_X1 U8444 ( .A(n6810), .ZN(n6801) );
  NAND2_X1 U8445 ( .A1(n7254), .A2(n7252), .ZN(n13859) );
  OAI21_X1 U8446 ( .B1(n7249), .B2(n6791), .A(n6789), .ZN(n11451) );
  INV_X1 U8447 ( .A(n6792), .ZN(n6791) );
  AND2_X1 U8448 ( .A1(n6790), .A2(n7277), .ZN(n6789) );
  AOI21_X1 U8449 ( .B1(n7280), .B2(n7278), .A(n6548), .ZN(n7277) );
  NAND2_X1 U8450 ( .A1(n10452), .A2(n11844), .ZN(n9262) );
  AOI21_X1 U8451 ( .B1(n7262), .B2(n7260), .A(n13720), .ZN(n7259) );
  INV_X1 U8452 ( .A(n13865), .ZN(n7260) );
  INV_X1 U8453 ( .A(n7262), .ZN(n7261) );
  OR2_X1 U8454 ( .A1(n10734), .A2(n10733), .ZN(n10891) );
  NOR2_X1 U8455 ( .A1(n10891), .A2(n10890), .ZN(n11037) );
  NAND2_X1 U8456 ( .A1(n7282), .A2(n7283), .ZN(n9804) );
  INV_X1 U8457 ( .A(n9535), .ZN(n7282) );
  INV_X1 U8458 ( .A(n10658), .ZN(n7251) );
  INV_X1 U8459 ( .A(n11743), .ZN(n11720) );
  AND4_X1 U8460 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(n11866)
         );
  INV_X1 U8461 ( .A(n7529), .ZN(n11653) );
  NAND2_X1 U8462 ( .A1(n11562), .A2(n14373), .ZN(n7529) );
  AOI21_X1 U8463 ( .B1(n10629), .B2(P1_REG2_REG_7__SCAN_IN), .A(n9325), .ZN(
        n9327) );
  AOI21_X1 U8464 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n10878), .A(n10353), .ZN(
        n10355) );
  AOI21_X1 U8465 ( .B1(n11034), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10539), .ZN(
        n10543) );
  NAND2_X1 U8466 ( .A1(n14557), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6728) );
  AND2_X1 U8467 ( .A1(n14564), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6730) );
  INV_X1 U8468 ( .A(n7169), .ZN(n7167) );
  NAND2_X1 U8469 ( .A1(n14270), .A2(n13923), .ZN(n7171) );
  NOR2_X1 U8470 ( .A1(n14070), .A2(n7170), .ZN(n7169) );
  INV_X1 U8471 ( .A(n11748), .ZN(n7170) );
  XNOR2_X1 U8472 ( .A(n14270), .B(n13923), .ZN(n14070) );
  AND2_X1 U8473 ( .A1(n11740), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11742) );
  INV_X1 U8474 ( .A(n7205), .ZN(n14117) );
  AOI21_X1 U8475 ( .B1(n14150), .B2(n7409), .A(n6559), .ZN(n7408) );
  INV_X1 U8476 ( .A(n11768), .ZN(n7409) );
  INV_X1 U8477 ( .A(n7207), .ZN(n14152) );
  INV_X1 U8478 ( .A(n7132), .ZN(n7131) );
  AOI21_X1 U8479 ( .B1(n7132), .B2(n7130), .A(n6571), .ZN(n7129) );
  NOR2_X1 U8480 ( .A1(n14181), .A2(n7133), .ZN(n7132) );
  AND2_X1 U8481 ( .A1(n9542), .A2(n14376), .ZN(n13898) );
  OR2_X1 U8482 ( .A1(n11518), .A2(n9172), .ZN(n11650) );
  INV_X1 U8483 ( .A(n7202), .ZN(n14230) );
  INV_X1 U8484 ( .A(n7127), .ZN(n7126) );
  AOI21_X1 U8485 ( .B1(n7127), .B2(n7125), .A(n6565), .ZN(n7124) );
  INV_X1 U8486 ( .A(n12083), .ZN(n7125) );
  NOR2_X1 U8487 ( .A1(n12083), .A2(n7423), .ZN(n7422) );
  INV_X1 U8488 ( .A(n11934), .ZN(n7423) );
  NOR2_X1 U8489 ( .A1(n11527), .A2(n13839), .ZN(n14245) );
  OR3_X1 U8490 ( .A1(n11150), .A2(n11149), .A3(n11148), .ZN(n11352) );
  NAND2_X1 U8491 ( .A1(n6745), .A2(n6744), .ZN(n11527) );
  INV_X1 U8492 ( .A(n11440), .ZN(n6745) );
  NAND2_X1 U8493 ( .A1(n6747), .A2(n6746), .ZN(n11440) );
  NOR2_X1 U8494 ( .A1(n7198), .A2(n14518), .ZN(n6747) );
  INV_X1 U8495 ( .A(n11047), .ZN(n6746) );
  NAND2_X1 U8496 ( .A1(n11037), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11150) );
  NOR3_X1 U8497 ( .A1(n11047), .A2(n14424), .A3(n14503), .ZN(n11160) );
  NOR2_X1 U8498 ( .A1(n11047), .A2(n14503), .ZN(n11127) );
  NAND2_X1 U8499 ( .A1(n10880), .A2(n10879), .ZN(n14471) );
  AOI21_X1 U8500 ( .B1(n6505), .B2(n10756), .A(n6533), .ZN(n7418) );
  AND2_X1 U8501 ( .A1(n7112), .A2(n10712), .ZN(n7110) );
  NAND2_X1 U8502 ( .A1(n7421), .A2(n10729), .ZN(n10730) );
  NAND2_X1 U8503 ( .A1(n7421), .A2(n6505), .ZN(n10882) );
  AND2_X1 U8504 ( .A1(n10457), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U8505 ( .A1(n7203), .A2(n10236), .ZN(n10034) );
  INV_X1 U8506 ( .A(n11549), .ZN(n6749) );
  OR2_X1 U8507 ( .A1(n11844), .A2(n14660), .ZN(n12061) );
  AND2_X1 U8508 ( .A1(n12015), .A2(n12014), .ZN(n14261) );
  AND3_X1 U8509 ( .A1(n7401), .A2(n7399), .A3(n6601), .ZN(n11780) );
  INV_X1 U8510 ( .A(n14691), .ZN(n14698) );
  INV_X1 U8511 ( .A(n10236), .ZN(n11857) );
  OR2_X1 U8512 ( .A1(n12011), .A2(n7524), .ZN(n9577) );
  OR3_X1 U8513 ( .A1(n8250), .A2(n8184), .A3(n8182), .ZN(n8193) );
  AND2_X1 U8514 ( .A1(n6541), .A2(n6820), .ZN(n6826) );
  NAND2_X1 U8515 ( .A1(n8235), .A2(n8250), .ZN(n13629) );
  AND2_X1 U8516 ( .A1(n9061), .A2(n9062), .ZN(n7415) );
  AND3_X1 U8517 ( .A1(n7274), .A2(n9056), .A3(n6827), .ZN(n9061) );
  INV_X1 U8518 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8519 ( .A1(n6816), .A2(n6819), .ZN(n12031) );
  NOR2_X1 U8520 ( .A1(n6818), .A2(n6817), .ZN(n6816) );
  OAI21_X1 U8521 ( .B1(n9150), .B2(P1_IR_REG_21__SCAN_IN), .A(n6576), .ZN(
        n6819) );
  NOR2_X1 U8522 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6817) );
  NAND2_X1 U8523 ( .A1(n9287), .A2(n7243), .ZN(n10805) );
  INV_X1 U8524 ( .A(n7244), .ZN(n7243) );
  NAND2_X1 U8525 ( .A1(n9287), .A2(n7246), .ZN(n10301) );
  AND2_X1 U8526 ( .A1(n15253), .A2(n9288), .ZN(n7246) );
  NAND2_X1 U8527 ( .A1(n7304), .A2(n7305), .ZN(n7925) );
  NAND2_X1 U8528 ( .A1(n7582), .A2(n6502), .ZN(n7305) );
  NAND2_X1 U8529 ( .A1(n7299), .A2(n15172), .ZN(n7304) );
  NAND2_X1 U8530 ( .A1(n6961), .A2(n7559), .ZN(n7812) );
  INV_X1 U8531 ( .A(n7788), .ZN(n7557) );
  OR2_X1 U8532 ( .A1(n9112), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9139) );
  INV_X1 U8533 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U8534 ( .A1(n9092), .A2(n9051), .ZN(n9107) );
  NAND2_X1 U8535 ( .A1(n8341), .A2(n7094), .ZN(n8369) );
  NAND2_X1 U8536 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7095), .ZN(n7094) );
  XNOR2_X1 U8537 ( .A(n8366), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n8367) );
  INV_X1 U8538 ( .A(n6895), .ZN(n8384) );
  OAI21_X1 U8539 ( .B1(n15238), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6562), .ZN(
        n6895) );
  NAND2_X1 U8540 ( .A1(n8349), .A2(n8348), .ZN(n8386) );
  NAND2_X1 U8541 ( .A1(n8381), .A2(n9306), .ZN(n8348) );
  OAI21_X1 U8542 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n8358), .A(n8357), .ZN(
        n8400) );
  OAI22_X1 U8543 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14915), .B1(n8407), .B2(
        n8406), .ZN(n8412) );
  NAND2_X1 U8544 ( .A1(n6884), .A2(n6883), .ZN(n8421) );
  INV_X1 U8545 ( .A(n14543), .ZN(n6883) );
  OR2_X1 U8546 ( .A1(n14542), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8547 ( .A1(n7359), .A2(n6518), .ZN(n12193) );
  OR2_X1 U8548 ( .A1(n10942), .A2(n10943), .ZN(n11081) );
  NAND2_X1 U8549 ( .A1(n11081), .A2(n6908), .ZN(n11327) );
  INV_X1 U8550 ( .A(n10216), .ZN(n14965) );
  NAND2_X1 U8551 ( .A1(n12281), .A2(n12139), .ZN(n12184) );
  OAI21_X1 U8552 ( .B1(n7366), .B2(n7358), .A(n7356), .ZN(n7355) );
  OAI21_X1 U8553 ( .B1(n7366), .B2(n7362), .A(n7358), .ZN(n7356) );
  NAND2_X1 U8554 ( .A1(n7358), .A2(n12195), .ZN(n7357) );
  NAND2_X1 U8555 ( .A1(n7378), .A2(n8559), .ZN(n10129) );
  INV_X1 U8556 ( .A(n9982), .ZN(n7378) );
  NAND2_X1 U8557 ( .A1(n8574), .A2(n9079), .ZN(n8540) );
  AND4_X1 U8558 ( .A1(n8697), .A2(n8696), .A3(n8695), .A4(n8694), .ZN(n12380)
         );
  AND2_X1 U8559 ( .A1(n12223), .A2(n12130), .ZN(n7380) );
  AND2_X1 U8560 ( .A1(n7381), .A2(n12130), .ZN(n12224) );
  NAND2_X1 U8561 ( .A1(n10166), .A2(n10165), .ZN(n10288) );
  NAND2_X1 U8562 ( .A1(n10155), .A2(n10143), .ZN(n10145) );
  NOR2_X1 U8563 ( .A1(n12251), .A2(n6910), .ZN(n6909) );
  INV_X1 U8564 ( .A(n12142), .ZN(n6910) );
  NAND2_X1 U8565 ( .A1(n12182), .A2(n12142), .ZN(n12252) );
  NAND2_X1 U8566 ( .A1(n9977), .A2(n9976), .ZN(n12257) );
  INV_X1 U8567 ( .A(n10294), .ZN(n6731) );
  NAND2_X1 U8568 ( .A1(n12127), .A2(n12126), .ZN(n12302) );
  NOR2_X1 U8569 ( .A1(n6698), .A2(n6641), .ZN(n6640) );
  NOR2_X1 U8570 ( .A1(n6699), .A2(n14938), .ZN(n6698) );
  INV_X1 U8571 ( .A(n12541), .ZN(n6699) );
  OAI21_X1 U8572 ( .B1(n12541), .B2(n12490), .A(n6697), .ZN(n6696) );
  OR2_X1 U8573 ( .A1(n12537), .A2(n12538), .ZN(n6697) );
  INV_X1 U8574 ( .A(n12851), .ZN(n12552) );
  INV_X1 U8575 ( .A(n12264), .ZN(n12553) );
  INV_X1 U8576 ( .A(n12380), .ZN(n12554) );
  INV_X1 U8577 ( .A(n11085), .ZN(n12556) );
  CLKBUF_X1 U8578 ( .A(n12563), .Z(n6655) );
  OR2_X1 U8579 ( .A1(n12481), .A2(n8548), .ZN(n8554) );
  INV_X1 U8580 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U8581 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n8548), .ZN(n10207) );
  NOR2_X1 U8582 ( .A1(n10199), .A2(n9673), .ZN(n9892) );
  AOI21_X1 U8583 ( .B1(n9890), .B2(n9658), .A(n9657), .ZN(n10010) );
  INV_X1 U8584 ( .A(n6768), .ZN(n10013) );
  INV_X1 U8585 ( .A(n7179), .ZN(n9844) );
  AOI21_X1 U8586 ( .B1(n10007), .B2(n9840), .A(n9839), .ZN(n9842) );
  INV_X1 U8587 ( .A(n7186), .ZN(n9701) );
  INV_X1 U8588 ( .A(n6767), .ZN(n9858) );
  AOI21_X1 U8589 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n10315) );
  INV_X1 U8590 ( .A(n6650), .ZN(n10473) );
  INV_X1 U8591 ( .A(n10475), .ZN(n7080) );
  INV_X1 U8592 ( .A(n7081), .ZN(n10476) );
  INV_X1 U8593 ( .A(n11177), .ZN(n6670) );
  OR2_X1 U8594 ( .A1(n12575), .A2(n12572), .ZN(n7184) );
  NOR2_X1 U8595 ( .A1(n14925), .A2(n8731), .ZN(n14924) );
  NAND2_X1 U8596 ( .A1(n7087), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7086) );
  INV_X1 U8597 ( .A(n12586), .ZN(n7087) );
  NOR2_X1 U8598 ( .A1(n12612), .A2(n12886), .ZN(n12618) );
  NAND2_X1 U8599 ( .A1(n7191), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U8600 ( .A1(n12619), .A2(n7191), .ZN(n6766) );
  INV_X1 U8601 ( .A(n12620), .ZN(n7191) );
  NAND2_X1 U8602 ( .A1(n12704), .A2(n12703), .ZN(n7195) );
  NAND2_X1 U8603 ( .A1(n12700), .A2(n12701), .ZN(n7194) );
  OAI21_X1 U8604 ( .B1(n12771), .B2(n12327), .A(n7052), .ZN(n12743) );
  AND2_X1 U8605 ( .A1(n7322), .A2(n7323), .ZN(n12809) );
  NAND2_X1 U8606 ( .A1(n8831), .A2(n8830), .ZN(n12937) );
  INV_X1 U8607 ( .A(n14448), .ZN(n12379) );
  NAND2_X1 U8608 ( .A1(n11020), .A2(n8691), .ZN(n11273) );
  NAND2_X1 U8609 ( .A1(n10776), .A2(n8648), .ZN(n10957) );
  NAND2_X1 U8610 ( .A1(n10839), .A2(n12360), .ZN(n10775) );
  AND3_X1 U8611 ( .A1(n8647), .A2(n8646), .A3(n8645), .ZN(n14988) );
  NAND2_X1 U8612 ( .A1(n10111), .A2(n7346), .ZN(n10867) );
  AND2_X1 U8613 ( .A1(n9035), .A2(n14940), .ZN(n14955) );
  INV_X1 U8614 ( .A(n12903), .ZN(n12889) );
  AND2_X1 U8615 ( .A1(n9995), .A2(n9032), .ZN(n12888) );
  INV_X1 U8616 ( .A(n12200), .ZN(n12965) );
  AND2_X1 U8617 ( .A1(n12766), .A2(n12765), .ZN(n12974) );
  NAND2_X1 U8618 ( .A1(n7342), .A2(n8876), .ZN(n12776) );
  NAND2_X1 U8619 ( .A1(n12789), .A2(n12788), .ZN(n7342) );
  NAND2_X1 U8620 ( .A1(n8855), .A2(n8854), .ZN(n12991) );
  NAND2_X1 U8621 ( .A1(n7056), .A2(n8997), .ZN(n12797) );
  NAND2_X1 U8622 ( .A1(n12807), .A2(n8996), .ZN(n7056) );
  NAND2_X1 U8623 ( .A1(n12846), .A2(n8811), .ZN(n12832) );
  NAND2_X1 U8624 ( .A1(n8995), .A2(n12416), .ZN(n12843) );
  NAND2_X1 U8625 ( .A1(n8790), .A2(n8789), .ZN(n13015) );
  NAND2_X1 U8626 ( .A1(n7324), .A2(n7326), .ZN(n12862) );
  NAND2_X1 U8627 ( .A1(n7329), .A2(n8768), .ZN(n12872) );
  NAND2_X1 U8628 ( .A1(n12882), .A2(n12879), .ZN(n7329) );
  NAND2_X1 U8629 ( .A1(n8760), .A2(n8759), .ZN(n13027) );
  NAND2_X1 U8630 ( .A1(n8744), .A2(n8743), .ZN(n13038) );
  AND2_X1 U8631 ( .A1(n9966), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13041) );
  NAND2_X1 U8632 ( .A1(n6654), .A2(n8456), .ZN(n13045) );
  INV_X1 U8633 ( .A(n8455), .ZN(n6654) );
  NAND2_X1 U8634 ( .A1(n7023), .A2(n7021), .ZN(n12476) );
  NAND2_X1 U8635 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n7022), .ZN(n7021) );
  NAND2_X1 U8636 ( .A1(n8510), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8512) );
  INV_X1 U8637 ( .A(n7039), .ZN(n7032) );
  AND2_X1 U8638 ( .A1(n7031), .A2(n7044), .ZN(n8889) );
  NAND2_X1 U8639 ( .A1(n13044), .A2(n7390), .ZN(n7389) );
  OR2_X1 U8640 ( .A1(n8943), .A2(n7388), .ZN(n7387) );
  INV_X1 U8641 ( .A(SI_13_), .ZN(n14403) );
  INV_X1 U8642 ( .A(n7017), .ZN(n8719) );
  AOI21_X1 U8643 ( .B1(n8702), .B2(n8701), .A(n7019), .ZN(n7017) );
  OAI21_X1 U8644 ( .B1(n6751), .B2(n6938), .A(n6936), .ZN(n8671) );
  OAI21_X1 U8645 ( .B1(n6751), .B2(n8640), .A(n8480), .ZN(n8658) );
  NAND2_X1 U8646 ( .A1(n6929), .A2(n8476), .ZN(n8611) );
  NAND2_X1 U8647 ( .A1(n8601), .A2(n8600), .ZN(n6929) );
  INV_X1 U8648 ( .A(n9729), .ZN(n9857) );
  OR3_X1 U8649 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8585) );
  INV_X1 U8650 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8569) );
  INV_X1 U8651 ( .A(n9675), .ZN(n9906) );
  OR2_X1 U8652 ( .A1(n11397), .A2(n11396), .ZN(n11398) );
  XNOR2_X1 U8653 ( .A(n11596), .B(n11597), .ZN(n7474) );
  NOR2_X1 U8654 ( .A1(n10913), .A2(n7459), .ZN(n7458) );
  INV_X1 U8655 ( .A(n10909), .ZN(n7459) );
  NAND2_X1 U8656 ( .A1(n10910), .A2(n10909), .ZN(n10912) );
  NAND2_X1 U8657 ( .A1(n7794), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U8658 ( .A1(n7683), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7695) );
  AND2_X1 U8659 ( .A1(n7693), .A2(n7692), .ZN(n6752) );
  NAND2_X1 U8660 ( .A1(n13159), .A2(n10054), .ZN(n10070) );
  NAND2_X2 U8661 ( .A1(n7894), .A2(n7893), .ZN(n11255) );
  CLKBUF_X1 U8662 ( .A(n13096), .Z(n13098) );
  OAI21_X1 U8663 ( .B1(n6753), .B2(n7488), .A(n7485), .ZN(n7490) );
  AOI21_X1 U8664 ( .B1(n6753), .B2(n7489), .A(n7488), .ZN(n13107) );
  NAND2_X1 U8665 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  NAND2_X1 U8666 ( .A1(n10102), .A2(n10103), .ZN(n10249) );
  NAND2_X1 U8667 ( .A1(n7484), .A2(n11574), .ZN(n7483) );
  INV_X1 U8668 ( .A(n7488), .ZN(n7484) );
  NAND2_X1 U8669 ( .A1(n7989), .A2(n7988), .ZN(n13581) );
  OR2_X1 U8670 ( .A1(n8254), .A2(n9132), .ZN(n6721) );
  OR2_X1 U8671 ( .A1(n8255), .A2(n7524), .ZN(n7703) );
  OR2_X1 U8672 ( .A1(n10250), .A2(n10251), .ZN(n10252) );
  NAND2_X1 U8673 ( .A1(n10249), .A2(n10248), .ZN(n10388) );
  NAND2_X1 U8674 ( .A1(n7469), .A2(n7470), .ZN(n13179) );
  XNOR2_X1 U8675 ( .A(n6753), .B(n11569), .ZN(n11571) );
  CLKBUF_X2 U8676 ( .A(n13213), .Z(n6748) );
  OAI21_X1 U8677 ( .B1(n13223), .B2(n13221), .A(n13220), .ZN(n13237) );
  INV_X1 U8678 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7908) );
  XNOR2_X1 U8679 ( .A(n13274), .B(n13273), .ZN(n14804) );
  OR2_X1 U8680 ( .A1(n14831), .A2(n14830), .ZN(n14834) );
  OAI22_X1 U8681 ( .A1(n13278), .A2(n14816), .B1(n14810), .B2(n13277), .ZN(
        n14829) );
  NAND2_X1 U8682 ( .A1(n6991), .A2(n10055), .ZN(n13510) );
  XNOR2_X1 U8683 ( .A(n13296), .B(n6992), .ZN(n6991) );
  INV_X1 U8684 ( .A(n8307), .ZN(n13513) );
  NOR2_X1 U8685 ( .A1(n13308), .A2(n13307), .ZN(n13522) );
  AOI211_X1 U8686 ( .C1(n13304), .C2(n13303), .A(n13451), .B(n6546), .ZN(
        n13308) );
  NAND2_X1 U8687 ( .A1(n7142), .A2(n7146), .ZN(n13303) );
  OR2_X1 U8688 ( .A1(n13312), .A2(n13473), .ZN(n6718) );
  NAND2_X1 U8689 ( .A1(n13631), .A2(n8236), .ZN(n8202) );
  INV_X1 U8690 ( .A(n7144), .ZN(n13316) );
  NAND2_X1 U8691 ( .A1(n13635), .A2(n8236), .ZN(n8158) );
  AND2_X1 U8692 ( .A1(n7437), .A2(n7435), .ZN(n13404) );
  NAND2_X1 U8693 ( .A1(n7153), .A2(n11796), .ZN(n13394) );
  NAND2_X1 U8694 ( .A1(n13414), .A2(n11795), .ZN(n7153) );
  OR2_X1 U8695 ( .A1(n11672), .A2(n8255), .ZN(n7625) );
  NAND2_X1 U8696 ( .A1(n7967), .A2(n7966), .ZN(n13587) );
  NAND2_X1 U8697 ( .A1(n7946), .A2(n7945), .ZN(n13593) );
  NAND2_X1 U8698 ( .A1(n11311), .A2(n11310), .ZN(n11415) );
  NAND2_X1 U8699 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  NAND2_X1 U8700 ( .A1(n10687), .A2(n10686), .ZN(n10689) );
  NAND2_X1 U8701 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  NAND2_X1 U8702 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  NAND2_X1 U8703 ( .A1(n10266), .A2(n10265), .ZN(n10268) );
  NAND2_X1 U8704 ( .A1(n13476), .A2(n10188), .ZN(n13498) );
  XNOR2_X1 U8705 ( .A(n6667), .B(n10377), .ZN(n14850) );
  INV_X2 U8706 ( .A(n14893), .ZN(n14895) );
  NAND2_X1 U8707 ( .A1(n13510), .A2(n6988), .ZN(n13606) );
  NOR2_X1 U8708 ( .A1(n6990), .A2(n6989), .ZN(n6988) );
  INV_X1 U8709 ( .A(n13511), .ZN(n6989) );
  NOR2_X1 U8710 ( .A1(n6992), .A2(n14859), .ZN(n6990) );
  AND2_X1 U8711 ( .A1(n13517), .A2(n13516), .ZN(n6758) );
  AND2_X1 U8712 ( .A1(n10079), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14843) );
  CLKBUF_X1 U8713 ( .A(n11800), .Z(n6719) );
  INV_X1 U8714 ( .A(n9497), .ZN(n10924) );
  AND2_X1 U8715 ( .A1(n7889), .A2(n6848), .ZN(n6847) );
  INV_X1 U8716 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9429) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9314) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9207) );
  INV_X1 U8719 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9131) );
  INV_X1 U8720 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9129) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n15157) );
  INV_X1 U8722 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9127) );
  INV_X1 U8723 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U8724 ( .A1(n10797), .A2(n10796), .ZN(n10973) );
  AND2_X1 U8725 ( .A1(n11827), .A2(n9814), .ZN(n9821) );
  NAND2_X1 U8726 ( .A1(n13885), .A2(n6778), .ZN(n13789) );
  AND2_X1 U8727 ( .A1(n13790), .A2(n13788), .ZN(n6778) );
  NOR2_X1 U8728 ( .A1(n6784), .A2(n13803), .ZN(n6783) );
  OAI22_X1 U8729 ( .A1(n6784), .A2(n6781), .B1(n13803), .B2(n6787), .ZN(n6780)
         );
  NOR2_X1 U8730 ( .A1(n13803), .A2(n13772), .ZN(n6781) );
  OR2_X1 U8731 ( .A1(n6788), .A2(n6786), .ZN(n6609) );
  INV_X1 U8732 ( .A(n13803), .ZN(n6786) );
  NAND2_X1 U8733 ( .A1(n10973), .A2(n10972), .ZN(n10974) );
  INV_X1 U8734 ( .A(n7283), .ZN(n9536) );
  AND2_X1 U8735 ( .A1(n7263), .A2(n6540), .ZN(n13813) );
  NAND2_X1 U8736 ( .A1(n6797), .A2(n6796), .ZN(n13653) );
  INV_X1 U8737 ( .A(n11473), .ZN(n6796) );
  OAI21_X1 U8738 ( .B1(n7254), .B2(n6803), .A(n6805), .ZN(n13829) );
  NAND2_X1 U8739 ( .A1(n10446), .A2(n10445), .ZN(n10659) );
  AND2_X1 U8740 ( .A1(n7270), .A2(n6525), .ZN(n13845) );
  XNOR2_X1 U8741 ( .A(n11451), .B(n11449), .ZN(n11448) );
  NAND2_X1 U8742 ( .A1(n7256), .A2(n7257), .ZN(n13877) );
  INV_X1 U8743 ( .A(n7258), .ZN(n7257) );
  OR2_X1 U8744 ( .A1(n13866), .A2(n6526), .ZN(n7256) );
  CLKBUF_X1 U8745 ( .A(n14473), .Z(n14498) );
  NAND2_X1 U8746 ( .A1(n9804), .A2(n9803), .ZN(n11828) );
  NAND2_X1 U8747 ( .A1(n11828), .A2(n11829), .ZN(n11827) );
  NAND2_X1 U8748 ( .A1(n7264), .A2(n7267), .ZN(n13886) );
  OR2_X1 U8749 ( .A1(n13908), .A2(n7268), .ZN(n7264) );
  NAND2_X1 U8750 ( .A1(n7249), .A2(n6794), .ZN(n10792) );
  OAI21_X1 U8751 ( .B1(n10446), .B2(n7251), .A(n7250), .ZN(n10666) );
  AND2_X1 U8752 ( .A1(n14480), .A2(n14691), .ZN(n14502) );
  INV_X1 U8753 ( .A(n12059), .ZN(n12098) );
  CLKBUF_X1 U8754 ( .A(n13950), .Z(n6678) );
  AOI21_X1 U8755 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10622), .A(n9241), .ZN(
        n9223) );
  AOI21_X1 U8756 ( .B1(n10714), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9928), .ZN(
        n9931) );
  INV_X1 U8757 ( .A(n6729), .ZN(n14552) );
  AND2_X1 U8758 ( .A1(n14028), .A2(n14579), .ZN(n14593) );
  INV_X1 U8759 ( .A(n14261), .ZN(n14064) );
  XOR2_X1 U8760 ( .A(n12089), .B(n11749), .Z(n14269) );
  OAI21_X1 U8761 ( .B1(n14082), .B2(n7168), .A(n7166), .ZN(n11749) );
  NAND2_X1 U8762 ( .A1(n14085), .A2(n7171), .ZN(n7168) );
  NAND2_X1 U8763 ( .A1(n7167), .A2(n7171), .ZN(n7166) );
  NAND2_X1 U8764 ( .A1(n14147), .A2(n11702), .ZN(n14138) );
  NAND2_X1 U8765 ( .A1(n14161), .A2(n11768), .ZN(n14146) );
  NAND2_X1 U8766 ( .A1(n14203), .A2(n11671), .ZN(n14178) );
  AND2_X1 U8767 ( .A1(n14215), .A2(n11763), .ZN(n14196) );
  NAND2_X1 U8768 ( .A1(n11633), .A2(n11632), .ZN(n14238) );
  NAND2_X1 U8769 ( .A1(n11512), .A2(n11934), .ZN(n11759) );
  NAND2_X1 U8770 ( .A1(n7159), .A2(n11424), .ZN(n11522) );
  NAND2_X1 U8771 ( .A1(n7394), .A2(n11144), .ZN(n11349) );
  NAND2_X1 U8772 ( .A1(n11142), .A2(n11141), .ZN(n7394) );
  NAND2_X1 U8773 ( .A1(n7173), .A2(n11113), .ZN(n11165) );
  NAND2_X1 U8774 ( .A1(n7113), .A2(n10707), .ZN(n10755) );
  NAND2_X1 U8775 ( .A1(n10706), .A2(n10705), .ZN(n7113) );
  AND2_X1 U8776 ( .A1(n14671), .A2(n10228), .ZN(n14647) );
  OAI211_X1 U8777 ( .C1(n14677), .C2(n14275), .A(n14274), .B(n14273), .ZN(
        n14351) );
  AND2_X1 U8778 ( .A1(n14278), .A2(n6762), .ZN(n6761) );
  AND2_X1 U8779 ( .A1(n14277), .A2(n14279), .ZN(n6762) );
  NAND2_X1 U8780 ( .A1(n7272), .A2(n6821), .ZN(n14367) );
  AND3_X1 U8781 ( .A1(n7416), .A2(n6541), .A3(n6822), .ZN(n6821) );
  NOR2_X1 U8782 ( .A1(n9087), .A2(n6823), .ZN(n6822) );
  NAND2_X1 U8783 ( .A1(n6824), .A2(n9174), .ZN(n6823) );
  XNOR2_X1 U8784 ( .A(n7284), .B(P1_IR_REG_25__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U8785 ( .A1(n9059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7284) );
  MUX2_X1 U8786 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9058), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9060) );
  NAND2_X1 U8787 ( .A1(n6966), .A2(n6972), .ZN(n8121) );
  NAND2_X1 U8788 ( .A1(n6969), .A2(n6972), .ZN(n8104) );
  OR2_X1 U8789 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  INV_X1 U8790 ( .A(n12019), .ZN(n12037) );
  INV_X1 U8791 ( .A(n12036), .ZN(n12030) );
  NAND2_X1 U8792 ( .A1(n8041), .A2(n8040), .ZN(n11659) );
  INV_X1 U8793 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9316) );
  INV_X1 U8794 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9199) );
  OR2_X1 U8795 ( .A1(n9198), .A2(n9197), .ZN(n9936) );
  INV_X1 U8796 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9168) );
  INV_X1 U8797 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9111) );
  AND2_X1 U8798 ( .A1(n9105), .A2(n9112), .ZN(n10448) );
  NAND2_X1 U8799 ( .A1(n6886), .A2(n8373), .ZN(n14393) );
  NAND2_X1 U8800 ( .A1(n15245), .A2(n15244), .ZN(n6886) );
  NAND2_X1 U8801 ( .A1(n8378), .A2(n6891), .ZN(n15236) );
  NAND2_X1 U8802 ( .A1(n15243), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n6891) );
  INV_X1 U8803 ( .A(n6892), .ZN(n8377) );
  XNOR2_X1 U8804 ( .A(n8383), .B(n8382), .ZN(n15238) );
  XNOR2_X1 U8805 ( .A(n8384), .B(n7100), .ZN(n14408) );
  INV_X1 U8806 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7100) );
  XNOR2_X1 U8807 ( .A(n8389), .B(n7098), .ZN(n15241) );
  INV_X1 U8808 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U8809 ( .A1(n7096), .A2(n8398), .ZN(n14420) );
  NAND2_X1 U8810 ( .A1(n14418), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7096) );
  OAI21_X1 U8811 ( .B1(n14420), .B2(n14421), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6651) );
  NAND2_X1 U8812 ( .A1(n6888), .A2(n6512), .ZN(n14539) );
  NOR2_X1 U8813 ( .A1(n8415), .A2(n8416), .ZN(n14542) );
  AND2_X1 U8814 ( .A1(n8415), .A2(n8416), .ZN(n14543) );
  NOR2_X1 U8815 ( .A1(n8421), .A2(n8420), .ZN(n14545) );
  AND2_X1 U8816 ( .A1(n8421), .A2(n8420), .ZN(n14546) );
  XNOR2_X1 U8817 ( .A(n6904), .B(n12290), .ZN(n12298) );
  INV_X1 U8818 ( .A(n12677), .ZN(n12670) );
  INV_X1 U8819 ( .A(n6773), .ZN(n6772) );
  OAI21_X1 U8820 ( .B1(n12697), .B2(n6771), .A(n12592), .ZN(n6770) );
  OAI21_X1 U8821 ( .B1(n9041), .B2(n12892), .A(n9040), .ZN(n9042) );
  INV_X1 U8822 ( .A(n6710), .ZN(n6709) );
  OAI22_X1 U8823 ( .A1(n12968), .A2(n12961), .B1(n15025), .B2(n12914), .ZN(
        n6710) );
  INV_X1 U8824 ( .A(n6713), .ZN(n6712) );
  OAI22_X1 U8825 ( .A1(n12968), .A2(n13039), .B1(n15010), .B2(n12967), .ZN(
        n6713) );
  NAND2_X1 U8826 ( .A1(n10672), .A2(n10671), .ZN(n10675) );
  AND2_X1 U8827 ( .A1(n7457), .A2(n7456), .ZN(n13088) );
  NAND2_X1 U8828 ( .A1(n10087), .A2(n10086), .ZN(n10090) );
  NAND2_X1 U8829 ( .A1(n6867), .A2(n8320), .ZN(n6865) );
  OAI21_X1 U8830 ( .B1(n13214), .B2(n7455), .A(n7454), .ZN(P2_U3531) );
  INV_X1 U8831 ( .A(n6667), .ZN(n7455) );
  NAND2_X1 U8832 ( .A1(n13214), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7454) );
  INV_X1 U8833 ( .A(n7448), .ZN(n11826) );
  OAI21_X1 U8834 ( .B1(n13518), .B2(n13504), .A(n7449), .ZN(n7448) );
  AOI21_X1 U8835 ( .B1(n13514), .B2(n13507), .A(n11825), .ZN(n7449) );
  INV_X1 U8836 ( .A(n6985), .ZN(P2_U3530) );
  AOI21_X1 U8837 ( .B1(n13606), .B2(n14895), .A(n6986), .ZN(n6985) );
  NOR2_X1 U8838 ( .A1(n14895), .A2(n6987), .ZN(n6986) );
  INV_X1 U8839 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6987) );
  INV_X1 U8840 ( .A(n6707), .ZN(n6706) );
  OAI21_X1 U8841 ( .B1(n14279), .B2(n13779), .A(n13778), .ZN(n6707) );
  NOR2_X1 U8842 ( .A1(n14536), .A2(n14535), .ZN(n14534) );
  AND2_X1 U8843 ( .A1(n6890), .A2(n6527), .ZN(n14536) );
  XNOR2_X1 U8844 ( .A(n6532), .B(n8435), .ZN(n7101) );
  AND2_X1 U8845 ( .A1(n9497), .A2(n14855), .ZN(n6517) );
  NOR2_X1 U8846 ( .A1(n8782), .A2(n7328), .ZN(n6501) );
  AND2_X1 U8847 ( .A1(n7581), .A2(SI_14_), .ZN(n6502) );
  INV_X1 U8848 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13044) );
  INV_X1 U8849 ( .A(n9526), .ZN(n13690) );
  AND2_X2 U8850 ( .A1(n9822), .A2(n11845), .ZN(n9526) );
  NAND2_X2 U8851 ( .A1(n8202), .A2(n8201), .ZN(n13520) );
  OR2_X1 U8852 ( .A1(n8311), .A2(n6687), .ZN(n6503) );
  INV_X2 U8853 ( .A(n11846), .ZN(n12026) );
  AND2_X1 U8854 ( .A1(n6488), .A2(n7403), .ZN(n6504) );
  AND2_X1 U8855 ( .A1(n7420), .A2(n10729), .ZN(n6505) );
  AND2_X1 U8856 ( .A1(n7070), .A2(n12416), .ZN(n6506) );
  NAND2_X1 U8857 ( .A1(n13687), .A2(n13842), .ZN(n6507) );
  XNOR2_X1 U8858 ( .A(n6691), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U8859 ( .A1(n11948), .A2(n11947), .ZN(n6508) );
  NAND2_X1 U8860 ( .A1(n12753), .A2(n12218), .ZN(n6509) );
  AND2_X1 U8861 ( .A1(n6727), .A2(n13206), .ZN(n6510) );
  AND2_X1 U8862 ( .A1(n12080), .A2(n11924), .ZN(n6511) );
  NAND2_X1 U8863 ( .A1(n14535), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6512) );
  INV_X1 U8864 ( .A(n7924), .ZN(n7303) );
  OR2_X1 U8865 ( .A1(n7958), .A2(n7957), .ZN(n6513) );
  OR2_X1 U8866 ( .A1(n7765), .A2(n7764), .ZN(n6514) );
  NOR2_X1 U8867 ( .A1(n13565), .A2(n13195), .ZN(n6515) );
  INV_X1 U8868 ( .A(n11873), .ZN(n7213) );
  AOI21_X1 U8869 ( .B1(n7020), .B2(n8487), .A(n6627), .ZN(n7018) );
  INV_X1 U8870 ( .A(n14204), .ZN(n7130) );
  INV_X1 U8871 ( .A(n12879), .ZN(n7327) );
  XNOR2_X1 U8872 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8600) );
  INV_X1 U8873 ( .A(n8600), .ZN(n6931) );
  NAND2_X1 U8874 ( .A1(n8043), .A2(n8042), .ZN(n13565) );
  INV_X1 U8875 ( .A(n13565), .ZN(n7004) );
  NAND2_X1 U8876 ( .A1(n11237), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U8877 ( .A1(n7010), .A2(n7009), .ZN(n11317) );
  INV_X1 U8878 ( .A(n11317), .ZN(n7008) );
  INV_X2 U8879 ( .A(n8214), .ZN(n8215) );
  INV_X1 U8880 ( .A(n9726), .ZN(n7180) );
  XNOR2_X1 U8881 ( .A(n12937), .B(n12811), .ZN(n12821) );
  INV_X1 U8882 ( .A(n12821), .ZN(n7318) );
  NAND2_X1 U8883 ( .A1(n7410), .A2(n9092), .ZN(n9087) );
  AND2_X1 U8884 ( .A1(n7365), .A2(n7367), .ZN(n6518) );
  OR2_X1 U8885 ( .A1(n12753), .A2(n12218), .ZN(n12453) );
  NOR2_X1 U8886 ( .A1(n8015), .A2(n8012), .ZN(n6519) );
  AND2_X1 U8887 ( .A1(n7050), .A2(n7049), .ZN(n6520) );
  AND2_X1 U8888 ( .A1(n6643), .A2(n6642), .ZN(n6521) );
  AND2_X1 U8889 ( .A1(n7937), .A2(n7936), .ZN(n6522) );
  AND3_X1 U8890 ( .A1(n7513), .A2(n7511), .A3(n7515), .ZN(n6523) );
  AND4_X1 U8891 ( .A1(n13334), .A2(n8303), .A3(n13363), .A4(n13353), .ZN(n6524) );
  NAND2_X1 U8892 ( .A1(n13680), .A2(n13679), .ZN(n6525) );
  OR2_X1 U8893 ( .A1(n7261), .A2(n13873), .ZN(n6526) );
  OR2_X1 U8894 ( .A1(n8404), .A2(n8405), .ZN(n6527) );
  NAND2_X1 U8895 ( .A1(n13532), .A2(n13100), .ZN(n6528) );
  NOR2_X1 U8896 ( .A1(n6913), .A2(n8597), .ZN(n8612) );
  OR2_X1 U8897 ( .A1(n12697), .A2(n12696), .ZN(n6529) );
  AND2_X1 U8898 ( .A1(n10158), .A2(n14937), .ZN(n6530) );
  OR2_X1 U8899 ( .A1(n13352), .A2(n13180), .ZN(n6531) );
  NAND2_X1 U8900 ( .A1(n8195), .A2(n8194), .ZN(n8247) );
  INV_X1 U8901 ( .A(n8247), .ZN(n6992) );
  INV_X1 U8902 ( .A(n9757), .ZN(n7084) );
  XOR2_X1 U8903 ( .A(n8439), .B(P3_ADDR_REG_19__SCAN_IN), .Z(n6532) );
  INV_X1 U8904 ( .A(n12375), .ZN(n7073) );
  INV_X1 U8905 ( .A(n13772), .ZN(n6788) );
  AND2_X1 U8906 ( .A1(n11893), .A2(n10881), .ZN(n6533) );
  INV_X1 U8907 ( .A(n13081), .ZN(n9504) );
  OR2_X1 U8908 ( .A1(n14503), .A2(n13939), .ZN(n6534) );
  INV_X1 U8909 ( .A(n13571), .ZN(n7006) );
  OR2_X1 U8910 ( .A1(n6520), .A2(n6924), .ZN(n6535) );
  OR2_X1 U8911 ( .A1(n8266), .A2(n8267), .ZN(n6536) );
  AND2_X1 U8912 ( .A1(n10112), .A2(n8621), .ZN(n6537) );
  AND2_X1 U8913 ( .A1(n13598), .A2(n11539), .ZN(n6538) );
  OR2_X1 U8914 ( .A1(n8393), .A2(n8392), .ZN(n6539) );
  NAND2_X1 U8915 ( .A1(n13712), .A2(n13711), .ZN(n6540) );
  AND2_X1 U8916 ( .A1(n6825), .A2(n9055), .ZN(n6541) );
  AND2_X1 U8917 ( .A1(n12191), .A2(n12197), .ZN(n6542) );
  OR2_X1 U8918 ( .A1(n12991), .A2(n12551), .ZN(n6543) );
  AND2_X1 U8919 ( .A1(n11926), .A2(n11999), .ZN(n6544) );
  OR2_X1 U8920 ( .A1(n13581), .A2(n13169), .ZN(n6545) );
  AND2_X1 U8921 ( .A1(n7141), .A2(n7142), .ZN(n6546) );
  AND2_X1 U8922 ( .A1(n13839), .A2(n13847), .ZN(n6547) );
  AND2_X1 U8923 ( .A1(n11216), .A2(n11215), .ZN(n6548) );
  AND2_X1 U8924 ( .A1(n7865), .A2(n7864), .ZN(n6549) );
  AND2_X1 U8925 ( .A1(n7976), .A2(n7975), .ZN(n6550) );
  NOR2_X1 U8926 ( .A1(n12618), .A2(n12619), .ZN(n6551) );
  AND2_X1 U8927 ( .A1(n6646), .A2(n6645), .ZN(n6552) );
  AND2_X1 U8928 ( .A1(n8997), .A2(n7058), .ZN(n6553) );
  XNOR2_X1 U8929 ( .A(n7538), .B(n9077), .ZN(n7696) );
  INV_X1 U8930 ( .A(n7696), .ZN(n6666) );
  NOR2_X1 U8931 ( .A1(n14327), .A2(n13932), .ZN(n6554) );
  OR2_X1 U8932 ( .A1(n10491), .A2(n10472), .ZN(n6555) );
  OR2_X1 U8933 ( .A1(n7921), .A2(n7923), .ZN(n6556) );
  AND2_X1 U8934 ( .A1(n11975), .A2(n11974), .ZN(n6557) );
  OR2_X1 U8935 ( .A1(n12645), .A2(n6765), .ZN(n6764) );
  AND2_X1 U8936 ( .A1(n8441), .A2(n7386), .ZN(n7385) );
  OR2_X1 U8937 ( .A1(n7905), .A2(n7904), .ZN(n6558) );
  AND2_X1 U8938 ( .A1(n14156), .A2(n11769), .ZN(n6559) );
  INV_X1 U8939 ( .A(n6957), .ZN(n6956) );
  NAND2_X1 U8940 ( .A1(n7592), .A2(SI_17_), .ZN(n6957) );
  NAND2_X1 U8941 ( .A1(n13565), .A2(n13195), .ZN(n6560) );
  INV_X1 U8942 ( .A(n7147), .ZN(n7146) );
  AND2_X1 U8943 ( .A1(n13557), .A2(n13375), .ZN(n6561) );
  INV_X1 U8944 ( .A(n6795), .ZN(n6794) );
  OR2_X1 U8945 ( .A1(n8383), .A2(n8382), .ZN(n6562) );
  NOR2_X1 U8946 ( .A1(n13598), .A2(n11539), .ZN(n6563) );
  NOR2_X1 U8947 ( .A1(n13557), .A2(n13091), .ZN(n6564) );
  NOR2_X1 U8948 ( .A1(n14246), .A2(n13681), .ZN(n6565) );
  NOR2_X1 U8949 ( .A1(n14492), .A2(n11914), .ZN(n6566) );
  OR2_X1 U8950 ( .A1(n7006), .A2(n13170), .ZN(n6567) );
  AND2_X1 U8951 ( .A1(n12968), .A2(n12197), .ZN(n6568) );
  INV_X1 U8952 ( .A(n8055), .ZN(n7503) );
  INV_X1 U8953 ( .A(n12314), .ZN(n6921) );
  INV_X1 U8954 ( .A(n7340), .ZN(n7339) );
  OR2_X1 U8955 ( .A1(n8887), .A2(n7341), .ZN(n7340) );
  AND2_X1 U8956 ( .A1(n14093), .A2(n11776), .ZN(n6569) );
  INV_X1 U8957 ( .A(n7866), .ZN(n7518) );
  INV_X1 U8958 ( .A(n7297), .ZN(n7296) );
  OAI21_X1 U8959 ( .B1(n7572), .B2(n7298), .A(n7528), .ZN(n7297) );
  AND2_X1 U8960 ( .A1(n12152), .A2(n12791), .ZN(n6570) );
  NOR2_X1 U8961 ( .A1(n14314), .A2(n13930), .ZN(n6571) );
  AND2_X1 U8962 ( .A1(n8054), .A2(n8053), .ZN(n6572) );
  AND2_X1 U8963 ( .A1(n7705), .A2(n7704), .ZN(n6573) );
  NOR2_X1 U8964 ( .A1(n7494), .A2(n7922), .ZN(n6574) );
  AND2_X1 U8965 ( .A1(n9129), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6575) );
  AND2_X1 U8966 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6576) );
  AND2_X1 U8967 ( .A1(n8481), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6577) );
  AND2_X1 U8968 ( .A1(n11934), .A2(n11925), .ZN(n12080) );
  OR2_X1 U8969 ( .A1(n9980), .A2(n10826), .ZN(n6578) );
  AND2_X1 U8970 ( .A1(n6920), .A2(n12313), .ZN(n6579) );
  NAND2_X1 U8971 ( .A1(n7520), .A2(n6874), .ZN(n6580) );
  INV_X1 U8972 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8973 ( .A1(n14083), .A2(n7169), .ZN(n6581) );
  NAND2_X1 U8974 ( .A1(n13688), .A2(n6525), .ZN(n6582) );
  OR2_X1 U8975 ( .A1(n8076), .A2(n8075), .ZN(n6583) );
  AND2_X1 U8976 ( .A1(n12771), .A2(n12321), .ZN(n6584) );
  OR2_X1 U8977 ( .A1(n7180), .A2(n9693), .ZN(n6585) );
  OR2_X1 U8978 ( .A1(n7978), .A2(n6550), .ZN(n6586) );
  AND2_X1 U8979 ( .A1(n13764), .A2(n13943), .ZN(n6587) );
  AND2_X1 U8980 ( .A1(n7366), .A2(n7362), .ZN(n6588) );
  INV_X1 U8981 ( .A(n7745), .ZN(n7746) );
  AND2_X1 U8982 ( .A1(n7829), .A2(n7828), .ZN(n6589) );
  INV_X1 U8983 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6824) );
  AND2_X1 U8984 ( .A1(n11949), .A2(n11950), .ZN(n14224) );
  INV_X1 U8985 ( .A(n14224), .ZN(n6837) );
  NOR2_X1 U8986 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n6590) );
  OR2_X1 U8987 ( .A1(n13388), .A2(n13194), .ZN(n6591) );
  AND2_X1 U8988 ( .A1(n11523), .A2(n11424), .ZN(n6592) );
  AND2_X1 U8989 ( .A1(n11908), .A2(n6828), .ZN(n6593) );
  AND2_X1 U8990 ( .A1(n7560), .A2(SI_8_), .ZN(n6594) );
  AND2_X1 U8991 ( .A1(n7330), .A2(n7326), .ZN(n6595) );
  AND2_X1 U8992 ( .A1(n6504), .A2(n11779), .ZN(n6596) );
  AND2_X1 U8993 ( .A1(n10673), .A2(n10671), .ZN(n6597) );
  INV_X1 U8994 ( .A(n10707), .ZN(n7114) );
  AND2_X1 U8995 ( .A1(n8661), .A2(n8648), .ZN(n6598) );
  AND2_X1 U8996 ( .A1(n6848), .A2(n7626), .ZN(n6599) );
  OR2_X1 U8997 ( .A1(n7785), .A2(n7787), .ZN(n6600) );
  NAND2_X1 U8998 ( .A1(n14270), .A2(n11778), .ZN(n6601) );
  OR2_X1 U8999 ( .A1(n12965), .A2(n8926), .ZN(n6602) );
  OR2_X1 U9000 ( .A1(n7786), .A2(n7508), .ZN(n6603) );
  AND2_X1 U9001 ( .A1(n6527), .A2(n6889), .ZN(n6604) );
  AND2_X1 U9002 ( .A1(n8452), .A2(n8513), .ZN(n6605) );
  NAND2_X1 U9003 ( .A1(n7228), .A2(n11912), .ZN(n6606) );
  OR2_X1 U9004 ( .A1(n7748), .A2(n7746), .ZN(n6607) );
  INV_X1 U9005 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9174) );
  INV_X1 U9006 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7390) );
  INV_X1 U9007 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7274) );
  INV_X1 U9008 ( .A(n7075), .ZN(n7074) );
  NAND2_X1 U9009 ( .A1(n12382), .A2(n7076), .ZN(n7075) );
  OR2_X1 U9010 ( .A1(n7213), .A2(n11874), .ZN(n6608) );
  INV_X1 U9011 ( .A(n7775), .ZN(n8257) );
  INV_X1 U9012 ( .A(n12842), .ZN(n7070) );
  AND2_X1 U9013 ( .A1(n7597), .A2(n9774), .ZN(n6610) );
  NAND2_X1 U9014 ( .A1(n11727), .A2(n11726), .ZN(n14283) );
  INV_X1 U9015 ( .A(n14283), .ZN(n7204) );
  AND2_X1 U9016 ( .A1(n11064), .A2(n7157), .ZN(n6611) );
  INV_X1 U9017 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6726) );
  INV_X1 U9018 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7027) );
  INV_X1 U9019 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6734) );
  XOR2_X1 U9020 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .Z(n6612) );
  XOR2_X1 U9021 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .Z(n6613) );
  NAND2_X1 U9022 ( .A1(n11427), .A2(n11426), .ZN(n14345) );
  INV_X1 U9023 ( .A(n14345), .ZN(n6744) );
  AND2_X1 U9024 ( .A1(n11597), .A2(n13066), .ZN(n6614) );
  AND2_X1 U9025 ( .A1(n8092), .A2(n8091), .ZN(n13126) );
  INV_X1 U9026 ( .A(n14295), .ZN(n7206) );
  INV_X1 U9027 ( .A(n8701), .ZN(n7020) );
  NAND2_X1 U9028 ( .A1(n7007), .A2(n7006), .ZN(n13457) );
  INV_X1 U9029 ( .A(n13457), .ZN(n7005) );
  NOR2_X1 U9030 ( .A1(n14924), .A2(n12568), .ZN(n6615) );
  AND2_X1 U9031 ( .A1(n14222), .A2(n11949), .ZN(n6616) );
  INV_X1 U9032 ( .A(SI_14_), .ZN(n15172) );
  AND2_X1 U9033 ( .A1(n6911), .A2(n12139), .ZN(n6617) );
  AND2_X1 U9034 ( .A1(n7613), .A2(n7889), .ZN(n6618) );
  AND2_X1 U9035 ( .A1(n11430), .A2(n11924), .ZN(n6619) );
  AND2_X1 U9036 ( .A1(n12522), .A2(n12851), .ZN(n6620) );
  AND2_X1 U9037 ( .A1(n12554), .A2(n12379), .ZN(n6621) );
  AND2_X1 U9038 ( .A1(n12230), .A2(n12406), .ZN(n6622) );
  NAND2_X1 U9039 ( .A1(n9287), .A2(n15253), .ZN(n6623) );
  NAND2_X1 U9040 ( .A1(n12160), .A2(n12292), .ZN(n7368) );
  OR2_X1 U9041 ( .A1(n12965), .A2(n12961), .ZN(n6624) );
  AND2_X1 U9042 ( .A1(n10452), .A2(n13939), .ZN(n6625) );
  NOR2_X1 U9043 ( .A1(n11328), .A2(n7377), .ZN(n6626) );
  INV_X1 U9044 ( .A(n8839), .ZN(n7323) );
  INV_X1 U9045 ( .A(n10429), .ZN(n7443) );
  INV_X1 U9046 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7013) );
  INV_X1 U9047 ( .A(n14503), .ZN(n7200) );
  XOR2_X1 U9048 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .Z(n6627) );
  INV_X1 U9049 ( .A(n12079), .ZN(n6755) );
  NAND2_X1 U9050 ( .A1(n7928), .A2(n7927), .ZN(n13598) );
  INV_X1 U9051 ( .A(n13598), .ZN(n7011) );
  INV_X1 U9052 ( .A(n14327), .ZN(n7201) );
  INV_X1 U9053 ( .A(n8174), .ZN(n7312) );
  OAI21_X1 U9054 ( .B1(n9170), .B2(P3_D_REG_0__SCAN_IN), .A(n8954), .ZN(n7369)
         );
  NOR2_X1 U9055 ( .A1(n10492), .A2(n10493), .ZN(n6628) );
  AND2_X1 U9056 ( .A1(n10249), .A2(n7479), .ZN(n6629) );
  AND2_X1 U9057 ( .A1(n7444), .A2(n10590), .ZN(n6630) );
  AND2_X1 U9058 ( .A1(n10973), .A2(n7280), .ZN(n6631) );
  INV_X1 U9059 ( .A(n7197), .ZN(n11361) );
  NOR2_X1 U9060 ( .A1(n11047), .A2(n7198), .ZN(n7197) );
  INV_X1 U9061 ( .A(n8038), .ZN(n7604) );
  INV_X1 U9062 ( .A(n6700), .ZN(n11388) );
  AOI21_X1 U9063 ( .B1(n8948), .B2(P3_IR_REG_25__SCAN_IN), .A(n6701), .ZN(
        n6700) );
  AND2_X1 U9064 ( .A1(n12572), .A2(n12575), .ZN(n6632) );
  NOR2_X1 U9065 ( .A1(n12702), .A2(n7194), .ZN(n6633) );
  AND2_X1 U9066 ( .A1(n10111), .A2(n8604), .ZN(n6634) );
  AND2_X1 U9067 ( .A1(n11081), .A2(n11080), .ZN(n6635) );
  INV_X1 U9068 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7022) );
  INV_X1 U9069 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7036) );
  INV_X1 U9070 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7043) );
  INV_X1 U9071 ( .A(n14868), .ZN(n6997) );
  NAND2_X1 U9072 ( .A1(n7913), .A2(n7912), .ZN(n13603) );
  INV_X1 U9073 ( .A(n13603), .ZN(n7009) );
  INV_X1 U9074 ( .A(n10036), .ZN(n7203) );
  OR2_X1 U9075 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7036), .ZN(n6636) );
  NAND2_X1 U9076 ( .A1(n8502), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6637) );
  INV_X1 U9077 ( .A(n7044), .ZN(n7041) );
  NAND2_X1 U9078 ( .A1(n11715), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7044) );
  INV_X1 U9079 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6738) );
  INV_X1 U9080 ( .A(SI_24_), .ZN(n6970) );
  INV_X1 U9081 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7095) );
  INV_X1 U9082 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7092) );
  AOI21_X1 U9083 ( .B1(n11805), .B2(n13488), .A(n11804), .ZN(n13517) );
  NAND2_X1 U9084 ( .A1(n11781), .A2(n14643), .ZN(n14267) );
  AOI21_X1 U9085 ( .B1(n14069), .B2(n14643), .A(n14068), .ZN(n14274) );
  INV_X2 U9086 ( .A(n13633), .ZN(n13636) );
  NOR2_X2 U9087 ( .A1(n12761), .A2(n6638), .ZN(n12745) );
  OR2_X2 U9088 ( .A1(n6499), .A2(n8543), .ZN(n8546) );
  NAND2_X1 U9089 ( .A1(n12716), .A2(n6602), .ZN(n6704) );
  NAND2_X1 U9090 ( .A1(n12316), .A2(n12463), .ZN(n6643) );
  NAND2_X1 U9091 ( .A1(n6741), .A2(n8473), .ZN(n8584) );
  NAND2_X1 U9092 ( .A1(n6927), .A2(n6928), .ZN(n8630) );
  NAND2_X1 U9093 ( .A1(n11736), .A2(n11735), .ZN(n14082) );
  NAND3_X1 U9094 ( .A1(n7120), .A2(n7415), .A3(n9147), .ZN(n6644) );
  NAND2_X1 U9095 ( .A1(n11643), .A2(n11642), .ZN(n14209) );
  NAND2_X1 U9096 ( .A1(n14071), .A2(n14070), .ZN(n6647) );
  NAND2_X1 U9097 ( .A1(n6750), .A2(n6749), .ZN(n11551) );
  NAND2_X1 U9098 ( .A1(n14111), .A2(n14113), .ZN(n14110) );
  NAND3_X1 U9099 ( .A1(n7532), .A2(n14048), .A3(n7531), .ZN(n6668) );
  NAND2_X1 U9100 ( .A1(n6736), .A2(n7604), .ZN(n8041) );
  NAND2_X1 U9101 ( .A1(n7940), .A2(n7939), .ZN(n7942) );
  AOI21_X1 U9102 ( .B1(n6962), .B2(n6963), .A(n6594), .ZN(n6960) );
  INV_X1 U9103 ( .A(n7603), .ZN(n6648) );
  NAND2_X1 U9104 ( .A1(n6768), .A2(n6585), .ZN(n7179) );
  NOR2_X2 U9105 ( .A1(n14913), .A2(n12576), .ZN(n12610) );
  XNOR2_X1 U9106 ( .A(n11187), .B(n11188), .ZN(n14898) );
  NAND2_X1 U9107 ( .A1(n9675), .A2(n7182), .ZN(n7181) );
  NAND2_X1 U9108 ( .A1(n7181), .A2(n9665), .ZN(n9894) );
  NAND2_X1 U9109 ( .A1(n12573), .A2(n6632), .ZN(n6715) );
  INV_X1 U9110 ( .A(n8039), .ZN(n6736) );
  NAND2_X1 U9111 ( .A1(n8041), .A2(n7601), .ZN(n7609) );
  OAI21_X1 U9112 ( .B1(n12612), .B2(n7190), .A(n6766), .ZN(n12645) );
  AOI21_X1 U9113 ( .B1(n12664), .B2(n6764), .A(n12663), .ZN(n12666) );
  XNOR2_X1 U9114 ( .A(n6529), .B(n12699), .ZN(n7196) );
  INV_X1 U9115 ( .A(n13333), .ZN(n11820) );
  OAI21_X2 U9116 ( .B1(n13354), .B2(n11817), .A(n6531), .ZN(n13333) );
  OR2_X2 U9117 ( .A1(n10326), .A2(n10308), .ZN(n6650) );
  NAND2_X1 U9118 ( .A1(n6671), .A2(n6670), .ZN(n12566) );
  NAND2_X1 U9119 ( .A1(n12568), .A2(n7087), .ZN(n7085) );
  NAND2_X1 U9120 ( .A1(n8425), .A2(n14434), .ZN(n6881) );
  NAND2_X1 U9121 ( .A1(n6881), .A2(n6882), .ZN(n6880) );
  NAND2_X1 U9122 ( .A1(n7404), .A2(n7403), .ZN(n6652) );
  AOI21_X2 U9123 ( .B1(n10507), .B2(n10506), .A(n10505), .ZN(n10508) );
  INV_X1 U9124 ( .A(n7275), .ZN(n7120) );
  AND3_X2 U9125 ( .A1(n9802), .A2(n9801), .A3(n9800), .ZN(n10236) );
  NAND2_X1 U9126 ( .A1(n10029), .A2(n11854), .ZN(n10028) );
  NAND2_X1 U9127 ( .A1(n14110), .A2(n11725), .ZN(n14098) );
  NAND2_X1 U9128 ( .A1(n11169), .A2(n11168), .ZN(n11345) );
  AOI21_X1 U9129 ( .B1(n11658), .B2(n11657), .A(n6554), .ZN(n14205) );
  OR2_X2 U9130 ( .A1(n14082), .A2(n6488), .ZN(n14083) );
  AOI21_X2 U9131 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10157) );
  NAND2_X1 U9132 ( .A1(n6732), .A2(n6731), .ZN(n10559) );
  AOI21_X1 U9133 ( .B1(n7379), .B2(n9981), .A(n6684), .ZN(n6683) );
  NAND2_X1 U9134 ( .A1(n8913), .A2(n8912), .ZN(n8922) );
  INV_X1 U9135 ( .A(n8922), .ZN(n8921) );
  NAND2_X1 U9136 ( .A1(n7789), .A2(n7557), .ZN(n6961) );
  NAND2_X1 U9137 ( .A1(n10940), .A2(n10939), .ZN(n10942) );
  NAND2_X1 U9138 ( .A1(n11369), .A2(n7376), .ZN(n12116) );
  NAND2_X1 U9139 ( .A1(n12123), .A2(n12122), .ZN(n12168) );
  NAND2_X1 U9140 ( .A1(n10858), .A2(n10859), .ZN(n10910) );
  NAND2_X1 U9141 ( .A1(n11235), .A2(n11234), .ZN(n11237) );
  NAND2_X1 U9142 ( .A1(n11536), .A2(n11535), .ZN(n11568) );
  NAND2_X1 U9143 ( .A1(n10260), .A2(n10259), .ZN(n10672) );
  AND2_X1 U9144 ( .A1(n10088), .A2(n10086), .ZN(n7481) );
  AOI21_X1 U9145 ( .B1(n13135), .B2(n13131), .A(n13133), .ZN(n13090) );
  OAI22_X1 U9146 ( .A1(n11568), .A2(n7483), .B1(n7485), .B2(n11575), .ZN(
        n13116) );
  NAND2_X1 U9147 ( .A1(n12911), .A2(n6624), .ZN(P3_U3487) );
  NAND2_X2 U9148 ( .A1(n12785), .A2(n12784), .ZN(n12787) );
  OAI21_X2 U9149 ( .B1(n8995), .B2(n7069), .A(n7067), .ZN(n12818) );
  OAI21_X2 U9150 ( .B1(n12901), .B2(n8992), .A(n12402), .ZN(n12880) );
  NAND2_X1 U9151 ( .A1(n6922), .A2(n7050), .ZN(n12729) );
  OAI211_X1 U9152 ( .C1(n8317), .C2(n6865), .A(n6656), .B(n8340), .ZN(P2_U3328) );
  NAND2_X1 U9153 ( .A1(n8317), .A2(n6864), .ZN(n6656) );
  NAND2_X1 U9154 ( .A1(n6971), .A2(n6970), .ZN(n6969) );
  NAND2_X1 U9155 ( .A1(n7568), .A2(n7567), .ZN(n7868) );
  NAND2_X1 U9156 ( .A1(n6692), .A2(n7548), .ZN(n6979) );
  NAND2_X1 U9157 ( .A1(n6980), .A2(n6982), .ZN(n6981) );
  INV_X1 U9158 ( .A(n6876), .ZN(n7306) );
  OAI211_X1 U9159 ( .C1(n8268), .C2(n7309), .A(n8273), .B(n7306), .ZN(n8279)
         );
  NAND2_X1 U9160 ( .A1(n11957), .A2(n11956), .ZN(n11960) );
  INV_X1 U9161 ( .A(n11976), .ZN(n6660) );
  NAND2_X2 U9162 ( .A1(n11511), .A2(n11510), .ZN(n13839) );
  AOI21_X2 U9163 ( .B1(n7677), .B2(n7676), .A(n7537), .ZN(n7697) );
  OAI22_X1 U9164 ( .A1(n11982), .A2(n6845), .B1(n11983), .B2(n6844), .ZN(
        n11987) );
  NAND2_X1 U9165 ( .A1(n7543), .A2(n7542), .ZN(n7730) );
  NOR3_X1 U9166 ( .A1(n11933), .A2(n11932), .A3(n11938), .ZN(n7530) );
  NAND2_X1 U9167 ( .A1(n11973), .A2(n11972), .ZN(n11976) );
  NAND2_X1 U9168 ( .A1(n11992), .A2(n11991), .ZN(n11994) );
  NAND2_X1 U9169 ( .A1(n10727), .A2(n10726), .ZN(n10750) );
  AOI21_X2 U9170 ( .B1(n10030), .B2(n12064), .A(n9914), .ZN(n10507) );
  NAND4_X1 U9171 ( .A1(n8310), .A2(n8308), .A3(n8309), .A4(n10924), .ZN(n8311)
         );
  NAND2_X2 U9172 ( .A1(n14114), .A2(n11773), .ZN(n14101) );
  XNOR2_X1 U9173 ( .A(n7697), .B(n6666), .ZN(n7524) );
  INV_X1 U9174 ( .A(n8062), .ZN(n6980) );
  INV_X1 U9175 ( .A(n9808), .ZN(n11848) );
  NAND3_X1 U9176 ( .A1(n9577), .A2(n9575), .A3(n9576), .ZN(n9808) );
  NOR2_X1 U9177 ( .A1(n12866), .A2(n12646), .ZN(n12663) );
  NOR2_X1 U9178 ( .A1(n12665), .A2(n12666), .ZN(n12697) );
  INV_X1 U9179 ( .A(n10207), .ZN(n7182) );
  NOR2_X1 U9180 ( .A1(n9692), .A2(n6769), .ZN(n9693) );
  NOR2_X2 U9181 ( .A1(n6777), .A2(n6776), .ZN(n11187) );
  OAI21_X2 U9182 ( .B1(n12610), .B2(n12609), .A(n12611), .ZN(n12617) );
  AOI21_X1 U9183 ( .B1(n9666), .B2(P3_REG2_REG_0__SCAN_IN), .A(n9893), .ZN(
        n9669) );
  AND2_X4 U9184 ( .A1(n11566), .A2(n13630), .ZN(n8027) );
  XNOR2_X2 U9185 ( .A(n7652), .B(n7651), .ZN(n11566) );
  OAI21_X2 U9186 ( .B1(n11400), .B2(n11399), .A(n11398), .ZN(n11402) );
  NAND2_X1 U9187 ( .A1(n13082), .A2(n10050), .ZN(n13160) );
  NOR2_X1 U9188 ( .A1(n13116), .A2(n13115), .ZN(n13114) );
  AOI21_X1 U9189 ( .B1(n13123), .B2(n13124), .A(n11601), .ZN(n13096) );
  NAND2_X1 U9190 ( .A1(n7135), .A2(n6528), .ZN(n7144) );
  NAND2_X1 U9191 ( .A1(n7469), .A2(n7467), .ZN(n13176) );
  INV_X1 U9192 ( .A(n11178), .ZN(n6671) );
  NOR2_X2 U9193 ( .A1(n14904), .A2(n11174), .ZN(n11178) );
  AND2_X2 U9194 ( .A1(n10325), .A2(n10324), .ZN(n10472) );
  NAND2_X1 U9195 ( .A1(n7627), .A2(n6673), .ZN(n6680) );
  NAND3_X1 U9196 ( .A1(n6981), .A2(n6984), .A3(n6983), .ZN(n8077) );
  NAND2_X1 U9197 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  NAND3_X1 U9198 ( .A1(n7134), .A2(n6675), .A3(n6674), .ZN(n11799) );
  NAND3_X1 U9199 ( .A1(n6676), .A2(n9984), .A3(n10129), .ZN(n10130) );
  XNOR2_X1 U9200 ( .A(n6704), .B(n12533), .ZN(n8936) );
  AND2_X1 U9201 ( .A1(n9383), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U9202 ( .A1(n8702), .A2(n7018), .ZN(n6940) );
  NAND2_X1 U9203 ( .A1(n12222), .A2(n12133), .ZN(n12233) );
  NAND2_X1 U9204 ( .A1(n10768), .A2(n10767), .ZN(n10770) );
  INV_X1 U9205 ( .A(n7031), .ZN(n7033) );
  INV_X1 U9206 ( .A(n7349), .ZN(n7348) );
  XNOR2_X2 U9207 ( .A(n12739), .B(n12746), .ZN(n6924) );
  NAND3_X1 U9208 ( .A1(n6826), .A2(n7416), .A3(n7272), .ZN(n9178) );
  NAND2_X1 U9209 ( .A1(n11551), .A2(n9574), .ZN(n9579) );
  XNOR2_X1 U9210 ( .A(n9179), .B(n6824), .ZN(n9180) );
  NAND2_X1 U9211 ( .A1(n14083), .A2(n11748), .ZN(n14071) );
  NAND2_X1 U9212 ( .A1(n13176), .A2(n11607), .ZN(n13060) );
  INV_X1 U9213 ( .A(n7479), .ZN(n7478) );
  NAND2_X1 U9214 ( .A1(n13160), .A2(n13161), .ZN(n13159) );
  NAND2_X1 U9215 ( .A1(n7381), .A2(n7380), .ZN(n12222) );
  NAND2_X1 U9216 ( .A1(n10560), .A2(n10765), .ZN(n10768) );
  NAND2_X1 U9217 ( .A1(n6578), .A2(n6683), .ZN(n9982) );
  NOR2_X1 U9218 ( .A1(n13361), .A2(n6685), .ZN(n13354) );
  NOR2_X2 U9219 ( .A1(n13362), .A2(n13363), .ZN(n13361) );
  OR2_X2 U9220 ( .A1(n13096), .A2(n13097), .ZN(n7469) );
  NAND3_X1 U9221 ( .A1(n6847), .A2(n6492), .A3(n6999), .ZN(n7630) );
  AOI21_X2 U9222 ( .B1(n11820), .B2(n11819), .A(n11818), .ZN(n13321) );
  XNOR2_X1 U9223 ( .A(n10336), .B(n13210), .ZN(n9949) );
  NAND2_X1 U9224 ( .A1(n13083), .A2(n13084), .ZN(n13082) );
  NAND2_X1 U9225 ( .A1(n11003), .A2(n11002), .ZN(n11235) );
  OAI22_X1 U9226 ( .A1(n13090), .A2(n13089), .B1(n11590), .B2(n11589), .ZN(
        n11591) );
  NAND2_X1 U9227 ( .A1(n7160), .A2(n14147), .ZN(n14140) );
  NAND2_X1 U9228 ( .A1(n9579), .A2(n9578), .ZN(n9910) );
  INV_X2 U9229 ( .A(n11682), .ZN(n9068) );
  NAND2_X1 U9230 ( .A1(n8485), .A2(n8484), .ZN(n8702) );
  NAND2_X1 U9231 ( .A1(n8498), .A2(n8497), .ZN(n8842) );
  INV_X1 U9232 ( .A(n6696), .ZN(n6695) );
  NAND2_X1 U9233 ( .A1(n7730), .A2(n7546), .ZN(n6692) );
  NAND2_X1 U9234 ( .A1(n7832), .A2(n7561), .ZN(n7564) );
  NAND2_X1 U9235 ( .A1(n6959), .A2(n6960), .ZN(n7832) );
  MUX2_X1 U9236 ( .A(n13934), .B(n13839), .S(n11953), .Z(n11944) );
  NAND2_X1 U9237 ( .A1(n10150), .A2(n10168), .ZN(n12355) );
  NAND2_X1 U9238 ( .A1(n7325), .A2(n6501), .ZN(n7324) );
  AOI21_X1 U9239 ( .B1(n6924), .B2(n12731), .A(n12730), .ZN(n12735) );
  AOI21_X1 U9240 ( .B1(n15009), .B2(n12913), .A(n12912), .ZN(n12966) );
  NOR2_X2 U9241 ( .A1(n12759), .A2(n12758), .ZN(n12761) );
  INV_X1 U9242 ( .A(n6916), .ZN(n6915) );
  NAND2_X1 U9243 ( .A1(n8842), .A2(n8840), .ZN(n8499) );
  INV_X1 U9244 ( .A(n14942), .ZN(n12337) );
  NAND2_X1 U9245 ( .A1(n8981), .A2(n12343), .ZN(n10209) );
  NAND2_X1 U9246 ( .A1(n8986), .A2(n12369), .ZN(n10983) );
  NAND2_X1 U9247 ( .A1(n8479), .A2(n8478), .ZN(n8641) );
  OAI21_X1 U9248 ( .B1(n6917), .B2(n6915), .A(n12494), .ZN(n12498) );
  INV_X1 U9249 ( .A(n7369), .ZN(n13042) );
  AND2_X4 U9250 ( .A1(n9981), .A2(n9980), .ZN(n12153) );
  NAND2_X1 U9251 ( .A1(n12127), .A2(n7382), .ZN(n7381) );
  INV_X1 U9252 ( .A(n10295), .ZN(n6732) );
  NAND2_X1 U9253 ( .A1(n13321), .A2(n13320), .ZN(n13524) );
  NAND2_X1 U9254 ( .A1(n8369), .A2(n8368), .ZN(n7093) );
  AOI21_X1 U9255 ( .B1(n15193), .B2(n8409), .A(n14538), .ZN(n8410) );
  NAND2_X1 U9256 ( .A1(n10028), .A2(n9911), .ZN(n10501) );
  NAND2_X1 U9257 ( .A1(n10620), .A2(n10619), .ZN(n14639) );
  NAND2_X1 U9258 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  INV_X1 U9259 ( .A(n12063), .ZN(n6750) );
  NAND2_X1 U9260 ( .A1(n7324), .A2(n6595), .ZN(n12859) );
  NAND2_X1 U9261 ( .A1(n12338), .A2(n8979), .ZN(n10827) );
  NAND2_X1 U9262 ( .A1(n6705), .A2(n7338), .ZN(n12759) );
  NAND2_X1 U9263 ( .A1(n7523), .A2(n10211), .ZN(n10210) );
  NAND2_X1 U9264 ( .A1(n8864), .A2(n7336), .ZN(n6705) );
  NAND2_X1 U9265 ( .A1(n6708), .A2(n6706), .ZN(P1_U3214) );
  NAND2_X1 U9266 ( .A1(n13773), .A2(n14504), .ZN(n6708) );
  NAND2_X1 U9267 ( .A1(n6711), .A2(n6709), .ZN(P3_U3486) );
  OR2_X1 U9268 ( .A1(n12966), .A2(n15023), .ZN(n6711) );
  NAND2_X1 U9269 ( .A1(n6714), .A2(n6712), .ZN(P3_U3454) );
  OR2_X1 U9270 ( .A1(n12966), .A2(n15012), .ZN(n6714) );
  NAND2_X1 U9271 ( .A1(n13653), .A2(n13652), .ZN(n14489) );
  INV_X1 U9272 ( .A(n11474), .ZN(n6797) );
  NAND2_X1 U9273 ( .A1(n12859), .A2(n8797), .ZN(n12848) );
  NAND2_X1 U9274 ( .A1(n10841), .A2(n8633), .ZN(n10778) );
  NOR2_X1 U9275 ( .A1(n11322), .A2(n14383), .ZN(n7285) );
  INV_X1 U9276 ( .A(n12798), .ZN(n8862) );
  NAND2_X1 U9277 ( .A1(n8062), .A2(SI_22_), .ZN(n6984) );
  OR2_X2 U9278 ( .A1(n9863), .A2(n9862), .ZN(n10322) );
  NOR2_X1 U9279 ( .A1(n9859), .A2(n9860), .ZN(n9863) );
  XNOR2_X1 U9280 ( .A(n9693), .B(n7180), .ZN(n10014) );
  NAND2_X1 U9281 ( .A1(n7179), .A2(n7178), .ZN(n9846) );
  AOI21_X1 U9282 ( .B1(n7196), .B2(n12592), .A(n7193), .ZN(n7192) );
  NOR2_X1 U9283 ( .A1(n9755), .A2(n10869), .ZN(n9754) );
  NAND2_X1 U9284 ( .A1(n13412), .A2(n7435), .ZN(n7433) );
  INV_X1 U9285 ( .A(n13426), .ZN(n6717) );
  AOI21_X2 U9286 ( .B1(n6717), .B2(n6560), .A(n6515), .ZN(n13412) );
  OAI21_X2 U9287 ( .B1(n13444), .B2(n11816), .A(n6567), .ZN(n13426) );
  NAND2_X1 U9288 ( .A1(n7231), .A2(n7229), .ZN(n11962) );
  NAND2_X1 U9289 ( .A1(n6838), .A2(n7218), .ZN(n12000) );
  NAND2_X1 U9290 ( .A1(n11878), .A2(n11879), .ZN(n11877) );
  OAI21_X1 U9291 ( .B1(n6557), .B2(n7222), .A(n7220), .ZN(n11982) );
  NAND2_X1 U9292 ( .A1(n7176), .A2(n7174), .ZN(n11793) );
  NAND2_X1 U9293 ( .A1(n7105), .A2(n7104), .ZN(n11493) );
  NAND3_X1 U9294 ( .A1(n13522), .A2(n13311), .A3(n6718), .ZN(n13313) );
  NAND3_X2 U9295 ( .A1(n7702), .A2(n7703), .A3(n6721), .ZN(n13158) );
  INV_X4 U9296 ( .A(n7678), .ZN(n9332) );
  OAI21_X2 U9297 ( .B1(n10423), .B2(n7445), .A(n7442), .ZN(n10810) );
  OAI21_X1 U9298 ( .B1(n11380), .B2(n8991), .A(n12397), .ZN(n12901) );
  NAND4_X2 U9299 ( .A1(n8552), .A2(n8553), .A3(n8554), .A4(n8551), .ZN(n10830)
         );
  AND2_X2 U9300 ( .A1(n6729), .A2(n6728), .ZN(n14569) );
  NOR2_X2 U9301 ( .A1(n14619), .A2(n15192), .ZN(n14623) );
  AOI21_X2 U9302 ( .B1(n10448), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9307), .ZN(
        n9243) );
  NAND2_X1 U9303 ( .A1(n8061), .A2(n8060), .ZN(n8062) );
  NAND2_X1 U9304 ( .A1(n8081), .A2(n8080), .ZN(n8101) );
  NAND2_X1 U9305 ( .A1(n12204), .A2(n12147), .ZN(n12150) );
  OAI21_X1 U9306 ( .B1(n7998), .B2(n7291), .A(n7289), .ZN(n7608) );
  INV_X8 U9307 ( .A(n9068), .ZN(n9517) );
  AOI21_X1 U9308 ( .B1(n9949), .B2(n10265), .A(n10272), .ZN(n7429) );
  XNOR2_X1 U9309 ( .A(n7789), .B(n7788), .ZN(n10628) );
  XNOR2_X2 U9310 ( .A(n13213), .B(n13081), .ZN(n9495) );
  NAND2_X1 U9311 ( .A1(n10421), .A2(n10420), .ZN(n10522) );
  NAND2_X1 U9312 ( .A1(n11199), .A2(n11198), .ZN(n11201) );
  NAND2_X1 U9313 ( .A1(n13771), .A2(n13772), .ZN(n13797) );
  XNOR2_X1 U9314 ( .A(n6979), .B(n7749), .ZN(n10447) );
  NAND2_X1 U9315 ( .A1(n13384), .A2(n6591), .ZN(n13362) );
  OAI21_X2 U9316 ( .B1(n11682), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6739), .ZN(
        n7536) );
  NAND2_X1 U9317 ( .A1(n7426), .A2(n7429), .ZN(n10421) );
  NAND2_X1 U9318 ( .A1(n8739), .A2(n8738), .ZN(n6740) );
  NAND2_X1 U9319 ( .A1(n8573), .A2(n8571), .ZN(n6741) );
  XNOR2_X2 U9320 ( .A(n9155), .B(n9153), .ZN(n14378) );
  NAND2_X1 U9321 ( .A1(n15253), .A2(n7119), .ZN(n7275) );
  NAND2_X1 U9322 ( .A1(n7173), .A2(n7172), .ZN(n11167) );
  INV_X1 U9323 ( .A(n11112), .ZN(n6743) );
  NAND2_X1 U9324 ( .A1(n14168), .A2(n14167), .ZN(n14166) );
  INV_X1 U9325 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7531) );
  NAND2_X1 U9326 ( .A1(n7207), .A2(n7206), .ZN(n14132) );
  INV_X1 U9327 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U9328 ( .A1(n14245), .A2(n14246), .ZN(n14248) );
  NAND2_X1 U9329 ( .A1(n7202), .A2(n7201), .ZN(n14210) );
  NAND2_X1 U9330 ( .A1(n11345), .A2(n11344), .ZN(n11423) );
  NAND2_X1 U9331 ( .A1(n7205), .A2(n7204), .ZN(n14089) );
  NAND2_X2 U9333 ( .A1(n10984), .A2(n12388), .ZN(n11021) );
  NAND2_X1 U9334 ( .A1(n10210), .A2(n8591), .ZN(n10113) );
  NOR2_X1 U9335 ( .A1(n14905), .A2(n8693), .ZN(n14904) );
  XNOR2_X1 U9336 ( .A(n11173), .B(n11188), .ZN(n14905) );
  AOI21_X2 U9337 ( .B1(n12677), .B2(n12676), .A(n12675), .ZN(n12684) );
  XNOR2_X1 U9338 ( .A(n12672), .B(n12671), .ZN(n12644) );
  OAI21_X2 U9339 ( .B1(n11307), .B2(n11306), .A(n11308), .ZN(n11413) );
  NAND2_X1 U9340 ( .A1(n7433), .A2(n7431), .ZN(n13384) );
  INV_X1 U9341 ( .A(n11423), .ZN(n6756) );
  INV_X1 U9342 ( .A(n14149), .ZN(n6757) );
  NAND2_X1 U9343 ( .A1(n8539), .A2(n8555), .ZN(n8472) );
  INV_X1 U9344 ( .A(n8293), .ZN(n13212) );
  AND3_X2 U9345 ( .A1(n7695), .A2(n7694), .A3(n6752), .ZN(n8293) );
  NAND3_X2 U9346 ( .A1(n12787), .A2(n12775), .A3(n12772), .ZN(n12771) );
  NAND2_X1 U9347 ( .A1(n7063), .A2(n7061), .ZN(n10954) );
  INV_X1 U9348 ( .A(n6923), .ZN(n6922) );
  NAND2_X1 U9349 ( .A1(n8984), .A2(n8983), .ZN(n7048) );
  NOR3_X2 U9350 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .A3(
        P2_IR_REG_18__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U9351 ( .A1(n11265), .A2(n11264), .ZN(n11400) );
  OAI21_X2 U9352 ( .B1(n13076), .B2(n13072), .A(n13073), .ZN(n13135) );
  NAND2_X1 U9353 ( .A1(n6552), .A2(n6761), .ZN(n14352) );
  INV_X1 U9354 ( .A(n7445), .ZN(n7444) );
  OAI21_X1 U9355 ( .B1(n13518), .B2(n14875), .A(n6758), .ZN(n13608) );
  NAND2_X1 U9356 ( .A1(n7195), .A2(n6633), .ZN(n7193) );
  NOR2_X1 U9357 ( .A1(n12621), .A2(n6759), .ZN(n12652) );
  AND2_X1 U9358 ( .A1(n12622), .A2(n12628), .ZN(n6759) );
  OAI21_X2 U9359 ( .B1(n7582), .B2(n7302), .A(n7300), .ZN(n7940) );
  NAND4_X1 U9360 ( .A1(n6760), .A2(n8442), .A3(n7077), .A4(n8447), .ZN(n8939)
         );
  NOR2_X1 U9361 ( .A1(n10015), .A2(n9728), .ZN(n9848) );
  OAI21_X1 U9362 ( .B1(n12705), .B2(n14926), .A(n7192), .ZN(P3_U3201) );
  OR2_X2 U9363 ( .A1(n9882), .A2(n9881), .ZN(n10325) );
  NOR2_X1 U9364 ( .A1(n9679), .A2(n9680), .ZN(n9725) );
  NOR2_X2 U9365 ( .A1(n12597), .A2(n12952), .ZN(n12629) );
  OR2_X2 U9366 ( .A1(n14101), .A2(n11775), .ZN(n7404) );
  NAND2_X1 U9367 ( .A1(n7405), .A2(n7408), .ZN(n14128) );
  NAND2_X1 U9368 ( .A1(n7419), .A2(n7418), .ZN(n10883) );
  INV_X2 U9369 ( .A(n7275), .ZN(n7272) );
  OR2_X2 U9370 ( .A1(n14022), .A2(n14021), .ZN(n14619) );
  NAND2_X1 U9371 ( .A1(n6481), .A2(n10589), .ZN(n7445) );
  XNOR2_X1 U9372 ( .A(n7812), .B(n7811), .ZN(n10708) );
  OAI21_X1 U9373 ( .B1(n11413), .B2(n11412), .A(n11414), .ZN(n11484) );
  XNOR2_X1 U9374 ( .A(n6763), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14043) );
  OR2_X1 U9375 ( .A1(n14623), .A2(n14022), .ZN(n6763) );
  NOR2_X1 U9376 ( .A1(n14897), .A2(n11189), .ZN(n12571) );
  XNOR2_X2 U9377 ( .A(n6764), .B(n12664), .ZN(n12646) );
  NOR2_X2 U9378 ( .A1(n9777), .A2(n10783), .ZN(n9859) );
  NAND3_X1 U9379 ( .A1(n12680), .A2(n6772), .A3(n6770), .ZN(P3_U3200) );
  AND2_X1 U9380 ( .A1(n11186), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6776) );
  AOI21_X1 U9381 ( .B1(n6628), .B2(n10495), .A(n6777), .ZN(n10496) );
  OAI21_X2 U9382 ( .B1(n10323), .B2(n7188), .A(n7187), .ZN(n6777) );
  NAND2_X1 U9383 ( .A1(n13894), .A2(n13770), .ZN(n13771) );
  NAND3_X1 U9384 ( .A1(n6785), .A2(n6782), .A3(n6780), .ZN(n13811) );
  NAND2_X1 U9385 ( .A1(n13894), .A2(n6783), .ZN(n6782) );
  INV_X1 U9386 ( .A(n6787), .ZN(n6784) );
  OR2_X1 U9387 ( .A1(n13894), .A2(n6609), .ZN(n6785) );
  NAND2_X1 U9388 ( .A1(n10665), .A2(n7248), .ZN(n6795) );
  INV_X1 U9389 ( .A(n7254), .ZN(n6800) );
  NAND2_X1 U9390 ( .A1(n7254), .A2(n6801), .ZN(n6804) );
  INV_X1 U9391 ( .A(n9253), .ZN(n9148) );
  NAND3_X1 U9392 ( .A1(n15253), .A2(n6813), .A3(n6814), .ZN(n9253) );
  AND2_X2 U9393 ( .A1(n6815), .A2(n6814), .ZN(n9147) );
  NOR2_X1 U9394 ( .A1(n9087), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U9395 ( .A1(n6829), .A2(n6593), .ZN(n11907) );
  NAND2_X1 U9396 ( .A1(n11903), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U9397 ( .A1(n6835), .A2(n6833), .ZN(n11952) );
  INV_X1 U9398 ( .A(n6834), .ZN(n6833) );
  OAI21_X1 U9399 ( .B1(n7215), .B2(n6837), .A(n11951), .ZN(n6834) );
  NAND3_X1 U9400 ( .A1(n11923), .A2(n6836), .A3(n7214), .ZN(n6835) );
  NAND3_X1 U9401 ( .A1(n11562), .A2(n14373), .A3(P1_REG0_REG_0__SCAN_IN), .ZN(
        n9192) );
  XNOR2_X2 U9402 ( .A(n9177), .B(n9176), .ZN(n11562) );
  OAI211_X1 U9403 ( .C1(n11994), .C2(n11995), .A(n6839), .B(n7217), .ZN(n6838)
         );
  NAND2_X1 U9404 ( .A1(n6840), .A2(n11993), .ZN(n6839) );
  NAND2_X1 U9405 ( .A1(n11994), .A2(n11995), .ZN(n6840) );
  NAND2_X1 U9406 ( .A1(n6843), .A2(n11870), .ZN(n11871) );
  NAND2_X1 U9407 ( .A1(n7237), .A2(n7238), .ZN(n6843) );
  NAND2_X1 U9408 ( .A1(n11987), .A2(n11988), .ZN(n11986) );
  NAND2_X1 U9409 ( .A1(n6846), .A2(n6492), .ZN(n7627) );
  AND2_X2 U9410 ( .A1(n6999), .A2(n7889), .ZN(n7451) );
  NAND3_X1 U9411 ( .A1(n6851), .A2(n6558), .A3(n6850), .ZN(n6849) );
  INV_X1 U9412 ( .A(n7906), .ZN(n6851) );
  NAND3_X1 U9413 ( .A1(n6857), .A2(n6856), .A3(n6860), .ZN(n7848) );
  NAND3_X1 U9414 ( .A1(n6859), .A2(n6589), .A3(n6858), .ZN(n6856) );
  NAND3_X1 U9415 ( .A1(n6859), .A2(n6861), .A3(n6858), .ZN(n6857) );
  OAI21_X1 U9416 ( .B1(n8058), .B2(n8057), .A(n6583), .ZN(n6863) );
  NAND2_X1 U9417 ( .A1(n7519), .A2(n6871), .ZN(n6868) );
  NAND2_X1 U9418 ( .A1(n6868), .A2(n6869), .ZN(n7509) );
  NAND3_X1 U9419 ( .A1(n6536), .A2(n7307), .A3(n8304), .ZN(n6877) );
  XNOR2_X1 U9420 ( .A(n6878), .B(n7101), .ZN(SUB_1596_U4) );
  INV_X1 U9421 ( .A(n6880), .ZN(n8433) );
  INV_X1 U9422 ( .A(n8434), .ZN(n6879) );
  INV_X1 U9423 ( .A(n14431), .ZN(n6882) );
  NAND2_X1 U9424 ( .A1(n6890), .A2(n6604), .ZN(n6888) );
  AOI21_X1 U9425 ( .B1(n12272), .B2(n12812), .A(n12151), .ZN(n12241) );
  NAND2_X1 U9426 ( .A1(n12272), .A2(n6903), .ZN(n6902) );
  NAND2_X1 U9427 ( .A1(n10942), .A2(n6908), .ZN(n6907) );
  NAND2_X1 U9428 ( .A1(n8924), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U9429 ( .A1(n8921), .A2(n8914), .ZN(n8924) );
  INV_X1 U9430 ( .A(n7385), .ZN(n6913) );
  NOR2_X2 U9431 ( .A1(n8501), .A2(n6926), .ZN(n8866) );
  NAND2_X1 U9432 ( .A1(n8601), .A2(n6930), .ZN(n6927) );
  NAND2_X1 U9433 ( .A1(n8641), .A2(n6936), .ZN(n6933) );
  NAND2_X1 U9434 ( .A1(n6933), .A2(n6934), .ZN(n8483) );
  XNOR2_X2 U9435 ( .A(n8488), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U9436 ( .A1(n8813), .A2(n8812), .ZN(n6941) );
  NAND2_X1 U9437 ( .A1(n8800), .A2(n8798), .ZN(n6942) );
  NAND2_X1 U9438 ( .A1(n8771), .A2(n8769), .ZN(n6943) );
  NAND2_X1 U9439 ( .A1(n8756), .A2(n8754), .ZN(n6944) );
  NAND2_X1 U9440 ( .A1(n12327), .A2(n12324), .ZN(n6946) );
  OAI21_X1 U9441 ( .B1(n12327), .B2(n12321), .A(n12324), .ZN(n6945) );
  NAND2_X1 U9442 ( .A1(n7961), .A2(n6949), .ZN(n6948) );
  NAND2_X1 U9443 ( .A1(n7789), .A2(n6962), .ZN(n6959) );
  NAND2_X1 U9444 ( .A1(n7310), .A2(n7311), .ZN(n6964) );
  NAND2_X1 U9445 ( .A1(n6964), .A2(n15031), .ZN(n6965) );
  INV_X1 U9446 ( .A(n8102), .ZN(n6971) );
  OAI21_X1 U9447 ( .B1(n7697), .B2(n6666), .A(n7539), .ZN(n7286) );
  NAND2_X1 U9448 ( .A1(n6976), .A2(n6973), .ZN(n7543) );
  INV_X1 U9449 ( .A(n6974), .ZN(n6973) );
  OAI21_X1 U9450 ( .B1(n7696), .B2(n6975), .A(n7540), .ZN(n6974) );
  INV_X1 U9451 ( .A(n7539), .ZN(n6975) );
  NAND2_X1 U9452 ( .A1(n7697), .A2(n7539), .ZN(n6976) );
  XNOR2_X2 U9453 ( .A(n7536), .B(SI_1_), .ZN(n7677) );
  NAND2_X1 U9454 ( .A1(n7293), .A2(n7292), .ZN(n6977) );
  NAND2_X1 U9455 ( .A1(n6979), .A2(n7549), .ZN(n7552) );
  NAND2_X1 U9456 ( .A1(n6981), .A2(n6984), .ZN(n11683) );
  NAND2_X1 U9457 ( .A1(n8077), .A2(n6984), .ZN(n8081) );
  CLKBUF_X1 U9458 ( .A(n6995), .Z(n6993) );
  INV_X1 U9459 ( .A(n6996), .ZN(n10531) );
  NAND3_X1 U9460 ( .A1(n6999), .A2(n7889), .A3(n7622), .ZN(n6998) );
  AND2_X2 U9461 ( .A1(n7613), .A2(n7452), .ZN(n6999) );
  AND4_X2 U9462 ( .A1(n7612), .A2(n7769), .A3(n7610), .A4(n7611), .ZN(n7889)
         );
  NOR2_X2 U9463 ( .A1(n13515), .A2(n13309), .ZN(n13297) );
  NOR2_X2 U9464 ( .A1(n13490), .A2(n13576), .ZN(n7007) );
  NOR2_X2 U9465 ( .A1(n11417), .A2(n13593), .ZN(n11487) );
  NOR2_X2 U9466 ( .A1(n11102), .A2(n11255), .ZN(n7010) );
  NAND2_X1 U9467 ( .A1(n7048), .A2(n12506), .ZN(n8985) );
  XNOR2_X1 U9468 ( .A(n7048), .B(n8620), .ZN(n14979) );
  NAND2_X4 U9469 ( .A1(n13050), .A2(n12542), .ZN(n9646) );
  NAND2_X1 U9470 ( .A1(n12807), .A2(n7057), .ZN(n7053) );
  NAND2_X1 U9471 ( .A1(n7053), .A2(n7054), .ZN(n12785) );
  NAND2_X1 U9472 ( .A1(n10837), .A2(n7064), .ZN(n7063) );
  OAI21_X1 U9473 ( .B1(n12503), .B2(n7066), .A(n12507), .ZN(n7065) );
  OAI21_X1 U9474 ( .B1(n11024), .B2(n12383), .A(n12375), .ZN(n11272) );
  NAND2_X1 U9475 ( .A1(n12383), .A2(n12375), .ZN(n7076) );
  AND2_X2 U9476 ( .A1(n7081), .A2(n7080), .ZN(n11172) );
  NOR2_X2 U9477 ( .A1(n9792), .A2(n9779), .ZN(n9878) );
  XNOR2_X2 U9478 ( .A(n9876), .B(n9877), .ZN(n9792) );
  AND2_X2 U9479 ( .A1(n9790), .A2(n9789), .ZN(n9876) );
  NOR2_X2 U9480 ( .A1(n9750), .A2(n9712), .ZN(n9749) );
  XNOR2_X2 U9481 ( .A(n12567), .B(n12575), .ZN(n14925) );
  OR2_X2 U9482 ( .A1(n12644), .A2(n15058), .ZN(n12677) );
  NOR2_X2 U9483 ( .A1(n12643), .A2(n7088), .ZN(n12672) );
  INV_X1 U9484 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U9485 ( .A1(n7099), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U9486 ( .A1(n11206), .A2(n7106), .ZN(n7105) );
  AOI21_X1 U9487 ( .B1(n12068), .B2(n10707), .A(n12070), .ZN(n7109) );
  NAND2_X1 U9488 ( .A1(n10706), .A2(n7109), .ZN(n7111) );
  NAND2_X1 U9489 ( .A1(n7111), .A2(n7110), .ZN(n10874) );
  NAND2_X1 U9490 ( .A1(n10756), .A2(n7114), .ZN(n7112) );
  OAI21_X1 U9492 ( .B1(n6742), .B2(n7126), .A(n7124), .ZN(n14225) );
  NAND2_X1 U9493 ( .A1(n7123), .A2(n7121), .ZN(n11643) );
  NAND2_X1 U9494 ( .A1(n11526), .A2(n7124), .ZN(n7123) );
  NAND2_X1 U9495 ( .A1(n13330), .A2(n7136), .ZN(n7134) );
  NAND2_X1 U9496 ( .A1(n13330), .A2(n13334), .ZN(n7135) );
  NOR2_X1 U9497 ( .A1(n11821), .A2(n13191), .ZN(n7147) );
  NAND2_X1 U9498 ( .A1(n7159), .A2(n6592), .ZN(n11525) );
  NAND2_X2 U9499 ( .A1(n7678), .A2(n9517), .ZN(n8255) );
  NAND2_X2 U9500 ( .A1(n7165), .A2(n7161), .ZN(n13081) );
  NAND3_X1 U9501 ( .A1(n7678), .A2(n7163), .A3(n7162), .ZN(n7161) );
  NAND2_X1 U9502 ( .A1(n7620), .A2(n7451), .ZN(n8324) );
  NAND2_X1 U9503 ( .A1(n13468), .A2(n6516), .ZN(n7176) );
  NAND2_X1 U9504 ( .A1(n10271), .A2(n10270), .ZN(n10273) );
  NAND2_X1 U9505 ( .A1(n9947), .A2(n9946), .ZN(n10416) );
  NAND2_X1 U9506 ( .A1(n8982), .A2(n12345), .ZN(n10110) );
  OR2_X1 U9507 ( .A1(n12481), .A2(n10834), .ZN(n8544) );
  NAND2_X1 U9508 ( .A1(n11787), .A2(n11786), .ZN(n13486) );
  NAND2_X1 U9509 ( .A1(n8993), .A2(n12411), .ZN(n12870) );
  NAND2_X1 U9510 ( .A1(n8990), .A2(n12390), .ZN(n11380) );
  INV_X1 U9511 ( .A(n8510), .ZN(n8509) );
  NAND2_X1 U9512 ( .A1(n11496), .A2(n11495), .ZN(n11785) );
  INV_X1 U9513 ( .A(n9625), .ZN(n9629) );
  NAND2_X1 U9514 ( .A1(n9630), .A2(n9629), .ZN(n9947) );
  NAND2_X1 U9515 ( .A1(n10526), .A2(n10525), .ZN(n10524) );
  NAND2_X1 U9516 ( .A1(n8375), .A2(n13983), .ZN(n8343) );
  XNOR2_X2 U9517 ( .A(n8454), .B(n8453), .ZN(n8459) );
  NOR2_X2 U9518 ( .A1(n10830), .A2(n10024), .ZN(n12333) );
  XNOR2_X2 U9519 ( .A(n12560), .B(n10147), .ZN(n10112) );
  NOR2_X2 U9520 ( .A1(n14914), .A2(n11383), .ZN(n14913) );
  NAND2_X1 U9521 ( .A1(n10493), .A2(n7189), .ZN(n7187) );
  XNOR2_X2 U9522 ( .A(n9154), .B(n9174), .ZN(n9158) );
  NOR2_X2 U9523 ( .A1(n14248), .A2(n14232), .ZN(n7202) );
  NOR2_X2 U9524 ( .A1(n10034), .A2(n11862), .ZN(n10513) );
  NOR2_X2 U9525 ( .A1(n14132), .A2(n14290), .ZN(n7205) );
  NOR2_X2 U9526 ( .A1(n14151), .A2(n14156), .ZN(n7207) );
  NAND2_X1 U9527 ( .A1(n11838), .A2(n11848), .ZN(n7209) );
  AND2_X1 U9528 ( .A1(n11871), .A2(n6608), .ZN(n7210) );
  NAND2_X1 U9529 ( .A1(n11872), .A2(n7210), .ZN(n7211) );
  NAND2_X1 U9530 ( .A1(n7211), .A2(n7212), .ZN(n11878) );
  OR2_X1 U9531 ( .A1(n7219), .A2(n11997), .ZN(n7218) );
  INV_X1 U9532 ( .A(n11996), .ZN(n7219) );
  NAND2_X1 U9533 ( .A1(n11978), .A2(n7223), .ZN(n7222) );
  INV_X1 U9534 ( .A(n11979), .ZN(n7224) );
  NAND2_X1 U9535 ( .A1(n7225), .A2(n7226), .ZN(n11918) );
  NAND3_X1 U9536 ( .A1(n11910), .A2(n11909), .A3(n6606), .ZN(n7225) );
  NAND2_X1 U9537 ( .A1(n11960), .A2(n7232), .ZN(n7231) );
  AOI21_X1 U9538 ( .B1(n7234), .B2(n7232), .A(n7230), .ZN(n7229) );
  NAND2_X1 U9539 ( .A1(n7237), .A2(n7236), .ZN(n11869) );
  INV_X1 U9540 ( .A(n11864), .ZN(n7239) );
  NAND2_X1 U9541 ( .A1(n9287), .A2(n7242), .ZN(n7241) );
  OR2_X2 U9542 ( .A1(n14476), .A2(n14477), .ZN(n14473) );
  NAND2_X1 U9543 ( .A1(n7247), .A2(n11452), .ZN(n14476) );
  NAND2_X1 U9544 ( .A1(n11448), .A2(n11447), .ZN(n7247) );
  NAND2_X1 U9545 ( .A1(n10446), .A2(n7250), .ZN(n7249) );
  NAND2_X1 U9546 ( .A1(n7251), .A2(n10660), .ZN(n7248) );
  INV_X1 U9547 ( .A(n7270), .ZN(n13833) );
  NAND2_X1 U9548 ( .A1(n7272), .A2(n7271), .ZN(n9065) );
  NAND2_X2 U9549 ( .A1(n7285), .A2(n11506), .ZN(n9822) );
  XNOR2_X1 U9550 ( .A(n7286), .B(n7708), .ZN(n9799) );
  NAND3_X1 U9551 ( .A1(n7533), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7293) );
  NAND2_X1 U9552 ( .A1(n8156), .A2(n7313), .ZN(n7310) );
  OAI21_X2 U9553 ( .B1(n12822), .B2(n7319), .A(n7316), .ZN(n12798) );
  INV_X1 U9554 ( .A(n12881), .ZN(n7325) );
  NAND2_X1 U9555 ( .A1(n11021), .A2(n7333), .ZN(n7331) );
  NAND2_X1 U9556 ( .A1(n7331), .A2(n7332), .ZN(n11299) );
  NAND2_X1 U9557 ( .A1(n10776), .A2(n6598), .ZN(n10955) );
  OR2_X2 U9558 ( .A1(n12848), .A2(n7070), .ZN(n12846) );
  NAND2_X1 U9559 ( .A1(n10113), .A2(n6537), .ZN(n7345) );
  AOI21_X1 U9560 ( .B1(n12745), .B2(n7350), .A(n7348), .ZN(n12717) );
  OR2_X1 U9561 ( .A1(n12745), .A2(n8897), .ZN(n7352) );
  NAND2_X1 U9562 ( .A1(n12717), .A2(n12723), .ZN(n12716) );
  NAND2_X1 U9563 ( .A1(n8937), .A2(n6605), .ZN(n8510) );
  NAND2_X1 U9564 ( .A1(n12214), .A2(n6588), .ZN(n7354) );
  OAI211_X1 U9565 ( .C1(n12214), .C2(n7357), .A(n7355), .B(n7354), .ZN(n12203)
         );
  NAND2_X1 U9566 ( .A1(n12214), .A2(n7363), .ZN(n7359) );
  INV_X1 U9567 ( .A(n12195), .ZN(n7366) );
  NAND2_X1 U9568 ( .A1(n7372), .A2(n10165), .ZN(n7371) );
  OAI211_X1 U9569 ( .C1(n10155), .C2(n7373), .A(n7371), .B(n10287), .ZN(n10292) );
  NAND2_X1 U9570 ( .A1(n11368), .A2(n12554), .ZN(n7376) );
  NAND2_X1 U9571 ( .A1(n11327), .A2(n11326), .ZN(n11329) );
  XNOR2_X1 U9572 ( .A(n12150), .B(n12148), .ZN(n12272) );
  NAND3_X1 U9573 ( .A1(n8946), .A2(n7389), .A3(n7387), .ZN(n11343) );
  OAI21_X1 U9574 ( .B1(n12062), .B2(n7391), .A(n9913), .ZN(n9588) );
  NAND2_X1 U9575 ( .A1(n12062), .A2(n7391), .ZN(n9913) );
  AND2_X1 U9576 ( .A1(n11852), .A2(n11847), .ZN(n7391) );
  NAND2_X1 U9577 ( .A1(n11142), .A2(n7395), .ZN(n7392) );
  NAND2_X1 U9578 ( .A1(n14101), .A2(n6504), .ZN(n7398) );
  NAND2_X1 U9579 ( .A1(n14101), .A2(n6596), .ZN(n7401) );
  NAND2_X1 U9580 ( .A1(n14179), .A2(n7406), .ZN(n7405) );
  NOR2_X4 U9581 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9092) );
  NAND2_X1 U9582 ( .A1(n14215), .A2(n7411), .ZN(n14195) );
  NAND3_X1 U9583 ( .A1(n7272), .A2(n9147), .A3(n9061), .ZN(n9152) );
  NAND2_X1 U9584 ( .A1(n10750), .A2(n6505), .ZN(n7419) );
  NAND2_X1 U9586 ( .A1(n10403), .A2(n7427), .ZN(n7426) );
  AND2_X1 U9587 ( .A1(n7433), .A2(n7434), .ZN(n13386) );
  INV_X1 U9588 ( .A(n13561), .ZN(n7439) );
  NAND2_X1 U9589 ( .A1(n13477), .A2(n11815), .ZN(n13444) );
  AOI21_X1 U9590 ( .B1(n7444), .B2(n7443), .A(n6510), .ZN(n7442) );
  NAND3_X1 U9591 ( .A1(n7654), .A2(n7653), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n7447) );
  NAND2_X1 U9592 ( .A1(n10910), .A2(n7458), .ZN(n11003) );
  OAI21_X1 U9593 ( .B1(n13098), .B2(n7460), .A(n7461), .ZN(n11615) );
  XNOR2_X1 U9594 ( .A(n7474), .B(n13066), .ZN(n13071) );
  OAI21_X1 U9595 ( .B1(n10102), .B2(n7478), .A(n7475), .ZN(n10260) );
  NAND2_X1 U9596 ( .A1(n13626), .A2(n7650), .ZN(n13630) );
  NAND2_X1 U9597 ( .A1(n10087), .A2(n7481), .ZN(n10101) );
  NAND2_X1 U9598 ( .A1(n11237), .A2(n7482), .ZN(n11265) );
  INV_X1 U9599 ( .A(n7490), .ZN(n13106) );
  NAND2_X1 U9600 ( .A1(n10672), .A2(n6597), .ZN(n10862) );
  NAND2_X1 U9601 ( .A1(n10862), .A2(n10860), .ZN(n10858) );
  NAND2_X1 U9602 ( .A1(n7691), .A2(n7690), .ZN(n7492) );
  NAND2_X1 U9603 ( .A1(n8120), .A2(n7498), .ZN(n7495) );
  INV_X1 U9604 ( .A(n7886), .ZN(n7506) );
  NAND3_X1 U9605 ( .A1(n7766), .A2(n6514), .A3(n6603), .ZN(n7507) );
  NAND2_X1 U9606 ( .A1(n7507), .A2(n6600), .ZN(n7807) );
  INV_X1 U9607 ( .A(n7787), .ZN(n7508) );
  NAND2_X1 U9608 ( .A1(n7509), .A2(n7510), .ZN(n8036) );
  NAND2_X1 U9609 ( .A1(n7851), .A2(n7512), .ZN(n7511) );
  NAND2_X1 U9610 ( .A1(n7847), .A2(n7514), .ZN(n7513) );
  NAND3_X1 U9611 ( .A1(n7959), .A2(n6513), .A3(n6586), .ZN(n7519) );
  NAND2_X1 U9612 ( .A1(n7521), .A2(n7522), .ZN(n7765) );
  NAND3_X1 U9613 ( .A1(n7729), .A2(n7728), .A3(n6607), .ZN(n7521) );
  XNOR2_X1 U9614 ( .A(n11799), .B(n11798), .ZN(n11805) );
  NAND2_X1 U9615 ( .A1(n11901), .A2(n11900), .ZN(n11903) );
  NAND2_X1 U9616 ( .A1(n11743), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U9617 ( .A1(n8862), .A2(n6543), .ZN(n8864) );
  NAND2_X1 U9618 ( .A1(n13302), .A2(n13304), .ZN(n13301) );
  INV_X1 U9619 ( .A(n6486), .ZN(n8239) );
  XNOR2_X2 U9620 ( .A(n12563), .B(n14937), .ZN(n14942) );
  OR2_X1 U9621 ( .A1(n6499), .A2(n8904), .ZN(n12486) );
  NAND2_X2 U9622 ( .A1(n8828), .A2(n8827), .ZN(n12822) );
  NAND4_X2 U9623 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n13949)
         );
  XNOR2_X1 U9624 ( .A(n8156), .B(n8155), .ZN(n13635) );
  CLKBUF_X1 U9625 ( .A(n13123), .Z(n13125) );
  XNOR2_X1 U9626 ( .A(n10047), .B(n10048), .ZN(n13083) );
  NOR2_X2 U9627 ( .A1(n14199), .A2(n14314), .ZN(n14187) );
  AOI21_X1 U9628 ( .B1(n8099), .B2(n8098), .A(n8097), .ZN(n8120) );
  XNOR2_X2 U9629 ( .A(n13947), .B(n10236), .ZN(n11854) );
  NAND2_X1 U9630 ( .A1(n9618), .A2(n14842), .ZN(n14884) );
  XNOR2_X1 U9631 ( .A(n12500), .B(n12694), .ZN(n7525) );
  NAND2_X1 U9632 ( .A1(n8168), .A2(n8167), .ZN(n13192) );
  INV_X1 U9633 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10126) );
  INV_X1 U9634 ( .A(n6748), .ZN(n9622) );
  AND2_X1 U9635 ( .A1(n7581), .A2(n7580), .ZN(n7527) );
  INV_X1 U9636 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10128) );
  AND2_X1 U9637 ( .A1(n7577), .A2(n7576), .ZN(n7528) );
  AOI21_X1 U9638 ( .B1(n6667), .B2(n14847), .A(n10183), .ZN(n7673) );
  INV_X1 U9639 ( .A(n7747), .ZN(n7748) );
  OAI21_X1 U9640 ( .B1(n11921), .B2(n12079), .A(n11925), .ZN(n11922) );
  NAND2_X1 U9641 ( .A1(n11946), .A2(n14246), .ZN(n11947) );
  INV_X1 U9642 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8443) );
  OAI21_X1 U9643 ( .B1(n13513), .B2(n8214), .A(n8265), .ZN(n8274) );
  INV_X1 U9644 ( .A(n12505), .ZN(n8661) );
  NAND2_X1 U9645 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  INV_X1 U9646 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9037) );
  INV_X1 U9647 ( .A(n8791), .ZN(n8805) );
  AND2_X1 U9648 ( .A1(n8124), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8140) );
  INV_X1 U9649 ( .A(n8110), .ZN(n8108) );
  INV_X1 U9650 ( .A(n8006), .ZN(n7642) );
  INV_X1 U9651 ( .A(n14860), .ZN(n10406) );
  INV_X1 U9652 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7646) );
  AND2_X1 U9653 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n11719), .ZN(n11718) );
  NOR2_X1 U9654 ( .A1(n11650), .A2(n11649), .ZN(n11663) );
  INV_X1 U9655 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9054) );
  INV_X1 U9656 ( .A(n7831), .ZN(n7561) );
  INV_X1 U9657 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7545) );
  OR2_X1 U9658 ( .A1(n14953), .A2(n9037), .ZN(n9038) );
  NOR2_X1 U9659 ( .A1(n8792), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8791) );
  OR2_X1 U9660 ( .A1(n9170), .A2(n8969), .ZN(n9009) );
  NAND2_X1 U9661 ( .A1(n8829), .A2(n11660), .ZN(n8498) );
  NAND2_X1 U9662 ( .A1(n8785), .A2(n8783), .ZN(n8494) );
  NAND2_X1 U9663 ( .A1(n11594), .A2(n11593), .ZN(n11595) );
  INV_X1 U9664 ( .A(n10676), .ZN(n10673) );
  INV_X1 U9665 ( .A(n10091), .ZN(n10088) );
  INV_X1 U9666 ( .A(n7895), .ZN(n7639) );
  OR2_X1 U9667 ( .A1(n8162), .A2(n8141), .ZN(n8204) );
  NAND2_X1 U9668 ( .A1(n8108), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8126) );
  OR2_X1 U9669 ( .A1(n8046), .A2(n7644), .ZN(n8067) );
  NAND2_X1 U9670 ( .A1(n7640), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9671 ( .A1(n6485), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7664) );
  NOR2_X1 U9672 ( .A1(n13532), .A2(n13192), .ZN(n11818) );
  NAND2_X1 U9673 ( .A1(n8085), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U9674 ( .A1(n7642), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8025) );
  INV_X1 U9675 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7962) );
  INV_X1 U9676 ( .A(n13704), .ZN(n13705) );
  AND2_X1 U9677 ( .A1(n11718), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11740) );
  INV_X1 U9678 ( .A(n11707), .ZN(n11719) );
  INV_X1 U9679 ( .A(n11697), .ZN(n11686) );
  INV_X1 U9680 ( .A(n14216), .ZN(n11657) );
  AND3_X1 U9681 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U9682 ( .A1(n9148), .A2(n9050), .ZN(n9150) );
  NAND2_X1 U9683 ( .A1(n7589), .A2(n7588), .ZN(n7592) );
  NAND2_X1 U9684 ( .A1(n7569), .A2(n8703), .ZN(n7573) );
  INV_X1 U9685 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U9686 ( .A1(n8364), .A2(n8365), .ZN(n8355) );
  INV_X1 U9687 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9751) );
  INV_X1 U9688 ( .A(n12763), .ZN(n12218) );
  AND4_X1 U9689 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8764), .ZN(n12299)
         );
  INV_X1 U9690 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9663) );
  INV_X1 U9691 ( .A(n14896), .ZN(n14916) );
  AND2_X1 U9692 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  INV_X1 U9693 ( .A(n12551), .ZN(n12812) );
  AND2_X1 U9694 ( .A1(n8762), .A2(n8761), .ZN(n8776) );
  NAND2_X1 U9695 ( .A1(n12556), .A2(n12385), .ZN(n12388) );
  AND2_X1 U9696 ( .A1(n9011), .A2(n12539), .ZN(n12861) );
  NAND2_X1 U9697 ( .A1(n8932), .A2(n12446), .ZN(n14944) );
  NAND2_X1 U9698 ( .A1(n9127), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8474) );
  AND2_X1 U9699 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  AND2_X1 U9700 ( .A1(n6682), .A2(n9497), .ZN(n10063) );
  OR2_X1 U9701 ( .A1(n8067), .A2(n13148), .ZN(n8086) );
  AND2_X1 U9702 ( .A1(n8160), .A2(n8127), .ZN(n13350) );
  OR2_X1 U9703 ( .A1(n8025), .A2(n8024), .ZN(n8044) );
  AND2_X1 U9704 ( .A1(n9344), .A2(n13632), .ZN(n9361) );
  INV_X1 U9705 ( .A(n13198), .ZN(n13117) );
  INV_X1 U9706 ( .A(n13437), .ZN(n13447) );
  INV_X1 U9707 ( .A(n11814), .ZN(n13480) );
  CLKBUF_X1 U9708 ( .A(n10043), .Z(n14849) );
  AND2_X1 U9709 ( .A1(n11686), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11708) );
  NOR2_X1 U9710 ( .A1(n10641), .A2(n10976), .ZN(n10717) );
  NAND2_X1 U9711 ( .A1(n13703), .A2(n13705), .ZN(n13706) );
  OR2_X1 U9712 ( .A1(n9298), .A2(n12102), .ZN(n14481) );
  NAND2_X1 U9713 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  AND3_X1 U9714 ( .A1(n9185), .A2(n9184), .A3(n9183), .ZN(n13849) );
  INV_X1 U9715 ( .A(n14647), .ZN(n14175) );
  OR2_X1 U9716 ( .A1(n9315), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9961) );
  OR2_X1 U9717 ( .A1(n12706), .A2(n8464), .ZN(n12724) );
  INV_X1 U9718 ( .A(n12311), .ZN(n12280) );
  AND4_X1 U9719 ( .A1(n12486), .A2(n12485), .A3(n12484), .A4(n12483), .ZN(
        n12709) );
  AND4_X1 U9720 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n12292)
         );
  AND4_X1 U9721 ( .A1(n8838), .A2(n8837), .A3(n8836), .A4(n8835), .ZN(n12811)
         );
  INV_X1 U9722 ( .A(n12888), .ZN(n14940) );
  AND3_X1 U9723 ( .A1(n9010), .A2(n8970), .A3(n9015), .ZN(n9031) );
  AND2_X1 U9724 ( .A1(n12417), .A2(n12416), .ZN(n12863) );
  OR2_X1 U9725 ( .A1(n14993), .A2(n15009), .ZN(n14959) );
  OR2_X1 U9726 ( .A1(n9335), .A2(n9334), .ZN(n9344) );
  OR2_X1 U9727 ( .A1(n13336), .A2(n8239), .ZN(n8168) );
  INV_X1 U9728 ( .A(n8027), .ZN(n8261) );
  NOR2_X1 U9729 ( .A1(n9763), .A2(n9762), .ZN(n13223) );
  AND2_X1 U9730 ( .A1(n14809), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15226) );
  NAND2_X1 U9731 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  INV_X1 U9732 ( .A(n11060), .ZN(n11066) );
  INV_X1 U9733 ( .A(n13498), .ZN(n13483) );
  AND2_X1 U9734 ( .A1(n14849), .A2(n14871), .ZN(n14875) );
  AND2_X1 U9735 ( .A1(n14844), .A2(n9485), .ZN(n9618) );
  AND2_X1 U9736 ( .A1(n7790), .A2(n7772), .ZN(n9355) );
  INV_X1 U9737 ( .A(n14481), .ZN(n14506) );
  AND2_X1 U9738 ( .A1(n11730), .A2(n11729), .ZN(n14099) );
  AND4_X1 U9739 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n13674) );
  INV_X1 U9740 ( .A(n14548), .ZN(n14617) );
  OAI21_X1 U9741 ( .B1(n14084), .B2(n14085), .A(n14083), .ZN(n14276) );
  INV_X1 U9742 ( .A(n12082), .ZN(n14241) );
  AND2_X1 U9743 ( .A1(n11916), .A2(n11924), .ZN(n12079) );
  AND2_X1 U9744 ( .A1(n14671), .A2(n14044), .ZN(n14654) );
  OR2_X1 U9745 ( .A1(n10226), .A2(n10225), .ZN(n14662) );
  AND2_X1 U9746 ( .A1(n14707), .A2(n14708), .ZN(n14677) );
  AND3_X1 U9747 ( .A1(n9565), .A2(n10222), .A3(n10226), .ZN(n9593) );
  AND2_X1 U9748 ( .A1(n9822), .A2(n9122), .ZN(n9297) );
  NAND2_X1 U9749 ( .A1(n7608), .A2(n7607), .ZN(n8061) );
  AND2_X1 U9750 ( .A1(n9614), .A2(n9435), .ZN(n14557) );
  AND2_X1 U9751 ( .A1(n9142), .A2(n9141), .ZN(n10709) );
  AND2_X1 U9752 ( .A1(n9662), .A2(n9661), .ZN(n14896) );
  INV_X1 U9753 ( .A(n9993), .ZN(n12288) );
  AND4_X1 U9754 ( .A1(n12486), .A2(n8911), .A3(n8910), .A4(n8909), .ZN(n12720)
         );
  INV_X1 U9755 ( .A(n12292), .ZN(n12778) );
  INV_X1 U9756 ( .A(n12850), .ZN(n12873) );
  INV_X1 U9757 ( .A(n11274), .ZN(n12555) );
  INV_X1 U9758 ( .A(P3_U3897), .ZN(n12562) );
  OR2_X1 U9759 ( .A1(n9672), .A2(n9664), .ZN(n14934) );
  OR2_X1 U9760 ( .A1(n9035), .A2(n9034), .ZN(n12903) );
  OR2_X1 U9761 ( .A1(n14955), .A2(n9033), .ZN(n12892) );
  INV_X1 U9762 ( .A(n15025), .ZN(n15023) );
  AND2_X2 U9763 ( .A1(n9031), .A2(n8977), .ZN(n15025) );
  OR2_X1 U9764 ( .A1(n15012), .A2(n14449), .ZN(n13033) );
  INV_X2 U9765 ( .A(n15012), .ZN(n15010) );
  AND2_X1 U9766 ( .A1(n9021), .A2(n9020), .ZN(n15012) );
  AND2_X1 U9767 ( .A1(n8952), .A2(n8951), .ZN(n13040) );
  INV_X1 U9768 ( .A(n12690), .ZN(n12694) );
  OR2_X1 U9769 ( .A1(n8718), .A2(n8717), .ZN(n12582) );
  INV_X1 U9770 ( .A(n13162), .ZN(n13187) );
  NAND2_X1 U9771 ( .A1(n8212), .A2(n8211), .ZN(n13190) );
  INV_X1 U9772 ( .A(n13126), .ZN(n13194) );
  INV_X1 U9773 ( .A(n13476), .ZN(n13392) );
  NAND2_X1 U9774 ( .A1(n9618), .A2(n9617), .ZN(n14893) );
  INV_X1 U9775 ( .A(n14839), .ZN(n14840) );
  INV_X1 U9776 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9965) );
  INV_X1 U9777 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9069) );
  INV_X1 U9778 ( .A(n14308), .ZN(n14174) );
  INV_X1 U9779 ( .A(n14502), .ZN(n13907) );
  CLKBUF_X1 U9780 ( .A(P1_U4016), .Z(n13948) );
  INV_X1 U9781 ( .A(n14753), .ZN(n14751) );
  AND3_X1 U9782 ( .A1(n14524), .A2(n14523), .A3(n14522), .ZN(n14527) );
  INV_X1 U9783 ( .A(n14742), .ZN(n14740) );
  AND2_X1 U9784 ( .A1(n9146), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9122) );
  BUF_X1 U9785 ( .A(n9180), .Z(n14373) );
  INV_X1 U9786 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9436) );
  AND2_X1 U9787 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9335), .ZN(P2_U3947) );
  INV_X1 U9788 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9518) );
  AND2_X1 U9789 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7534) );
  NAND2_X1 U9790 ( .A1(n9068), .A2(n7534), .ZN(n9258) );
  NAND3_X1 U9791 ( .A1(n11682), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n7535) );
  NAND2_X1 U9792 ( .A1(n9258), .A2(n7535), .ZN(n7676) );
  INV_X1 U9793 ( .A(SI_1_), .ZN(n9081) );
  NOR2_X1 U9794 ( .A1(n7536), .A2(n9081), .ZN(n7537) );
  INV_X1 U9795 ( .A(SI_2_), .ZN(n9077) );
  NAND2_X1 U9796 ( .A1(n7538), .A2(SI_2_), .ZN(n7539) );
  XNOR2_X1 U9797 ( .A(n7541), .B(SI_3_), .ZN(n7708) );
  INV_X1 U9798 ( .A(n7708), .ZN(n7540) );
  NAND2_X1 U9799 ( .A1(n7541), .A2(SI_3_), .ZN(n7542) );
  XNOR2_X1 U9800 ( .A(n7547), .B(SI_4_), .ZN(n7731) );
  INV_X1 U9801 ( .A(n7731), .ZN(n7546) );
  NAND2_X1 U9802 ( .A1(n7547), .A2(SI_4_), .ZN(n7548) );
  XNOR2_X1 U9803 ( .A(n7550), .B(SI_5_), .ZN(n7749) );
  INV_X1 U9804 ( .A(n7749), .ZN(n7549) );
  NAND2_X1 U9805 ( .A1(n7550), .A2(SI_5_), .ZN(n7551) );
  MUX2_X1 U9806 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9517), .Z(n7554) );
  NAND2_X1 U9807 ( .A1(n7768), .A2(n7553), .ZN(n7556) );
  NAND2_X1 U9808 ( .A1(n7554), .A2(SI_6_), .ZN(n7555) );
  NAND2_X1 U9809 ( .A1(n7558), .A2(SI_7_), .ZN(n7559) );
  MUX2_X1 U9810 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9517), .Z(n7560) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9517), .Z(n7562) );
  NAND2_X1 U9812 ( .A1(n7562), .A2(SI_9_), .ZN(n7563) );
  NAND2_X1 U9813 ( .A1(n7564), .A2(n7563), .ZN(n7853) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9517), .Z(n7566) );
  NAND2_X1 U9815 ( .A1(n7853), .A2(n7565), .ZN(n7568) );
  NAND2_X1 U9816 ( .A1(n7566), .A2(SI_10_), .ZN(n7567) );
  MUX2_X1 U9817 ( .A(n8486), .B(n9207), .S(n9517), .Z(n7569) );
  INV_X1 U9818 ( .A(SI_11_), .ZN(n8703) );
  INV_X1 U9819 ( .A(n7569), .ZN(n7570) );
  NAND2_X1 U9820 ( .A1(n7570), .A2(SI_11_), .ZN(n7571) );
  MUX2_X1 U9821 ( .A(n9316), .B(n9314), .S(n9517), .Z(n7574) );
  INV_X1 U9822 ( .A(SI_12_), .ZN(n9124) );
  INV_X1 U9823 ( .A(n7574), .ZN(n7575) );
  NAND2_X1 U9824 ( .A1(n7575), .A2(SI_12_), .ZN(n7576) );
  MUX2_X1 U9825 ( .A(n9436), .B(n9429), .S(n9517), .Z(n7578) );
  INV_X1 U9826 ( .A(n7578), .ZN(n7579) );
  NAND2_X1 U9827 ( .A1(n7579), .A2(SI_13_), .ZN(n7580) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9517), .Z(n7924) );
  MUX2_X1 U9829 ( .A(n7027), .B(n9965), .S(n9517), .Z(n7584) );
  INV_X1 U9830 ( .A(SI_15_), .ZN(n7583) );
  NAND2_X1 U9831 ( .A1(n7584), .A2(n7583), .ZN(n7587) );
  INV_X1 U9832 ( .A(n7584), .ZN(n7585) );
  NAND2_X1 U9833 ( .A1(n7585), .A2(SI_15_), .ZN(n7586) );
  MUX2_X1 U9834 ( .A(n10126), .B(n10128), .S(n9517), .Z(n7589) );
  INV_X1 U9835 ( .A(SI_16_), .ZN(n7588) );
  INV_X1 U9836 ( .A(n7589), .ZN(n7590) );
  NAND2_X1 U9837 ( .A1(n7590), .A2(SI_16_), .ZN(n7591) );
  INV_X1 U9838 ( .A(SI_17_), .ZN(n9549) );
  INV_X1 U9839 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10304) );
  INV_X1 U9840 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10306) );
  MUX2_X1 U9841 ( .A(n10304), .B(n10306), .S(n9517), .Z(n7979) );
  MUX2_X1 U9842 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9517), .Z(n8000) );
  NOR2_X1 U9843 ( .A1(n8000), .A2(SI_18_), .ZN(n7595) );
  MUX2_X1 U9844 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9517), .Z(n7596) );
  XNOR2_X1 U9845 ( .A(n7596), .B(SI_19_), .ZN(n8019) );
  INV_X1 U9846 ( .A(n8000), .ZN(n8017) );
  INV_X1 U9847 ( .A(SI_18_), .ZN(n9641) );
  NOR2_X1 U9848 ( .A1(n8017), .A2(n9641), .ZN(n7593) );
  NOR2_X1 U9849 ( .A1(n8019), .A2(n7593), .ZN(n7594) );
  INV_X1 U9850 ( .A(n7596), .ZN(n7597) );
  INV_X1 U9851 ( .A(SI_19_), .ZN(n9774) );
  INV_X1 U9852 ( .A(SI_20_), .ZN(n10384) );
  NAND2_X1 U9853 ( .A1(n7603), .A2(n10384), .ZN(n7598) );
  NAND2_X1 U9854 ( .A1(n7600), .A2(n7598), .ZN(n8039) );
  INV_X1 U9855 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11660) );
  INV_X1 U9856 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10923) );
  MUX2_X1 U9857 ( .A(n11660), .B(n10923), .S(n9517), .Z(n8038) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9517), .Z(n7599) );
  NAND2_X1 U9859 ( .A1(n7599), .A2(SI_21_), .ZN(n8060) );
  OAI21_X1 U9860 ( .B1(SI_21_), .B2(n7599), .A(n8060), .ZN(n7606) );
  AND2_X1 U9861 ( .A1(n7600), .A2(n7606), .ZN(n7601) );
  NAND2_X1 U9862 ( .A1(n7604), .A2(SI_20_), .ZN(n7602) );
  NOR2_X1 U9863 ( .A1(n7604), .A2(SI_20_), .ZN(n7605) );
  NOR2_X1 U9864 ( .A1(n7606), .A2(n7605), .ZN(n7607) );
  NAND2_X1 U9865 ( .A1(n7609), .A2(n8061), .ZN(n11672) );
  NOR2_X1 U9866 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7612) );
  NOR2_X2 U9867 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7611) );
  NOR2_X2 U9868 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7610) );
  NOR2_X1 U9869 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7619) );
  NOR2_X1 U9870 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7618) );
  NOR2_X1 U9871 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7617) );
  NOR2_X1 U9872 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7616) );
  INV_X1 U9873 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7622) );
  INV_X1 U9874 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15043) );
  OR2_X1 U9875 ( .A1(n6653), .A2(n15043), .ZN(n7624) );
  INV_X1 U9876 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7626) );
  INV_X1 U9877 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U9878 ( .A1(n7630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7631) );
  OR2_X1 U9879 ( .A1(n7632), .A2(n7709), .ZN(n7633) );
  XNOR2_X2 U9880 ( .A(n7633), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U9881 ( .A1(n13561), .A2(n8215), .ZN(n7661) );
  NAND2_X1 U9882 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7754) );
  INV_X1 U9883 ( .A(n7754), .ZN(n7634) );
  NAND2_X1 U9884 ( .A1(n7634), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7777) );
  INV_X1 U9885 ( .A(n7777), .ZN(n7635) );
  NAND2_X1 U9886 ( .A1(n7635), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7796) );
  INV_X1 U9887 ( .A(n7796), .ZN(n7636) );
  NAND2_X1 U9888 ( .A1(n7636), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7822) );
  INV_X1 U9889 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U9890 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7638) );
  INV_X1 U9891 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7929) );
  INV_X1 U9892 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11404) );
  INV_X1 U9893 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13118) );
  INV_X1 U9894 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8024) );
  INV_X1 U9895 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9896 ( .A1(n8046), .A2(n7644), .ZN(n7645) );
  NAND2_X1 U9897 ( .A1(n8067), .A2(n7645), .ZN(n13417) );
  NAND2_X1 U9898 ( .A1(n7648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7647) );
  MUX2_X1 U9899 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7647), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7650) );
  INV_X1 U9900 ( .A(n7649), .ZN(n13626) );
  INV_X1 U9901 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7651) );
  OR2_X1 U9902 ( .A1(n13417), .A2(n8239), .ZN(n7659) );
  INV_X1 U9903 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15185) );
  INV_X2 U9904 ( .A(n7969), .ZN(n8256) );
  NAND2_X1 U9905 ( .A1(n8256), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U9906 ( .A1(n8206), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7655) );
  OAI211_X1 U9907 ( .C1(n15185), .C2(n8261), .A(n7656), .B(n7655), .ZN(n7657)
         );
  INV_X1 U9908 ( .A(n7657), .ZN(n7658) );
  NAND2_X1 U9909 ( .A1(n7659), .A2(n7658), .ZN(n13438) );
  NAND2_X1 U9910 ( .A1(n13438), .A2(n8214), .ZN(n7660) );
  NAND2_X1 U9911 ( .A1(n7661), .A2(n7660), .ZN(n8057) );
  NAND2_X1 U9912 ( .A1(n7683), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7663) );
  NAND2_X1 U9913 ( .A1(n7682), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7662) );
  INV_X1 U9914 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U9915 ( .A1(n9517), .A2(SI_0_), .ZN(n7667) );
  INV_X1 U9916 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n15032) );
  XNOR2_X1 U9917 ( .A(n7667), .B(n15032), .ZN(n13639) );
  MUX2_X1 U9918 ( .A(n9460), .B(n13639), .S(n7678), .Z(n14847) );
  INV_X1 U9919 ( .A(n7673), .ZN(n7671) );
  NAND2_X1 U9920 ( .A1(n6667), .A2(n8093), .ZN(n7670) );
  NAND3_X1 U9921 ( .A1(n7671), .A2(n7670), .A3(n7669), .ZN(n7675) );
  NAND2_X1 U9922 ( .A1(n8263), .A2(n11500), .ZN(n7672) );
  NAND2_X1 U9923 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NAND2_X1 U9924 ( .A1(n7675), .A2(n7674), .ZN(n7689) );
  XNOR2_X1 U9925 ( .A(n7677), .B(n7676), .ZN(n9516) );
  NAND2_X1 U9926 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7679) );
  MUX2_X1 U9927 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7679), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7681) );
  INV_X1 U9928 ( .A(n7713), .ZN(n7680) );
  NAND2_X1 U9929 ( .A1(n7681), .A2(n7680), .ZN(n9458) );
  INV_X1 U9930 ( .A(n9458), .ZN(n9466) );
  NAND2_X1 U9931 ( .A1(n8027), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9932 ( .A1(n7682), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9933 ( .A1(n7683), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7684) );
  OAI22_X1 U9934 ( .A1(n9622), .A2(n8093), .B1(n9504), .B2(n6517), .ZN(n7687)
         );
  OAI21_X1 U9935 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7691) );
  NAND2_X1 U9936 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  NAND2_X1 U9937 ( .A1(n8143), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U9938 ( .A1(n8027), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9939 ( .A1(n8032), .A2(n13212), .ZN(n7705) );
  NOR2_X1 U9940 ( .A1(n7713), .A2(n7709), .ZN(n7698) );
  MUX2_X1 U9941 ( .A(n7709), .B(n7698), .S(P2_IR_REG_2__SCAN_IN), .Z(n7701) );
  INV_X1 U9942 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7699) );
  NAND2_X1 U9943 ( .A1(n7713), .A2(n7699), .ZN(n7710) );
  INV_X1 U9944 ( .A(n7710), .ZN(n7700) );
  NAND2_X1 U9945 ( .A1(n9332), .A2(n9383), .ZN(n7702) );
  NAND2_X1 U9946 ( .A1(n8093), .A2(n13158), .ZN(n7704) );
  INV_X1 U9947 ( .A(n13158), .ZN(n10397) );
  NAND2_X1 U9948 ( .A1(n13212), .A2(n8093), .ZN(n7706) );
  OAI21_X1 U9949 ( .B1(n8093), .B2(n10397), .A(n7706), .ZN(n7707) );
  NAND2_X1 U9950 ( .A1(n9799), .A2(n8236), .ZN(n7716) );
  NAND2_X1 U9951 ( .A1(n7710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7711) );
  MUX2_X1 U9952 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7711), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n7714) );
  NAND2_X1 U9953 ( .A1(n7713), .A2(n7712), .ZN(n7732) );
  AOI22_X1 U9954 ( .A1(n8021), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9332), .B2(
        n9351), .ZN(n7715) );
  AND2_X2 U9955 ( .A1(n7716), .A2(n7715), .ZN(n14860) );
  INV_X1 U9956 ( .A(n6517), .ZN(n8093) );
  NAND2_X1 U9957 ( .A1(n8257), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9958 ( .A1(n7794), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7719) );
  INV_X1 U9959 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U9960 ( .A1(n6485), .A2(n10411), .ZN(n7718) );
  NAND2_X1 U9961 ( .A1(n8027), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9962 ( .A1(n13211), .A2(n8093), .ZN(n7721) );
  OAI21_X1 U9963 ( .B1(n14860), .B2(n8093), .A(n7721), .ZN(n7725) );
  NAND2_X1 U9964 ( .A1(n7724), .A2(n7725), .ZN(n7723) );
  INV_X1 U9965 ( .A(n13211), .ZN(n9951) );
  OAI22_X1 U9966 ( .A1(n9951), .A2(n8214), .B1(n14860), .B2(n7820), .ZN(n7722)
         );
  NAND2_X1 U9967 ( .A1(n7723), .A2(n7722), .ZN(n7729) );
  INV_X1 U9968 ( .A(n7724), .ZN(n7727) );
  INV_X1 U9969 ( .A(n7725), .ZN(n7726) );
  NAND2_X1 U9970 ( .A1(n7727), .A2(n7726), .ZN(n7728) );
  XNOR2_X1 U9971 ( .A(n7730), .B(n7731), .ZN(n9907) );
  NAND2_X1 U9972 ( .A1(n9907), .A2(n8236), .ZN(n7737) );
  NAND2_X1 U9973 ( .A1(n7732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7733) );
  MUX2_X1 U9974 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7733), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7735) );
  AND2_X1 U9975 ( .A1(n7735), .A2(n7734), .ZN(n9352) );
  AOI22_X1 U9976 ( .A1(n8021), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9332), .B2(
        n9352), .ZN(n7736) );
  NAND2_X1 U9977 ( .A1(n7737), .A2(n7736), .ZN(n10336) );
  NAND2_X1 U9978 ( .A1(n10336), .A2(n8093), .ZN(n7744) );
  INV_X1 U9979 ( .A(n8093), .ZN(n8032) );
  NAND2_X1 U9980 ( .A1(n7683), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U9981 ( .A1(n7682), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7741) );
  OAI21_X1 U9982 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7754), .ZN(n10333) );
  INV_X1 U9983 ( .A(n10333), .ZN(n7738) );
  NAND2_X1 U9984 ( .A1(n6486), .A2(n7738), .ZN(n7740) );
  NAND2_X1 U9985 ( .A1(n8027), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7739) );
  NAND4_X1 U9986 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n13210)
         );
  NAND2_X1 U9987 ( .A1(n8032), .A2(n13210), .ZN(n7743) );
  NAND2_X1 U9988 ( .A1(n7744), .A2(n7743), .ZN(n7747) );
  AOI22_X1 U9989 ( .A1(n10336), .A2(n8032), .B1(n13210), .B2(n8093), .ZN(n7745) );
  NAND2_X1 U9990 ( .A1(n10447), .A2(n8236), .ZN(n7752) );
  OR2_X1 U9991 ( .A1(n6492), .A2(n7709), .ZN(n7750) );
  XNOR2_X1 U9992 ( .A(n7750), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9374) );
  AOI22_X1 U9993 ( .A1(n8021), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9332), .B2(
        n9374), .ZN(n7751) );
  NAND2_X1 U9994 ( .A1(n7752), .A2(n7751), .ZN(n14868) );
  NAND2_X1 U9995 ( .A1(n14868), .A2(n8032), .ZN(n7761) );
  NAND2_X1 U9996 ( .A1(n7683), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U9997 ( .A1(n7794), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7758) );
  INV_X1 U9998 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U9999 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  AND2_X1 U10000 ( .A1(n7777), .A2(n7755), .ZN(n10279) );
  NAND2_X1 U10001 ( .A1(n6485), .A2(n10279), .ZN(n7757) );
  NAND2_X1 U10002 ( .A1(n8027), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10003 ( .A1(n13209), .A2(n8214), .ZN(n7760) );
  NAND2_X1 U10004 ( .A1(n7761), .A2(n7760), .ZN(n7764) );
  AOI22_X1 U10005 ( .A1(n14868), .A2(n8214), .B1(n8032), .B2(n13209), .ZN(
        n7762) );
  AOI21_X1 U10006 ( .B1(n7765), .B2(n7764), .A(n7762), .ZN(n7763) );
  INV_X1 U10007 ( .A(n7763), .ZN(n7766) );
  XNOR2_X1 U10008 ( .A(n7768), .B(n7767), .ZN(n10621) );
  NAND2_X1 U10009 ( .A1(n10621), .A2(n8236), .ZN(n7774) );
  NAND2_X1 U10010 ( .A1(n6492), .A2(n7769), .ZN(n7813) );
  NAND2_X1 U10011 ( .A1(n7813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7771) );
  INV_X1 U10012 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10013 ( .A1(n7771), .A2(n7770), .ZN(n7790) );
  OR2_X1 U10014 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  AOI22_X1 U10015 ( .A1(n8021), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9332), .B2(
        n9355), .ZN(n7773) );
  NAND2_X1 U10016 ( .A1(n10567), .A2(n8214), .ZN(n7784) );
  INV_X2 U10017 ( .A(n7775), .ZN(n8206) );
  NAND2_X1 U10018 ( .A1(n8206), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U10019 ( .A1(n7794), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7781) );
  INV_X1 U10020 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10021 ( .A1(n7777), .A2(n7776), .ZN(n7778) );
  AND2_X1 U10022 ( .A1(n7796), .A2(n7778), .ZN(n10533) );
  NAND2_X1 U10023 ( .A1(n6486), .A2(n10533), .ZN(n7780) );
  NAND2_X1 U10024 ( .A1(n8027), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7779) );
  NAND4_X1 U10025 ( .A1(n7782), .A2(n7781), .A3(n7780), .A4(n7779), .ZN(n13208) );
  NAND2_X1 U10026 ( .A1(n8215), .A2(n13208), .ZN(n7783) );
  NAND2_X1 U10027 ( .A1(n7784), .A2(n7783), .ZN(n7787) );
  AOI22_X1 U10028 ( .A1(n10567), .A2(n8032), .B1(n13208), .B2(n8214), .ZN(
        n7785) );
  INV_X1 U10029 ( .A(n7785), .ZN(n7786) );
  NAND2_X1 U10030 ( .A1(n10628), .A2(n8236), .ZN(n7793) );
  NAND2_X1 U10031 ( .A1(n7790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7791) );
  XNOR2_X1 U10032 ( .A(n7791), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9418) );
  AOI22_X1 U10033 ( .A1(n8021), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9332), .B2(
        n9418), .ZN(n7792) );
  NAND2_X1 U10034 ( .A1(n14878), .A2(n8032), .ZN(n7803) );
  NAND2_X1 U10035 ( .A1(n8206), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10036 ( .A1(n7794), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7800) );
  INV_X1 U10037 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10038 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  AND2_X1 U10039 ( .A1(n7822), .A2(n7797), .ZN(n10434) );
  NAND2_X1 U10040 ( .A1(n6486), .A2(n10434), .ZN(n7799) );
  NAND2_X1 U10041 ( .A1(n8027), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7798) );
  NAND4_X1 U10042 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n13207) );
  NAND2_X1 U10043 ( .A1(n13207), .A2(n8214), .ZN(n7802) );
  NAND2_X1 U10044 ( .A1(n7803), .A2(n7802), .ZN(n7808) );
  NAND2_X1 U10045 ( .A1(n7807), .A2(n7808), .ZN(n7806) );
  NAND2_X1 U10046 ( .A1(n14878), .A2(n8214), .ZN(n7804) );
  OAI21_X1 U10047 ( .B1(n10597), .B2(n8214), .A(n7804), .ZN(n7805) );
  INV_X1 U10048 ( .A(n7807), .ZN(n7810) );
  INV_X1 U10049 ( .A(n7808), .ZN(n7809) );
  NAND2_X1 U10050 ( .A1(n7815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7814) );
  MUX2_X1 U10051 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7814), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7818) );
  INV_X1 U10052 ( .A(n7815), .ZN(n7817) );
  INV_X1 U10053 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10054 ( .A1(n7817), .A2(n7816), .ZN(n7854) );
  NAND2_X1 U10055 ( .A1(n7818), .A2(n7854), .ZN(n9419) );
  INV_X1 U10056 ( .A(n9419), .ZN(n9444) );
  AOI22_X1 U10057 ( .A1(n8021), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9332), .B2(
        n9444), .ZN(n7819) );
  NAND2_X1 U10058 ( .A1(n6727), .A2(n8214), .ZN(n7829) );
  NAND2_X1 U10059 ( .A1(n8206), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10060 ( .A1(n8256), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U10061 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  AND2_X1 U10062 ( .A1(n7837), .A2(n7823), .ZN(n10677) );
  NAND2_X1 U10063 ( .A1(n6485), .A2(n10677), .ZN(n7825) );
  NAND2_X1 U10064 ( .A1(n8027), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7824) );
  NAND4_X1 U10065 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7824), .ZN(n13206) );
  NAND2_X1 U10066 ( .A1(n8215), .A2(n13206), .ZN(n7828) );
  AOI22_X1 U10067 ( .A1(n6727), .A2(n8215), .B1(n13206), .B2(n8214), .ZN(n7830) );
  XNOR2_X1 U10068 ( .A(n7832), .B(n7831), .ZN(n10713) );
  NAND2_X1 U10069 ( .A1(n10713), .A2(n8236), .ZN(n7835) );
  NAND2_X1 U10070 ( .A1(n7854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10071 ( .A(n7833), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9765) );
  AOI22_X1 U10072 ( .A1(n8021), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9332), .B2(
        n9765), .ZN(n7834) );
  NAND2_X1 U10073 ( .A1(n10927), .A2(n8215), .ZN(n7844) );
  NAND2_X1 U10074 ( .A1(n8256), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10075 ( .A1(n8206), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7841) );
  INV_X1 U10076 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10077 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  AND2_X1 U10078 ( .A1(n7877), .A2(n7838), .ZN(n10852) );
  NAND2_X1 U10079 ( .A1(n6485), .A2(n10852), .ZN(n7840) );
  NAND2_X1 U10080 ( .A1(n8027), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7839) );
  NAND4_X1 U10081 ( .A1(n7842), .A2(n7841), .A3(n7840), .A4(n7839), .ZN(n13205) );
  NAND2_X1 U10082 ( .A1(n13205), .A2(n8214), .ZN(n7843) );
  NAND2_X1 U10083 ( .A1(n7844), .A2(n7843), .ZN(n7849) );
  NAND2_X1 U10084 ( .A1(n7848), .A2(n7849), .ZN(n7847) );
  INV_X1 U10085 ( .A(n13205), .ZN(n10813) );
  NAND2_X1 U10086 ( .A1(n10927), .A2(n8214), .ZN(n7845) );
  OAI21_X1 U10087 ( .B1(n10813), .B2(n8214), .A(n7845), .ZN(n7846) );
  INV_X1 U10088 ( .A(n7848), .ZN(n7851) );
  INV_X1 U10089 ( .A(n7849), .ZN(n7850) );
  XNOR2_X1 U10090 ( .A(n7853), .B(n7852), .ZN(n10877) );
  NAND2_X1 U10091 ( .A1(n10877), .A2(n8236), .ZN(n7859) );
  INV_X1 U10092 ( .A(n7854), .ZN(n7856) );
  INV_X1 U10093 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10094 ( .A1(n7856), .A2(n7855), .ZN(n7871) );
  NAND2_X1 U10095 ( .A1(n7871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7857) );
  XNOR2_X1 U10096 ( .A(n7857), .B(P2_IR_REG_10__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U10097 ( .A1(n8021), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n13226), 
        .B2(n9332), .ZN(n7858) );
  NAND2_X1 U10098 ( .A1(n11062), .A2(n8214), .ZN(n7865) );
  NAND2_X1 U10099 ( .A1(n8206), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10100 ( .A1(n8256), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U10101 ( .A(n7877), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U10102 ( .A1(n6486), .A2(n10918), .ZN(n7861) );
  NAND2_X1 U10103 ( .A1(n8027), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7860) );
  NAND4_X1 U10104 ( .A1(n7863), .A2(n7862), .A3(n7861), .A4(n7860), .ZN(n13204) );
  NAND2_X1 U10105 ( .A1(n8215), .A2(n13204), .ZN(n7864) );
  AOI22_X1 U10106 ( .A1(n11062), .A2(n8215), .B1(n13204), .B2(n8214), .ZN(
        n7866) );
  NAND2_X1 U10107 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  NAND2_X1 U10108 ( .A1(n7870), .A2(n7869), .ZN(n11033) );
  NAND2_X1 U10109 ( .A1(n11033), .A2(n8236), .ZN(n7874) );
  OAI21_X1 U10110 ( .B1(n7871), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7872) );
  XNOR2_X1 U10111 ( .A(n7872), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U10112 ( .A1(n13234), .A2(n9332), .B1(n8021), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U10113 ( .A1(n11291), .A2(n8215), .ZN(n7884) );
  NAND2_X1 U10114 ( .A1(n8206), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10115 ( .A1(n8256), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7881) );
  INV_X1 U10116 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7876) );
  INV_X1 U10117 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7875) );
  OAI21_X1 U10118 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7878) );
  AND2_X1 U10119 ( .A1(n7878), .A2(n7895), .ZN(n11073) );
  NAND2_X1 U10120 ( .A1(n6485), .A2(n11073), .ZN(n7880) );
  NAND2_X1 U10121 ( .A1(n8027), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7879) );
  NAND4_X1 U10122 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n13203) );
  NAND2_X1 U10123 ( .A1(n13203), .A2(n8214), .ZN(n7883) );
  NAND2_X1 U10124 ( .A1(n7884), .A2(n7883), .ZN(n7887) );
  INV_X1 U10125 ( .A(n13203), .ZN(n11095) );
  NAND2_X1 U10126 ( .A1(n11291), .A2(n8214), .ZN(n7885) );
  OAI21_X1 U10127 ( .B1(n11095), .B2(n8214), .A(n7885), .ZN(n7886) );
  NAND2_X1 U10128 ( .A1(n11114), .A2(n8236), .ZN(n7894) );
  NAND2_X1 U10129 ( .A1(n6492), .A2(n7889), .ZN(n7891) );
  NAND2_X1 U10130 ( .A1(n7891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7890) );
  MUX2_X1 U10131 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7890), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7892) );
  OR2_X1 U10132 ( .A1(n7891), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7910) );
  AND2_X1 U10133 ( .A1(n7892), .A2(n7910), .ZN(n13270) );
  AOI22_X1 U10134 ( .A1(n8021), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9332), 
        .B2(n13270), .ZN(n7893) );
  NAND2_X1 U10135 ( .A1(n11255), .A2(n8214), .ZN(n7902) );
  NAND2_X1 U10136 ( .A1(n8206), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10137 ( .A1(n8256), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7899) );
  INV_X1 U10138 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n13240) );
  NAND2_X1 U10139 ( .A1(n7895), .A2(n13240), .ZN(n7896) );
  AND2_X1 U10140 ( .A1(n7930), .A2(n7896), .ZN(n11244) );
  NAND2_X1 U10141 ( .A1(n6486), .A2(n11244), .ZN(n7898) );
  NAND2_X1 U10142 ( .A1(n8027), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7897) );
  NAND4_X1 U10143 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n13202) );
  NAND2_X1 U10144 ( .A1(n8215), .A2(n13202), .ZN(n7901) );
  NAND2_X1 U10145 ( .A1(n7902), .A2(n7901), .ZN(n7904) );
  AOI22_X1 U10146 ( .A1(n11255), .A2(n8215), .B1(n13202), .B2(n8214), .ZN(
        n7903) );
  AOI21_X1 U10147 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7906) );
  XNOR2_X1 U10148 ( .A(n7907), .B(n7527), .ZN(n11145) );
  NAND2_X1 U10149 ( .A1(n11145), .A2(n8236), .ZN(n7913) );
  NAND2_X1 U10150 ( .A1(n7910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7909) );
  MUX2_X1 U10151 ( .A(n7909), .B(P2_IR_REG_31__SCAN_IN), .S(n7908), .Z(n7911)
         );
  OR2_X1 U10152 ( .A1(n7910), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7943) );
  AND2_X1 U10153 ( .A1(n7911), .A2(n7943), .ZN(n14778) );
  AOI22_X1 U10154 ( .A1(n8021), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9332), 
        .B2(n14778), .ZN(n7912) );
  NAND2_X1 U10155 ( .A1(n13603), .A2(n8215), .ZN(n7919) );
  NAND2_X1 U10156 ( .A1(n8206), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10157 ( .A1(n8256), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7916) );
  XNOR2_X1 U10158 ( .A(n7930), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U10159 ( .A1(n6485), .A2(n11268), .ZN(n7915) );
  NAND2_X1 U10160 ( .A1(n8027), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7914) );
  NAND4_X1 U10161 ( .A1(n7917), .A2(n7916), .A3(n7915), .A4(n7914), .ZN(n13201) );
  NAND2_X1 U10162 ( .A1(n13201), .A2(n8214), .ZN(n7918) );
  NAND2_X1 U10163 ( .A1(n7919), .A2(n7918), .ZN(n7922) );
  INV_X1 U10164 ( .A(n13201), .ZN(n11309) );
  NAND2_X1 U10165 ( .A1(n13603), .A2(n8214), .ZN(n7920) );
  OAI21_X1 U10166 ( .B1(n11309), .B2(n8093), .A(n7920), .ZN(n7921) );
  INV_X1 U10167 ( .A(n7922), .ZN(n7923) );
  XNOR2_X1 U10168 ( .A(n7925), .B(n7924), .ZN(n11346) );
  NAND2_X1 U10169 ( .A1(n11346), .A2(n8236), .ZN(n7928) );
  NAND2_X1 U10170 ( .A1(n7943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  XNOR2_X1 U10171 ( .A(n7926), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14790) );
  AOI22_X1 U10172 ( .A1(n8021), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9332), 
        .B2(n14790), .ZN(n7927) );
  NAND2_X1 U10173 ( .A1(n13598), .A2(n8214), .ZN(n7937) );
  NAND2_X1 U10174 ( .A1(n8256), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10175 ( .A1(n8027), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7934) );
  OAI21_X1 U10176 ( .B1(n7930), .B2(n7929), .A(n11404), .ZN(n7931) );
  AND2_X1 U10177 ( .A1(n7931), .A2(n7947), .ZN(n11407) );
  NAND2_X1 U10178 ( .A1(n6485), .A2(n11407), .ZN(n7933) );
  NAND2_X1 U10179 ( .A1(n8206), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7932) );
  NAND4_X1 U10180 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n13200) );
  NAND2_X1 U10181 ( .A1(n8215), .A2(n13200), .ZN(n7936) );
  AOI22_X1 U10182 ( .A1(n13598), .A2(n7820), .B1(n13200), .B2(n8214), .ZN(
        n7938) );
  OR2_X1 U10183 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  NAND2_X1 U10184 ( .A1(n7942), .A2(n7941), .ZN(n11425) );
  NAND2_X1 U10185 ( .A1(n11425), .A2(n8236), .ZN(n7946) );
  OAI21_X1 U10186 ( .B1(n7943), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7944) );
  XNOR2_X1 U10187 ( .A(n7944), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U10188 ( .A1(n8021), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n14800), 
        .B2(n9332), .ZN(n7945) );
  NAND2_X1 U10189 ( .A1(n13593), .A2(n7820), .ZN(n7954) );
  NAND2_X1 U10190 ( .A1(n8256), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10191 ( .A1(n8027), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7951) );
  INV_X1 U10192 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U10193 ( .A1(n7947), .A2(n11537), .ZN(n7948) );
  AND2_X1 U10194 ( .A1(n7971), .A2(n7948), .ZN(n11418) );
  NAND2_X1 U10195 ( .A1(n6485), .A2(n11418), .ZN(n7950) );
  NAND2_X1 U10196 ( .A1(n8206), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7949) );
  NAND4_X1 U10197 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n13199) );
  NAND2_X1 U10198 ( .A1(n13199), .A2(n8214), .ZN(n7953) );
  NAND2_X1 U10199 ( .A1(n7954), .A2(n7953), .ZN(n7957) );
  AOI22_X1 U10200 ( .A1(n13593), .A2(n8214), .B1(n7820), .B2(n13199), .ZN(
        n7955) );
  AOI21_X1 U10201 ( .B1(n7958), .B2(n7957), .A(n7955), .ZN(n7956) );
  INV_X1 U10202 ( .A(n7956), .ZN(n7959) );
  NAND2_X1 U10203 ( .A1(n11509), .A2(n8236), .ZN(n7967) );
  NAND2_X1 U10204 ( .A1(n6492), .A2(n6618), .ZN(n7964) );
  NAND2_X1 U10205 ( .A1(n7964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7963) );
  MUX2_X1 U10206 ( .A(n7963), .B(P2_IR_REG_31__SCAN_IN), .S(n7962), .Z(n7965)
         );
  OR2_X1 U10207 ( .A1(n7964), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7983) );
  AND2_X1 U10208 ( .A1(n7965), .A2(n7983), .ZN(n13276) );
  AOI22_X1 U10209 ( .A1(n8021), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9332), 
        .B2(n13276), .ZN(n7966) );
  NAND2_X1 U10210 ( .A1(n13587), .A2(n8214), .ZN(n7976) );
  INV_X1 U10211 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U10212 ( .A1(n8027), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7968) );
  OAI21_X1 U10213 ( .B1(n13277), .B2(n7969), .A(n7968), .ZN(n7974) );
  INV_X1 U10214 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10215 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  NAND2_X1 U10216 ( .A1(n7990), .A2(n7972), .ZN(n13110) );
  INV_X1 U10217 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13263) );
  OAI22_X1 U10218 ( .A1(n13110), .A2(n8239), .B1(n7775), .B2(n13263), .ZN(
        n7973) );
  OR2_X1 U10219 ( .A1(n7974), .A2(n7973), .ZN(n13198) );
  NAND2_X1 U10220 ( .A1(n7820), .A2(n13198), .ZN(n7975) );
  NAND2_X1 U10221 ( .A1(n13587), .A2(n7820), .ZN(n7977) );
  OAI21_X1 U10222 ( .B1(n13117), .B2(n7820), .A(n7977), .ZN(n7978) );
  XNOR2_X1 U10223 ( .A(n7979), .B(SI_17_), .ZN(n7980) );
  XNOR2_X1 U10224 ( .A(n7981), .B(n7980), .ZN(n11634) );
  NAND2_X1 U10225 ( .A1(n11634), .A2(n8236), .ZN(n7989) );
  NAND2_X1 U10226 ( .A1(n7983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7982) );
  MUX2_X1 U10227 ( .A(n7982), .B(P2_IR_REG_31__SCAN_IN), .S(n7984), .Z(n7986)
         );
  INV_X1 U10228 ( .A(n7983), .ZN(n7985) );
  NAND2_X1 U10229 ( .A1(n7985), .A2(n7984), .ZN(n8001) );
  NAND2_X1 U10230 ( .A1(n7986), .A2(n8001), .ZN(n14823) );
  INV_X1 U10231 ( .A(n14823), .ZN(n7987) );
  AOI22_X1 U10232 ( .A1(n8021), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9332), 
        .B2(n7987), .ZN(n7988) );
  NAND2_X1 U10233 ( .A1(n13581), .A2(n8032), .ZN(n7995) );
  NAND2_X1 U10234 ( .A1(n7990), .A2(n13118), .ZN(n7991) );
  NAND2_X1 U10235 ( .A1(n8006), .A2(n7991), .ZN(n13494) );
  AOI22_X1 U10236 ( .A1(n8256), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8206), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10237 ( .A1(n8027), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7992) );
  OAI211_X1 U10238 ( .C1(n13494), .C2(n8239), .A(n7993), .B(n7992), .ZN(n13197) );
  NAND2_X1 U10239 ( .A1(n13197), .A2(n8214), .ZN(n7994) );
  NAND2_X1 U10240 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  AOI22_X1 U10241 ( .A1(n13581), .A2(n8214), .B1(n8215), .B2(n13197), .ZN(
        n7996) );
  NAND2_X1 U10242 ( .A1(n7998), .A2(n9641), .ZN(n7999) );
  NAND2_X1 U10243 ( .A1(n11638), .A2(n8236), .ZN(n8004) );
  NAND2_X1 U10244 ( .A1(n8001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8002) );
  XNOR2_X1 U10245 ( .A(n8002), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15225) );
  AOI22_X1 U10246 ( .A1(n8021), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9332), 
        .B2(n15225), .ZN(n8003) );
  INV_X1 U10247 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8010) );
  INV_X1 U10248 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10249 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  NAND2_X1 U10250 ( .A1(n8025), .A2(n8007), .ZN(n13474) );
  OR2_X1 U10251 ( .A1(n13474), .A2(n8239), .ZN(n8009) );
  AOI22_X1 U10252 ( .A1(n8256), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8206), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n8008) );
  OAI211_X1 U10253 ( .C1(n8261), .C2(n8010), .A(n8009), .B(n8008), .ZN(n13196)
         );
  AND2_X1 U10254 ( .A1(n13196), .A2(n8215), .ZN(n8011) );
  AOI21_X1 U10255 ( .B1(n13576), .B2(n8214), .A(n8011), .ZN(n8012) );
  NAND2_X1 U10256 ( .A1(n13576), .A2(n8032), .ZN(n8014) );
  NAND2_X1 U10257 ( .A1(n13196), .A2(n8214), .ZN(n8013) );
  NAND2_X1 U10258 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  OAI21_X1 U10259 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8020) );
  XNOR2_X1 U10260 ( .A(n8020), .B(n8019), .ZN(n11644) );
  NAND2_X1 U10261 ( .A1(n11644), .A2(n8236), .ZN(n8023) );
  AOI22_X1 U10262 ( .A1(n8021), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9332), 
        .B2(n11500), .ZN(n8022) );
  NAND2_X1 U10263 ( .A1(n13571), .A2(n8215), .ZN(n8031) );
  NAND2_X1 U10264 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U10265 ( .A1(n8044), .A2(n8026), .ZN(n13458) );
  AOI22_X1 U10266 ( .A1(n8256), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8206), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10267 ( .A1(n8027), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8028) );
  OAI211_X1 U10268 ( .C1(n13458), .C2(n8239), .A(n8029), .B(n8028), .ZN(n13436) );
  NAND2_X1 U10269 ( .A1(n13436), .A2(n8214), .ZN(n8030) );
  NAND2_X1 U10270 ( .A1(n8031), .A2(n8030), .ZN(n8035) );
  AOI22_X1 U10271 ( .A1(n13571), .A2(n8214), .B1(n8032), .B2(n13436), .ZN(
        n8033) );
  AOI21_X1 U10272 ( .B1(n8036), .B2(n8035), .A(n8033), .ZN(n8034) );
  NOR2_X1 U10273 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  NAND2_X1 U10274 ( .A1(n8039), .A2(n8038), .ZN(n8040) );
  OR2_X1 U10275 ( .A1(n6653), .A2(n10923), .ZN(n8042) );
  NAND2_X1 U10276 ( .A1(n13565), .A2(n8214), .ZN(n8054) );
  INV_X1 U10277 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13136) );
  NAND2_X1 U10278 ( .A1(n8044), .A2(n13136), .ZN(n8045) );
  NAND2_X1 U10279 ( .A1(n8046), .A2(n8045), .ZN(n13428) );
  OR2_X1 U10280 ( .A1(n13428), .A2(n8239), .ZN(n8052) );
  INV_X1 U10281 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10282 ( .A1(n8256), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10283 ( .A1(n8206), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8047) );
  OAI211_X1 U10284 ( .C1(n8049), .C2(n8261), .A(n8048), .B(n8047), .ZN(n8050)
         );
  INV_X1 U10285 ( .A(n8050), .ZN(n8051) );
  NAND2_X1 U10286 ( .A1(n8052), .A2(n8051), .ZN(n13195) );
  NAND2_X1 U10287 ( .A1(n13195), .A2(n8215), .ZN(n8053) );
  AOI22_X1 U10288 ( .A1(n13565), .A2(n8215), .B1(n13195), .B2(n8214), .ZN(
        n8055) );
  AOI22_X1 U10289 ( .A1(n13561), .A2(n8214), .B1(n8032), .B2(n13438), .ZN(
        n8056) );
  AOI21_X1 U10290 ( .B1(n8058), .B2(n8057), .A(n8056), .ZN(n8059) );
  INV_X1 U10291 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8500) );
  INV_X1 U10292 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10953) );
  MUX2_X1 U10293 ( .A(n8500), .B(n10953), .S(n9517), .Z(n8063) );
  NAND2_X1 U10294 ( .A1(n11683), .A2(n8063), .ZN(n8064) );
  NAND2_X1 U10295 ( .A1(n8077), .A2(n8064), .ZN(n10952) );
  OR2_X1 U10296 ( .A1(n6653), .A2(n10953), .ZN(n8065) );
  INV_X1 U10297 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U10298 ( .A1(n8067), .A2(n13148), .ZN(n8068) );
  AND2_X1 U10299 ( .A1(n8086), .A2(n8068), .ZN(n13400) );
  NAND2_X1 U10300 ( .A1(n13400), .A2(n6486), .ZN(n8074) );
  INV_X1 U10301 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10302 ( .A1(n8256), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10303 ( .A1(n8206), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8069) );
  OAI211_X1 U10304 ( .C1(n8071), .C2(n8261), .A(n8070), .B(n8069), .ZN(n8072)
         );
  INV_X1 U10305 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U10306 ( .A1(n8074), .A2(n8073), .ZN(n13375) );
  AOI22_X1 U10307 ( .A1(n13557), .A2(n8214), .B1(n8215), .B2(n13375), .ZN(
        n8076) );
  INV_X1 U10308 ( .A(n13557), .ZN(n13403) );
  INV_X1 U10309 ( .A(n13375), .ZN(n13091) );
  OAI22_X1 U10310 ( .A1(n13403), .A2(n8214), .B1(n13091), .B2(n7820), .ZN(
        n8075) );
  INV_X1 U10311 ( .A(n8096), .ZN(n8099) );
  MUX2_X1 U10312 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9517), .Z(n8078) );
  NAND2_X1 U10313 ( .A1(n8078), .A2(SI_23_), .ZN(n8100) );
  OAI21_X1 U10314 ( .B1(SI_23_), .B2(n8078), .A(n8100), .ZN(n8079) );
  INV_X1 U10315 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U10316 ( .A1(n8101), .A2(n8082), .ZN(n11693) );
  OR2_X1 U10317 ( .A1(n11693), .A2(n8255), .ZN(n8084) );
  INV_X1 U10318 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8502) );
  OR2_X1 U10319 ( .A1(n6653), .A2(n8502), .ZN(n8083) );
  INV_X1 U10320 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U10321 ( .A1(n8086), .A2(n13067), .ZN(n8087) );
  NAND2_X1 U10322 ( .A1(n8110), .A2(n8087), .ZN(n13378) );
  OR2_X1 U10323 ( .A1(n13378), .A2(n8239), .ZN(n8092) );
  INV_X1 U10324 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15160) );
  NAND2_X1 U10325 ( .A1(n8256), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10326 ( .A1(n8206), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8088) );
  OAI211_X1 U10327 ( .C1(n15160), .C2(n8261), .A(n8089), .B(n8088), .ZN(n8090)
         );
  INV_X1 U10328 ( .A(n8090), .ZN(n8091) );
  OAI22_X1 U10329 ( .A1(n13549), .A2(n8093), .B1(n13126), .B2(n7820), .ZN(
        n8095) );
  INV_X1 U10330 ( .A(n8095), .ZN(n8098) );
  AOI22_X1 U10331 ( .A1(n13388), .A2(n8214), .B1(n8215), .B2(n13194), .ZN(
        n8094) );
  INV_X1 U10332 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11704) );
  INV_X1 U10333 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11323) );
  MUX2_X1 U10334 ( .A(n11704), .B(n11323), .S(n9517), .Z(n8103) );
  NAND2_X1 U10335 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  NAND2_X1 U10336 ( .A1(n8121), .A2(n8105), .ZN(n11703) );
  OR2_X1 U10337 ( .A1(n6653), .A2(n11323), .ZN(n8106) );
  INV_X1 U10338 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10339 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  NAND2_X1 U10340 ( .A1(n8126), .A2(n8111), .ZN(n13366) );
  OR2_X1 U10341 ( .A1(n13366), .A2(n8239), .ZN(n8117) );
  INV_X1 U10342 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10343 ( .A1(n8256), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10344 ( .A1(n8257), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8112) );
  OAI211_X1 U10345 ( .C1(n8114), .C2(n8261), .A(n8113), .B(n8112), .ZN(n8115)
         );
  INV_X1 U10346 ( .A(n8115), .ZN(n8116) );
  NAND2_X1 U10347 ( .A1(n8117), .A2(n8116), .ZN(n13377) );
  AOI22_X1 U10348 ( .A1(n13369), .A2(n8214), .B1(n8215), .B2(n13377), .ZN(
        n8119) );
  INV_X1 U10349 ( .A(n13369), .ZN(n13543) );
  INV_X1 U10350 ( .A(n13377), .ZN(n13099) );
  OAI22_X1 U10351 ( .A1(n13543), .A2(n8093), .B1(n13099), .B2(n7820), .ZN(
        n8118) );
  MUX2_X1 U10352 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9517), .Z(n8132) );
  XNOR2_X1 U10353 ( .A(n8132), .B(SI_25_), .ZN(n8135) );
  XNOR2_X1 U10354 ( .A(n8136), .B(n8135), .ZN(n11714) );
  NAND2_X1 U10355 ( .A1(n11714), .A2(n8236), .ZN(n8123) );
  INV_X1 U10356 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15202) );
  OR2_X1 U10357 ( .A1(n6653), .A2(n15202), .ZN(n8122) );
  INV_X1 U10358 ( .A(n8126), .ZN(n8124) );
  INV_X1 U10359 ( .A(n8140), .ZN(n8160) );
  INV_X1 U10360 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U10361 ( .A1(n8126), .A2(n8125), .ZN(n8127) );
  INV_X1 U10362 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10363 ( .A1(n8256), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10364 ( .A1(n8206), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8128) );
  OAI211_X1 U10365 ( .C1(n8130), .C2(n8261), .A(n8129), .B(n8128), .ZN(n8131)
         );
  AOI21_X1 U10366 ( .B1(n13350), .B2(n6486), .A(n8131), .ZN(n13180) );
  INV_X1 U10367 ( .A(n13180), .ZN(n13193) );
  AOI22_X1 U10368 ( .A1(n13537), .A2(n8214), .B1(n8215), .B2(n13193), .ZN(
        n8220) );
  OAI22_X1 U10369 ( .A1(n13352), .A2(n8214), .B1(n13180), .B2(n7820), .ZN(
        n8219) );
  INV_X1 U10370 ( .A(n8132), .ZN(n8133) );
  INV_X1 U10371 ( .A(SI_25_), .ZN(n11390) );
  NAND2_X1 U10372 ( .A1(n8133), .A2(n11390), .ZN(n8134) );
  INV_X1 U10373 ( .A(SI_26_), .ZN(n13055) );
  MUX2_X1 U10374 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9517), .Z(n8153) );
  MUX2_X1 U10375 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9517), .Z(n8174) );
  XNOR2_X1 U10376 ( .A(n8174), .B(SI_27_), .ZN(n8137) );
  INV_X1 U10377 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11563) );
  OR2_X1 U10378 ( .A1(n6653), .A2(n11563), .ZN(n8138) );
  NAND2_X1 U10379 ( .A1(n8140), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8162) );
  INV_X1 U10380 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10381 ( .A1(n8162), .A2(n8141), .ZN(n8142) );
  NAND2_X1 U10382 ( .A1(n13324), .A2(n6485), .ZN(n8149) );
  INV_X1 U10383 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10384 ( .A1(n8256), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10385 ( .A1(n8206), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8144) );
  OAI211_X1 U10386 ( .C1(n8146), .C2(n8261), .A(n8145), .B(n8144), .ZN(n8147)
         );
  INV_X1 U10387 ( .A(n8147), .ZN(n8148) );
  NAND2_X1 U10388 ( .A1(n8149), .A2(n8148), .ZN(n13191) );
  AND2_X1 U10389 ( .A1(n13191), .A2(n8215), .ZN(n8150) );
  AOI21_X1 U10390 ( .B1(n13526), .B2(n8214), .A(n8150), .ZN(n8232) );
  NAND2_X1 U10391 ( .A1(n13526), .A2(n8215), .ZN(n8152) );
  NAND2_X1 U10392 ( .A1(n13191), .A2(n8214), .ZN(n8151) );
  NAND2_X1 U10393 ( .A1(n8152), .A2(n8151), .ZN(n8231) );
  NAND2_X1 U10394 ( .A1(n8232), .A2(n8231), .ZN(n8228) );
  INV_X1 U10395 ( .A(n8153), .ZN(n8154) );
  XNOR2_X1 U10396 ( .A(n8154), .B(SI_26_), .ZN(n8155) );
  OR2_X1 U10397 ( .A1(n6653), .A2(n7043), .ZN(n8157) );
  INV_X1 U10398 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10399 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U10400 ( .A1(n8162), .A2(n8161), .ZN(n13336) );
  INV_X1 U10401 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10402 ( .A1(n8256), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10403 ( .A1(n8257), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U10404 ( .C1(n8165), .C2(n8261), .A(n8164), .B(n8163), .ZN(n8166)
         );
  INV_X1 U10405 ( .A(n8166), .ZN(n8167) );
  AND2_X1 U10406 ( .A1(n13192), .A2(n8215), .ZN(n8169) );
  AOI21_X1 U10407 ( .B1(n13532), .B2(n8214), .A(n8169), .ZN(n8225) );
  NAND2_X1 U10408 ( .A1(n13532), .A2(n8215), .ZN(n8171) );
  NAND2_X1 U10409 ( .A1(n13192), .A2(n8214), .ZN(n8170) );
  NAND2_X1 U10410 ( .A1(n8171), .A2(n8170), .ZN(n8224) );
  NAND2_X1 U10411 ( .A1(n8225), .A2(n8224), .ZN(n8172) );
  NAND2_X1 U10412 ( .A1(n8228), .A2(n8172), .ZN(n8218) );
  AOI21_X1 U10413 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8173) );
  INV_X1 U10414 ( .A(SI_27_), .ZN(n15031) );
  MUX2_X1 U10415 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9517), .Z(n8176) );
  XNOR2_X1 U10416 ( .A(n8176), .B(n15044), .ZN(n8199) );
  NAND2_X1 U10417 ( .A1(n8200), .A2(n8199), .ZN(n8179) );
  INV_X1 U10418 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U10419 ( .A1(n8177), .A2(n15044), .ZN(n8178) );
  NAND2_X1 U10420 ( .A1(n8179), .A2(n8178), .ZN(n8234) );
  INV_X1 U10421 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11622) );
  INV_X1 U10422 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8237) );
  MUX2_X1 U10423 ( .A(n11622), .B(n8237), .S(n9517), .Z(n8183) );
  XNOR2_X1 U10424 ( .A(n8183), .B(SI_29_), .ZN(n8233) );
  INV_X1 U10425 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12472) );
  MUX2_X1 U10426 ( .A(n12472), .B(n7022), .S(n9517), .Z(n8181) );
  INV_X1 U10427 ( .A(SI_30_), .ZN(n12114) );
  NOR2_X1 U10428 ( .A1(n8181), .A2(n12114), .ZN(n8184) );
  MUX2_X1 U10429 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9517), .Z(n8180) );
  XNOR2_X1 U10430 ( .A(n8180), .B(SI_31_), .ZN(n8182) );
  INV_X1 U10431 ( .A(n8182), .ZN(n8189) );
  INV_X1 U10432 ( .A(n8181), .ZN(n8251) );
  OAI21_X1 U10433 ( .B1(n8189), .B2(n12114), .A(n8251), .ZN(n8187) );
  OAI21_X1 U10434 ( .B1(n8182), .B2(SI_30_), .A(n8181), .ZN(n8186) );
  INV_X1 U10435 ( .A(SI_29_), .ZN(n12110) );
  NAND2_X1 U10436 ( .A1(n8183), .A2(n12110), .ZN(n8249) );
  NOR2_X1 U10437 ( .A1(n8184), .A2(n8249), .ZN(n8185) );
  AOI22_X1 U10438 ( .A1(n8187), .A2(n8186), .B1(n8185), .B2(n8189), .ZN(n8192)
         );
  OAI21_X1 U10439 ( .B1(n8251), .B2(SI_30_), .A(n8249), .ZN(n8188) );
  NOR2_X1 U10440 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  NAND2_X1 U10441 ( .A1(n8250), .A2(n8190), .ZN(n8191) );
  NAND2_X1 U10442 ( .A1(n13625), .A2(n8236), .ZN(n8195) );
  INV_X1 U10443 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12474) );
  OR2_X1 U10444 ( .A1(n6653), .A2(n12474), .ZN(n8194) );
  INV_X1 U10445 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10446 ( .A1(n8256), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10447 ( .A1(n8206), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10448 ( .C1(n8261), .C2(n8198), .A(n8197), .B(n8196), .ZN(n13292)
         );
  INV_X1 U10449 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8898) );
  OR2_X1 U10450 ( .A1(n6653), .A2(n8898), .ZN(n8201) );
  INV_X1 U10451 ( .A(n8204), .ZN(n8203) );
  NAND2_X1 U10452 ( .A1(n8203), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11806) );
  INV_X1 U10453 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11617) );
  NAND2_X1 U10454 ( .A1(n8204), .A2(n11617), .ZN(n8205) );
  NAND2_X1 U10455 ( .A1(n11806), .A2(n8205), .ZN(n13312) );
  OR2_X1 U10456 ( .A1(n13312), .A2(n8239), .ZN(n8212) );
  INV_X1 U10457 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U10458 ( .A1(n8256), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10459 ( .A1(n8206), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8207) );
  OAI211_X1 U10460 ( .C1(n8209), .C2(n8261), .A(n8208), .B(n8207), .ZN(n8210)
         );
  INV_X1 U10461 ( .A(n8210), .ZN(n8211) );
  AND2_X1 U10462 ( .A1(n13190), .A2(n8214), .ZN(n8213) );
  AOI21_X1 U10463 ( .B1(n13520), .B2(n7820), .A(n8213), .ZN(n8270) );
  NAND2_X1 U10464 ( .A1(n13520), .A2(n8214), .ZN(n8217) );
  NAND2_X1 U10465 ( .A1(n13190), .A2(n8215), .ZN(n8216) );
  NAND2_X1 U10466 ( .A1(n8217), .A2(n8216), .ZN(n8269) );
  INV_X1 U10467 ( .A(n8218), .ZN(n8223) );
  INV_X1 U10468 ( .A(n8219), .ZN(n8222) );
  INV_X1 U10469 ( .A(n8220), .ZN(n8221) );
  NAND3_X1 U10470 ( .A1(n8223), .A2(n8222), .A3(n8221), .ZN(n8230) );
  INV_X1 U10471 ( .A(n8224), .ZN(n8227) );
  INV_X1 U10472 ( .A(n8225), .ZN(n8226) );
  NAND3_X1 U10473 ( .A1(n8228), .A2(n8227), .A3(n8226), .ZN(n8229) );
  OAI211_X1 U10474 ( .C1(n8232), .C2(n8231), .A(n8230), .B(n8229), .ZN(n8246)
         );
  OR2_X1 U10475 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  OR2_X1 U10476 ( .A1(n6653), .A2(n8237), .ZN(n8238) );
  OR2_X1 U10477 ( .A1(n11806), .A2(n8239), .ZN(n8245) );
  INV_X1 U10478 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10479 ( .A1(n8256), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10480 ( .A1(n8206), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8240) );
  OAI211_X1 U10481 ( .C1(n8242), .C2(n8261), .A(n8241), .B(n8240), .ZN(n8243)
         );
  INV_X1 U10482 ( .A(n8243), .ZN(n8244) );
  OAI22_X1 U10483 ( .A1(n11809), .A2(n8214), .B1(n13305), .B2(n8215), .ZN(
        n8266) );
  INV_X1 U10484 ( .A(n13305), .ZN(n10345) );
  AOI22_X1 U10485 ( .A1(n13515), .A2(n8214), .B1(n8215), .B2(n10345), .ZN(
        n8267) );
  INV_X1 U10486 ( .A(n13292), .ZN(n8262) );
  MUX2_X1 U10487 ( .A(n8262), .B(n8214), .S(n8247), .Z(n8248) );
  NAND2_X1 U10488 ( .A1(n8250), .A2(n8249), .ZN(n8253) );
  XNOR2_X1 U10489 ( .A(n8251), .B(SI_30_), .ZN(n8252) );
  INV_X1 U10490 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10491 ( .A1(n8256), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10492 ( .A1(n8257), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8258) );
  OAI211_X1 U10493 ( .C1(n8261), .C2(n8260), .A(n8259), .B(n8258), .ZN(n13189)
         );
  AOI22_X1 U10494 ( .A1(n8307), .A2(n8214), .B1(n7820), .B2(n13189), .ZN(n8275) );
  NOR2_X1 U10495 ( .A1(n8262), .A2(n8215), .ZN(n8280) );
  NAND2_X1 U10496 ( .A1(n6682), .A2(n11500), .ZN(n9499) );
  INV_X1 U10497 ( .A(n10922), .ZN(n10072) );
  NAND2_X1 U10498 ( .A1(n10922), .A2(n6754), .ZN(n10075) );
  OAI211_X1 U10499 ( .C1(n9499), .C2(n10072), .A(n9497), .B(n10075), .ZN(n8264) );
  OAI21_X1 U10500 ( .B1(n8280), .B2(n8264), .A(n13189), .ZN(n8265) );
  AOI22_X1 U10501 ( .A1(n8275), .A2(n8274), .B1(n8267), .B2(n8266), .ZN(n8268)
         );
  INV_X1 U10502 ( .A(n8269), .ZN(n8272) );
  INV_X1 U10503 ( .A(n8270), .ZN(n8271) );
  NAND4_X1 U10504 ( .A1(n6536), .A2(n8304), .A3(n8272), .A4(n8271), .ZN(n8273)
         );
  INV_X1 U10505 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U10506 ( .A1(n8279), .A2(n8278), .ZN(n8285) );
  NAND2_X1 U10507 ( .A1(n7820), .A2(n13292), .ZN(n8283) );
  INV_X1 U10508 ( .A(n8280), .ZN(n8281) );
  NAND2_X1 U10509 ( .A1(n8281), .A2(n8214), .ZN(n8282) );
  MUX2_X1 U10510 ( .A(n8283), .B(n8282), .S(n8247), .Z(n8284) );
  NAND2_X1 U10511 ( .A1(n8285), .A2(n8284), .ZN(n8317) );
  INV_X1 U10512 ( .A(n10183), .ZN(n8286) );
  AND2_X1 U10513 ( .A1(n8286), .A2(n8263), .ZN(n9493) );
  OAI22_X1 U10514 ( .A1(n9493), .A2(n6754), .B1(n9497), .B2(n10922), .ZN(n8287) );
  INV_X1 U10515 ( .A(n13189), .ZN(n8306) );
  NAND2_X1 U10516 ( .A1(n13520), .A2(n13190), .ZN(n11823) );
  XNOR2_X1 U10517 ( .A(n13388), .B(n13126), .ZN(n13385) );
  INV_X1 U10518 ( .A(n13436), .ZN(n13170) );
  NAND2_X1 U10519 ( .A1(n13571), .A2(n13170), .ZN(n13431) );
  OR2_X1 U10520 ( .A1(n13571), .A2(n13170), .ZN(n8289) );
  INV_X1 U10521 ( .A(n13196), .ZN(n13446) );
  XNOR2_X1 U10522 ( .A(n13576), .B(n13446), .ZN(n11814) );
  INV_X1 U10523 ( .A(n13197), .ZN(n13169) );
  XNOR2_X1 U10524 ( .A(n13581), .B(n13169), .ZN(n13500) );
  XNOR2_X1 U10525 ( .A(n13587), .B(n13117), .ZN(n11497) );
  INV_X1 U10526 ( .A(n13199), .ZN(n11494) );
  XNOR2_X1 U10527 ( .A(n13593), .B(n11494), .ZN(n11483) );
  OR2_X1 U10528 ( .A1(n13598), .A2(n13200), .ZN(n11414) );
  NAND2_X1 U10529 ( .A1(n13598), .A2(n13200), .ZN(n11411) );
  AND2_X1 U10530 ( .A1(n11414), .A2(n11411), .ZN(n11312) );
  XNOR2_X1 U10531 ( .A(n13603), .B(n11309), .ZN(n11202) );
  INV_X1 U10532 ( .A(n13204), .ZN(n11061) );
  XNOR2_X1 U10533 ( .A(n11062), .B(n11061), .ZN(n11056) );
  INV_X1 U10534 ( .A(n13202), .ZN(n8290) );
  NAND2_X1 U10535 ( .A1(n11255), .A2(n8290), .ZN(n8291) );
  NAND2_X1 U10536 ( .A1(n11203), .A2(n8291), .ZN(n11198) );
  XNOR2_X1 U10537 ( .A(n11291), .B(n13203), .ZN(n11060) );
  XNOR2_X1 U10538 ( .A(n14878), .B(n10597), .ZN(n10429) );
  XNOR2_X1 U10539 ( .A(n10567), .B(n13208), .ZN(n10525) );
  INV_X1 U10540 ( .A(n14847), .ZN(n10377) );
  NAND4_X1 U10541 ( .A1(n14850), .A2(n9495), .A3(n9629), .A4(n10072), .ZN(
        n8294) );
  XNOR2_X1 U10542 ( .A(n13211), .B(n14860), .ZN(n10404) );
  NOR2_X1 U10543 ( .A1(n8294), .A2(n10404), .ZN(n8295) );
  XNOR2_X1 U10544 ( .A(n14868), .B(n13209), .ZN(n10272) );
  NAND4_X1 U10545 ( .A1(n10525), .A2(n8295), .A3(n10272), .A4(n9949), .ZN(
        n8296) );
  NOR2_X1 U10546 ( .A1(n10429), .A2(n8296), .ZN(n8297) );
  XNOR2_X1 U10547 ( .A(n10927), .B(n13205), .ZN(n10688) );
  NAND4_X1 U10548 ( .A1(n11060), .A2(n8297), .A3(n10688), .A4(n7118), .ZN(
        n8298) );
  OR4_X1 U10549 ( .A1(n13449), .A2(n11814), .A3(n13500), .A4(n8300), .ZN(n8301) );
  XNOR2_X1 U10550 ( .A(n13557), .B(n13091), .ZN(n13393) );
  INV_X1 U10551 ( .A(n13438), .ZN(n13137) );
  XNOR2_X1 U10552 ( .A(n13561), .B(n13137), .ZN(n13411) );
  INV_X1 U10553 ( .A(n13195), .ZN(n13448) );
  XNOR2_X1 U10554 ( .A(n13565), .B(n13448), .ZN(n13432) );
  NOR2_X1 U10555 ( .A1(n13385), .A2(n8302), .ZN(n8303) );
  XNOR2_X1 U10556 ( .A(n13369), .B(n13377), .ZN(n13363) );
  XNOR2_X1 U10557 ( .A(n13537), .B(n13193), .ZN(n13353) );
  NAND2_X1 U10558 ( .A1(n8312), .A2(n6754), .ZN(n8310) );
  INV_X1 U10559 ( .A(n8305), .ZN(n8309) );
  NAND3_X1 U10560 ( .A1(n8307), .A2(n8306), .A3(n6754), .ZN(n8308) );
  INV_X1 U10561 ( .A(n8312), .ZN(n8315) );
  NAND2_X1 U10562 ( .A1(n10924), .A2(n11500), .ZN(n8314) );
  MUX2_X1 U10563 ( .A(n8263), .B(n10924), .S(n10072), .Z(n8313) );
  OAI22_X1 U10564 ( .A1(n8315), .A2(n8314), .B1(n8313), .B2(n6754), .ZN(n8316)
         );
  INV_X1 U10565 ( .A(n8322), .ZN(n8319) );
  NAND2_X1 U10566 ( .A1(n8319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8331) );
  INV_X1 U10567 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8330) );
  XNOR2_X1 U10568 ( .A(n8331), .B(n8330), .ZN(n9333) );
  OR2_X1 U10569 ( .A1(n9333), .A2(P2_U3088), .ZN(n11110) );
  INV_X1 U10570 ( .A(n11110), .ZN(n8320) );
  NOR2_X1 U10571 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8321) );
  NAND2_X1 U10572 ( .A1(n8322), .A2(n8321), .ZN(n8326) );
  NAND2_X1 U10573 ( .A1(n8328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8323) );
  MUX2_X1 U10574 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8323), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8325) );
  NAND2_X1 U10575 ( .A1(n8325), .A2(n8324), .ZN(n13638) );
  INV_X1 U10576 ( .A(n13638), .ZN(n9472) );
  NAND2_X1 U10577 ( .A1(n8326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8327) );
  MUX2_X1 U10578 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8327), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8329) );
  NAND2_X1 U10579 ( .A1(n8329), .A2(n8328), .ZN(n11505) );
  NAND2_X1 U10580 ( .A1(n8331), .A2(n8330), .ZN(n8332) );
  NAND2_X1 U10581 ( .A1(n8332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8334) );
  INV_X1 U10582 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10583 ( .A(n8334), .B(n8333), .ZN(n11324) );
  NOR2_X1 U10584 ( .A1(n11505), .A2(n11324), .ZN(n8335) );
  NAND2_X1 U10585 ( .A1(n9472), .A2(n8335), .ZN(n9046) );
  AND2_X1 U10586 ( .A1(n9046), .A2(n9333), .ZN(n10079) );
  INV_X1 U10587 ( .A(n14843), .ZN(n14845) );
  INV_X1 U10588 ( .A(n9494), .ZN(n8337) );
  NAND2_X1 U10589 ( .A1(n10063), .A2(n8337), .ZN(n13445) );
  NOR4_X1 U10590 ( .A1(n14845), .A2(n6719), .A3(n10075), .A4(n13445), .ZN(
        n8339) );
  OAI21_X1 U10591 ( .B1(n11110), .B2(n6682), .A(P2_B_REG_SCAN_IN), .ZN(n8338)
         );
  OR2_X1 U10592 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  INV_X1 U10593 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14434) );
  INV_X1 U10594 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15193) );
  INV_X1 U10595 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14775) );
  INV_X1 U10596 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15069) );
  INV_X1 U10597 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10352) );
  INV_X1 U10598 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9603) );
  INV_X1 U10599 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U10600 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8364) );
  INV_X1 U10601 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9249) );
  XNOR2_X1 U10602 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n8368) );
  NAND2_X1 U10603 ( .A1(n8371), .A2(n8370), .ZN(n8341) );
  NAND2_X1 U10604 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8342), .ZN(n8344) );
  NAND2_X1 U10605 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8345), .ZN(n8346) );
  NAND2_X1 U10606 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8347), .ZN(n8349) );
  INV_X1 U10607 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9306) );
  OR2_X1 U10608 ( .A1(n9249), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n8350) );
  INV_X1 U10609 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10610 ( .A1(n8352), .A2(n8351), .ZN(n8354) );
  XOR2_X1 U10611 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8352), .Z(n8388) );
  INV_X1 U10612 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9237) );
  XNOR2_X1 U10613 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n9603), .ZN(n8394) );
  NOR2_X1 U10614 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8362), .ZN(n8358) );
  NAND2_X1 U10615 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8362), .ZN(n8357) );
  XOR2_X1 U10616 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n8399) );
  INV_X1 U10617 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15047) );
  AOI22_X1 U10618 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .B1(n15069), .B2(n15047), .ZN(n8402) );
  XOR2_X1 U10619 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n8361) );
  XNOR2_X1 U10620 ( .A(n8407), .B(n8361), .ZN(n14535) );
  INV_X1 U10621 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14531) );
  XNOR2_X1 U10622 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n8363) );
  XOR2_X1 U10623 ( .A(n8363), .B(n8362), .Z(n14421) );
  XOR2_X1 U10624 ( .A(n8365), .B(n8364), .Z(n8393) );
  NOR2_X1 U10625 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n8367), .ZN(n8380) );
  XNOR2_X1 U10626 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8367), .ZN(n15237) );
  INV_X1 U10627 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14394) );
  XNOR2_X1 U10628 ( .A(n8369), .B(n8368), .ZN(n14392) );
  NAND2_X1 U10629 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n8372), .ZN(n8373) );
  AOI21_X1 U10630 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n10198), .A(n8371), .ZN(
        n15240) );
  INV_X1 U10631 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15239) );
  NOR2_X1 U10632 ( .A1(n15240), .A2(n15239), .ZN(n15244) );
  NAND2_X1 U10633 ( .A1(n14392), .A2(n14393), .ZN(n8374) );
  NOR2_X1 U10634 ( .A1(n14392), .A2(n14393), .ZN(n14391) );
  XNOR2_X1 U10635 ( .A(n13983), .B(n8375), .ZN(n8376) );
  NAND2_X1 U10636 ( .A1(n8377), .A2(n8376), .ZN(n8378) );
  NOR2_X1 U10637 ( .A1(n15237), .A2(n15236), .ZN(n8379) );
  NAND2_X1 U10638 ( .A1(n8384), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8387) );
  XOR2_X1 U10639 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n8385) );
  XOR2_X1 U10640 ( .A(n8386), .B(n8385), .Z(n14407) );
  XNOR2_X1 U10641 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8388), .ZN(n15242) );
  NAND2_X1 U10642 ( .A1(n15241), .A2(n15242), .ZN(n8391) );
  NAND2_X1 U10643 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n8389), .ZN(n8390) );
  XNOR2_X1 U10644 ( .A(n8395), .B(n8394), .ZN(n8397) );
  NAND2_X1 U10645 ( .A1(n8396), .A2(n8397), .ZN(n8398) );
  NAND2_X1 U10646 ( .A1(n14421), .A2(n14420), .ZN(n14419) );
  XNOR2_X1 U10647 ( .A(n8400), .B(n8399), .ZN(n14530) );
  NAND2_X1 U10648 ( .A1(n14529), .A2(n14530), .ZN(n8401) );
  AOI21_X2 U10649 ( .B1(n14531), .B2(n8401), .A(n14528), .ZN(n8404) );
  XNOR2_X1 U10650 ( .A(n8403), .B(n8402), .ZN(n8405) );
  XNOR2_X1 U10651 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8408) );
  INV_X1 U10652 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14915) );
  INV_X1 U10653 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14560) );
  NOR2_X1 U10654 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14560), .ZN(n8406) );
  XNOR2_X1 U10655 ( .A(n8408), .B(n8412), .ZN(n14540) );
  NAND2_X1 U10656 ( .A1(n14539), .A2(n14540), .ZN(n8409) );
  NOR2_X1 U10657 ( .A1(n14539), .A2(n14540), .ZN(n14538) );
  INV_X1 U10658 ( .A(n8410), .ZN(n8415) );
  INV_X1 U10659 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8411) );
  NOR2_X1 U10660 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n8411), .ZN(n8413) );
  INV_X1 U10661 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14575) );
  OAI22_X1 U10662 ( .A1(n8413), .A2(n8412), .B1(P3_ADDR_REG_14__SCAN_IN), .B2(
        n14575), .ZN(n8417) );
  XOR2_X1 U10663 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n8414) );
  XOR2_X1 U10664 ( .A(n8417), .B(n8414), .Z(n8416) );
  XNOR2_X1 U10665 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .ZN(n8419) );
  INV_X1 U10666 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14587) );
  NOR2_X1 U10667 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14587), .ZN(n8418) );
  INV_X1 U10668 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12599) );
  OAI22_X1 U10669 ( .A1(n8418), .A2(n8417), .B1(P1_ADDR_REG_15__SCAN_IN), .B2(
        n12599), .ZN(n8423) );
  XOR2_X1 U10670 ( .A(n8419), .B(n8423), .Z(n8420) );
  NOR2_X1 U10671 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14545), .ZN(n8422) );
  INV_X1 U10672 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n8428) );
  INV_X1 U10673 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14600) );
  INV_X1 U10674 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12637) );
  NOR2_X1 U10675 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12637), .ZN(n8424) );
  OAI22_X1 U10676 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14600), .B1(n8424), 
        .B2(n8423), .ZN(n8426) );
  XNOR2_X1 U10677 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8426), .ZN(n8427) );
  XNOR2_X1 U10678 ( .A(n8428), .B(n8427), .ZN(n14432) );
  NAND2_X1 U10679 ( .A1(n14433), .A2(n14432), .ZN(n8425) );
  NOR2_X1 U10680 ( .A1(n14433), .A2(n14432), .ZN(n14431) );
  NOR2_X1 U10681 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8426), .ZN(n8430) );
  NOR2_X1 U10682 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  NOR2_X1 U10683 ( .A1(n8430), .A2(n8429), .ZN(n8437) );
  INV_X1 U10684 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8438) );
  NOR2_X1 U10685 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8438), .ZN(n8431) );
  AOI21_X1 U10686 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8438), .A(n8431), .ZN(
        n8432) );
  XOR2_X1 U10687 ( .A(n8437), .B(n8432), .Z(n8434) );
  XNOR2_X1 U10688 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8435) );
  INV_X1 U10689 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14634) );
  NOR2_X1 U10690 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14634), .ZN(n8436) );
  OAI22_X1 U10691 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8438), .B1(n8437), .B2(
        n8436), .ZN(n8439) );
  NAND2_X1 U10692 ( .A1(n9666), .A2(n8440), .ZN(n8597) );
  NAND4_X1 U10693 ( .A1(n8450), .A2(n8449), .A3(n8448), .A4(n8912), .ZN(n8942)
         );
  INV_X1 U10694 ( .A(n8942), .ZN(n8451) );
  NAND2_X1 U10695 ( .A1(n8451), .A2(n7390), .ZN(n8944) );
  NAND2_X1 U10696 ( .A1(n8509), .A2(n8511), .ZN(n8455) );
  INV_X1 U10697 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10698 ( .A1(n8455), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8457) );
  INV_X1 U10699 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8456) );
  INV_X1 U10700 ( .A(n6694), .ZN(n8458) );
  NAND2_X1 U10701 ( .A1(n8458), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8469) );
  INV_X1 U10702 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12910) );
  OR2_X1 U10703 ( .A1(n6484), .A2(n12910), .ZN(n8468) );
  NAND2_X4 U10704 ( .A1(n8461), .A2(n8460), .ZN(n8905) );
  NAND2_X1 U10705 ( .A1(n8605), .A2(n9751), .ZN(n8622) );
  OR2_X1 U10706 ( .A1(n8622), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8634) );
  NOR2_X1 U10707 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_8__SCAN_IN), 
        .ZN(n8462) );
  INV_X1 U10708 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12169) );
  INV_X1 U10709 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8761) );
  INV_X1 U10710 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8775) );
  INV_X1 U10711 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10712 ( .A1(n8821), .A2(n8820), .ZN(n8833) );
  INV_X1 U10713 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12273) );
  INV_X1 U10714 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15199) );
  INV_X1 U10715 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15029) );
  INV_X1 U10716 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U10717 ( .A1(n15029), .A2(n15182), .ZN(n8463) );
  INV_X1 U10718 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12196) );
  NOR2_X1 U10719 ( .A1(n8523), .A2(n12196), .ZN(n8464) );
  INV_X1 U10720 ( .A(n12724), .ZN(n8465) );
  OR2_X1 U10721 ( .A1(n6499), .A2(n8465), .ZN(n8467) );
  INV_X1 U10722 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12963) );
  OR2_X1 U10723 ( .A1(n8908), .A2(n12963), .ZN(n8466) );
  INV_X1 U10724 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14380) );
  INV_X1 U10725 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U10726 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n15204), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n15043), .ZN(n8840) );
  INV_X1 U10727 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9187) );
  AOI22_X1 U10728 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n9187), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7013), .ZN(n8798) );
  AOI22_X1 U10729 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n10126), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10128), .ZN(n8769) );
  NAND2_X1 U10730 ( .A1(n9069), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10731 ( .A1(n8472), .A2(n8471), .ZN(n8573) );
  NAND2_X1 U10732 ( .A1(n8584), .A2(n8582), .ZN(n8475) );
  NAND2_X1 U10733 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n9111), .ZN(n8477) );
  NAND2_X1 U10734 ( .A1(n8630), .A2(n8477), .ZN(n8479) );
  NAND2_X1 U10735 ( .A1(n9131), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10736 ( .A1(n6691), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U10737 ( .A1(n9168), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10738 ( .A1(n8684), .A2(n8683), .ZN(n8485) );
  NAND2_X1 U10739 ( .A1(n9199), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8484) );
  XNOR2_X1 U10740 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8701) );
  NAND2_X1 U10741 ( .A1(n8486), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U10742 ( .A1(n8724), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10743 ( .A1(n9436), .A2(n8488), .ZN(n8489) );
  XNOR2_X1 U10744 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8738) );
  INV_X1 U10745 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10746 ( .A1(n8491), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8492) );
  XNOR2_X1 U10747 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8754) );
  AOI22_X1 U10748 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10306), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10304), .ZN(n8783) );
  INV_X1 U10749 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10905) );
  INV_X1 U10750 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U10751 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10905), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n10950), .ZN(n8812) );
  NAND2_X1 U10752 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8496), .ZN(n8497) );
  AOI22_X1 U10753 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n10953), .B2(n8500), .ZN(n8852) );
  INV_X1 U10754 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U10755 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n8502), .B2(n11694), .ZN(n8865) );
  NAND2_X1 U10756 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8503), .ZN(n8504) );
  NAND2_X1 U10757 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n15202), .ZN(n8506) );
  INV_X1 U10758 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U10759 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n7043), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14380), .ZN(n8888) );
  INV_X1 U10760 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14374) );
  AOI22_X1 U10761 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8898), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14374), .ZN(n8507) );
  INV_X1 U10762 ( .A(n8507), .ZN(n8508) );
  XNOR2_X2 U10763 ( .A(n8512), .B(n8511), .ZN(n12542) );
  NAND2_X1 U10764 ( .A1(n8939), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8514) );
  INV_X1 U10765 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8513) );
  BUF_X4 U10766 ( .A(n8574), .Z(n12477) );
  NAND2_X1 U10767 ( .A1(n11564), .A2(n12477), .ZN(n8517) );
  NAND2_X1 U10768 ( .A1(n6483), .A2(SI_28_), .ZN(n8516) );
  AOI22_X1 U10769 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n11563), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n7036), .ZN(n8518) );
  XNOR2_X1 U10770 ( .A(n8519), .B(n8518), .ZN(n13049) );
  NAND2_X1 U10771 ( .A1(n13049), .A2(n12477), .ZN(n8521) );
  OR2_X1 U10772 ( .A1(n8515), .A2(n15031), .ZN(n8520) );
  NAND2_X2 U10773 ( .A1(n8521), .A2(n8520), .ZN(n12739) );
  INV_X1 U10774 ( .A(n12739), .ZN(n12968) );
  NAND2_X1 U10775 ( .A1(n8847), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8528) );
  OAI21_X1 U10776 ( .B1(n8892), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n8522) );
  INV_X1 U10777 ( .A(n8522), .ZN(n8524) );
  NOR2_X1 U10778 ( .A1(n8524), .A2(n8523), .ZN(n12736) );
  OR2_X1 U10779 ( .A1(n8905), .A2(n12736), .ZN(n8527) );
  NAND2_X1 U10780 ( .A1(n8458), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10781 ( .A1(n6495), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10782 ( .A1(n8847), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8534) );
  INV_X1 U10783 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12767) );
  OR2_X1 U10784 ( .A1(n6694), .A2(n12767), .ZN(n8533) );
  NAND2_X1 U10785 ( .A1(n8882), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U10786 ( .A1(n8892), .A2(n8529), .ZN(n12768) );
  INV_X1 U10787 ( .A(n12768), .ZN(n8530) );
  OR2_X1 U10788 ( .A1(n8905), .A2(n8530), .ZN(n8532) );
  INV_X1 U10789 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12919) );
  OR2_X1 U10790 ( .A1(n6484), .A2(n12919), .ZN(n8531) );
  AOI22_X1 U10791 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(
        P2_DATAO_REG_25__SCAN_IN), .B1(n11715), .B2(n15202), .ZN(n8535) );
  XNOR2_X1 U10792 ( .A(n8536), .B(n8535), .ZN(n11387) );
  NAND2_X1 U10793 ( .A1(n11387), .A2(n12477), .ZN(n8538) );
  NAND2_X1 U10794 ( .A1(n6483), .A2(SI_25_), .ZN(n8537) );
  NAND2_X2 U10795 ( .A1(n8538), .A2(n8537), .ZN(n12975) );
  NAND2_X1 U10796 ( .A1(n8575), .A2(SI_1_), .ZN(n8541) );
  XNOR2_X1 U10797 ( .A(n8539), .B(n8555), .ZN(n9079) );
  OAI211_X2 U10798 ( .C1(n9646), .C2(n9906), .A(n8541), .B(n8540), .ZN(n10826)
         );
  INV_X1 U10799 ( .A(n10826), .ZN(n8560) );
  INV_X1 U10800 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8542) );
  INV_X1 U10801 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10802 ( .A1(n8564), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8545) );
  INV_X1 U10803 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U10804 ( .A1(n8560), .A2(n12564), .ZN(n12338) );
  INV_X1 U10805 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8548) );
  INV_X1 U10806 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n8549) );
  INV_X1 U10807 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8550) );
  OR2_X1 U10808 ( .A1(n6494), .A2(n8550), .ZN(n8552) );
  NAND2_X1 U10809 ( .A1(n6498), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8551) );
  INV_X1 U10810 ( .A(n8555), .ZN(n8557) );
  INV_X1 U10811 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U10812 ( .A1(n9255), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10813 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  MUX2_X1 U10814 ( .A(n8558), .B(SI_0_), .S(n9517), .Z(n13059) );
  MUX2_X1 U10815 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13059), .S(n9646), .Z(n10655)
         );
  NAND2_X1 U10816 ( .A1(n10830), .A2(n10655), .ZN(n10828) );
  NAND2_X1 U10817 ( .A1(n10827), .A2(n10828), .ZN(n8562) );
  NAND2_X1 U10818 ( .A1(n8559), .A2(n8560), .ZN(n8561) );
  NAND2_X1 U10819 ( .A1(n8562), .A2(n8561), .ZN(n14941) );
  INV_X1 U10820 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9652) );
  INV_X1 U10821 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n8563) );
  INV_X1 U10822 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U10823 ( .A1(n6498), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8565) );
  INV_X1 U10824 ( .A(n6500), .ZN(n9653) );
  INV_X1 U10825 ( .A(n8571), .ZN(n8572) );
  XNOR2_X1 U10826 ( .A(n8573), .B(n8572), .ZN(n9078) );
  NAND2_X1 U10827 ( .A1(n8574), .A2(n9078), .ZN(n8577) );
  NAND2_X1 U10828 ( .A1(n8575), .A2(n9077), .ZN(n8576) );
  OAI211_X1 U10829 ( .C1(n9653), .C2(n9646), .A(n8577), .B(n8576), .ZN(n14937)
         );
  INV_X1 U10830 ( .A(n12563), .ZN(n10158) );
  NAND2_X1 U10831 ( .A1(n6497), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8581) );
  INV_X1 U10832 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9704) );
  OR2_X1 U10833 ( .A1(n6490), .A2(n9704), .ZN(n8580) );
  OR2_X1 U10834 ( .A1(n8905), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8579) );
  INV_X1 U10835 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9703) );
  OR2_X1 U10836 ( .A1(n6494), .A2(n9703), .ZN(n8578) );
  AND4_X2 U10837 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n14945)
         );
  INV_X1 U10838 ( .A(SI_3_), .ZN(n9070) );
  NAND2_X1 U10839 ( .A1(n12478), .A2(n9070), .ZN(n8590) );
  INV_X1 U10840 ( .A(n8582), .ZN(n8583) );
  XNOR2_X1 U10841 ( .A(n8584), .B(n8583), .ZN(n9071) );
  NAND2_X1 U10842 ( .A1(n12477), .A2(n9071), .ZN(n8589) );
  INV_X1 U10843 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U10844 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8585), .ZN(n8586) );
  XNOR2_X1 U10845 ( .A(n8587), .B(n8586), .ZN(n9726) );
  OR2_X1 U10846 ( .A1(n9646), .A2(n7180), .ZN(n8588) );
  NAND2_X1 U10847 ( .A1(n14945), .A2(n10216), .ZN(n12345) );
  AND2_X2 U10848 ( .A1(n12345), .A2(n12347), .ZN(n12502) );
  INV_X1 U10849 ( .A(n12502), .ZN(n10211) );
  NAND2_X1 U10850 ( .A1(n12561), .A2(n10216), .ZN(n8591) );
  INV_X1 U10851 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10117) );
  OR2_X1 U10852 ( .A1(n6490), .A2(n10117), .ZN(n8596) );
  AND2_X1 U10853 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8592) );
  NOR2_X1 U10854 ( .A1(n8605), .A2(n8592), .ZN(n10118) );
  OR2_X1 U10855 ( .A1(n8905), .A2(n10118), .ZN(n8595) );
  INV_X1 U10856 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15016) );
  OR2_X1 U10857 ( .A1(n6494), .A2(n15016), .ZN(n8594) );
  NAND2_X1 U10858 ( .A1(n6498), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8593) );
  NAND4_X1 U10859 ( .A1(n8596), .A2(n8595), .A3(n8594), .A4(n8593), .ZN(n12560) );
  NAND2_X1 U10860 ( .A1(n8597), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8598) );
  MUX2_X1 U10861 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8598), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8599) );
  AND2_X1 U10862 ( .A1(n8599), .A2(n8613), .ZN(n9729) );
  XNOR2_X1 U10863 ( .A(n8601), .B(n6931), .ZN(n9075) );
  NAND2_X1 U10864 ( .A1(n12477), .A2(n9075), .ZN(n8603) );
  INV_X1 U10865 ( .A(SI_4_), .ZN(n9074) );
  NAND2_X1 U10866 ( .A1(n12478), .A2(n9074), .ZN(n8602) );
  OAI211_X1 U10867 ( .C1(n9729), .C2(n9646), .A(n8603), .B(n8602), .ZN(n10147)
         );
  NAND2_X1 U10868 ( .A1(n12560), .A2(n6914), .ZN(n8604) );
  NAND2_X1 U10869 ( .A1(n6498), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8610) );
  INV_X1 U10870 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10869) );
  OR2_X1 U10871 ( .A1(n6490), .A2(n10869), .ZN(n8609) );
  OR2_X1 U10872 ( .A1(n8605), .A2(n9751), .ZN(n8606) );
  AND2_X1 U10873 ( .A1(n8622), .A2(n8606), .ZN(n10870) );
  OR2_X1 U10874 ( .A1(n8905), .A2(n10870), .ZN(n8608) );
  INV_X1 U10875 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9712) );
  OR2_X1 U10876 ( .A1(n6494), .A2(n9712), .ZN(n8607) );
  INV_X1 U10877 ( .A(SI_5_), .ZN(n9085) );
  NAND2_X1 U10878 ( .A1(n6483), .A2(n9085), .ZN(n8619) );
  XNOR2_X1 U10879 ( .A(n8611), .B(n6612), .ZN(n9086) );
  NAND2_X1 U10880 ( .A1(n12477), .A2(n9086), .ZN(n8618) );
  INV_X1 U10881 ( .A(n8612), .ZN(n8616) );
  NAND2_X1 U10882 ( .A1(n8613), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8614) );
  MUX2_X1 U10883 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8614), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8615) );
  NAND2_X1 U10884 ( .A1(n8616), .A2(n8615), .ZN(n9757) );
  OR2_X1 U10885 ( .A1(n9646), .A2(n7084), .ZN(n8617) );
  NAND2_X1 U10886 ( .A1(n10844), .A2(n14976), .ZN(n12356) );
  INV_X1 U10887 ( .A(n10844), .ZN(n10150) );
  INV_X1 U10888 ( .A(n14976), .ZN(n10168) );
  NAND2_X1 U10889 ( .A1(n10844), .A2(n10168), .ZN(n8621) );
  NAND2_X1 U10890 ( .A1(n8847), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8627) );
  INV_X1 U10891 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9716) );
  OR2_X1 U10892 ( .A1(n6490), .A2(n9716), .ZN(n8626) );
  NAND2_X1 U10893 ( .A1(n8622), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8623) );
  AND2_X1 U10894 ( .A1(n8634), .A2(n8623), .ZN(n10840) );
  OR2_X1 U10895 ( .A1(n8905), .A2(n10840), .ZN(n8625) );
  INV_X1 U10896 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15019) );
  OR2_X1 U10897 ( .A1(n6484), .A2(n15019), .ZN(n8624) );
  OR2_X1 U10898 ( .A1(n8612), .A2(n13044), .ZN(n8628) );
  XNOR2_X1 U10899 ( .A(n8628), .B(n8642), .ZN(n9739) );
  NAND2_X1 U10900 ( .A1(n6483), .A2(SI_6_), .ZN(n8632) );
  XNOR2_X1 U10901 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8629) );
  XNOR2_X1 U10902 ( .A(n8630), .B(n8629), .ZN(n9082) );
  NAND2_X1 U10903 ( .A1(n12477), .A2(n9082), .ZN(n8631) );
  OAI211_X1 U10904 ( .C1(n9646), .C2(n9739), .A(n8632), .B(n8631), .ZN(n10293)
         );
  NAND2_X1 U10905 ( .A1(n10779), .A2(n10293), .ZN(n12360) );
  INV_X2 U10906 ( .A(n10779), .ZN(n12559) );
  INV_X1 U10907 ( .A(n10293), .ZN(n14983) );
  NAND2_X1 U10908 ( .A1(n12559), .A2(n14983), .ZN(n12359) );
  NAND2_X1 U10909 ( .A1(n12360), .A2(n12359), .ZN(n10842) );
  NAND2_X1 U10910 ( .A1(n12559), .A2(n10293), .ZN(n8633) );
  NAND2_X1 U10911 ( .A1(n8847), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8639) );
  INV_X1 U10912 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10783) );
  OR2_X1 U10913 ( .A1(n6490), .A2(n10783), .ZN(n8638) );
  AND2_X1 U10914 ( .A1(n8634), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8635) );
  NOR2_X1 U10915 ( .A1(n8663), .A2(n8635), .ZN(n10784) );
  OR2_X1 U10916 ( .A1(n8905), .A2(n10784), .ZN(n8637) );
  INV_X1 U10917 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9779) );
  OR2_X1 U10918 ( .A1(n6494), .A2(n9779), .ZN(n8636) );
  INV_X1 U10919 ( .A(SI_7_), .ZN(n9072) );
  NAND2_X1 U10920 ( .A1(n6483), .A2(n9072), .ZN(n8647) );
  XNOR2_X1 U10921 ( .A(n6751), .B(n8640), .ZN(n9073) );
  NAND2_X1 U10922 ( .A1(n12477), .A2(n9073), .ZN(n8646) );
  NAND2_X1 U10923 ( .A1(n8612), .A2(n8642), .ZN(n8653) );
  NAND2_X1 U10924 ( .A1(n8653), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8644) );
  INV_X1 U10925 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8643) );
  XNOR2_X1 U10926 ( .A(n8644), .B(n8643), .ZN(n9791) );
  INV_X1 U10927 ( .A(n9791), .ZN(n9877) );
  OR2_X1 U10928 ( .A1(n9646), .A2(n9877), .ZN(n8645) );
  NAND2_X1 U10929 ( .A1(n10959), .A2(n14988), .ZN(n12364) );
  INV_X1 U10930 ( .A(n14988), .ZN(n10561) );
  NAND2_X1 U10931 ( .A1(n12558), .A2(n10561), .ZN(n12365) );
  NAND2_X2 U10932 ( .A1(n12364), .A2(n12365), .ZN(n10777) );
  NAND2_X1 U10933 ( .A1(n12558), .A2(n14988), .ZN(n8648) );
  NAND2_X1 U10934 ( .A1(n8847), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8652) );
  INV_X1 U10935 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n9865) );
  OR2_X1 U10936 ( .A1(n6490), .A2(n9865), .ZN(n8651) );
  XNOR2_X1 U10937 ( .A(n8663), .B(P3_REG3_REG_8__SCAN_IN), .ZN(n10960) );
  OR2_X1 U10938 ( .A1(n8905), .A2(n10960), .ZN(n8650) );
  INV_X1 U10939 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9864) );
  OR2_X1 U10940 ( .A1(n6484), .A2(n9864), .ZN(n8649) );
  INV_X1 U10941 ( .A(n8686), .ZN(n8657) );
  NAND2_X1 U10942 ( .A1(n8654), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8655) );
  MUX2_X1 U10943 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8655), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8656) );
  NAND2_X1 U10944 ( .A1(n8657), .A2(n8656), .ZN(n9880) );
  NAND2_X1 U10945 ( .A1(n6483), .A2(SI_8_), .ZN(n8660) );
  XNOR2_X1 U10946 ( .A(n8658), .B(n6613), .ZN(n9096) );
  NAND2_X1 U10947 ( .A1(n12477), .A2(n9096), .ZN(n8659) );
  OAI211_X1 U10948 ( .C1(n9646), .C2(n9880), .A(n8660), .B(n8659), .ZN(n15000)
         );
  NAND2_X1 U10949 ( .A1(n10986), .A2(n15000), .ZN(n12369) );
  INV_X1 U10950 ( .A(n10986), .ZN(n12557) );
  INV_X1 U10951 ( .A(n15000), .ZN(n10961) );
  NAND2_X1 U10952 ( .A1(n12557), .A2(n10961), .ZN(n12370) );
  NAND2_X1 U10953 ( .A1(n10986), .A2(n10961), .ZN(n8662) );
  AND2_X2 U10954 ( .A1(n10955), .A2(n8662), .ZN(n10985) );
  NAND2_X1 U10955 ( .A1(n8847), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8668) );
  INV_X1 U10956 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10309) );
  OR2_X1 U10957 ( .A1(n6490), .A2(n10309), .ZN(n8667) );
  INV_X1 U10958 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10308) );
  OR2_X1 U10959 ( .A1(n6484), .A2(n10308), .ZN(n8666) );
  INV_X1 U10960 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9873) );
  INV_X1 U10961 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10318) );
  AOI21_X1 U10962 ( .B1(n8663), .B2(n9873), .A(n10318), .ZN(n8664) );
  OR2_X1 U10963 ( .A1(n8677), .A2(n8664), .ZN(n10946) );
  INV_X1 U10964 ( .A(n10946), .ZN(n10990) );
  OR2_X1 U10965 ( .A1(n8905), .A2(n10990), .ZN(n8665) );
  OR2_X1 U10966 ( .A1(n8686), .A2(n13044), .ZN(n8669) );
  INV_X1 U10967 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8685) );
  XNOR2_X1 U10968 ( .A(n8669), .B(n8685), .ZN(n14399) );
  XNOR2_X1 U10969 ( .A(n8671), .B(n8670), .ZN(n14396) );
  NAND2_X1 U10970 ( .A1(n12477), .A2(n14396), .ZN(n8674) );
  INV_X1 U10971 ( .A(SI_9_), .ZN(n8672) );
  NAND2_X1 U10972 ( .A1(n6483), .A2(n8672), .ZN(n8673) );
  OAI211_X1 U10973 ( .C1(n10491), .C2(n9646), .A(n8674), .B(n8673), .ZN(n15005) );
  NAND2_X1 U10974 ( .A1(n11085), .A2(n15005), .ZN(n8675) );
  INV_X1 U10975 ( .A(n15005), .ZN(n12385) );
  NAND2_X1 U10976 ( .A1(n8847), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8682) );
  INV_X1 U10977 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11025) );
  OR2_X1 U10978 ( .A1(n6490), .A2(n11025), .ZN(n8681) );
  OR2_X1 U10979 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  AND2_X1 U10980 ( .A1(n8707), .A2(n8678), .ZN(n11086) );
  OR2_X1 U10981 ( .A1(n8905), .A2(n11086), .ZN(n8680) );
  INV_X1 U10982 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10478) );
  OR2_X1 U10983 ( .A1(n6484), .A2(n10478), .ZN(n8679) );
  XNOR2_X1 U10984 ( .A(n8684), .B(n8683), .ZN(n9091) );
  NAND2_X1 U10985 ( .A1(n12477), .A2(n9091), .ZN(n8690) );
  INV_X1 U10986 ( .A(SI_10_), .ZN(n9090) );
  NAND2_X1 U10987 ( .A1(n6483), .A2(n9090), .ZN(n8689) );
  NAND2_X1 U10988 ( .A1(n8686), .A2(n8685), .ZN(n8698) );
  NAND2_X1 U10989 ( .A1(n8698), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8687) );
  XNOR2_X1 U10990 ( .A(n8687), .B(n15098), .ZN(n11186) );
  INV_X1 U10991 ( .A(n11186), .ZN(n10489) );
  OR2_X1 U10992 ( .A1(n9646), .A2(n10489), .ZN(n8688) );
  NAND2_X1 U10993 ( .A1(n11274), .A2(n11089), .ZN(n12375) );
  INV_X1 U10994 ( .A(n11089), .ZN(n11254) );
  NAND2_X1 U10995 ( .A1(n12555), .A2(n11254), .ZN(n8989) );
  NAND2_X1 U10996 ( .A1(n12375), .A2(n8989), .ZN(n12511) );
  NAND2_X1 U10997 ( .A1(n12555), .A2(n11089), .ZN(n8691) );
  NAND2_X1 U10998 ( .A1(n8847), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8697) );
  INV_X1 U10999 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8692) );
  OR2_X1 U11000 ( .A1(n6490), .A2(n8692), .ZN(n8696) );
  INV_X1 U11001 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11331) );
  XNOR2_X1 U11002 ( .A(n8707), .B(n11331), .ZN(n11332) );
  OR2_X1 U11003 ( .A1(n8905), .A2(n11332), .ZN(n8695) );
  INV_X1 U11004 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8693) );
  OR2_X1 U11005 ( .A1(n6484), .A2(n8693), .ZN(n8694) );
  OAI21_X1 U11006 ( .B1(n8698), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8700) );
  INV_X1 U11007 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11008 ( .A(n8700), .B(n8699), .ZN(n14900) );
  XNOR2_X1 U11009 ( .A(n8702), .B(n8701), .ZN(n14400) );
  NAND2_X1 U11010 ( .A1(n12477), .A2(n14400), .ZN(n8705) );
  NAND2_X1 U11011 ( .A1(n6483), .A2(n8703), .ZN(n8704) );
  OAI211_X1 U11012 ( .C1(n11188), .C2(n9646), .A(n8705), .B(n8704), .ZN(n14448) );
  NAND2_X1 U11013 ( .A1(n12380), .A2(n14448), .ZN(n8706) );
  NAND2_X1 U11014 ( .A1(n8847), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8712) );
  INV_X1 U11015 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11302) );
  OR2_X1 U11016 ( .A1(n6490), .A2(n11302), .ZN(n8711) );
  OAI21_X1 U11017 ( .B1(n8707), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8708) );
  AND2_X1 U11018 ( .A1(n8708), .A2(n8729), .ZN(n11371) );
  OR2_X1 U11019 ( .A1(n8905), .A2(n11371), .ZN(n8710) );
  INV_X1 U11020 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11175) );
  OR2_X1 U11021 ( .A1(n6484), .A2(n11175), .ZN(n8709) );
  AND2_X1 U11022 ( .A1(n8713), .A2(n8612), .ZN(n8716) );
  NOR2_X1 U11023 ( .A1(n8716), .A2(n13044), .ZN(n8714) );
  MUX2_X1 U11024 ( .A(n13044), .B(n8714), .S(P3_IR_REG_12__SCAN_IN), .Z(n8718)
         );
  NAND2_X1 U11025 ( .A1(n8716), .A2(n8715), .ZN(n8740) );
  INV_X1 U11026 ( .A(n8740), .ZN(n8717) );
  NAND2_X1 U11027 ( .A1(n6483), .A2(SI_12_), .ZN(n8721) );
  XNOR2_X1 U11028 ( .A(n8719), .B(n6627), .ZN(n9123) );
  NAND2_X1 U11029 ( .A1(n12477), .A2(n9123), .ZN(n8720) );
  OAI211_X1 U11030 ( .C1(n9646), .C2(n12582), .A(n8721), .B(n8720), .ZN(n11377) );
  NAND2_X1 U11031 ( .A1(n12264), .A2(n11377), .ZN(n12390) );
  INV_X1 U11032 ( .A(n11377), .ZN(n14444) );
  NAND2_X1 U11033 ( .A1(n12553), .A2(n14444), .ZN(n12391) );
  NAND2_X1 U11034 ( .A1(n12390), .A2(n12391), .ZN(n11300) );
  NAND2_X1 U11035 ( .A1(n11299), .A2(n11300), .ZN(n8723) );
  NAND2_X1 U11036 ( .A1(n12553), .A2(n11377), .ZN(n8722) );
  NAND2_X1 U11037 ( .A1(n8723), .A2(n8722), .ZN(n11381) );
  XNOR2_X1 U11038 ( .A(n8724), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U11039 ( .A1(n14404), .A2(n12477), .ZN(n8728) );
  INV_X1 U11040 ( .A(n9646), .ZN(n8817) );
  NAND2_X1 U11041 ( .A1(n8740), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8726) );
  XNOR2_X1 U11042 ( .A(n8726), .B(n8725), .ZN(n14917) );
  AOI22_X1 U11043 ( .A1(n6483), .A2(n14403), .B1(n8817), .B2(n14917), .ZN(
        n8727) );
  NAND2_X1 U11044 ( .A1(n8728), .A2(n8727), .ZN(n14440) );
  INV_X1 U11045 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11383) );
  OR2_X1 U11046 ( .A1(n6490), .A2(n11383), .ZN(n8735) );
  AND2_X1 U11047 ( .A1(n8729), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8730) );
  NOR2_X1 U11048 ( .A1(n8746), .A2(n8730), .ZN(n12267) );
  OR2_X1 U11049 ( .A1(n8905), .A2(n12267), .ZN(n8734) );
  INV_X1 U11050 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8731) );
  OR2_X1 U11051 ( .A1(n6484), .A2(n8731), .ZN(n8733) );
  NAND2_X1 U11052 ( .A1(n6497), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8732) );
  NAND4_X1 U11053 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n12899) );
  OR2_X1 U11054 ( .A1(n14440), .A2(n12899), .ZN(n12398) );
  NAND2_X1 U11055 ( .A1(n14440), .A2(n12899), .ZN(n12397) );
  NAND2_X1 U11056 ( .A1(n12398), .A2(n12397), .ZN(n12395) );
  NAND2_X1 U11057 ( .A1(n11381), .A2(n12395), .ZN(n8737) );
  INV_X1 U11058 ( .A(n12899), .ZN(n12171) );
  OR2_X1 U11059 ( .A1(n14440), .A2(n12171), .ZN(n8736) );
  NAND2_X1 U11060 ( .A1(n8737), .A2(n8736), .ZN(n12893) );
  XNOR2_X1 U11061 ( .A(n8739), .B(n8738), .ZN(n9171) );
  NAND2_X1 U11062 ( .A1(n9171), .A2(n12477), .ZN(n8744) );
  OR2_X1 U11063 ( .A1(n8740), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11064 ( .A1(n8757), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U11065 ( .A(n8742), .B(n8741), .ZN(n12580) );
  AOI22_X1 U11066 ( .A1(n6483), .A2(n15172), .B1(n8817), .B2(n12580), .ZN(
        n8743) );
  INV_X1 U11067 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11068 ( .A1(n6694), .A2(n8745), .ZN(n8751) );
  INV_X1 U11069 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12956) );
  OR2_X1 U11070 ( .A1(n6484), .A2(n12956), .ZN(n8750) );
  NOR2_X1 U11071 ( .A1(n8746), .A2(n12169), .ZN(n8747) );
  OR2_X1 U11072 ( .A1(n8762), .A2(n8747), .ZN(n12174) );
  INV_X1 U11073 ( .A(n12174), .ZN(n12902) );
  OR2_X1 U11074 ( .A1(n6499), .A2(n12902), .ZN(n8749) );
  NAND2_X1 U11075 ( .A1(n8847), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8748) );
  NAND4_X1 U11076 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n12885) );
  OR2_X1 U11077 ( .A1(n13038), .A2(n12885), .ZN(n12402) );
  NAND2_X1 U11078 ( .A1(n13038), .A2(n12885), .ZN(n12401) );
  NAND2_X1 U11079 ( .A1(n12402), .A2(n12401), .ZN(n12900) );
  NAND2_X1 U11080 ( .A1(n12893), .A2(n12900), .ZN(n8753) );
  INV_X1 U11081 ( .A(n12885), .ZN(n12124) );
  OR2_X1 U11082 ( .A1(n13038), .A2(n12124), .ZN(n8752) );
  NAND2_X1 U11083 ( .A1(n8753), .A2(n8752), .ZN(n12881) );
  INV_X1 U11084 ( .A(n8754), .ZN(n8755) );
  XNOR2_X1 U11085 ( .A(n8756), .B(n8755), .ZN(n14409) );
  NAND2_X1 U11086 ( .A1(n14409), .A2(n12477), .ZN(n8760) );
  OAI21_X1 U11087 ( .B1(n8757), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8758) );
  XNOR2_X1 U11088 ( .A(n8758), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U11089 ( .A1(n6483), .A2(SI_15_), .B1(n8817), .B2(n12628), .ZN(
        n8759) );
  NAND2_X1 U11090 ( .A1(n6498), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8767) );
  INV_X1 U11091 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12886) );
  OR2_X1 U11092 ( .A1(n6694), .A2(n12886), .ZN(n8766) );
  INV_X1 U11093 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12952) );
  OR2_X1 U11094 ( .A1(n6494), .A2(n12952), .ZN(n8765) );
  NOR2_X1 U11095 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  OR2_X1 U11096 ( .A1(n8776), .A2(n8763), .ZN(n12887) );
  INV_X1 U11097 ( .A(n12887), .ZN(n12308) );
  OR2_X1 U11098 ( .A1(n8905), .A2(n12308), .ZN(n8764) );
  OR2_X1 U11099 ( .A1(n13027), .A2(n12299), .ZN(n12405) );
  NAND2_X1 U11100 ( .A1(n13027), .A2(n12299), .ZN(n12411) );
  NAND2_X1 U11101 ( .A1(n12405), .A2(n12411), .ZN(n12879) );
  NAND2_X1 U11102 ( .A1(n13027), .A2(n12897), .ZN(n8768) );
  INV_X1 U11103 ( .A(n8769), .ZN(n8770) );
  XNOR2_X1 U11104 ( .A(n8771), .B(n8770), .ZN(n14414) );
  NAND2_X1 U11105 ( .A1(n14414), .A2(n12477), .ZN(n8774) );
  NAND2_X1 U11106 ( .A1(n8786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8772) );
  XNOR2_X1 U11107 ( .A(n8772), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U11108 ( .A1(n6483), .A2(SI_16_), .B1(n8817), .B2(n12634), .ZN(
        n8773) );
  INV_X1 U11109 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12875) );
  OR2_X1 U11110 ( .A1(n6694), .A2(n12875), .ZN(n8781) );
  INV_X1 U11111 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12949) );
  OR2_X1 U11112 ( .A1(n6494), .A2(n12949), .ZN(n8780) );
  OR2_X1 U11113 ( .A1(n8776), .A2(n8775), .ZN(n8777) );
  AND2_X1 U11114 ( .A1(n8792), .A2(n8777), .ZN(n12225) );
  OR2_X1 U11115 ( .A1(n8905), .A2(n12225), .ZN(n8779) );
  NAND2_X1 U11116 ( .A1(n8847), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8778) );
  NAND4_X1 U11117 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(n12884) );
  AND2_X1 U11118 ( .A1(n13021), .A2(n12884), .ZN(n8782) );
  INV_X1 U11119 ( .A(n13021), .ZN(n12230) );
  INV_X1 U11120 ( .A(n12884), .ZN(n12406) );
  INV_X1 U11121 ( .A(n8783), .ZN(n8784) );
  XNOR2_X1 U11122 ( .A(n8785), .B(n8784), .ZN(n9548) );
  NAND2_X1 U11123 ( .A1(n9548), .A2(n12477), .ZN(n8790) );
  NAND2_X1 U11124 ( .A1(n8945), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8787) );
  MUX2_X1 U11125 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8787), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8788) );
  NAND2_X1 U11126 ( .A1(n8788), .A2(n8814), .ZN(n12664) );
  INV_X1 U11127 ( .A(n12664), .ZN(n12671) );
  AOI22_X1 U11128 ( .A1(n6483), .A2(SI_17_), .B1(n8817), .B2(n12671), .ZN(
        n8789) );
  NAND2_X1 U11129 ( .A1(n8847), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8796) );
  INV_X1 U11130 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12866) );
  OR2_X1 U11131 ( .A1(n6694), .A2(n12866), .ZN(n8795) );
  AOI21_X1 U11132 ( .B1(n8792), .B2(P3_REG3_REG_17__SCAN_IN), .A(n8791), .ZN(
        n12234) );
  OR2_X1 U11133 ( .A1(n6499), .A2(n12234), .ZN(n8794) );
  INV_X1 U11134 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n15058) );
  OR2_X1 U11135 ( .A1(n6484), .A2(n15058), .ZN(n8793) );
  OR2_X1 U11136 ( .A1(n13015), .A2(n12850), .ZN(n12417) );
  NAND2_X1 U11137 ( .A1(n13015), .A2(n12850), .ZN(n12416) );
  NAND2_X1 U11138 ( .A1(n13015), .A2(n12873), .ZN(n8797) );
  INV_X1 U11139 ( .A(n8798), .ZN(n8799) );
  XNOR2_X1 U11140 ( .A(n8800), .B(n8799), .ZN(n9640) );
  NAND2_X1 U11141 ( .A1(n9640), .A2(n12477), .ZN(n8803) );
  NAND2_X1 U11142 ( .A1(n8814), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8801) );
  XNOR2_X1 U11143 ( .A(n8801), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U11144 ( .A1(n6483), .A2(SI_18_), .B1(n8817), .B2(n12688), .ZN(
        n8802) );
  NAND2_X1 U11145 ( .A1(n8847), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8810) );
  INV_X1 U11146 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8804) );
  OR2_X1 U11147 ( .A1(n6694), .A2(n8804), .ZN(n8809) );
  AND2_X1 U11148 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(n8805), .ZN(n8806) );
  NOR2_X1 U11149 ( .A1(n8821), .A2(n8806), .ZN(n12853) );
  OR2_X1 U11150 ( .A1(n8905), .A2(n12853), .ZN(n8808) );
  INV_X1 U11151 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12945) );
  OR2_X1 U11152 ( .A1(n6484), .A2(n12945), .ZN(n8807) );
  NAND2_X1 U11153 ( .A1(n12944), .A2(n12858), .ZN(n12423) );
  NAND2_X1 U11154 ( .A1(n12830), .A2(n12423), .ZN(n12842) );
  OR2_X1 U11155 ( .A1(n12944), .A2(n12834), .ZN(n8811) );
  XNOR2_X1 U11156 ( .A(n8813), .B(n8812), .ZN(n9773) );
  NAND2_X1 U11157 ( .A1(n9773), .A2(n12477), .ZN(n8819) );
  INV_X1 U11158 ( .A(n8913), .ZN(n8815) );
  NAND2_X1 U11159 ( .A1(n8815), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8816) );
  AOI22_X1 U11160 ( .A1(n6483), .A2(n9774), .B1(n8817), .B2(n12694), .ZN(n8818) );
  NAND2_X1 U11161 ( .A1(n6497), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8826) );
  INV_X1 U11162 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12837) );
  OR2_X1 U11163 ( .A1(n6694), .A2(n12837), .ZN(n8825) );
  OR2_X1 U11164 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  AND2_X1 U11165 ( .A1(n8822), .A2(n8833), .ZN(n12838) );
  OR2_X1 U11166 ( .A1(n8905), .A2(n12838), .ZN(n8824) );
  INV_X1 U11167 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12940) );
  OR2_X1 U11168 ( .A1(n6494), .A2(n12940), .ZN(n8823) );
  INV_X1 U11169 ( .A(n12522), .ZN(n13005) );
  NAND2_X1 U11170 ( .A1(n13005), .A2(n12552), .ZN(n8827) );
  XNOR2_X1 U11171 ( .A(n8829), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10383) );
  NAND2_X1 U11172 ( .A1(n10383), .A2(n12477), .ZN(n8831) );
  NAND2_X1 U11173 ( .A1(n6483), .A2(SI_20_), .ZN(n8830) );
  NAND2_X1 U11174 ( .A1(n8847), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8838) );
  INV_X1 U11175 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n8832) );
  OR2_X1 U11176 ( .A1(n6694), .A2(n8832), .ZN(n8837) );
  NAND2_X1 U11177 ( .A1(n8833), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8834) );
  AND2_X1 U11178 ( .A1(n8845), .A2(n8834), .ZN(n12826) );
  OR2_X1 U11179 ( .A1(n6499), .A2(n12826), .ZN(n8836) );
  INV_X1 U11180 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12938) );
  OR2_X1 U11181 ( .A1(n6484), .A2(n12938), .ZN(n8835) );
  INV_X1 U11182 ( .A(n12811), .ZN(n12835) );
  AND2_X1 U11183 ( .A1(n12937), .A2(n12835), .ZN(n8839) );
  INV_X1 U11184 ( .A(n8840), .ZN(n8841) );
  XNOR2_X1 U11185 ( .A(n8842), .B(n8841), .ZN(n10576) );
  NAND2_X1 U11186 ( .A1(n10576), .A2(n12477), .ZN(n8844) );
  NAND2_X1 U11187 ( .A1(n6483), .A2(SI_21_), .ZN(n8843) );
  INV_X1 U11188 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12814) );
  OR2_X1 U11189 ( .A1(n6694), .A2(n12814), .ZN(n8851) );
  AND2_X1 U11190 ( .A1(n8845), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8846) );
  NOR2_X1 U11191 ( .A1(n8856), .A2(n8846), .ZN(n12813) );
  OR2_X1 U11192 ( .A1(n6499), .A2(n12813), .ZN(n8850) );
  INV_X1 U11193 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12934) );
  OR2_X1 U11194 ( .A1(n6484), .A2(n12934), .ZN(n8849) );
  NAND2_X1 U11195 ( .A1(n8847), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8848) );
  NAND4_X1 U11196 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(n12800) );
  NAND2_X1 U11197 ( .A1(n12933), .A2(n12800), .ZN(n12434) );
  OR2_X1 U11198 ( .A1(n12933), .A2(n12800), .ZN(n12435) );
  XNOR2_X1 U11199 ( .A(n8853), .B(n8852), .ZN(n10701) );
  NAND2_X1 U11200 ( .A1(n10701), .A2(n12477), .ZN(n8855) );
  NAND2_X1 U11201 ( .A1(n6483), .A2(SI_22_), .ZN(n8854) );
  INV_X1 U11202 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12803) );
  OR2_X1 U11203 ( .A1(n6694), .A2(n12803), .ZN(n8861) );
  NOR2_X1 U11204 ( .A1(n8856), .A2(n12273), .ZN(n8857) );
  OR2_X1 U11205 ( .A1(n8869), .A2(n8857), .ZN(n12804) );
  INV_X1 U11206 ( .A(n12804), .ZN(n12276) );
  OR2_X1 U11207 ( .A1(n8905), .A2(n12276), .ZN(n8860) );
  INV_X1 U11208 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12929) );
  OR2_X1 U11209 ( .A1(n6494), .A2(n12929), .ZN(n8859) );
  NAND2_X1 U11210 ( .A1(n6497), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8858) );
  NAND4_X1 U11211 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n12551) );
  NAND2_X1 U11212 ( .A1(n12991), .A2(n12551), .ZN(n8863) );
  XNOR2_X1 U11213 ( .A(n8866), .B(n8865), .ZN(n10935) );
  NAND2_X1 U11214 ( .A1(n10935), .A2(n12477), .ZN(n8868) );
  NAND2_X1 U11215 ( .A1(n6483), .A2(SI_23_), .ZN(n8867) );
  INV_X1 U11216 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12793) );
  OR2_X1 U11217 ( .A1(n6694), .A2(n12793), .ZN(n8874) );
  INV_X1 U11218 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12927) );
  OR2_X1 U11219 ( .A1(n6494), .A2(n12927), .ZN(n8873) );
  OR2_X1 U11220 ( .A1(n8869), .A2(n15199), .ZN(n8870) );
  AND2_X1 U11221 ( .A1(n8880), .A2(n8870), .ZN(n12792) );
  OR2_X1 U11222 ( .A1(n8905), .A2(n12792), .ZN(n8872) );
  NAND2_X1 U11223 ( .A1(n6498), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8871) );
  NAND4_X1 U11224 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8871), .ZN(n12801) );
  NAND2_X1 U11225 ( .A1(n12154), .A2(n12801), .ZN(n12772) );
  INV_X1 U11226 ( .A(n12801), .ZN(n12447) );
  NAND2_X1 U11227 ( .A1(n12926), .A2(n12447), .ZN(n8875) );
  NAND2_X1 U11228 ( .A1(n12772), .A2(n8875), .ZN(n12788) );
  NAND2_X1 U11229 ( .A1(n12926), .A2(n12801), .ZN(n8876) );
  XNOR2_X1 U11230 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8877), .ZN(n11341) );
  NAND2_X1 U11231 ( .A1(n11341), .A2(n12477), .ZN(n8879) );
  NAND2_X1 U11232 ( .A1(n6483), .A2(SI_24_), .ZN(n8878) );
  INV_X2 U11233 ( .A(n12152), .ZN(n12981) );
  INV_X1 U11234 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12779) );
  OR2_X1 U11235 ( .A1(n6694), .A2(n12779), .ZN(n8886) );
  NAND2_X1 U11236 ( .A1(n8880), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8881) );
  AND2_X1 U11237 ( .A1(n8882), .A2(n8881), .ZN(n12780) );
  OR2_X1 U11238 ( .A1(n6499), .A2(n12780), .ZN(n8885) );
  INV_X1 U11239 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12922) );
  OR2_X1 U11240 ( .A1(n6484), .A2(n12922), .ZN(n8884) );
  NAND2_X1 U11241 ( .A1(n6498), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8883) );
  NAND4_X1 U11242 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n12764) );
  AND2_X1 U11243 ( .A1(n12981), .A2(n12764), .ZN(n8887) );
  NAND2_X1 U11244 ( .A1(n12975), .A2(n12292), .ZN(n12324) );
  NAND2_X1 U11245 ( .A1(n13053), .A2(n12477), .ZN(n8891) );
  NAND2_X1 U11246 ( .A1(n6483), .A2(SI_26_), .ZN(n8890) );
  NAND2_X2 U11247 ( .A1(n8891), .A2(n8890), .ZN(n12753) );
  INV_X1 U11248 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12751) );
  OR2_X1 U11249 ( .A1(n6694), .A2(n12751), .ZN(n8896) );
  INV_X1 U11250 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12917) );
  OR2_X1 U11251 ( .A1(n6494), .A2(n12917), .ZN(n8895) );
  XNOR2_X1 U11252 ( .A(n8892), .B(n15029), .ZN(n12750) );
  OR2_X1 U11253 ( .A1(n8905), .A2(n12750), .ZN(n8894) );
  NAND2_X1 U11254 ( .A1(n6497), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8893) );
  NAND4_X1 U11255 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n12763) );
  NOR2_X1 U11256 ( .A1(n12753), .A2(n12763), .ZN(n8897) );
  INV_X1 U11257 ( .A(n12753), .ZN(n12972) );
  NAND2_X1 U11258 ( .A1(n12200), .A2(n8926), .ZN(n8998) );
  NAND2_X1 U11259 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8898), .ZN(n8900) );
  AOI22_X1 U11260 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8237), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n11622), .ZN(n12112) );
  XNOR2_X1 U11261 ( .A(n12111), .B(n12112), .ZN(n12107) );
  NAND2_X1 U11262 ( .A1(n12107), .A2(n12477), .ZN(n8903) );
  NAND2_X1 U11263 ( .A1(n6483), .A2(SI_29_), .ZN(n8902) );
  INV_X1 U11264 ( .A(n12706), .ZN(n8904) );
  OR2_X1 U11265 ( .A1(n6694), .A2(n9037), .ZN(n8911) );
  INV_X1 U11266 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8906) );
  OR2_X1 U11267 ( .A1(n6484), .A2(n8906), .ZN(n8910) );
  INV_X1 U11268 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8907) );
  OR2_X1 U11269 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  NAND2_X1 U11270 ( .A1(n9036), .A2(n12720), .ZN(n12461) );
  INV_X1 U11271 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11272 ( .A1(n8955), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8916) );
  INV_X1 U11273 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11274 ( .A1(n12544), .A2(n12690), .ZN(n9011) );
  MUX2_X1 U11275 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8919), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8920) );
  NAND2_X2 U11276 ( .A1(n8920), .A2(n8955), .ZN(n12332) );
  NAND2_X1 U11277 ( .A1(n8922), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8923) );
  MUX2_X1 U11278 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8923), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8925) );
  NAND2_X1 U11279 ( .A1(n8925), .A2(n8924), .ZN(n10386) );
  NAND2_X1 U11280 ( .A1(n12329), .A2(n9012), .ZN(n12539) );
  INV_X1 U11281 ( .A(n12542), .ZN(n9648) );
  NAND2_X1 U11282 ( .A1(n9648), .A2(n9671), .ZN(n9664) );
  INV_X1 U11283 ( .A(n8926), .ZN(n12732) );
  INV_X1 U11284 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8927) );
  OR2_X1 U11285 ( .A1(n6694), .A2(n8927), .ZN(n8931) );
  INV_X1 U11286 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14439) );
  OR2_X1 U11287 ( .A1(n6484), .A2(n14439), .ZN(n8930) );
  NAND2_X1 U11288 ( .A1(n6498), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8929) );
  NAND4_X1 U11289 ( .A1(n12486), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(
        n12550) );
  NAND2_X1 U11290 ( .A1(n9664), .A2(n9646), .ZN(n8932) );
  INV_X1 U11291 ( .A(P3_B_REG_SCAN_IN), .ZN(n8933) );
  NOR2_X1 U11292 ( .A1(n12542), .A2(n8933), .ZN(n8934) );
  NOR2_X1 U11293 ( .A1(n14944), .A2(n8934), .ZN(n12707) );
  AOI22_X1 U11294 ( .A1(n12898), .A2(n12732), .B1(n12550), .B2(n12707), .ZN(
        n8935) );
  OAI21_X1 U11295 ( .B1(n8936), .B2(n12861), .A(n8935), .ZN(n9027) );
  NOR2_X1 U11296 ( .A1(n8937), .A2(n13044), .ZN(n8938) );
  MUX2_X1 U11297 ( .A(n13044), .B(n8938), .S(P3_IR_REG_26__SCAN_IN), .Z(n8941)
         );
  INV_X1 U11298 ( .A(n8939), .ZN(n8940) );
  NOR2_X1 U11299 ( .A1(n8945), .A2(n8944), .ZN(n8947) );
  INV_X1 U11300 ( .A(n8947), .ZN(n8946) );
  XNOR2_X1 U11301 ( .A(n11343), .B(P3_B_REG_SCAN_IN), .ZN(n8950) );
  NOR2_X1 U11302 ( .A1(n8947), .A2(n13044), .ZN(n8948) );
  INV_X1 U11303 ( .A(n8937), .ZN(n8949) );
  OR2_X1 U11304 ( .A1(n9170), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8952) );
  OR2_X1 U11305 ( .A1(n13052), .A2(n6700), .ZN(n8951) );
  INV_X1 U11306 ( .A(n11343), .ZN(n8953) );
  OR2_X1 U11307 ( .A1(n13052), .A2(n8953), .ZN(n8954) );
  NAND2_X1 U11308 ( .A1(n13040), .A2(n13042), .ZN(n9010) );
  OAI21_X1 U11309 ( .B1(n8955), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8957) );
  INV_X1 U11310 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8956) );
  XNOR2_X1 U11311 ( .A(n8957), .B(n8956), .ZN(n9966) );
  NOR2_X1 U11312 ( .A1(n11388), .A2(n11343), .ZN(n8958) );
  NAND2_X1 U11313 ( .A1(n13052), .A2(n8958), .ZN(n9967) );
  NOR2_X1 U11314 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8962) );
  NOR4_X1 U11315 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8961) );
  NOR4_X1 U11316 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8960) );
  NOR4_X1 U11317 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8959) );
  NAND4_X1 U11318 ( .A1(n8962), .A2(n8961), .A3(n8960), .A4(n8959), .ZN(n8968)
         );
  NOR4_X1 U11319 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8966) );
  NOR4_X1 U11320 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8965) );
  NOR4_X1 U11321 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8964) );
  NOR4_X1 U11322 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8963) );
  NAND4_X1 U11323 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n8967)
         );
  NOR2_X1 U11324 ( .A1(n8968), .A2(n8967), .ZN(n8969) );
  AND2_X1 U11325 ( .A1(n9995), .A2(n9009), .ZN(n8970) );
  INV_X1 U11326 ( .A(n13040), .ZN(n9029) );
  NAND2_X1 U11327 ( .A1(n9029), .A2(n7369), .ZN(n9015) );
  OAI22_X1 U11328 ( .A1(n15004), .A2(n9012), .B1(n12690), .B2(n9005), .ZN(
        n8971) );
  NAND2_X1 U11329 ( .A1(n10386), .A2(n12694), .ZN(n12490) );
  AOI21_X1 U11330 ( .B1(n8971), .B2(n12490), .A(n12446), .ZN(n8975) );
  NAND2_X1 U11331 ( .A1(n12446), .A2(n12490), .ZN(n9968) );
  NAND2_X1 U11332 ( .A1(n9012), .A2(n12694), .ZN(n8972) );
  OR2_X1 U11333 ( .A1(n9005), .A2(n8972), .ZN(n9003) );
  NAND2_X1 U11334 ( .A1(n12463), .A2(n9003), .ZN(n9028) );
  NAND2_X1 U11335 ( .A1(n9968), .A2(n9028), .ZN(n8973) );
  NAND2_X1 U11336 ( .A1(n13040), .A2(n8973), .ZN(n8974) );
  OAI21_X1 U11337 ( .B1(n13040), .B2(n8975), .A(n8974), .ZN(n8976) );
  INV_X1 U11338 ( .A(n8976), .ZN(n8977) );
  MUX2_X1 U11339 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n9027), .S(n15025), .Z(
        n8978) );
  INV_X1 U11340 ( .A(n8978), .ZN(n9008) );
  INV_X1 U11341 ( .A(n10655), .ZN(n10024) );
  NAND2_X1 U11342 ( .A1(n12333), .A2(n12338), .ZN(n8980) );
  NAND2_X1 U11343 ( .A1(n14936), .A2(n12337), .ZN(n8981) );
  INV_X1 U11344 ( .A(n14937), .ZN(n10134) );
  NAND2_X1 U11345 ( .A1(n10158), .A2(n10134), .ZN(n12343) );
  NAND2_X1 U11346 ( .A1(n10209), .A2(n12502), .ZN(n8982) );
  NAND2_X1 U11347 ( .A1(n10110), .A2(n12514), .ZN(n8984) );
  INV_X1 U11348 ( .A(n12560), .ZN(n12350) );
  NAND2_X1 U11349 ( .A1(n12350), .A2(n6914), .ZN(n8983) );
  INV_X1 U11350 ( .A(n10842), .ZN(n12503) );
  INV_X1 U11351 ( .A(n10777), .ZN(n12507) );
  NAND2_X1 U11352 ( .A1(n10954), .A2(n12505), .ZN(n8986) );
  NOR2_X1 U11353 ( .A1(n12556), .A2(n15005), .ZN(n8987) );
  NAND2_X1 U11354 ( .A1(n12556), .A2(n15005), .ZN(n8988) );
  INV_X1 U11355 ( .A(n8989), .ZN(n12383) );
  XNOR2_X1 U11356 ( .A(n12554), .B(n12379), .ZN(n12382) );
  NAND2_X1 U11357 ( .A1(n12380), .A2(n12379), .ZN(n12376) );
  INV_X1 U11358 ( .A(n11300), .ZN(n12513) );
  NAND2_X1 U11359 ( .A1(n11298), .A2(n12513), .ZN(n8990) );
  INV_X1 U11360 ( .A(n12398), .ZN(n8991) );
  INV_X1 U11361 ( .A(n12401), .ZN(n8992) );
  NAND2_X1 U11362 ( .A1(n12880), .A2(n7327), .ZN(n8993) );
  XNOR2_X1 U11363 ( .A(n13021), .B(n12884), .ZN(n12871) );
  NAND2_X1 U11364 ( .A1(n12870), .A2(n12871), .ZN(n8994) );
  NAND2_X1 U11365 ( .A1(n13021), .A2(n12406), .ZN(n12412) );
  NAND2_X1 U11366 ( .A1(n8994), .A2(n12412), .ZN(n12857) );
  NAND2_X1 U11367 ( .A1(n12857), .A2(n12863), .ZN(n8995) );
  NAND2_X1 U11368 ( .A1(n12522), .A2(n12552), .ZN(n12428) );
  AND2_X1 U11369 ( .A1(n12428), .A2(n12830), .ZN(n12420) );
  OR2_X1 U11370 ( .A1(n12522), .A2(n12552), .ZN(n12429) );
  OR2_X2 U11371 ( .A1(n12818), .A2(n12821), .ZN(n12820) );
  INV_X1 U11372 ( .A(n12937), .ZN(n12261) );
  NAND2_X1 U11373 ( .A1(n12261), .A2(n12835), .ZN(n12433) );
  INV_X1 U11374 ( .A(n12800), .ZN(n12824) );
  NAND2_X1 U11375 ( .A1(n12933), .A2(n12824), .ZN(n8996) );
  INV_X1 U11376 ( .A(n12933), .ZN(n12213) );
  NAND2_X1 U11377 ( .A1(n12213), .A2(n12800), .ZN(n8997) );
  NAND2_X1 U11378 ( .A1(n12991), .A2(n12812), .ZN(n12438) );
  INV_X1 U11379 ( .A(n12788), .ZN(n12784) );
  NAND2_X1 U11380 ( .A1(n12152), .A2(n12764), .ZN(n12319) );
  NAND2_X1 U11381 ( .A1(n12981), .A2(n12791), .ZN(n12321) );
  NAND2_X1 U11382 ( .A1(n12739), .A2(n12197), .ZN(n12721) );
  NAND2_X1 U11383 ( .A1(n8998), .A2(n12721), .ZN(n12314) );
  XOR2_X1 U11384 ( .A(n12533), .B(n12495), .Z(n9041) );
  OAI21_X1 U11385 ( .B1(n9005), .B2(n9012), .A(n12690), .ZN(n8999) );
  NAND2_X1 U11386 ( .A1(n8999), .A2(n12332), .ZN(n9001) );
  OAI21_X1 U11387 ( .B1(n12329), .B2(n9012), .A(n9005), .ZN(n9000) );
  NAND2_X1 U11388 ( .A1(n9001), .A2(n9000), .ZN(n9971) );
  INV_X1 U11389 ( .A(n12490), .ZN(n9994) );
  AND2_X1 U11390 ( .A1(n15004), .A2(n9994), .ZN(n9002) );
  NAND2_X1 U11391 ( .A1(n9971), .A2(n9002), .ZN(n9004) );
  NAND2_X1 U11392 ( .A1(n9004), .A2(n9003), .ZN(n14993) );
  NAND2_X1 U11393 ( .A1(n10386), .A2(n12690), .ZN(n14938) );
  INV_X1 U11394 ( .A(n14938), .ZN(n12540) );
  AND2_X1 U11395 ( .A1(n9005), .A2(n12540), .ZN(n15009) );
  NAND2_X1 U11396 ( .A1(n15025), .A2(n14959), .ZN(n12957) );
  INV_X1 U11397 ( .A(n9036), .ZN(n9023) );
  NAND2_X1 U11398 ( .A1(n15025), .A2(n15001), .ZN(n12961) );
  OAI22_X1 U11399 ( .A1(n9041), .A2(n12957), .B1(n9023), .B2(n12961), .ZN(
        n9006) );
  INV_X1 U11400 ( .A(n9006), .ZN(n9007) );
  NAND2_X1 U11401 ( .A1(n9008), .A2(n9007), .ZN(P3_U3488) );
  INV_X1 U11402 ( .A(n9009), .ZN(n9014) );
  OR2_X1 U11403 ( .A1(n9010), .A2(n9014), .ZN(n9992) );
  INV_X1 U11404 ( .A(n9011), .ZN(n9013) );
  NAND2_X1 U11405 ( .A1(n12332), .A2(n9012), .ZN(n12538) );
  NAND2_X1 U11406 ( .A1(n9013), .A2(n9978), .ZN(n9986) );
  INV_X1 U11407 ( .A(n9971), .ZN(n9016) );
  OAI22_X1 U11408 ( .A1(n9992), .A2(n9986), .B1(n9996), .B2(n9016), .ZN(n9017)
         );
  NAND2_X1 U11409 ( .A1(n9017), .A2(n9995), .ZN(n9021) );
  INV_X1 U11410 ( .A(n9992), .ZN(n9019) );
  NOR2_X1 U11411 ( .A1(n12463), .A2(n12490), .ZN(n9018) );
  AND2_X1 U11412 ( .A1(n9995), .A2(n9018), .ZN(n9975) );
  NAND2_X1 U11413 ( .A1(n9019), .A2(n9975), .ZN(n9020) );
  MUX2_X1 U11414 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9027), .S(n15010), .Z(
        n9022) );
  INV_X1 U11415 ( .A(n9022), .ZN(n9026) );
  INV_X1 U11416 ( .A(n14959), .ZN(n14449) );
  OAI22_X1 U11417 ( .A1(n9041), .A2(n13033), .B1(n9023), .B2(n13039), .ZN(
        n9024) );
  INV_X1 U11418 ( .A(n9024), .ZN(n9025) );
  NAND2_X1 U11419 ( .A1(n9026), .A2(n9025), .ZN(P3_U3456) );
  XNOR2_X1 U11420 ( .A(n9029), .B(n9028), .ZN(n9030) );
  NAND3_X1 U11421 ( .A1(n9031), .A2(n9968), .A3(n9030), .ZN(n9035) );
  NOR2_X1 U11422 ( .A1(n15004), .A2(n14938), .ZN(n9032) );
  INV_X2 U11423 ( .A(n14955), .ZN(n14953) );
  NAND2_X1 U11424 ( .A1(n9027), .A2(n14953), .ZN(n9044) );
  NOR2_X1 U11425 ( .A1(n12332), .A2(n14938), .ZN(n14952) );
  NOR2_X1 U11426 ( .A1(n14993), .A2(n14952), .ZN(n9033) );
  NAND2_X1 U11427 ( .A1(n15001), .A2(n14938), .ZN(n9034) );
  AOI22_X1 U11428 ( .A1(n9036), .A2(n12889), .B1(n12706), .B2(n12888), .ZN(
        n9039) );
  INV_X1 U11429 ( .A(n9042), .ZN(n9043) );
  NAND2_X1 U11430 ( .A1(n9044), .A2(n9043), .ZN(P3_U3204) );
  INV_X1 U11431 ( .A(n9333), .ZN(n9045) );
  NOR2_X1 U11432 ( .A1(n9046), .A2(n9045), .ZN(n9335) );
  INV_X1 U11435 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9050) );
  INV_X1 U11436 ( .A(n9065), .ZN(n9057) );
  INV_X1 U11437 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11438 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  NAND2_X1 U11439 ( .A1(n9065), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U11440 ( .A1(n9152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9063) );
  INV_X1 U11441 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9062) );
  XNOR2_X1 U11442 ( .A(n9063), .B(n9062), .ZN(n14383) );
  NAND2_X1 U11443 ( .A1(n9149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9064) );
  MUX2_X1 U11444 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9064), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9066) );
  NAND2_X1 U11445 ( .A1(n9066), .A2(n9065), .ZN(n9146) );
  INV_X1 U11446 ( .A(n9122), .ZN(n9118) );
  INV_X1 U11447 ( .A(n9967), .ZN(n9067) );
  AND2_X2 U11448 ( .A1(n9067), .A2(n13041), .ZN(P3_U3897) );
  AND2_X1 U11449 ( .A1(n9068), .A2(P2_U3088), .ZN(n13633) );
  OAI222_X1 U11450 ( .A1(n13636), .A2(n9069), .B1(n13637), .B2(n9516), .C1(
        P2_U3088), .C2(n9458), .ZN(P2_U3326) );
  OAI222_X1 U11451 ( .A1(n9726), .A2(P3_U3151), .B1(n13057), .B2(n9071), .C1(
        n9070), .C2(n13054), .ZN(P3_U3292) );
  OAI222_X1 U11452 ( .A1(n9791), .A2(P3_U3151), .B1(n13057), .B2(n9073), .C1(
        n9072), .C2(n13054), .ZN(P3_U3288) );
  OAI222_X1 U11453 ( .A1(n9857), .A2(P3_U3151), .B1(n13057), .B2(n9075), .C1(
        n9074), .C2(n13054), .ZN(P3_U3291) );
  OAI222_X1 U11454 ( .A1(n6500), .A2(P3_U3151), .B1(n13057), .B2(n9078), .C1(
        n9077), .C2(n13054), .ZN(P3_U3293) );
  INV_X1 U11455 ( .A(n9079), .ZN(n9080) );
  OAI222_X1 U11456 ( .A1(P3_U3151), .A2(n9906), .B1(n13054), .B2(n9081), .C1(
        n13057), .C2(n9080), .ZN(P3_U3294) );
  INV_X1 U11457 ( .A(n9082), .ZN(n9084) );
  INV_X1 U11458 ( .A(SI_6_), .ZN(n9083) );
  OAI222_X1 U11459 ( .A1(n9739), .A2(P3_U3151), .B1(n13057), .B2(n9084), .C1(
        n9083), .C2(n13054), .ZN(P3_U3289) );
  OAI222_X1 U11460 ( .A1(n9757), .A2(P3_U3151), .B1(n13057), .B2(n9086), .C1(
        n9085), .C2(n13054), .ZN(P3_U3290) );
  INV_X1 U11461 ( .A(n9907), .ZN(n9133) );
  NAND2_X1 U11462 ( .A1(n9087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9088) );
  XNOR2_X1 U11463 ( .A(n9088), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13999) );
  INV_X1 U11464 ( .A(n13999), .ZN(n9089) );
  OAI222_X1 U11465 ( .A1(n14379), .A2(n7545), .B1(n14382), .B2(n9133), .C1(
        n9089), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U11466 ( .A1(n13057), .A2(n9091), .B1(n13054), .B2(n9090), .C1(
        n11186), .C2(P3_U3151), .ZN(P3_U3285) );
  NOR2_X1 U11467 ( .A1(n9092), .A2(n6493), .ZN(n9093) );
  MUX2_X1 U11468 ( .A(n14366), .B(n9093), .S(P1_IR_REG_2__SCAN_IN), .Z(n9094)
         );
  INV_X1 U11469 ( .A(n9094), .ZN(n9095) );
  OAI222_X1 U11470 ( .A1(n13968), .A2(P1_U3086), .B1(n14382), .B2(n7524), .C1(
        n6726), .C2(n14379), .ZN(P1_U3353) );
  INV_X1 U11471 ( .A(SI_8_), .ZN(n9098) );
  INV_X1 U11472 ( .A(n9096), .ZN(n9097) );
  OAI222_X1 U11473 ( .A1(P3_U3151), .A2(n9880), .B1(n13054), .B2(n9098), .C1(
        n13057), .C2(n9097), .ZN(P3_U3287) );
  INV_X1 U11474 ( .A(n9087), .ZN(n9100) );
  NAND2_X1 U11475 ( .A1(n9100), .A2(n9099), .ZN(n9102) );
  NAND2_X1 U11476 ( .A1(n9102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U11477 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9101), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9105) );
  INV_X1 U11478 ( .A(n9102), .ZN(n9104) );
  INV_X1 U11479 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11480 ( .A1(n9104), .A2(n9103), .ZN(n9112) );
  INV_X1 U11481 ( .A(n10448), .ZN(n9106) );
  INV_X1 U11482 ( .A(n10447), .ZN(n9128) );
  OAI222_X1 U11483 ( .A1(n9106), .A2(P1_U3086), .B1(n14382), .B2(n9128), .C1(
        n6738), .C2(n14379), .ZN(P1_U3350) );
  INV_X1 U11484 ( .A(n9799), .ZN(n9126) );
  NAND2_X1 U11485 ( .A1(n9107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U11486 ( .A(n9108), .B(n9052), .ZN(n13981) );
  OAI222_X1 U11487 ( .A1(n14379), .A2(n6734), .B1(n14382), .B2(n9126), .C1(
        n13981), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U11488 ( .A(n10621), .ZN(n9130) );
  NAND2_X1 U11489 ( .A1(n9112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9109) );
  XNOR2_X1 U11490 ( .A(n9109), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10622) );
  INV_X1 U11491 ( .A(n10622), .ZN(n9110) );
  OAI222_X1 U11492 ( .A1(n14379), .A2(n9111), .B1(n14382), .B2(n9130), .C1(
        n9110), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U11493 ( .A(n10628), .ZN(n9134) );
  NAND2_X1 U11494 ( .A1(n9139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9113) );
  XNOR2_X1 U11495 ( .A(n9113), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10629) );
  INV_X1 U11496 ( .A(n14379), .ZN(n14369) );
  AOI22_X1 U11497 ( .A1(n10629), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14369), .ZN(n9114) );
  OAI21_X1 U11498 ( .B1(n9134), .B2(n14382), .A(n9114), .ZN(P1_U3348) );
  NAND2_X1 U11499 ( .A1(n11322), .A2(P1_B_REG_SCAN_IN), .ZN(n9117) );
  INV_X1 U11500 ( .A(n14383), .ZN(n9269) );
  OAI21_X1 U11501 ( .B1(n11322), .B2(P1_B_REG_SCAN_IN), .A(n9269), .ZN(n9115)
         );
  INV_X1 U11502 ( .A(n9115), .ZN(n9116) );
  OAI21_X1 U11503 ( .B1(n11506), .B2(n9117), .A(n9116), .ZN(n9569) );
  NAND2_X1 U11504 ( .A1(n9297), .A2(n9569), .ZN(n14674) );
  INV_X1 U11505 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9120) );
  NOR3_X1 U11506 ( .A1(n11506), .A2(n9118), .A3(n9269), .ZN(n9119) );
  AOI21_X1 U11507 ( .B1(n14674), .B2(n9120), .A(n9119), .ZN(P1_U3446) );
  INV_X1 U11508 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11509 ( .A1(n11322), .A2(n14383), .ZN(n9566) );
  INV_X1 U11510 ( .A(n9566), .ZN(n9121) );
  AOI22_X1 U11511 ( .A1(n14674), .A2(n9282), .B1(n9122), .B2(n9121), .ZN(
        P1_U3445) );
  INV_X1 U11512 ( .A(n9123), .ZN(n9125) );
  OAI222_X1 U11513 ( .A1(n13057), .A2(n9125), .B1(n13054), .B2(n9124), .C1(
        n12582), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U11514 ( .A(n9351), .ZN(n14761) );
  OAI222_X1 U11515 ( .A1(n13636), .A2(n9127), .B1(n13637), .B2(n9126), .C1(
        P2_U3088), .C2(n14761), .ZN(P2_U3324) );
  INV_X1 U11516 ( .A(n9374), .ZN(n9380) );
  OAI222_X1 U11517 ( .A1(n13636), .A2(n9129), .B1(n13637), .B2(n9128), .C1(
        P2_U3088), .C2(n9380), .ZN(P2_U3322) );
  INV_X1 U11518 ( .A(n9355), .ZN(n9411) );
  OAI222_X1 U11519 ( .A1(n13636), .A2(n9131), .B1(n13637), .B2(n9130), .C1(
        P2_U3088), .C2(n9411), .ZN(P2_U3321) );
  INV_X1 U11520 ( .A(n9383), .ZN(n9396) );
  OAI222_X1 U11521 ( .A1(n13636), .A2(n9132), .B1(n13637), .B2(n7524), .C1(
        P2_U3088), .C2(n9396), .ZN(P2_U3325) );
  INV_X1 U11522 ( .A(n9352), .ZN(n9564) );
  OAI222_X1 U11523 ( .A1(n13636), .A2(n15157), .B1(n13637), .B2(n9133), .C1(
        P2_U3088), .C2(n9564), .ZN(P2_U3323) );
  INV_X1 U11524 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9135) );
  INV_X1 U11525 ( .A(n9418), .ZN(n9366) );
  OAI222_X1 U11526 ( .A1(n13636), .A2(n9135), .B1(n13637), .B2(n9134), .C1(
        P2_U3088), .C2(n9366), .ZN(P2_U3320) );
  NAND2_X1 U11527 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9136) );
  MUX2_X1 U11528 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9136), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9138) );
  INV_X1 U11529 ( .A(n9092), .ZN(n9137) );
  OAI222_X1 U11530 ( .A1(n9519), .A2(P1_U3086), .B1(n14382), .B2(n9516), .C1(
        n9518), .C2(n14379), .ZN(P1_U3354) );
  INV_X1 U11531 ( .A(n10708), .ZN(n9144) );
  OAI21_X1 U11532 ( .B1(n9139), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9140) );
  MUX2_X1 U11533 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9140), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9142) );
  INV_X1 U11534 ( .A(n9287), .ZN(n9141) );
  AOI22_X1 U11535 ( .A1(n10709), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n14369), .ZN(n9143) );
  OAI21_X1 U11536 ( .B1(n9144), .B2(n14382), .A(n9143), .ZN(P1_U3347) );
  INV_X1 U11537 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9145) );
  OAI222_X1 U11538 ( .A1(n13636), .A2(n9145), .B1(n13637), .B2(n9144), .C1(
        P2_U3088), .C2(n9419), .ZN(P2_U3319) );
  INV_X1 U11539 ( .A(n9297), .ZN(n10225) );
  INV_X1 U11540 ( .A(n9146), .ZN(n9156) );
  NAND2_X1 U11541 ( .A1(n9156), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12105) );
  NAND2_X1 U11542 ( .A1(n10225), .A2(n12105), .ZN(n9161) );
  NAND2_X1 U11543 ( .A1(n9150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11544 ( .A1(n14385), .A2(n12019), .ZN(n12033) );
  INV_X1 U11545 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9153) );
  OAI21_X1 U11546 ( .B1(n12033), .B2(n9156), .A(n11685), .ZN(n9160) );
  INV_X1 U11547 ( .A(n9160), .ZN(n9157) );
  NAND2_X1 U11548 ( .A1(n9161), .A2(n9157), .ZN(n9233) );
  INV_X1 U11549 ( .A(n14378), .ZN(n11750) );
  INV_X1 U11550 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n14670) );
  INV_X1 U11551 ( .A(n9158), .ZN(n13964) );
  INV_X1 U11552 ( .A(n13964), .ZN(n14376) );
  AOI21_X1 U11553 ( .B1(n11750), .B2(n14670), .A(n14376), .ZN(n13967) );
  OAI21_X1 U11554 ( .B1(n11750), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13967), .ZN(
        n9159) );
  INV_X1 U11555 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9259) );
  XNOR2_X1 U11556 ( .A(n9159), .B(n9259), .ZN(n9163) );
  NAND2_X1 U11557 ( .A1(n9161), .A2(n9160), .ZN(n14633) );
  INV_X1 U11558 ( .A(n14633), .ZN(n10549) );
  AOI22_X1 U11559 ( .A1(n10549), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9162) );
  OAI21_X1 U11560 ( .B1(n9233), .B2(n9163), .A(n9162), .ZN(P1_U3243) );
  NOR2_X1 U11561 ( .A1(n10549), .A2(n13948), .ZN(P1_U3085) );
  INV_X1 U11562 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9164) );
  INV_X1 U11563 ( .A(n10713), .ZN(n9169) );
  INV_X1 U11564 ( .A(n9765), .ZN(n9450) );
  OAI222_X1 U11565 ( .A1(n13636), .A2(n9164), .B1(n13637), .B2(n9169), .C1(
        P2_U3088), .C2(n9450), .ZN(P2_U3318) );
  NOR2_X1 U11566 ( .A1(n9287), .A2(n14366), .ZN(n9165) );
  MUX2_X1 U11567 ( .A(n14366), .B(n9165), .S(P1_IR_REG_9__SCAN_IN), .Z(n9167)
         );
  AND2_X1 U11568 ( .A1(n9287), .A2(n9166), .ZN(n9196) );
  OR2_X1 U11569 ( .A1(n9167), .A2(n9196), .ZN(n9605) );
  OAI222_X1 U11570 ( .A1(n9605), .A2(P1_U3086), .B1(n14382), .B2(n9169), .C1(
        n9168), .C2(n14379), .ZN(P1_U3346) );
  NAND2_X1 U11571 ( .A1(n13041), .A2(n9170), .ZN(n9204) );
  AND2_X1 U11572 ( .A1(n9204), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11573 ( .A1(n9204), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11574 ( .A1(n9204), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11575 ( .A1(n9204), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11576 ( .A1(n9204), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11577 ( .A1(n9204), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11578 ( .A1(n9204), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11579 ( .A1(n9204), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11580 ( .A1(n9204), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11581 ( .A1(n9204), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11582 ( .A1(n9204), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11583 ( .A1(n9204), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11584 ( .A1(n9204), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11585 ( .A1(n9204), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11586 ( .A1(n9204), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11587 ( .A1(n9204), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11588 ( .A1(n9204), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11589 ( .A1(n9204), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11590 ( .A1(n9204), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11591 ( .A1(n9204), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11592 ( .A1(n9204), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11593 ( .A1(n9204), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11594 ( .A1(n9204), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11595 ( .A1(n9204), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11596 ( .A1(n9204), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11597 ( .A1(n9204), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11598 ( .A1(n9204), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  OAI222_X1 U11599 ( .A1(n13057), .A2(n9171), .B1(n13054), .B2(n15172), .C1(
        n12580), .C2(P3_U3151), .ZN(P3_U3281) );
  NAND2_X1 U11600 ( .A1(n10632), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10641) );
  INV_X1 U11601 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U11602 ( .A1(n10717), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10734) );
  INV_X1 U11603 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10733) );
  INV_X1 U11604 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10890) );
  INV_X1 U11605 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11149) );
  INV_X1 U11606 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11148) );
  INV_X1 U11607 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U11608 ( .A1(n11431), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11518) );
  INV_X1 U11609 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11610 ( .A1(n11518), .A2(n9172), .ZN(n9173) );
  NAND2_X1 U11611 ( .A1(n11650), .A2(n9173), .ZN(n13889) );
  INV_X1 U11612 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9176) );
  INV_X1 U11613 ( .A(n11562), .ZN(n9181) );
  NAND2_X1 U11614 ( .A1(n9178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9179) );
  INV_X1 U11615 ( .A(n9180), .ZN(n9182) );
  OR2_X1 U11616 ( .A1(n13889), .A2(n11720), .ZN(n9185) );
  AOI22_X1 U11617 ( .A1(n6491), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n11653), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n9184) );
  AND2_X2 U11618 ( .A1(n11562), .A2(n9182), .ZN(n9188) );
  NAND2_X1 U11619 ( .A1(n11039), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9183) );
  INV_X1 U11620 ( .A(n13849), .ZN(n13691) );
  NAND2_X1 U11621 ( .A1(n13691), .A2(P1_U4016), .ZN(n9186) );
  OAI21_X1 U11622 ( .B1(n13948), .B2(n9187), .A(n9186), .ZN(P1_U3578) );
  NAND2_X1 U11623 ( .A1(n11743), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U11624 ( .A1(n9188), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11625 ( .A1(n11152), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U11626 ( .A1(n11844), .A2(P1_U4016), .ZN(n9193) );
  OAI21_X1 U11627 ( .B1(n13948), .B2(n15032), .A(n9193), .ZN(P1_U3560) );
  INV_X1 U11628 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14366) );
  NOR2_X1 U11629 ( .A1(n9196), .A2(n6493), .ZN(n9194) );
  MUX2_X1 U11630 ( .A(n14366), .B(n9194), .S(P1_IR_REG_10__SCAN_IN), .Z(n9198)
         );
  INV_X1 U11631 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11632 ( .A1(n9196), .A2(n9195), .ZN(n9315) );
  INV_X1 U11633 ( .A(n9315), .ZN(n9197) );
  INV_X1 U11634 ( .A(n10877), .ZN(n9200) );
  OAI222_X1 U11635 ( .A1(n9936), .A2(P1_U3086), .B1(n14382), .B2(n9200), .C1(
        n9199), .C2(n14379), .ZN(P1_U3345) );
  INV_X1 U11636 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9201) );
  INV_X1 U11637 ( .A(n13226), .ZN(n13216) );
  OAI222_X1 U11638 ( .A1(n13636), .A2(n9201), .B1(n13637), .B2(n9200), .C1(
        P2_U3088), .C2(n13216), .ZN(P2_U3317) );
  INV_X1 U11639 ( .A(n11033), .ZN(n9206) );
  NAND2_X1 U11640 ( .A1(n9315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11641 ( .A(n9202), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U11642 ( .A1(n11034), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n14369), .ZN(n9203) );
  OAI21_X1 U11643 ( .B1(n9206), .B2(n14382), .A(n9203), .ZN(P1_U3344) );
  INV_X1 U11644 ( .A(n9204), .ZN(n9205) );
  INV_X1 U11645 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15053) );
  NOR2_X1 U11646 ( .A1(n9205), .A2(n15053), .ZN(P3_U3243) );
  INV_X1 U11647 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15071) );
  NOR2_X1 U11648 ( .A1(n9205), .A2(n15071), .ZN(P3_U3250) );
  INV_X1 U11649 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15162) );
  NOR2_X1 U11650 ( .A1(n9205), .A2(n15162), .ZN(P3_U3260) );
  INV_X1 U11651 ( .A(n13234), .ZN(n13243) );
  OAI222_X1 U11652 ( .A1(n13636), .A2(n9207), .B1(n13637), .B2(n9206), .C1(
        P2_U3088), .C2(n13243), .ZN(P2_U3316) );
  INV_X1 U11653 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n15056) );
  NAND2_X1 U11654 ( .A1(n10830), .A2(P3_U3897), .ZN(n9208) );
  OAI21_X1 U11655 ( .B1(P3_U3897), .B2(n15056), .A(n9208), .ZN(P3_U3491) );
  INV_X1 U11656 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U11657 ( .A1(n10150), .A2(P3_U3897), .ZN(n9209) );
  OAI21_X1 U11658 ( .B1(P3_U3897), .B2(n15194), .A(n9209), .ZN(P3_U3496) );
  INV_X1 U11659 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15183) );
  NAND2_X1 U11660 ( .A1(n12897), .A2(P3_U3897), .ZN(n9210) );
  OAI21_X1 U11661 ( .B1(P3_U3897), .B2(n15183), .A(n9210), .ZN(P3_U3506) );
  INV_X1 U11662 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9211) );
  INV_X1 U11663 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9212) );
  MUX2_X1 U11664 ( .A(n9212), .B(P1_REG2_REG_1__SCAN_IN), .S(n9519), .Z(n13958) );
  AND2_X1 U11665 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13963) );
  NAND2_X1 U11666 ( .A1(n13958), .A2(n13963), .ZN(n13957) );
  INV_X1 U11667 ( .A(n9519), .ZN(n13953) );
  NAND2_X1 U11668 ( .A1(n13953), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U11669 ( .A1(n13957), .A2(n9213), .ZN(n13973) );
  NAND2_X1 U11670 ( .A1(n13974), .A2(n13973), .ZN(n13972) );
  OR2_X1 U11671 ( .A1(n13968), .A2(n9211), .ZN(n9214) );
  NAND2_X1 U11672 ( .A1(n13972), .A2(n9214), .ZN(n13987) );
  XNOR2_X1 U11673 ( .A(n13981), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n13988) );
  NAND2_X1 U11674 ( .A1(n13987), .A2(n13988), .ZN(n13986) );
  INV_X1 U11675 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10237) );
  OR2_X1 U11676 ( .A1(n13981), .A2(n10237), .ZN(n9215) );
  NAND2_X1 U11677 ( .A1(n13986), .A2(n9215), .ZN(n14006) );
  INV_X1 U11678 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9216) );
  XNOR2_X1 U11679 ( .A(n13999), .B(n9216), .ZN(n14007) );
  INV_X1 U11680 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9217) );
  MUX2_X1 U11681 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9217), .S(n10448), .Z(n9218) );
  INV_X1 U11682 ( .A(n9218), .ZN(n9308) );
  NOR2_X1 U11683 ( .A1(n9309), .A2(n9308), .ZN(n9307) );
  XNOR2_X1 U11684 ( .A(n10622), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9242) );
  NOR2_X1 U11685 ( .A1(n9243), .A2(n9242), .ZN(n9241) );
  INV_X1 U11686 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9219) );
  MUX2_X1 U11687 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9219), .S(n10629), .Z(n9220) );
  INV_X1 U11688 ( .A(n9220), .ZN(n9222) );
  OR2_X1 U11689 ( .A1(n14376), .A2(n14378), .ZN(n9221) );
  OR2_X1 U11690 ( .A1(n9233), .A2(n9221), .ZN(n14566) );
  NOR2_X1 U11691 ( .A1(n9223), .A2(n9222), .ZN(n9325) );
  AOI211_X1 U11692 ( .C1(n9223), .C2(n9222), .A(n14566), .B(n9325), .ZN(n9240)
         );
  INV_X1 U11693 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9596) );
  MUX2_X1 U11694 ( .A(n9596), .B(P1_REG1_REG_2__SCAN_IN), .S(n13968), .Z(
        n13977) );
  INV_X1 U11695 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14744) );
  MUX2_X1 U11696 ( .A(n14744), .B(P1_REG1_REG_1__SCAN_IN), .S(n9519), .Z(
        n13956) );
  AND2_X1 U11697 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13955) );
  NAND2_X1 U11698 ( .A1(n13956), .A2(n13955), .ZN(n13954) );
  NAND2_X1 U11699 ( .A1(n13953), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11700 ( .A1(n13954), .A2(n9224), .ZN(n13976) );
  NAND2_X1 U11701 ( .A1(n13977), .A2(n13976), .ZN(n13975) );
  OR2_X1 U11702 ( .A1(n13968), .A2(n9596), .ZN(n9225) );
  NAND2_X1 U11703 ( .A1(n13975), .A2(n9225), .ZN(n13990) );
  XNOR2_X1 U11704 ( .A(n13981), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n13991) );
  NAND2_X1 U11705 ( .A1(n13990), .A2(n13991), .ZN(n13989) );
  INV_X1 U11706 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9226) );
  OR2_X1 U11707 ( .A1(n13981), .A2(n9226), .ZN(n9227) );
  NAND2_X1 U11708 ( .A1(n13989), .A2(n9227), .ZN(n14002) );
  INV_X1 U11709 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9228) );
  XNOR2_X1 U11710 ( .A(n13999), .B(n9228), .ZN(n14003) );
  AND2_X1 U11711 ( .A1(n14002), .A2(n14003), .ZN(n14000) );
  AOI21_X1 U11712 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n13999), .A(n14000), .ZN(
        n9304) );
  INV_X1 U11713 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9916) );
  MUX2_X1 U11714 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9916), .S(n10448), .Z(n9303) );
  NAND2_X1 U11715 ( .A1(n9304), .A2(n9303), .ZN(n9302) );
  OAI21_X1 U11716 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10448), .A(n9302), .ZN(
        n9245) );
  INV_X1 U11717 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9229) );
  MUX2_X1 U11718 ( .A(n9229), .B(P1_REG1_REG_6__SCAN_IN), .S(n10622), .Z(n9246) );
  NOR2_X1 U11719 ( .A1(n9245), .A2(n9246), .ZN(n9244) );
  AOI21_X1 U11720 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10622), .A(n9244), .ZN(
        n9232) );
  INV_X1 U11721 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9230) );
  MUX2_X1 U11722 ( .A(n9230), .B(P1_REG1_REG_7__SCAN_IN), .S(n10629), .Z(n9231) );
  OR2_X1 U11723 ( .A1(n9233), .A2(n11750), .ZN(n14548) );
  NOR2_X1 U11724 ( .A1(n9232), .A2(n9231), .ZN(n9318) );
  AOI211_X1 U11725 ( .C1(n9232), .C2(n9231), .A(n14548), .B(n9318), .ZN(n9239)
         );
  INV_X1 U11726 ( .A(n9233), .ZN(n9234) );
  AND2_X1 U11727 ( .A1(n9234), .A2(n14376), .ZN(n14625) );
  NAND2_X1 U11728 ( .A1(n14625), .A2(n10629), .ZN(n9236) );
  NAND2_X1 U11729 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9235) );
  OAI211_X1 U11730 ( .C1(n9237), .C2(n14633), .A(n9236), .B(n9235), .ZN(n9238)
         );
  OR3_X1 U11731 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(P1_U3250) );
  AOI211_X1 U11732 ( .C1(n9243), .C2(n9242), .A(n14566), .B(n9241), .ZN(n9252)
         );
  AOI211_X1 U11733 ( .C1(n9246), .C2(n9245), .A(n14548), .B(n9244), .ZN(n9251)
         );
  NAND2_X1 U11734 ( .A1(n14625), .A2(n10622), .ZN(n9248) );
  NAND2_X1 U11735 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9247) );
  OAI211_X1 U11736 ( .C1(n9249), .C2(n14633), .A(n9248), .B(n9247), .ZN(n9250)
         );
  OR3_X1 U11737 ( .A1(n9252), .A2(n9251), .A3(n9250), .ZN(P1_U3249) );
  NAND2_X1 U11738 ( .A1(n9253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9254) );
  XNOR2_X1 U11739 ( .A(n9254), .B(P1_IR_REG_20__SCAN_IN), .ZN(n12036) );
  INV_X4 U11740 ( .A(n13682), .ZN(n13800) );
  NAND2_X2 U11741 ( .A1(n14658), .A2(n12030), .ZN(n14683) );
  AND2_X2 U11742 ( .A1(n13800), .A2(n14683), .ZN(n10452) );
  INV_X1 U11743 ( .A(SI_0_), .ZN(n9256) );
  OAI21_X1 U11744 ( .B1(n9517), .B2(n9256), .A(n9255), .ZN(n9257) );
  NAND2_X1 U11745 ( .A1(n9258), .A2(n9257), .ZN(n14386) );
  MUX2_X1 U11746 ( .A(n9259), .B(n14386), .S(n11685), .Z(n14660) );
  OAI22_X1 U11748 ( .A1(n14660), .A2(n13690), .B1(n9822), .B2(n9259), .ZN(
        n9260) );
  INV_X1 U11749 ( .A(n9260), .ZN(n9261) );
  AND2_X1 U11750 ( .A1(n9262), .A2(n9261), .ZN(n9267) );
  NAND2_X1 U11751 ( .A1(n11844), .A2(n9526), .ZN(n9266) );
  INV_X1 U11752 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9263) );
  OAI22_X1 U11753 ( .A1(n14660), .A2(n13682), .B1(n9822), .B2(n9263), .ZN(
        n9264) );
  INV_X1 U11754 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U11755 ( .A1(n9266), .A2(n9265), .ZN(n9512) );
  NAND2_X1 U11756 ( .A1(n9267), .A2(n9512), .ZN(n9514) );
  OAI21_X1 U11757 ( .B1(n9267), .B2(n9512), .A(n9514), .ZN(n9268) );
  INV_X1 U11758 ( .A(n9268), .ZN(n13962) );
  OR2_X1 U11759 ( .A1(n9569), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9271) );
  OR2_X1 U11760 ( .A1(n11506), .A2(n9269), .ZN(n9270) );
  NAND2_X1 U11761 ( .A1(n9271), .A2(n9270), .ZN(n10222) );
  INV_X1 U11762 ( .A(n10222), .ZN(n9285) );
  NOR4_X1 U11763 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9275) );
  NOR4_X1 U11764 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9274) );
  NOR4_X1 U11765 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9273) );
  NOR4_X1 U11766 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9272) );
  AND4_X1 U11767 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n9281)
         );
  NOR2_X1 U11768 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .ZN(
        n9279) );
  NOR4_X1 U11769 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9278) );
  NOR4_X1 U11770 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9277) );
  NOR4_X1 U11771 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9276) );
  AND4_X1 U11772 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n9280)
         );
  NAND2_X1 U11773 ( .A1(n9281), .A2(n9280), .ZN(n9567) );
  NOR2_X1 U11774 ( .A1(n9567), .A2(n9282), .ZN(n9283) );
  OR2_X1 U11775 ( .A1(n9569), .A2(n9283), .ZN(n9284) );
  AND2_X1 U11776 ( .A1(n9284), .A2(n9566), .ZN(n9592) );
  NAND2_X1 U11777 ( .A1(n9285), .A2(n9592), .ZN(n9298) );
  INV_X1 U11778 ( .A(n9298), .ZN(n9291) );
  XNOR2_X2 U11779 ( .A(n9289), .B(P1_IR_REG_19__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U11780 ( .A1(n14044), .A2(n12030), .ZN(n9296) );
  AND2_X2 U11781 ( .A1(n9296), .A2(n14658), .ZN(n14691) );
  AND3_X1 U11782 ( .A1(n9297), .A2(n14698), .A3(n12033), .ZN(n9290) );
  NAND2_X1 U11783 ( .A1(n9291), .A2(n9290), .ZN(n14475) );
  OR2_X1 U11784 ( .A1(n14683), .A2(n14044), .ZN(n10226) );
  NAND2_X1 U11785 ( .A1(n9298), .A2(n10226), .ZN(n9824) );
  AND2_X1 U11786 ( .A1(n9824), .A2(n9297), .ZN(n14480) );
  INV_X1 U11787 ( .A(n14660), .ZN(n9573) );
  INV_X1 U11788 ( .A(n12033), .ZN(n9542) );
  NAND2_X1 U11789 ( .A1(n6678), .A2(n13898), .ZN(n14663) );
  NAND2_X1 U11790 ( .A1(n9296), .A2(n9542), .ZN(n9823) );
  NAND2_X1 U11791 ( .A1(n9297), .A2(n9823), .ZN(n12102) );
  INV_X1 U11792 ( .A(n12102), .ZN(n9565) );
  NAND2_X1 U11793 ( .A1(n9824), .A2(n9565), .ZN(n11831) );
  NAND2_X1 U11794 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n11831), .ZN(n9299) );
  OAI21_X1 U11795 ( .B1(n14663), .B2(n14481), .A(n9299), .ZN(n9300) );
  AOI21_X1 U11796 ( .B1(n14502), .B2(n9573), .A(n9300), .ZN(n9301) );
  OAI21_X1 U11797 ( .B1(n13962), .B2(n14475), .A(n9301), .ZN(P1_U3232) );
  OAI21_X1 U11798 ( .B1(n9304), .B2(n9303), .A(n9302), .ZN(n9312) );
  NAND2_X1 U11799 ( .A1(n14625), .A2(n10448), .ZN(n9305) );
  NAND2_X1 U11800 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10465) );
  OAI211_X1 U11801 ( .C1(n9306), .C2(n14633), .A(n9305), .B(n10465), .ZN(n9311) );
  AOI211_X1 U11802 ( .C1(n9309), .C2(n9308), .A(n9307), .B(n14566), .ZN(n9310)
         );
  AOI211_X1 U11803 ( .C1(n14617), .C2(n9312), .A(n9311), .B(n9310), .ZN(n9313)
         );
  INV_X1 U11804 ( .A(n9313), .ZN(P1_U3248) );
  INV_X1 U11805 ( .A(n11114), .ZN(n9317) );
  INV_X1 U11806 ( .A(n13270), .ZN(n13254) );
  OAI222_X1 U11807 ( .A1(n13636), .A2(n9314), .B1(n13637), .B2(n9317), .C1(
        n13254), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U11808 ( .A1(n9961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9431) );
  XNOR2_X1 U11809 ( .A(n9431), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14025) );
  INV_X1 U11810 ( .A(n14025), .ZN(n10551) );
  OAI222_X1 U11811 ( .A1(P1_U3086), .A2(n10551), .B1(n14382), .B2(n9317), .C1(
        n9316), .C2(n14379), .ZN(P1_U3343) );
  AOI21_X1 U11812 ( .B1(n10629), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9318), .ZN(
        n9321) );
  INV_X1 U11813 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9319) );
  MUX2_X1 U11814 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9319), .S(n10709), .Z(n9320) );
  NAND2_X1 U11815 ( .A1(n9321), .A2(n9320), .ZN(n9598) );
  OAI21_X1 U11816 ( .B1(n9321), .B2(n9320), .A(n9598), .ZN(n9330) );
  NAND2_X1 U11817 ( .A1(n14625), .A2(n10709), .ZN(n9323) );
  NAND2_X1 U11818 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9322) );
  OAI211_X1 U11819 ( .C1(n9324), .C2(n14633), .A(n9323), .B(n9322), .ZN(n9329)
         );
  XNOR2_X1 U11820 ( .A(n10709), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9326) );
  NOR2_X1 U11821 ( .A1(n9327), .A2(n9326), .ZN(n9604) );
  AOI211_X1 U11822 ( .C1(n9327), .C2(n9326), .A(n14566), .B(n9604), .ZN(n9328)
         );
  AOI211_X1 U11823 ( .C1(n14617), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9331)
         );
  INV_X1 U11824 ( .A(n9331), .ZN(P1_U3251) );
  AOI21_X1 U11825 ( .B1(n10063), .B2(n9333), .A(n9332), .ZN(n9334) );
  AND2_X1 U11826 ( .A1(n9494), .A2(n9344), .ZN(n14809) );
  INV_X1 U11827 ( .A(n15226), .ZN(n14824) );
  NOR2_X2 U11828 ( .A1(n9344), .A2(P2_U3088), .ZN(n15233) );
  AND2_X1 U11829 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10262) );
  INV_X1 U11830 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9336) );
  MUX2_X1 U11831 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9336), .S(n9383), .Z(n9339)
         );
  INV_X1 U11832 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9621) );
  MUX2_X1 U11833 ( .A(n9621), .B(P2_REG1_REG_1__SCAN_IN), .S(n9458), .Z(n9338)
         );
  AND2_X1 U11834 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9337) );
  NAND2_X1 U11835 ( .A1(n9338), .A2(n9337), .ZN(n9462) );
  OAI21_X1 U11836 ( .B1(n9621), .B2(n9458), .A(n9462), .ZN(n9382) );
  INV_X1 U11837 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n14889) );
  MUX2_X1 U11838 ( .A(n14889), .B(P2_REG1_REG_3__SCAN_IN), .S(n9351), .Z(
        n14764) );
  AOI21_X1 U11839 ( .B1(n9351), .B2(P2_REG1_REG_3__SCAN_IN), .A(n14763), .ZN(
        n9553) );
  INV_X1 U11840 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9340) );
  MUX2_X1 U11841 ( .A(n9340), .B(P2_REG1_REG_4__SCAN_IN), .S(n9352), .Z(n9552)
         );
  NOR2_X1 U11842 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  INV_X1 U11843 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14891) );
  MUX2_X1 U11844 ( .A(n14891), .B(P2_REG1_REG_5__SCAN_IN), .S(n9374), .Z(n9368) );
  NOR2_X1 U11845 ( .A1(n9369), .A2(n9368), .ZN(n9367) );
  AOI21_X1 U11846 ( .B1(n9374), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9367), .ZN(
        n9405) );
  INV_X1 U11847 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10575) );
  MUX2_X1 U11848 ( .A(n10575), .B(P2_REG1_REG_6__SCAN_IN), .S(n9355), .Z(n9404) );
  NOR2_X1 U11849 ( .A1(n9405), .A2(n9404), .ZN(n9403) );
  NOR2_X1 U11850 ( .A1(n9411), .A2(n10575), .ZN(n9343) );
  INV_X1 U11851 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11852 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9341), .S(n9418), .Z(n9342)
         );
  INV_X1 U11853 ( .A(n9414), .ZN(n9346) );
  NOR3_X1 U11854 ( .A1(n9403), .A2(n9343), .A3(n9342), .ZN(n9345) );
  NOR2_X1 U11855 ( .A1(n9494), .A2(P2_U3088), .ZN(n13632) );
  NAND2_X1 U11856 ( .A1(n9361), .A2(n6719), .ZN(n14780) );
  NOR3_X1 U11857 ( .A1(n9346), .A2(n9345), .A3(n14780), .ZN(n9347) );
  AOI211_X1 U11858 ( .C1(n15233), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10262), .B(
        n9347), .ZN(n9365) );
  INV_X1 U11859 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9348) );
  MUX2_X1 U11860 ( .A(n9348), .B(P2_REG2_REG_1__SCAN_IN), .S(n9458), .Z(n9456)
         );
  NAND3_X1 U11861 ( .A1(n9456), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n9457) );
  OR2_X1 U11862 ( .A1(n9458), .A2(n9348), .ZN(n9390) );
  INV_X1 U11863 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9349) );
  MUX2_X1 U11864 ( .A(n9349), .B(P2_REG2_REG_2__SCAN_IN), .S(n9383), .Z(n9391)
         );
  AOI21_X1 U11865 ( .B1(n9457), .B2(n9390), .A(n9391), .ZN(n9389) );
  AOI21_X1 U11866 ( .B1(n9383), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9389), .ZN(
        n14769) );
  INV_X1 U11867 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9350) );
  MUX2_X1 U11868 ( .A(n9350), .B(P2_REG2_REG_3__SCAN_IN), .S(n9351), .Z(n14768) );
  NOR2_X1 U11869 ( .A1(n14769), .A2(n14768), .ZN(n14767) );
  AOI21_X1 U11870 ( .B1(n9351), .B2(P2_REG2_REG_3__SCAN_IN), .A(n14767), .ZN(
        n9557) );
  INV_X1 U11871 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9353) );
  MUX2_X1 U11872 ( .A(n9353), .B(P2_REG2_REG_4__SCAN_IN), .S(n9352), .Z(n9556)
         );
  NOR2_X1 U11873 ( .A1(n9557), .A2(n9556), .ZN(n9555) );
  NOR2_X1 U11874 ( .A1(n9564), .A2(n9353), .ZN(n9373) );
  INV_X1 U11875 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10278) );
  MUX2_X1 U11876 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10278), .S(n9374), .Z(n9354) );
  OAI21_X1 U11877 ( .B1(n9555), .B2(n9373), .A(n9354), .ZN(n9400) );
  NAND2_X1 U11878 ( .A1(n9374), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9399) );
  INV_X1 U11879 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9356) );
  MUX2_X1 U11880 ( .A(n9356), .B(P2_REG2_REG_6__SCAN_IN), .S(n9355), .Z(n9398)
         );
  AOI21_X1 U11881 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9397) );
  INV_X1 U11882 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n15159) );
  MUX2_X1 U11883 ( .A(n15159), .B(P2_REG2_REG_7__SCAN_IN), .S(n9418), .Z(n9358) );
  NOR2_X1 U11884 ( .A1(n9411), .A2(n9356), .ZN(n9360) );
  INV_X1 U11885 ( .A(n9360), .ZN(n9357) );
  NAND2_X1 U11886 ( .A1(n9358), .A2(n9357), .ZN(n9363) );
  MUX2_X1 U11887 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n15159), .S(n9418), .Z(n9359) );
  OAI21_X1 U11888 ( .B1(n9397), .B2(n9360), .A(n9359), .ZN(n9423) );
  INV_X1 U11889 ( .A(n9361), .ZN(n9362) );
  NOR2_X2 U11890 ( .A1(n9362), .A2(n6719), .ZN(n14833) );
  OAI211_X1 U11891 ( .C1(n9397), .C2(n9363), .A(n9423), .B(n14833), .ZN(n9364)
         );
  OAI211_X1 U11892 ( .C1(n14824), .C2(n9366), .A(n9365), .B(n9364), .ZN(
        P2_U3221) );
  NAND2_X1 U11893 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10105) );
  AOI211_X1 U11894 ( .C1(n9369), .C2(n9368), .A(n9367), .B(n14780), .ZN(n9370)
         );
  INV_X1 U11895 ( .A(n9370), .ZN(n9371) );
  NAND2_X1 U11896 ( .A1(n10105), .A2(n9371), .ZN(n9372) );
  AOI21_X1 U11897 ( .B1(n15233), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9372), .ZN(
        n9379) );
  INV_X1 U11898 ( .A(n9373), .ZN(n9376) );
  MUX2_X1 U11899 ( .A(n10278), .B(P2_REG2_REG_5__SCAN_IN), .S(n9374), .Z(n9375) );
  NAND2_X1 U11900 ( .A1(n9376), .A2(n9375), .ZN(n9377) );
  OAI211_X1 U11901 ( .C1(n9555), .C2(n9377), .A(n14833), .B(n9400), .ZN(n9378)
         );
  OAI211_X1 U11902 ( .C1(n14824), .C2(n9380), .A(n9379), .B(n9378), .ZN(
        P2_U3219) );
  INV_X1 U11903 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9381) );
  NOR2_X1 U11904 ( .A1(n9381), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9388) );
  INV_X1 U11905 ( .A(n9382), .ZN(n9386) );
  MUX2_X1 U11906 ( .A(n9336), .B(P2_REG1_REG_2__SCAN_IN), .S(n9383), .Z(n9385)
         );
  AOI211_X1 U11907 ( .C1(n9386), .C2(n9385), .A(n9384), .B(n14780), .ZN(n9387)
         );
  AOI211_X1 U11908 ( .C1(n15233), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9388), .B(
        n9387), .ZN(n9395) );
  INV_X1 U11909 ( .A(n9389), .ZN(n9393) );
  NAND3_X1 U11910 ( .A1(n9391), .A2(n9457), .A3(n9390), .ZN(n9392) );
  NAND3_X1 U11911 ( .A1(n14833), .A2(n9393), .A3(n9392), .ZN(n9394) );
  OAI211_X1 U11912 ( .C1(n14824), .C2(n9396), .A(n9395), .B(n9394), .ZN(
        P2_U3216) );
  INV_X1 U11913 ( .A(n9397), .ZN(n9402) );
  NAND3_X1 U11914 ( .A1(n9400), .A2(n9399), .A3(n9398), .ZN(n9401) );
  NAND3_X1 U11915 ( .A1(n9402), .A2(n14833), .A3(n9401), .ZN(n9410) );
  NAND2_X1 U11916 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10391) );
  AOI211_X1 U11917 ( .C1(n9405), .C2(n9404), .A(n9403), .B(n14780), .ZN(n9406)
         );
  INV_X1 U11918 ( .A(n9406), .ZN(n9407) );
  NAND2_X1 U11919 ( .A1(n10391), .A2(n9407), .ZN(n9408) );
  AOI21_X1 U11920 ( .B1(n15233), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9408), .ZN(
        n9409) );
  OAI211_X1 U11921 ( .C1(n14824), .C2(n9411), .A(n9410), .B(n9409), .ZN(
        P2_U3220) );
  NAND2_X1 U11922 ( .A1(n9418), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9413) );
  INV_X1 U11923 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10615) );
  MUX2_X1 U11924 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10615), .S(n9419), .Z(n9412) );
  AOI21_X1 U11925 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(n9439) );
  NAND3_X1 U11926 ( .A1(n9414), .A2(n9413), .A3(n9412), .ZN(n9415) );
  INV_X1 U11927 ( .A(n14780), .ZN(n15223) );
  NAND2_X1 U11928 ( .A1(n9415), .A2(n15223), .ZN(n9428) );
  INV_X1 U11929 ( .A(n15233), .ZN(n14774) );
  INV_X1 U11930 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11931 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10679) );
  OAI21_X1 U11932 ( .B1(n14774), .B2(n9416), .A(n10679), .ZN(n9417) );
  AOI21_X1 U11933 ( .B1(n9444), .B2(n15226), .A(n9417), .ZN(n9427) );
  NAND2_X1 U11934 ( .A1(n9418), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9422) );
  INV_X1 U11935 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9420) );
  MUX2_X1 U11936 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9420), .S(n9419), .Z(n9421)
         );
  AOI21_X1 U11937 ( .B1(n9423), .B2(n9422), .A(n9421), .ZN(n9443) );
  INV_X1 U11938 ( .A(n9443), .ZN(n9425) );
  NAND3_X1 U11939 ( .A1(n9423), .A2(n9422), .A3(n9421), .ZN(n9424) );
  NAND3_X1 U11940 ( .A1(n9425), .A2(n14833), .A3(n9424), .ZN(n9426) );
  OAI211_X1 U11941 ( .C1(n9439), .C2(n9428), .A(n9427), .B(n9426), .ZN(
        P2_U3222) );
  INV_X1 U11942 ( .A(n11145), .ZN(n9437) );
  INV_X1 U11943 ( .A(n14778), .ZN(n13257) );
  OAI222_X1 U11944 ( .A1(n13636), .A2(n9429), .B1(n13637), .B2(n9437), .C1(
        n13257), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U11945 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U11946 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  NAND2_X1 U11947 ( .A1(n9432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9434) );
  INV_X1 U11948 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11949 ( .A1(n9434), .A2(n9433), .ZN(n9614) );
  OR2_X1 U11950 ( .A1(n9434), .A2(n9433), .ZN(n9435) );
  INV_X1 U11951 ( .A(n14557), .ZN(n9438) );
  OAI222_X1 U11952 ( .A1(P1_U3086), .A2(n9438), .B1(n14382), .B2(n9437), .C1(
        n9436), .C2(n14379), .ZN(P1_U3342) );
  INV_X1 U11953 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10934) );
  MUX2_X1 U11954 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10934), .S(n9765), .Z(n9440) );
  NAND2_X1 U11955 ( .A1(n9441), .A2(n9440), .ZN(n9761) );
  OAI21_X1 U11956 ( .B1(n9441), .B2(n9440), .A(n9761), .ZN(n9442) );
  NAND2_X1 U11957 ( .A1(n9442), .A2(n15223), .ZN(n9454) );
  AOI21_X1 U11958 ( .B1(n9444), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9443), .ZN(
        n9447) );
  INV_X1 U11959 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U11960 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9445), .S(n9765), .Z(n9446)
         );
  NAND2_X1 U11961 ( .A1(n9447), .A2(n9446), .ZN(n9764) );
  OAI21_X1 U11962 ( .B1(n9447), .B2(n9446), .A(n9764), .ZN(n9452) );
  NAND2_X1 U11963 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n9449) );
  NAND2_X1 U11964 ( .A1(n15233), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9448) );
  OAI211_X1 U11965 ( .C1(n14824), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9451)
         );
  AOI21_X1 U11966 ( .B1(n9452), .B2(n14833), .A(n9451), .ZN(n9453) );
  NAND2_X1 U11967 ( .A1(n9454), .A2(n9453), .ZN(P2_U3223) );
  INV_X1 U11968 ( .A(n14833), .ZN(n15230) );
  INV_X1 U11969 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9455) );
  NOR2_X1 U11970 ( .A1(n15230), .A2(n9455), .ZN(n14754) );
  AOI22_X1 U11971 ( .A1(n14754), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14833), .B2(
        n9456), .ZN(n9469) );
  INV_X1 U11972 ( .A(n9457), .ZN(n9468) );
  INV_X1 U11973 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14887) );
  MUX2_X1 U11974 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9621), .S(n9458), .Z(n9459)
         );
  OAI21_X1 U11975 ( .B1(n14887), .B2(n9460), .A(n9459), .ZN(n9461) );
  NAND3_X1 U11976 ( .A1(n15223), .A2(n9462), .A3(n9461), .ZN(n9464) );
  AOI22_X1 U11977 ( .A1(n15233), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n9463) );
  NAND2_X1 U11978 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  AOI21_X1 U11979 ( .B1(n9466), .B2(n15226), .A(n9465), .ZN(n9467) );
  OAI21_X1 U11980 ( .B1(n9469), .B2(n9468), .A(n9467), .ZN(P2_U3215) );
  XNOR2_X1 U11981 ( .A(n11324), .B(P2_B_REG_SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11982 ( .A1(n9470), .A2(n11505), .ZN(n9471) );
  INV_X1 U11983 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14846) );
  AND2_X1 U11984 ( .A1(n13638), .A2(n11505), .ZN(n9473) );
  AOI21_X1 U11985 ( .B1(n14838), .B2(n14846), .A(n9473), .ZN(n10062) );
  INV_X1 U11986 ( .A(n10062), .ZN(n9474) );
  AND2_X1 U11987 ( .A1(n9474), .A2(n14843), .ZN(n14844) );
  NOR2_X1 U11988 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n9478) );
  NOR4_X1 U11989 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n9477) );
  NOR4_X1 U11990 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9476) );
  NOR4_X1 U11991 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9475) );
  NAND4_X1 U11992 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(n9484)
         );
  NOR4_X1 U11993 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9482) );
  NOR4_X1 U11994 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9481) );
  NOR4_X1 U11995 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9480) );
  NOR4_X1 U11996 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9479) );
  NAND4_X1 U11997 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9483)
         );
  OAI21_X1 U11998 ( .B1(n9484), .B2(n9483), .A(n14838), .ZN(n10061) );
  NAND2_X1 U11999 ( .A1(n10924), .A2(n8263), .ZN(n14848) );
  NAND2_X1 U12000 ( .A1(n10055), .A2(n11500), .ZN(n10077) );
  NAND2_X1 U12001 ( .A1(n10063), .A2(n10075), .ZN(n10180) );
  AND3_X1 U12002 ( .A1(n10061), .A2(n10077), .A3(n10180), .ZN(n9485) );
  INV_X1 U12003 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14841) );
  NAND2_X1 U12004 ( .A1(n14838), .A2(n14841), .ZN(n9487) );
  NAND2_X1 U12005 ( .A1(n13638), .A2(n11324), .ZN(n9486) );
  NAND2_X1 U12006 ( .A1(n9487), .A2(n9486), .ZN(n14842) );
  INV_X1 U12007 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9509) );
  INV_X1 U12008 ( .A(n9495), .ZN(n9489) );
  NAND2_X1 U12009 ( .A1(n9489), .A2(n9488), .ZN(n9624) );
  NAND2_X1 U12010 ( .A1(n9495), .A2(n10044), .ZN(n9490) );
  AND2_X1 U12011 ( .A1(n9624), .A2(n9490), .ZN(n10185) );
  INV_X1 U12012 ( .A(n14855), .ZN(n14871) );
  NAND2_X1 U12013 ( .A1(n9495), .A2(n9496), .ZN(n9628) );
  OAI21_X1 U12014 ( .B1(n9496), .B2(n9495), .A(n9628), .ZN(n9500) );
  NAND2_X1 U12015 ( .A1(n9497), .A2(n10072), .ZN(n9498) );
  NAND2_X1 U12016 ( .A1(n9499), .A2(n9498), .ZN(n13488) );
  NAND2_X1 U12017 ( .A1(n9500), .A2(n13488), .ZN(n9501) );
  OAI211_X1 U12018 ( .C1(n10185), .C2(n14849), .A(n9502), .B(n9501), .ZN(
        n10186) );
  INV_X1 U12019 ( .A(n10186), .ZN(n9507) );
  INV_X1 U12020 ( .A(n10075), .ZN(n9503) );
  OR2_X1 U12021 ( .A1(n14848), .A2(n9503), .ZN(n14859) );
  NAND2_X1 U12022 ( .A1(n9504), .A2(n14847), .ZN(n9632) );
  NAND2_X1 U12023 ( .A1(n10377), .A2(n13081), .ZN(n9505) );
  AND3_X1 U12024 ( .A1(n10055), .A2(n9632), .A3(n9505), .ZN(n10191) );
  AOI21_X1 U12025 ( .B1(n14877), .B2(n13081), .A(n10191), .ZN(n9506) );
  OAI211_X1 U12026 ( .C1(n10185), .C2(n14871), .A(n9507), .B(n9506), .ZN(n9619) );
  NAND2_X1 U12027 ( .A1(n14886), .A2(n9619), .ZN(n9508) );
  OAI21_X1 U12028 ( .B1(n14886), .B2(n9509), .A(n9508), .ZN(P2_U3433) );
  OR2_X1 U12029 ( .A1(n12031), .A2(n11835), .ZN(n9511) );
  NAND2_X2 U12030 ( .A1(n9511), .A2(n9510), .ZN(n13798) );
  OR2_X1 U12031 ( .A1(n9512), .A2(n13752), .ZN(n9513) );
  NAND2_X1 U12032 ( .A1(n6678), .A2(n9526), .ZN(n9524) );
  OR2_X1 U12033 ( .A1(n12011), .A2(n9516), .ZN(n9522) );
  OR2_X1 U12034 ( .A1(n11685), .A2(n9519), .ZN(n9520) );
  OR2_X1 U12035 ( .A1(n11544), .A2(n13682), .ZN(n9523) );
  NAND2_X1 U12036 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  XNOR2_X1 U12037 ( .A(n9525), .B(n13752), .ZN(n9529) );
  NAND2_X1 U12038 ( .A1(n6678), .A2(n10452), .ZN(n9528) );
  NAND2_X1 U12039 ( .A1(n11555), .A2(n9526), .ZN(n9527) );
  AND2_X1 U12040 ( .A1(n9528), .A2(n9527), .ZN(n9530) );
  NAND2_X1 U12041 ( .A1(n9529), .A2(n9530), .ZN(n9803) );
  INV_X1 U12042 ( .A(n9529), .ZN(n9532) );
  INV_X1 U12043 ( .A(n9530), .ZN(n9531) );
  NAND2_X1 U12044 ( .A1(n9532), .A2(n9531), .ZN(n9533) );
  NAND2_X1 U12045 ( .A1(n9803), .A2(n9533), .ZN(n9535) );
  INV_X1 U12046 ( .A(n9804), .ZN(n9534) );
  AOI21_X1 U12047 ( .B1(n9536), .B2(n9535), .A(n9534), .ZN(n9547) );
  NAND2_X1 U12048 ( .A1(n11555), .A2(n14691), .ZN(n14682) );
  INV_X1 U12049 ( .A(n14682), .ZN(n9537) );
  AOI22_X1 U12050 ( .A1(n14480), .A2(n9537), .B1(n11831), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9546) );
  OR2_X1 U12051 ( .A1(n11656), .A2(n9596), .ZN(n9540) );
  INV_X1 U12052 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9591) );
  OR2_X1 U12053 ( .A1(n7529), .A2(n9591), .ZN(n9539) );
  NAND2_X1 U12054 ( .A1(n11152), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12055 ( .A1(n13949), .A2(n13898), .ZN(n9544) );
  NAND2_X1 U12056 ( .A1(n9542), .A2(n13964), .ZN(n13846) );
  INV_X2 U12057 ( .A(n13846), .ZN(n13899) );
  NAND2_X1 U12058 ( .A1(n11844), .A2(n13899), .ZN(n9543) );
  NAND2_X1 U12059 ( .A1(n9544), .A2(n9543), .ZN(n11552) );
  NAND2_X1 U12060 ( .A1(n11552), .A2(n14506), .ZN(n9545) );
  OAI211_X1 U12061 ( .C1(n9547), .C2(n14475), .A(n9546), .B(n9545), .ZN(
        P1_U3222) );
  INV_X1 U12062 ( .A(n9548), .ZN(n9550) );
  OAI222_X1 U12063 ( .A1(n13057), .A2(n9550), .B1(n13054), .B2(n9549), .C1(
        n12664), .C2(P3_U3151), .ZN(P3_U3278) );
  AOI211_X1 U12064 ( .C1(n9553), .C2(n9552), .A(n9551), .B(n14780), .ZN(n9554)
         );
  INV_X1 U12065 ( .A(n9554), .ZN(n9560) );
  AOI211_X1 U12066 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n15230), .ZN(n9558)
         );
  INV_X1 U12067 ( .A(n9558), .ZN(n9559) );
  NAND2_X1 U12068 ( .A1(n9560), .A2(n9559), .ZN(n9562) );
  NAND2_X1 U12069 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10092) );
  INV_X1 U12070 ( .A(n10092), .ZN(n9561) );
  AOI211_X1 U12071 ( .C1(n15233), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9562), .B(
        n9561), .ZN(n9563) );
  OAI21_X1 U12072 ( .B1(n14824), .B2(n9564), .A(n9563), .ZN(P2_U3218) );
  OAI21_X1 U12073 ( .B1(n9569), .B2(P1_D_REG_0__SCAN_IN), .A(n9566), .ZN(n9571) );
  INV_X1 U12074 ( .A(n9567), .ZN(n9568) );
  OR2_X1 U12075 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  AND2_X1 U12076 ( .A1(n9571), .A2(n9570), .ZN(n10223) );
  AND2_X2 U12077 ( .A1(n9593), .A2(n10223), .ZN(n14742) );
  NAND2_X1 U12078 ( .A1(n11845), .A2(n14385), .ZN(n9572) );
  AND2_X1 U12079 ( .A1(n13798), .A2(n9572), .ZN(n10582) );
  NAND2_X1 U12080 ( .A1(n10582), .A2(n14044), .ZN(n14707) );
  NAND2_X1 U12081 ( .A1(n11835), .A2(n12030), .ZN(n14665) );
  OR2_X1 U12082 ( .A1(n14665), .A2(n14385), .ZN(n14708) );
  AND2_X1 U12083 ( .A1(n11844), .A2(n9573), .ZN(n11549) );
  OR2_X1 U12084 ( .A1(n13950), .A2(n11555), .ZN(n9574) );
  OR2_X1 U12085 ( .A1(n12023), .A2(n6726), .ZN(n9576) );
  OR2_X1 U12086 ( .A1(n11685), .A2(n13968), .ZN(n9575) );
  OR2_X1 U12087 ( .A1(n13949), .A2(n9808), .ZN(n11849) );
  NAND2_X1 U12088 ( .A1(n13949), .A2(n9808), .ZN(n11839) );
  NAND2_X1 U12089 ( .A1(n11849), .A2(n11839), .ZN(n12062) );
  INV_X1 U12090 ( .A(n12062), .ZN(n9578) );
  OAI21_X1 U12091 ( .B1(n9579), .B2(n9578), .A(n9910), .ZN(n9580) );
  INV_X1 U12092 ( .A(n9580), .ZN(n10235) );
  AND2_X1 U12093 ( .A1(n11544), .A2(n14660), .ZN(n11546) );
  INV_X1 U12094 ( .A(n11546), .ZN(n9581) );
  NAND2_X1 U12095 ( .A1(n11546), .A2(n11848), .ZN(n10036) );
  AOI211_X1 U12096 ( .C1(n9808), .C2(n9581), .A(n14683), .B(n7203), .ZN(n10233) );
  AOI21_X1 U12097 ( .B1(n14691), .B2(n9808), .A(n10233), .ZN(n9589) );
  AND2_X1 U12098 ( .A1(n13950), .A2(n11544), .ZN(n11840) );
  INV_X1 U12099 ( .A(n11840), .ZN(n11847) );
  OR2_X1 U12100 ( .A1(n13950), .A2(n11544), .ZN(n9582) );
  NAND2_X1 U12101 ( .A1(n12061), .A2(n9582), .ZN(n11852) );
  NAND2_X1 U12102 ( .A1(n11835), .A2(n14385), .ZN(n11837) );
  NAND2_X1 U12103 ( .A1(n12019), .A2(n12036), .ZN(n12010) );
  NAND2_X1 U12104 ( .A1(n11837), .A2(n12010), .ZN(n14643) );
  INV_X1 U12105 ( .A(n6678), .ZN(n11547) );
  INV_X1 U12106 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12107 ( .A1(n11743), .A2(n9834), .ZN(n9586) );
  NAND2_X1 U12108 ( .A1(n11152), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U12109 ( .A1(n11039), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U12110 ( .A1(n11653), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9583) );
  INV_X1 U12111 ( .A(n13947), .ZN(n9587) );
  INV_X1 U12112 ( .A(n13898), .ZN(n13848) );
  OAI22_X1 U12113 ( .A1(n11547), .A2(n13846), .B1(n9587), .B2(n13848), .ZN(
        n11832) );
  AOI21_X1 U12114 ( .B1(n9588), .B2(n14643), .A(n11832), .ZN(n10230) );
  OAI211_X1 U12115 ( .C1(n14677), .C2(n10235), .A(n9589), .B(n10230), .ZN(
        n9594) );
  NAND2_X1 U12116 ( .A1(n9594), .A2(n14742), .ZN(n9590) );
  OAI21_X1 U12117 ( .B1(n14742), .B2(n9591), .A(n9590), .ZN(P1_U3465) );
  AND2_X2 U12118 ( .A1(n9593), .A2(n9592), .ZN(n14753) );
  NAND2_X1 U12119 ( .A1(n9594), .A2(n14753), .ZN(n9595) );
  OAI21_X1 U12120 ( .B1(n14753), .B2(n9596), .A(n9595), .ZN(P1_U3530) );
  INV_X1 U12121 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9597) );
  MUX2_X1 U12122 ( .A(n9597), .B(P1_REG1_REG_9__SCAN_IN), .S(n9605), .Z(n9600)
         );
  OAI21_X1 U12123 ( .B1(n10709), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9598), .ZN(
        n9599) );
  NAND2_X1 U12124 ( .A1(n9599), .A2(n9600), .ZN(n9933) );
  OAI21_X1 U12125 ( .B1(n9600), .B2(n9599), .A(n9933), .ZN(n9612) );
  INV_X1 U12126 ( .A(n9605), .ZN(n10714) );
  NAND2_X1 U12127 ( .A1(n14625), .A2(n10714), .ZN(n9602) );
  NAND2_X1 U12128 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9601) );
  OAI211_X1 U12129 ( .C1(n9603), .C2(n14633), .A(n9602), .B(n9601), .ZN(n9611)
         );
  INV_X1 U12130 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9606) );
  MUX2_X1 U12131 ( .A(n9606), .B(P1_REG2_REG_9__SCAN_IN), .S(n9605), .Z(n9607)
         );
  INV_X1 U12132 ( .A(n9607), .ZN(n9608) );
  NOR2_X1 U12133 ( .A1(n9609), .A2(n9608), .ZN(n9928) );
  AOI211_X1 U12134 ( .C1(n9609), .C2(n9608), .A(n14566), .B(n9928), .ZN(n9610)
         );
  AOI211_X1 U12135 ( .C1(n14617), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9613)
         );
  INV_X1 U12136 ( .A(n9613), .ZN(P1_U3252) );
  INV_X1 U12137 ( .A(n11346), .ZN(n9643) );
  NAND2_X1 U12138 ( .A1(n9614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9615) );
  XNOR2_X1 U12139 ( .A(n9615), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U12140 ( .A1(n14564), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14369), .ZN(n9616) );
  OAI21_X1 U12141 ( .B1(n9643), .B2(n14382), .A(n9616), .ZN(P1_U3341) );
  INV_X1 U12142 ( .A(n14842), .ZN(n9617) );
  NAND2_X1 U12143 ( .A1(n14895), .A2(n9619), .ZN(n9620) );
  OAI21_X1 U12144 ( .B1(n14895), .B2(n9621), .A(n9620), .ZN(P2_U3500) );
  INV_X2 U12145 ( .A(n14884), .ZN(n14886) );
  INV_X1 U12146 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12147 ( .A1(n9622), .A2(n9504), .ZN(n9623) );
  NAND2_X1 U12148 ( .A1(n9624), .A2(n9623), .ZN(n9626) );
  OAI21_X1 U12149 ( .B1(n9626), .B2(n9625), .A(n9942), .ZN(n10399) );
  INV_X1 U12150 ( .A(n10399), .ZN(n9635) );
  NAND2_X1 U12151 ( .A1(n9622), .A2(n13081), .ZN(n9627) );
  NAND2_X1 U12152 ( .A1(n9628), .A2(n9627), .ZN(n9630) );
  OAI21_X1 U12153 ( .B1(n9630), .B2(n9629), .A(n9947), .ZN(n9631) );
  AOI222_X1 U12154 ( .A1(n13488), .A2(n9631), .B1(n13211), .B2(n13437), .C1(
        n6748), .C2(n13435), .ZN(n10400) );
  AOI21_X1 U12155 ( .B1(n9632), .B2(n13158), .A(n13492), .ZN(n9633) );
  OR2_X1 U12156 ( .A1(n9632), .A2(n13158), .ZN(n10407) );
  AND2_X1 U12157 ( .A1(n9633), .A2(n10407), .ZN(n10395) );
  AOI21_X1 U12158 ( .B1(n14877), .B2(n13158), .A(n10395), .ZN(n9634) );
  OAI211_X1 U12159 ( .C1(n14875), .C2(n9635), .A(n10400), .B(n9634), .ZN(n9638) );
  NAND2_X1 U12160 ( .A1(n9638), .A2(n14886), .ZN(n9636) );
  OAI21_X1 U12161 ( .B1(n14886), .B2(n9637), .A(n9636), .ZN(P2_U3436) );
  NAND2_X1 U12162 ( .A1(n9638), .A2(n14895), .ZN(n9639) );
  OAI21_X1 U12163 ( .B1(n14895), .B2(n9336), .A(n9639), .ZN(P2_U3501) );
  INV_X1 U12164 ( .A(n9640), .ZN(n9642) );
  INV_X1 U12165 ( .A(n12688), .ZN(n12673) );
  OAI222_X1 U12166 ( .A1(n13057), .A2(n9642), .B1(n13054), .B2(n9641), .C1(
        n12673), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U12167 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9644) );
  INV_X1 U12168 ( .A(n14790), .ZN(n13272) );
  OAI222_X1 U12169 ( .A1(n13636), .A2(n9644), .B1(n13637), .B2(n9643), .C1(
        n13272), .C2(P2_U3088), .ZN(P2_U3313) );
  OR2_X1 U12170 ( .A1(n9966), .A2(P3_U3151), .ZN(n12547) );
  INV_X1 U12171 ( .A(n12547), .ZN(n9645) );
  OR2_X1 U12172 ( .A1(n9995), .A2(n9645), .ZN(n9662) );
  NAND2_X1 U12173 ( .A1(n12446), .A2(n9966), .ZN(n9647) );
  AND2_X1 U12174 ( .A1(n9647), .A2(n9646), .ZN(n9660) );
  NAND2_X1 U12175 ( .A1(n9662), .A2(n9660), .ZN(n9672) );
  MUX2_X1 U12176 ( .A(n9672), .B(n12562), .S(n9648), .Z(n14918) );
  MUX2_X1 U12177 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13050), .Z(n9649) );
  NOR2_X1 U12178 ( .A1(n9649), .A2(n9906), .ZN(n9650) );
  AOI21_X1 U12179 ( .B1(n9649), .B2(n9906), .A(n9650), .ZN(n9891) );
  MUX2_X1 U12180 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13050), .Z(n10199) );
  INV_X1 U12181 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U12182 ( .A1(n9891), .A2(n9892), .ZN(n9890) );
  INV_X1 U12183 ( .A(n9650), .ZN(n9658) );
  MUX2_X1 U12184 ( .A(n9652), .B(n9651), .S(n13050), .Z(n9654) );
  NAND2_X1 U12185 ( .A1(n9654), .A2(n9653), .ZN(n9702) );
  INV_X1 U12186 ( .A(n9654), .ZN(n9655) );
  NAND2_X1 U12187 ( .A1(n9655), .A2(n6500), .ZN(n9656) );
  NAND2_X1 U12188 ( .A1(n9702), .A2(n9656), .ZN(n9657) );
  AND3_X1 U12189 ( .A1(n9890), .A2(n9658), .A3(n9657), .ZN(n9659) );
  AND2_X1 U12190 ( .A1(P3_U3897), .A2(n12542), .ZN(n12703) );
  OAI21_X1 U12191 ( .B1(n10010), .B2(n9659), .A(n12703), .ZN(n9686) );
  INV_X1 U12192 ( .A(n9660), .ZN(n9661) );
  OAI22_X1 U12193 ( .A1(n14916), .A2(n9663), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8563), .ZN(n9684) );
  NAND2_X1 U12194 ( .A1(n9666), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9665) );
  NOR2_X1 U12195 ( .A1(n10834), .A2(n9894), .ZN(n9893) );
  NAND2_X1 U12196 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n6500), .ZN(n9667) );
  OAI21_X1 U12197 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n6500), .A(n9667), .ZN(
        n9668) );
  NOR2_X1 U12198 ( .A1(n9669), .A2(n9668), .ZN(n9692) );
  AOI21_X1 U12199 ( .B1(n9669), .B2(n9668), .A(n9692), .ZN(n9670) );
  NOR2_X1 U12200 ( .A1(n14934), .A2(n9670), .ZN(n9683) );
  NAND2_X1 U12201 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9673), .ZN(n9674) );
  AOI21_X1 U12202 ( .B1(n9675), .B2(n9674), .A(n9677), .ZN(n9676) );
  INV_X1 U12203 ( .A(n9676), .ZN(n9897) );
  NOR2_X1 U12204 ( .A1(n8542), .A2(n9897), .ZN(n9896) );
  NOR2_X1 U12205 ( .A1(n9677), .A2(n9896), .ZN(n9680) );
  NAND2_X1 U12206 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n9076), .ZN(n9678) );
  OAI21_X1 U12207 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n6500), .A(n9678), .ZN(
        n9679) );
  AOI21_X1 U12208 ( .B1(n9680), .B2(n9679), .A(n9725), .ZN(n9681) );
  NOR2_X1 U12209 ( .A1(n14926), .A2(n9681), .ZN(n9682) );
  NOR3_X1 U12210 ( .A1(n9684), .A2(n9683), .A3(n9682), .ZN(n9685) );
  OAI211_X1 U12211 ( .C1(n14918), .C2(n6500), .A(n9686), .B(n9685), .ZN(
        P3_U3184) );
  NAND2_X1 U12212 ( .A1(n10830), .A2(n10024), .ZN(n12330) );
  INV_X1 U12213 ( .A(n12330), .ZN(n9687) );
  NOR2_X1 U12214 ( .A1(n12333), .A2(n9687), .ZN(n12504) );
  NAND2_X1 U12215 ( .A1(n9971), .A2(n15004), .ZN(n9987) );
  AND2_X1 U12216 ( .A1(n9987), .A2(n12861), .ZN(n9688) );
  OAI22_X1 U12217 ( .A1(n12504), .A2(n9688), .B1(n8559), .B2(n14944), .ZN(
        n10654) );
  INV_X1 U12218 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9689) );
  OAI22_X1 U12219 ( .A1(n10024), .A2(n13039), .B1(n15010), .B2(n9689), .ZN(
        n9690) );
  AOI21_X1 U12220 ( .B1(n10654), .B2(n15010), .A(n9690), .ZN(n9691) );
  INV_X1 U12221 ( .A(n9691), .ZN(P3_U3390) );
  NAND2_X1 U12222 ( .A1(n9857), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12223 ( .A1(n9729), .A2(n10117), .ZN(n9694) );
  NAND2_X1 U12224 ( .A1(n9695), .A2(n9694), .ZN(n9843) );
  NOR2_X1 U12225 ( .A1(n7084), .A2(n9696), .ZN(n9697) );
  NAND2_X1 U12226 ( .A1(n9739), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9775) );
  OR2_X1 U12227 ( .A1(n9739), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12228 ( .A1(n9775), .A2(n9698), .ZN(n9700) );
  INV_X1 U12229 ( .A(n9776), .ZN(n9699) );
  AOI21_X1 U12230 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9744) );
  INV_X1 U12231 ( .A(n9702), .ZN(n10009) );
  MUX2_X1 U12232 ( .A(n9704), .B(n9703), .S(n12623), .Z(n9705) );
  NAND2_X1 U12233 ( .A1(n9705), .A2(n7180), .ZN(n9840) );
  INV_X1 U12234 ( .A(n9705), .ZN(n9706) );
  NAND2_X1 U12235 ( .A1(n9706), .A2(n9726), .ZN(n9707) );
  AND2_X1 U12236 ( .A1(n9840), .A2(n9707), .ZN(n10008) );
  OAI21_X1 U12237 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10007) );
  MUX2_X1 U12238 ( .A(n10117), .B(n15016), .S(n12623), .Z(n9708) );
  NAND2_X1 U12239 ( .A1(n9708), .A2(n9729), .ZN(n9711) );
  INV_X1 U12240 ( .A(n9708), .ZN(n9709) );
  NAND2_X1 U12241 ( .A1(n9709), .A2(n9857), .ZN(n9710) );
  NAND2_X1 U12242 ( .A1(n9711), .A2(n9710), .ZN(n9839) );
  INV_X1 U12243 ( .A(n9711), .ZN(n9746) );
  MUX2_X1 U12244 ( .A(n10869), .B(n9712), .S(n12623), .Z(n9713) );
  NAND2_X1 U12245 ( .A1(n9713), .A2(n7084), .ZN(n9722) );
  INV_X1 U12246 ( .A(n9713), .ZN(n9714) );
  NAND2_X1 U12247 ( .A1(n9714), .A2(n9757), .ZN(n9715) );
  AND2_X1 U12248 ( .A1(n9722), .A2(n9715), .ZN(n9745) );
  OAI21_X1 U12249 ( .B1(n9842), .B2(n9746), .A(n9745), .ZN(n9748) );
  MUX2_X1 U12250 ( .A(n9716), .B(n15019), .S(n12623), .Z(n9718) );
  INV_X1 U12251 ( .A(n9739), .ZN(n9717) );
  NAND2_X1 U12252 ( .A1(n9718), .A2(n9717), .ZN(n9778) );
  INV_X1 U12253 ( .A(n9718), .ZN(n9719) );
  NAND2_X1 U12254 ( .A1(n9719), .A2(n9739), .ZN(n9720) );
  NAND2_X1 U12255 ( .A1(n9778), .A2(n9720), .ZN(n9721) );
  AOI21_X1 U12256 ( .B1(n9748), .B2(n9722), .A(n9721), .ZN(n9785) );
  AND3_X1 U12257 ( .A1(n9748), .A2(n9722), .A3(n9721), .ZN(n9723) );
  OAI21_X1 U12258 ( .B1(n9785), .B2(n9723), .A(n12703), .ZN(n9743) );
  NAND2_X1 U12259 ( .A1(n9739), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9789) );
  OR2_X1 U12260 ( .A1(n9739), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12261 ( .A1(n9789), .A2(n9724), .ZN(n9734) );
  INV_X1 U12262 ( .A(n9734), .ZN(n9737) );
  NOR2_X1 U12263 ( .A1(n7180), .A2(n9727), .ZN(n9728) );
  NAND2_X1 U12264 ( .A1(n9857), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U12265 ( .A1(n9729), .A2(n15016), .ZN(n9730) );
  NAND2_X1 U12266 ( .A1(n9731), .A2(n9730), .ZN(n9847) );
  NOR2_X1 U12267 ( .A1(n7084), .A2(n9732), .ZN(n9733) );
  INV_X1 U12268 ( .A(n9735), .ZN(n9736) );
  OAI21_X1 U12269 ( .B1(n9737), .B2(n9736), .A(n9790), .ZN(n9741) );
  INV_X1 U12270 ( .A(n14926), .ZN(n12678) );
  AND2_X1 U12271 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n10298) );
  AOI21_X1 U12272 ( .B1(n14896), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10298), .ZN(
        n9738) );
  OAI21_X1 U12273 ( .B1(n14918), .B2(n9739), .A(n9738), .ZN(n9740) );
  AOI21_X1 U12274 ( .B1(n9741), .B2(n12678), .A(n9740), .ZN(n9742) );
  OAI211_X1 U12275 ( .C1(n9744), .C2(n14934), .A(n9743), .B(n9742), .ZN(
        P3_U3188) );
  OR3_X1 U12276 ( .A1(n9842), .A2(n9746), .A3(n9745), .ZN(n9747) );
  INV_X1 U12277 ( .A(n12703), .ZN(n14928) );
  AOI21_X1 U12278 ( .B1(n9748), .B2(n9747), .A(n14928), .ZN(n9760) );
  AOI21_X1 U12279 ( .B1(n9712), .B2(n9750), .A(n9749), .ZN(n9753) );
  NOR2_X1 U12280 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9751), .ZN(n10170) );
  AOI21_X1 U12281 ( .B1(n14896), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10170), .ZN(
        n9752) );
  OAI21_X1 U12282 ( .B1(n14926), .B2(n9753), .A(n9752), .ZN(n9759) );
  AOI21_X1 U12283 ( .B1(n10869), .B2(n9755), .A(n9754), .ZN(n9756) );
  OAI22_X1 U12284 ( .A1(n14918), .A2(n9757), .B1(n9756), .B2(n14934), .ZN(
        n9758) );
  OR3_X1 U12285 ( .A1(n9760), .A2(n9759), .A3(n9758), .ZN(P3_U3187) );
  OAI21_X1 U12286 ( .B1(n9765), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9761), .ZN(
        n9763) );
  INV_X1 U12287 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n13215) );
  MUX2_X1 U12288 ( .A(n13215), .B(P2_REG1_REG_10__SCAN_IN), .S(n13226), .Z(
        n9762) );
  AOI211_X1 U12289 ( .C1(n9763), .C2(n9762), .A(n14780), .B(n13223), .ZN(n9772) );
  OAI21_X1 U12290 ( .B1(n9765), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9764), .ZN(
        n9768) );
  INV_X1 U12291 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9766) );
  MUX2_X1 U12292 ( .A(n9766), .B(P2_REG2_REG_10__SCAN_IN), .S(n13226), .Z(
        n9767) );
  NOR2_X1 U12293 ( .A1(n9768), .A2(n9767), .ZN(n13225) );
  AOI211_X1 U12294 ( .C1(n9768), .C2(n9767), .A(n15230), .B(n13225), .ZN(n9771) );
  NAND2_X1 U12295 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10915)
         );
  NAND2_X1 U12296 ( .A1(n15233), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9769) );
  OAI211_X1 U12297 ( .C1(n14824), .C2(n13216), .A(n10915), .B(n9769), .ZN(
        n9770) );
  OR3_X1 U12298 ( .A1(n9772), .A2(n9771), .A3(n9770), .ZN(P2_U3224) );
  OAI222_X1 U12299 ( .A1(P3_U3151), .A2(n12694), .B1(n13054), .B2(n9774), .C1(
        n13057), .C2(n9773), .ZN(P3_U3276) );
  AOI21_X1 U12300 ( .B1(n10783), .B2(n9777), .A(n9859), .ZN(n9798) );
  INV_X1 U12301 ( .A(n9778), .ZN(n9784) );
  MUX2_X1 U12302 ( .A(n10783), .B(n9779), .S(n12623), .Z(n9780) );
  NAND2_X1 U12303 ( .A1(n9780), .A2(n9877), .ZN(n9870) );
  INV_X1 U12304 ( .A(n9780), .ZN(n9781) );
  NAND2_X1 U12305 ( .A1(n9781), .A2(n9791), .ZN(n9782) );
  AND2_X1 U12306 ( .A1(n9870), .A2(n9782), .ZN(n9783) );
  OAI21_X1 U12307 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9871) );
  INV_X1 U12308 ( .A(n9871), .ZN(n9787) );
  NOR3_X1 U12309 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(n9786) );
  OAI21_X1 U12310 ( .B1(n9787), .B2(n9786), .A(n12703), .ZN(n9797) );
  INV_X1 U12311 ( .A(n14918), .ZN(n12669) );
  AND2_X1 U12312 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10563) );
  INV_X1 U12313 ( .A(n10563), .ZN(n9788) );
  OAI21_X1 U12314 ( .B1(n14916), .B2(n8351), .A(n9788), .ZN(n9795) );
  AOI21_X1 U12315 ( .B1(n9779), .B2(n9792), .A(n9878), .ZN(n9793) );
  NOR2_X1 U12316 ( .A1(n9793), .A2(n14926), .ZN(n9794) );
  AOI211_X1 U12317 ( .C1(n12669), .C2(n9877), .A(n9795), .B(n9794), .ZN(n9796)
         );
  OAI211_X1 U12318 ( .C1(n9798), .C2(n14934), .A(n9797), .B(n9796), .ZN(
        P3_U3189) );
  NAND2_X1 U12319 ( .A1(n6482), .A2(n9799), .ZN(n9802) );
  OR2_X1 U12320 ( .A1(n12023), .A2(n6734), .ZN(n9801) );
  OR2_X1 U12321 ( .A1(n11685), .A2(n13981), .ZN(n9800) );
  NAND2_X1 U12322 ( .A1(n13949), .A2(n9526), .ZN(n9806) );
  NAND2_X1 U12323 ( .A1(n9808), .A2(n13800), .ZN(n9805) );
  NAND2_X1 U12324 ( .A1(n9806), .A2(n9805), .ZN(n9807) );
  XNOR2_X1 U12325 ( .A(n9807), .B(n13752), .ZN(n9813) );
  NAND2_X1 U12326 ( .A1(n13949), .A2(n10452), .ZN(n9810) );
  NAND2_X1 U12327 ( .A1(n9808), .A2(n9526), .ZN(n9809) );
  NAND2_X1 U12328 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  XNOR2_X1 U12329 ( .A(n9813), .B(n9811), .ZN(n11829) );
  INV_X1 U12330 ( .A(n9811), .ZN(n9812) );
  NAND2_X1 U12331 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U12332 ( .A1(n13947), .A2(n9526), .ZN(n9816) );
  OR2_X1 U12333 ( .A1(n10236), .A2(n13682), .ZN(n9815) );
  NAND2_X1 U12334 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  XNOR2_X1 U12335 ( .A(n9817), .B(n13752), .ZN(n10363) );
  BUF_X2 U12336 ( .A(n10452), .Z(n13764) );
  NAND2_X1 U12337 ( .A1(n13947), .A2(n13764), .ZN(n9819) );
  OR2_X1 U12338 ( .A1(n10236), .A2(n13690), .ZN(n9818) );
  NAND2_X1 U12339 ( .A1(n9819), .A2(n9818), .ZN(n10364) );
  XNOR2_X1 U12340 ( .A(n10363), .B(n10364), .ZN(n9820) );
  OAI211_X1 U12341 ( .C1(n9821), .C2(n9820), .A(n10367), .B(n14504), .ZN(n9838) );
  NAND3_X1 U12342 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n9825) );
  NAND2_X1 U12343 ( .A1(n9825), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9826) );
  AND2_X1 U12344 ( .A1(n9826), .A2(n12105), .ZN(n14511) );
  INV_X1 U12345 ( .A(n14511), .ZN(n13904) );
  NAND2_X1 U12346 ( .A1(n13949), .A2(n13899), .ZN(n9833) );
  NAND2_X1 U12347 ( .A1(n12006), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12348 ( .A1(n6491), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9830) );
  INV_X1 U12349 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9827) );
  XNOR2_X1 U12350 ( .A(n9827), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10579) );
  NAND2_X1 U12351 ( .A1(n11743), .A2(n10579), .ZN(n9829) );
  NAND2_X1 U12352 ( .A1(n11039), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9828) );
  NAND2_X1 U12353 ( .A1(n13946), .A2(n13898), .ZN(n9832) );
  NAND2_X1 U12354 ( .A1(n9833), .A2(n9832), .ZN(n10033) );
  INV_X1 U12355 ( .A(n10033), .ZN(n9835) );
  OAI22_X1 U12356 ( .A1(n9835), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9834), .ZN(n9836) );
  AOI21_X1 U12357 ( .B1(n9834), .B2(n13904), .A(n9836), .ZN(n9837) );
  OAI211_X1 U12358 ( .C1(n10236), .C2(n13907), .A(n9838), .B(n9837), .ZN(
        P1_U3218) );
  AND3_X1 U12359 ( .A1(n10007), .A2(n9840), .A3(n9839), .ZN(n9841) );
  OAI21_X1 U12360 ( .B1(n9842), .B2(n9841), .A(n12703), .ZN(n9856) );
  NAND2_X1 U12361 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  AOI21_X1 U12362 ( .B1(n9846), .B2(n9845), .A(n14934), .ZN(n9854) );
  NAND2_X1 U12363 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  AOI21_X1 U12364 ( .B1(n9850), .B2(n9849), .A(n14926), .ZN(n9853) );
  INV_X1 U12365 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U12366 ( .A1(n14916), .A2(n9851), .ZN(n9852) );
  AND2_X1 U12367 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10149) );
  NOR4_X1 U12368 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n10149), .ZN(n9855)
         );
  OAI211_X1 U12369 ( .C1(n14918), .C2(n9857), .A(n9856), .B(n9855), .ZN(
        P3_U3186) );
  NOR2_X1 U12370 ( .A1(n9877), .A2(n9858), .ZN(n9860) );
  NAND2_X1 U12371 ( .A1(n9880), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10321) );
  OAI21_X1 U12372 ( .B1(n9880), .B2(P3_REG2_REG_8__SCAN_IN), .A(n10321), .ZN(
        n9862) );
  INV_X1 U12373 ( .A(n10322), .ZN(n9861) );
  AOI21_X1 U12374 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9889) );
  MUX2_X1 U12375 ( .A(n9865), .B(n9864), .S(n12623), .Z(n9866) );
  INV_X1 U12376 ( .A(n9880), .ZN(n9886) );
  NAND2_X1 U12377 ( .A1(n9866), .A2(n9886), .ZN(n10307) );
  INV_X1 U12378 ( .A(n9866), .ZN(n9867) );
  NAND2_X1 U12379 ( .A1(n9867), .A2(n9880), .ZN(n9868) );
  NAND2_X1 U12380 ( .A1(n10307), .A2(n9868), .ZN(n9869) );
  AND3_X1 U12381 ( .A1(n9871), .A2(n9870), .A3(n9869), .ZN(n9872) );
  OAI21_X1 U12382 ( .B1(n10315), .B2(n9872), .A(n12703), .ZN(n9888) );
  INV_X1 U12383 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n9875) );
  NOR2_X1 U12384 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9873), .ZN(n10772) );
  INV_X1 U12385 ( .A(n10772), .ZN(n9874) );
  OAI21_X1 U12386 ( .B1(n14916), .B2(n9875), .A(n9874), .ZN(n9885) );
  NOR2_X1 U12387 ( .A1(n9877), .A2(n9876), .ZN(n9879) );
  NAND2_X1 U12388 ( .A1(n9880), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10324) );
  OAI21_X1 U12389 ( .B1(n9880), .B2(P3_REG1_REG_8__SCAN_IN), .A(n10324), .ZN(
        n9881) );
  NAND2_X1 U12390 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  AOI21_X1 U12391 ( .B1(n10325), .B2(n9883), .A(n14926), .ZN(n9884) );
  AOI211_X1 U12392 ( .C1(n12669), .C2(n9886), .A(n9885), .B(n9884), .ZN(n9887)
         );
  OAI211_X1 U12393 ( .C1(n9889), .C2(n14934), .A(n9888), .B(n9887), .ZN(
        P3_U3190) );
  OAI21_X1 U12394 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9904) );
  AOI21_X1 U12395 ( .B1(n10834), .B2(n9894), .A(n9893), .ZN(n9902) );
  OAI22_X1 U12396 ( .A1(n14916), .A2(n9895), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8543), .ZN(n9900) );
  AOI21_X1 U12397 ( .B1(n8542), .B2(n9897), .A(n9896), .ZN(n9898) );
  NOR2_X1 U12398 ( .A1(n14926), .A2(n9898), .ZN(n9899) );
  NOR2_X1 U12399 ( .A1(n9900), .A2(n9899), .ZN(n9901) );
  OAI21_X1 U12400 ( .B1(n9902), .B2(n14934), .A(n9901), .ZN(n9903) );
  AOI21_X1 U12401 ( .B1(n12703), .B2(n9904), .A(n9903), .ZN(n9905) );
  OAI21_X1 U12402 ( .B1(n9906), .B2(n14918), .A(n9905), .ZN(P3_U3183) );
  INV_X1 U12403 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12404 ( .A1(n9907), .A2(n12025), .ZN(n9909) );
  INV_X2 U12405 ( .A(n12013), .ZN(n11646) );
  AOI22_X1 U12406 ( .A1(n11646), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11645), 
        .B2(n13999), .ZN(n9908) );
  INV_X1 U12407 ( .A(n11862), .ZN(n10581) );
  XNOR2_X1 U12408 ( .A(n13946), .B(n10581), .ZN(n12065) );
  NAND2_X1 U12409 ( .A1(n9910), .A2(n11849), .ZN(n10029) );
  OR2_X1 U12410 ( .A1(n13947), .A2(n11857), .ZN(n9911) );
  XOR2_X1 U12411 ( .A(n10501), .B(n12065), .Z(n10583) );
  OR2_X1 U12412 ( .A1(n13949), .A2(n11848), .ZN(n9912) );
  NAND2_X1 U12413 ( .A1(n9913), .A2(n9912), .ZN(n10030) );
  INV_X1 U12414 ( .A(n11854), .ZN(n12064) );
  NOR2_X1 U12415 ( .A1(n13947), .A2(n10236), .ZN(n9914) );
  XNOR2_X1 U12416 ( .A(n10507), .B(n12065), .ZN(n9922) );
  NAND2_X1 U12417 ( .A1(n6491), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12418 ( .A1(n11653), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9919) );
  AOI21_X1 U12419 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U12420 ( .A1(n9915), .A2(n10457), .ZN(n10456) );
  NAND2_X1 U12421 ( .A1(n11743), .A2(n10456), .ZN(n9918) );
  OR2_X1 U12422 ( .A1(n11656), .A2(n9916), .ZN(n9917) );
  NAND2_X1 U12423 ( .A1(n13947), .A2(n13899), .ZN(n9921) );
  OAI21_X1 U12424 ( .B1(n11866), .B2(n13848), .A(n9921), .ZN(n10368) );
  AOI21_X1 U12425 ( .B1(n9922), .B2(n14643), .A(n10368), .ZN(n10588) );
  AOI211_X1 U12426 ( .C1(n11862), .C2(n10034), .A(n14683), .B(n10513), .ZN(
        n10586) );
  AOI21_X1 U12427 ( .B1(n14691), .B2(n11862), .A(n10586), .ZN(n9923) );
  OAI211_X1 U12428 ( .C1(n10583), .C2(n14677), .A(n10588), .B(n9923), .ZN(
        n9926) );
  NAND2_X1 U12429 ( .A1(n9926), .A2(n14742), .ZN(n9924) );
  OAI21_X1 U12430 ( .B1(n14742), .B2(n9925), .A(n9924), .ZN(P1_U3471) );
  NAND2_X1 U12431 ( .A1(n9926), .A2(n14753), .ZN(n9927) );
  OAI21_X1 U12432 ( .B1(n14753), .B2(n9228), .A(n9927), .ZN(P1_U3532) );
  MUX2_X1 U12433 ( .A(n10899), .B(P1_REG2_REG_10__SCAN_IN), .S(n9936), .Z(
        n9929) );
  INV_X1 U12434 ( .A(n9929), .ZN(n9930) );
  NOR2_X1 U12435 ( .A1(n9931), .A2(n9930), .ZN(n10353) );
  AOI211_X1 U12436 ( .C1(n9931), .C2(n9930), .A(n14566), .B(n10353), .ZN(n9940) );
  INV_X1 U12437 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9932) );
  MUX2_X1 U12438 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9932), .S(n9936), .Z(n9935) );
  OAI21_X1 U12439 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10714), .A(n9933), .ZN(
        n9934) );
  NOR2_X1 U12440 ( .A1(n9934), .A2(n9935), .ZN(n10347) );
  AOI211_X1 U12441 ( .C1(n9935), .C2(n9934), .A(n14548), .B(n10347), .ZN(n9939) );
  INV_X1 U12442 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15046) );
  INV_X1 U12443 ( .A(n9936), .ZN(n10878) );
  NAND2_X1 U12444 ( .A1(n14625), .A2(n10878), .ZN(n9937) );
  NAND2_X1 U12445 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14472)
         );
  OAI211_X1 U12446 ( .C1(n15046), .C2(n14633), .A(n9937), .B(n14472), .ZN(
        n9938) );
  OR3_X1 U12447 ( .A1(n9940), .A2(n9939), .A3(n9938), .ZN(P1_U3253) );
  NAND2_X1 U12448 ( .A1(n8293), .A2(n10397), .ZN(n9941) );
  NAND2_X1 U12449 ( .A1(n9951), .A2(n14860), .ZN(n9943) );
  INV_X1 U12450 ( .A(n9949), .ZN(n9944) );
  OAI21_X1 U12451 ( .B1(n9945), .B2(n9944), .A(n10266), .ZN(n9956) );
  OAI211_X1 U12452 ( .C1(n10410), .C2(n10093), .A(n10280), .B(n10055), .ZN(
        n10334) );
  OAI21_X1 U12453 ( .B1(n10093), .B2(n14859), .A(n10334), .ZN(n9955) );
  INV_X1 U12454 ( .A(n9956), .ZN(n10339) );
  NAND2_X1 U12455 ( .A1(n8293), .A2(n13158), .ZN(n9946) );
  INV_X1 U12456 ( .A(n10404), .ZN(n10415) );
  NAND2_X1 U12457 ( .A1(n10416), .A2(n10415), .ZN(n10414) );
  NAND2_X1 U12458 ( .A1(n9951), .A2(n10406), .ZN(n9948) );
  NAND2_X1 U12459 ( .A1(n10414), .A2(n9948), .ZN(n9950) );
  NAND2_X1 U12460 ( .A1(n9950), .A2(n9949), .ZN(n10271) );
  OAI21_X1 U12461 ( .B1(n9950), .B2(n9949), .A(n10271), .ZN(n9953) );
  INV_X1 U12462 ( .A(n13209), .ZN(n10527) );
  OAI22_X1 U12463 ( .A1(n9951), .A2(n13445), .B1(n10527), .B2(n13447), .ZN(
        n9952) );
  AOI21_X1 U12464 ( .B1(n9953), .B2(n13488), .A(n9952), .ZN(n9954) );
  OAI21_X1 U12465 ( .B1(n10339), .B2(n14849), .A(n9954), .ZN(n10331) );
  AOI211_X1 U12466 ( .C1(n14855), .C2(n9956), .A(n9955), .B(n10331), .ZN(
        n10121) );
  NAND2_X1 U12467 ( .A1(n14893), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9957) );
  OAI21_X1 U12468 ( .B1(n10121), .B2(n14893), .A(n9957), .ZN(P2_U3503) );
  INV_X1 U12469 ( .A(n11425), .ZN(n9964) );
  INV_X1 U12470 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U12471 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  OAI21_X1 U12472 ( .B1(n9961), .B2(n9960), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9963) );
  INV_X1 U12473 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9962) );
  XNOR2_X1 U12474 ( .A(n9963), .B(n9962), .ZN(n14026) );
  OAI222_X1 U12475 ( .A1(n14379), .A2(n7027), .B1(n14382), .B2(n9964), .C1(
        n14026), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U12476 ( .A(n14800), .ZN(n13273) );
  OAI222_X1 U12477 ( .A1(n13636), .A2(n9965), .B1(n13637), .B2(n9964), .C1(
        P2_U3088), .C2(n13273), .ZN(P2_U3312) );
  INV_X1 U12478 ( .A(n9986), .ZN(n9970) );
  NAND3_X1 U12479 ( .A1(n9968), .A2(n9967), .A3(n9966), .ZN(n9969) );
  AOI21_X1 U12480 ( .B1(n9996), .B2(n9970), .A(n9969), .ZN(n9973) );
  NAND2_X1 U12481 ( .A1(n9992), .A2(n9971), .ZN(n9972) );
  NAND2_X1 U12482 ( .A1(n9973), .A2(n9972), .ZN(n9974) );
  NAND2_X1 U12483 ( .A1(n9974), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9977) );
  NAND2_X1 U12484 ( .A1(n9996), .A2(n9975), .ZN(n9976) );
  NOR2_X1 U12485 ( .A1(n12257), .A2(P3_U3151), .ZN(n10131) );
  INV_X1 U12486 ( .A(n10827), .ZN(n12501) );
  NAND2_X1 U12487 ( .A1(n12332), .A2(n12690), .ZN(n9979) );
  NAND2_X1 U12488 ( .A1(n9979), .A2(n10386), .ZN(n9980) );
  NAND2_X1 U12489 ( .A1(n12564), .A2(n9982), .ZN(n9983) );
  OAI21_X1 U12490 ( .B1(n12501), .B2(n9984), .A(n10130), .ZN(n9990) );
  NAND3_X1 U12491 ( .A1(n12564), .A2(n12153), .A3(n10826), .ZN(n9985) );
  AOI21_X1 U12492 ( .B1(n9985), .B2(n10129), .A(n10828), .ZN(n9989) );
  OAI22_X1 U12493 ( .A1(n9992), .A2(n9987), .B1(n9996), .B2(n9986), .ZN(n9988)
         );
  OAI21_X1 U12494 ( .B1(n9990), .B2(n9989), .A(n12280), .ZN(n10004) );
  NAND2_X1 U12495 ( .A1(n9995), .A2(n15001), .ZN(n9991) );
  INV_X1 U12496 ( .A(n10830), .ZN(n10001) );
  AND2_X1 U12497 ( .A1(n9995), .A2(n9994), .ZN(n9998) );
  NAND2_X1 U12498 ( .A1(n9998), .A2(n12898), .ZN(n12543) );
  INV_X1 U12499 ( .A(n12543), .ZN(n9997) );
  INV_X1 U12500 ( .A(n9996), .ZN(n10000) );
  NAND2_X1 U12501 ( .A1(n9997), .A2(n10000), .ZN(n12291) );
  AND2_X1 U12502 ( .A1(n12896), .A2(n9998), .ZN(n9999) );
  NAND2_X1 U12503 ( .A1(n10000), .A2(n9999), .ZN(n12303) );
  OAI22_X1 U12504 ( .A1(n10001), .A2(n12291), .B1(n10158), .B2(n12303), .ZN(
        n10002) );
  AOI21_X1 U12505 ( .B1(n10826), .B2(n9993), .A(n10002), .ZN(n10003) );
  OAI211_X1 U12506 ( .C1(n10131), .C2(n8543), .A(n10004), .B(n10003), .ZN(
        P3_U3162) );
  OAI22_X1 U12507 ( .A1(n12961), .A2(n10024), .B1(n15025), .B2(n8550), .ZN(
        n10005) );
  AOI21_X1 U12508 ( .B1(n10654), .B2(n15025), .A(n10005), .ZN(n10006) );
  INV_X1 U12509 ( .A(n10006), .ZN(P3_U3459) );
  INV_X1 U12510 ( .A(n10007), .ZN(n10012) );
  NOR3_X1 U12511 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(n10011) );
  OAI21_X1 U12512 ( .B1(n10012), .B2(n10011), .A(n12703), .ZN(n10023) );
  AOI21_X1 U12513 ( .B1(n9704), .B2(n10014), .A(n10013), .ZN(n10020) );
  INV_X1 U12514 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12515 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10215), .ZN(n10160) );
  AOI21_X1 U12516 ( .B1(n9703), .B2(n10016), .A(n10015), .ZN(n10017) );
  NOR2_X1 U12517 ( .A1(n14926), .A2(n10017), .ZN(n10018) );
  AOI211_X1 U12518 ( .C1(n14896), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10160), .B(
        n10018), .ZN(n10019) );
  OAI21_X1 U12519 ( .B1(n10020), .B2(n14934), .A(n10019), .ZN(n10021) );
  AOI21_X1 U12520 ( .B1(n7180), .B2(n12669), .A(n10021), .ZN(n10022) );
  NAND2_X1 U12521 ( .A1(n10023), .A2(n10022), .ZN(P3_U3185) );
  INV_X1 U12522 ( .A(n12504), .ZN(n10026) );
  OAI22_X1 U12523 ( .A1(n12288), .A2(n10024), .B1(n8559), .B2(n12303), .ZN(
        n10025) );
  AOI21_X1 U12524 ( .B1(n10026), .B2(n12280), .A(n10025), .ZN(n10027) );
  OAI21_X1 U12525 ( .B1(n10131), .B2(n8549), .A(n10027), .ZN(P3_U3172) );
  INV_X1 U12526 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10040) );
  OAI21_X1 U12527 ( .B1(n10029), .B2(n11854), .A(n10028), .ZN(n10241) );
  INV_X1 U12528 ( .A(n10241), .ZN(n10038) );
  INV_X1 U12529 ( .A(n14707), .ZN(n14723) );
  XNOR2_X1 U12530 ( .A(n11854), .B(n10030), .ZN(n10031) );
  INV_X1 U12531 ( .A(n14643), .ZN(n14676) );
  NOR2_X1 U12532 ( .A1(n10031), .A2(n14676), .ZN(n10032) );
  AOI211_X1 U12533 ( .C1(n14723), .C2(n10241), .A(n10033), .B(n10032), .ZN(
        n10244) );
  INV_X1 U12534 ( .A(n10034), .ZN(n10035) );
  AOI211_X1 U12535 ( .C1(n11857), .C2(n10036), .A(n14683), .B(n10035), .ZN(
        n10240) );
  AOI21_X1 U12536 ( .B1(n14691), .B2(n11857), .A(n10240), .ZN(n10037) );
  OAI211_X1 U12537 ( .C1(n10038), .C2(n14708), .A(n10244), .B(n10037), .ZN(
        n10041) );
  NAND2_X1 U12538 ( .A1(n10041), .A2(n14742), .ZN(n10039) );
  OAI21_X1 U12539 ( .B1(n14742), .B2(n10040), .A(n10039), .ZN(P1_U3468) );
  NAND2_X1 U12540 ( .A1(n10041), .A2(n14753), .ZN(n10042) );
  OAI21_X1 U12541 ( .B1(n14753), .B2(n9226), .A(n10042), .ZN(P1_U3531) );
  NAND2_X4 U12542 ( .A1(n10043), .A2(n10183), .ZN(n11612) );
  NAND2_X1 U12543 ( .A1(n6748), .A2(n10911), .ZN(n10048) );
  OR2_X1 U12544 ( .A1(n11612), .A2(n10377), .ZN(n10046) );
  NAND2_X1 U12545 ( .A1(n10044), .A2(n10911), .ZN(n10045) );
  INV_X1 U12546 ( .A(n10047), .ZN(n10049) );
  NAND2_X1 U12547 ( .A1(n10049), .A2(n10048), .ZN(n10050) );
  XNOR2_X1 U12548 ( .A(n11612), .B(n13158), .ZN(n10051) );
  NAND2_X1 U12549 ( .A1(n13212), .A2(n10911), .ZN(n10052) );
  XNOR2_X1 U12550 ( .A(n10051), .B(n10052), .ZN(n13161) );
  INV_X1 U12551 ( .A(n10051), .ZN(n10053) );
  NAND2_X1 U12552 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  XNOR2_X1 U12553 ( .A(n11612), .B(n10406), .ZN(n10056) );
  AND2_X1 U12554 ( .A1(n10911), .A2(n13211), .ZN(n10057) );
  NAND2_X1 U12555 ( .A1(n10056), .A2(n10057), .ZN(n10086) );
  INV_X1 U12556 ( .A(n10056), .ZN(n10059) );
  INV_X1 U12557 ( .A(n10057), .ZN(n10058) );
  NAND2_X1 U12558 ( .A1(n10059), .A2(n10058), .ZN(n10060) );
  NAND2_X1 U12559 ( .A1(n10086), .A2(n10060), .ZN(n10069) );
  NAND2_X1 U12560 ( .A1(n10062), .A2(n10061), .ZN(n10179) );
  OR2_X1 U12561 ( .A1(n10179), .A2(n14842), .ZN(n10078) );
  NOR2_X1 U12562 ( .A1(n10078), .A2(n14845), .ZN(n10071) );
  INV_X1 U12563 ( .A(n10063), .ZN(n10064) );
  AND2_X1 U12564 ( .A1(n14859), .A2(n10064), .ZN(n10065) );
  INV_X1 U12565 ( .A(n10070), .ZN(n10067) );
  INV_X1 U12566 ( .A(n10087), .ZN(n10068) );
  AOI211_X1 U12567 ( .C1(n10070), .C2(n10069), .A(n13187), .B(n10068), .ZN(
        n10085) );
  INV_X1 U12568 ( .A(n10071), .ZN(n10076) );
  INV_X1 U12569 ( .A(n14848), .ZN(n10073) );
  NAND2_X1 U12570 ( .A1(n10073), .A2(n10072), .ZN(n10187) );
  INV_X1 U12571 ( .A(n10077), .ZN(n10074) );
  INV_X1 U12572 ( .A(n13173), .ZN(n13154) );
  NAND2_X1 U12573 ( .A1(n13181), .A2(n13437), .ZN(n13138) );
  INV_X1 U12574 ( .A(n13210), .ZN(n10274) );
  OAI22_X1 U12575 ( .A1(n14860), .A2(n13154), .B1(n13138), .B2(n10274), .ZN(
        n10084) );
  NAND2_X1 U12576 ( .A1(n13181), .A2(n13435), .ZN(n13139) );
  NAND2_X1 U12577 ( .A1(n10078), .A2(n10077), .ZN(n10081) );
  AND2_X1 U12578 ( .A1(n10079), .A2(n10180), .ZN(n10080) );
  NAND2_X1 U12579 ( .A1(n10081), .A2(n10080), .ZN(n10380) );
  NAND2_X1 U12580 ( .A1(n10380), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13183) );
  INV_X1 U12581 ( .A(n13183), .ZN(n13151) );
  NOR2_X1 U12582 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10411), .ZN(n14759) );
  AOI21_X1 U12583 ( .B1(n13151), .B2(n10411), .A(n14759), .ZN(n10082) );
  OAI21_X1 U12584 ( .B1(n13139), .B2(n8293), .A(n10082), .ZN(n10083) );
  OR3_X1 U12585 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(P2_U3190) );
  XNOR2_X1 U12586 ( .A(n11612), .B(n10093), .ZN(n10099) );
  INV_X2 U12587 ( .A(n10055), .ZN(n13492) );
  NAND2_X1 U12588 ( .A1(n13210), .A2(n10911), .ZN(n10098) );
  XNOR2_X1 U12589 ( .A(n10099), .B(n10098), .ZN(n10091) );
  INV_X1 U12590 ( .A(n10101), .ZN(n10089) );
  AOI21_X1 U12591 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(n10097) );
  INV_X1 U12592 ( .A(n13139), .ZN(n13156) );
  OAI21_X1 U12593 ( .B1(n13183), .B2(n10333), .A(n10092), .ZN(n10095) );
  OAI22_X1 U12594 ( .A1(n10093), .A2(n13154), .B1(n13138), .B2(n10527), .ZN(
        n10094) );
  AOI211_X1 U12595 ( .C1(n13156), .C2(n13211), .A(n10095), .B(n10094), .ZN(
        n10096) );
  OAI21_X1 U12596 ( .B1(n10097), .B2(n13187), .A(n10096), .ZN(P2_U3202) );
  XNOR2_X1 U12597 ( .A(n14868), .B(n11612), .ZN(n10245) );
  NAND2_X1 U12598 ( .A1(n13209), .A2(n10911), .ZN(n10246) );
  XNOR2_X1 U12599 ( .A(n10245), .B(n10246), .ZN(n10103) );
  NAND2_X1 U12600 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  OAI21_X1 U12601 ( .B1(n10103), .B2(n10102), .A(n10249), .ZN(n10108) );
  INV_X1 U12602 ( .A(n13208), .ZN(n10427) );
  OAI22_X1 U12603 ( .A1(n6997), .A2(n13154), .B1(n13138), .B2(n10427), .ZN(
        n10107) );
  NAND2_X1 U12604 ( .A1(n13151), .A2(n10279), .ZN(n10104) );
  OAI211_X1 U12605 ( .C1(n13139), .C2(n10274), .A(n10105), .B(n10104), .ZN(
        n10106) );
  AOI211_X1 U12606 ( .C1(n10108), .C2(n13162), .A(n10107), .B(n10106), .ZN(
        n10109) );
  INV_X1 U12607 ( .A(n10109), .ZN(P2_U3199) );
  XNOR2_X1 U12608 ( .A(n10110), .B(n10112), .ZN(n14972) );
  OAI211_X1 U12609 ( .C1(n10113), .C2(n10112), .A(n10111), .B(n14947), .ZN(
        n10116) );
  OAI22_X1 U12610 ( .A1(n10844), .A2(n14944), .B1(n14945), .B2(n14943), .ZN(
        n10114) );
  INV_X1 U12611 ( .A(n10114), .ZN(n10115) );
  AND2_X1 U12612 ( .A1(n10116), .A2(n10115), .ZN(n14971) );
  MUX2_X1 U12613 ( .A(n14971), .B(n10117), .S(n14955), .Z(n10120) );
  INV_X1 U12614 ( .A(n10118), .ZN(n10151) );
  AOI22_X1 U12615 ( .A1(n12889), .A2(n6914), .B1(n12888), .B2(n10151), .ZN(
        n10119) );
  OAI211_X1 U12616 ( .C1(n12892), .C2(n14972), .A(n10120), .B(n10119), .ZN(
        P3_U3229) );
  INV_X1 U12617 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10123) );
  OR2_X1 U12618 ( .A1(n10121), .A2(n14884), .ZN(n10122) );
  OAI21_X1 U12619 ( .B1(n14886), .B2(n10123), .A(n10122), .ZN(P2_U3442) );
  NAND2_X1 U12620 ( .A1(n6623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U12621 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10124), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10125) );
  NAND2_X1 U12622 ( .A1(n10125), .A2(n10301), .ZN(n14596) );
  INV_X1 U12623 ( .A(n11509), .ZN(n10127) );
  OAI222_X1 U12624 ( .A1(P1_U3086), .A2(n14596), .B1(n14382), .B2(n10127), 
        .C1(n10126), .C2(n14379), .ZN(P1_U3339) );
  INV_X1 U12625 ( .A(n13276), .ZN(n14810) );
  OAI222_X1 U12626 ( .A1(n13636), .A2(n10128), .B1(n13637), .B2(n10127), .C1(
        n14810), .C2(P2_U3088), .ZN(P2_U3311) );
  XNOR2_X1 U12627 ( .A(n12153), .B(n14937), .ZN(n10137) );
  XNOR2_X1 U12628 ( .A(n10137), .B(n6655), .ZN(n10140) );
  NAND2_X1 U12629 ( .A1(n10130), .A2(n10129), .ZN(n10141) );
  XOR2_X1 U12630 ( .A(n10140), .B(n10141), .Z(n10136) );
  OAI22_X1 U12631 ( .A1(n8559), .A2(n12291), .B1(n14945), .B2(n12303), .ZN(
        n10133) );
  NOR2_X1 U12632 ( .A1(n10131), .A2(n8563), .ZN(n10132) );
  AOI211_X1 U12633 ( .C1(n10134), .C2(n9993), .A(n10133), .B(n10132), .ZN(
        n10135) );
  OAI21_X1 U12634 ( .B1(n12311), .B2(n10136), .A(n10135), .ZN(P3_U3177) );
  XNOR2_X1 U12635 ( .A(n10163), .B(n12560), .ZN(n10146) );
  INV_X1 U12636 ( .A(n10137), .ZN(n10138) );
  NOR2_X1 U12637 ( .A1(n10138), .A2(n6655), .ZN(n10139) );
  XNOR2_X1 U12638 ( .A(n10216), .B(n12153), .ZN(n10142) );
  XNOR2_X1 U12639 ( .A(n10142), .B(n14945), .ZN(n10156) );
  NAND2_X1 U12640 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  NAND2_X1 U12641 ( .A1(n12561), .A2(n10142), .ZN(n10143) );
  INV_X1 U12642 ( .A(n10166), .ZN(n10144) );
  AOI21_X1 U12643 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(n10154) );
  OAI22_X1 U12644 ( .A1(n12288), .A2(n10147), .B1(n14945), .B2(n12291), .ZN(
        n10148) );
  AOI211_X1 U12645 ( .C1(n12294), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        n10153) );
  NAND2_X1 U12646 ( .A1(n12257), .A2(n10151), .ZN(n10152) );
  OAI211_X1 U12647 ( .C1(n10154), .C2(n12311), .A(n10153), .B(n10152), .ZN(
        P3_U3170) );
  OAI211_X1 U12648 ( .C1(n10157), .C2(n10156), .A(n10155), .B(n12280), .ZN(
        n10162) );
  OAI22_X1 U12649 ( .A1(n12288), .A2(n14965), .B1(n10158), .B2(n12291), .ZN(
        n10159) );
  AOI211_X1 U12650 ( .C1(n12294), .C2(n12560), .A(n10160), .B(n10159), .ZN(
        n10161) );
  OAI211_X1 U12651 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12307), .A(n10162), .B(
        n10161), .ZN(P3_U3158) );
  INV_X1 U12652 ( .A(n10163), .ZN(n10164) );
  NAND2_X1 U12653 ( .A1(n10164), .A2(n12350), .ZN(n10165) );
  XNOR2_X1 U12654 ( .A(n14976), .B(n12153), .ZN(n10289) );
  XNOR2_X1 U12655 ( .A(n10289), .B(n10844), .ZN(n10287) );
  XNOR2_X1 U12656 ( .A(n10288), .B(n10287), .ZN(n10167) );
  NAND2_X1 U12657 ( .A1(n10167), .A2(n12280), .ZN(n10172) );
  OAI22_X1 U12658 ( .A1(n12288), .A2(n10168), .B1(n12350), .B2(n12291), .ZN(
        n10169) );
  AOI211_X1 U12659 ( .C1(n12294), .C2(n12559), .A(n10170), .B(n10169), .ZN(
        n10171) );
  OAI211_X1 U12660 ( .C1(n10870), .C2(n12307), .A(n10172), .B(n10171), .ZN(
        P3_U3167) );
  INV_X1 U12661 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11649) );
  NAND2_X1 U12662 ( .A1(n11675), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11687) );
  INV_X1 U12663 ( .A(n11687), .ZN(n10173) );
  NAND2_X1 U12664 ( .A1(n10173), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U12665 ( .A1(n11708), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11707) );
  NAND2_X1 U12666 ( .A1(n11742), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11753) );
  OR2_X1 U12667 ( .A1(n11720), .A2(n11753), .ZN(n10177) );
  NAND2_X1 U12668 ( .A1(n9188), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U12669 ( .A1(n6491), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U12670 ( .A1(n12006), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n10174) );
  NAND4_X1 U12671 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n13804) );
  NAND2_X1 U12672 ( .A1(n13804), .A2(P1_U4016), .ZN(n10178) );
  OAI21_X1 U12673 ( .B1(n8237), .B2(P1_U4016), .A(n10178), .ZN(P1_U3589) );
  INV_X1 U12674 ( .A(n10179), .ZN(n10182) );
  AND3_X1 U12675 ( .A1(n14843), .A2(n14842), .A3(n10180), .ZN(n10181) );
  NAND2_X1 U12676 ( .A1(n10182), .A2(n10181), .ZN(n10189) );
  NOR2_X1 U12677 ( .A1(n10183), .A2(n6754), .ZN(n10184) );
  NAND2_X1 U12678 ( .A1(n13476), .A2(n10184), .ZN(n13462) );
  INV_X1 U12679 ( .A(n13462), .ZN(n10196) );
  INV_X1 U12680 ( .A(n10185), .ZN(n10195) );
  MUX2_X1 U12681 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10186), .S(n13476), .Z(
        n10194) );
  INV_X1 U12682 ( .A(n10187), .ZN(n10188) );
  INV_X1 U12683 ( .A(n10189), .ZN(n10190) );
  INV_X1 U12684 ( .A(n13473), .ZN(n13495) );
  AOI22_X1 U12685 ( .A1(n13507), .A2(n10191), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13495), .ZN(n10192) );
  OAI21_X1 U12686 ( .B1(n9504), .B2(n13498), .A(n10192), .ZN(n10193) );
  AOI211_X1 U12687 ( .C1(n10196), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10197) );
  INV_X1 U12688 ( .A(n10197), .ZN(P2_U3264) );
  INV_X1 U12689 ( .A(n14934), .ZN(n12592) );
  OAI22_X1 U12690 ( .A1(n14916), .A2(n10198), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8549), .ZN(n10206) );
  NAND2_X1 U12691 ( .A1(n14926), .A2(n14928), .ZN(n10201) );
  AND2_X1 U12692 ( .A1(n10201), .A2(n10199), .ZN(n10204) );
  INV_X1 U12693 ( .A(n10199), .ZN(n10200) );
  OAI21_X1 U12694 ( .B1(n12592), .B2(n10201), .A(n10200), .ZN(n10202) );
  NAND2_X1 U12695 ( .A1(n10202), .A2(n14918), .ZN(n10203) );
  MUX2_X1 U12696 ( .A(n10204), .B(n10203), .S(P3_IR_REG_0__SCAN_IN), .Z(n10205) );
  AOI211_X1 U12697 ( .C1(n12592), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10208) );
  INV_X1 U12698 ( .A(n10208), .ZN(P3_U3182) );
  XOR2_X1 U12699 ( .A(n10209), .B(n12502), .Z(n14966) );
  INV_X1 U12700 ( .A(n14993), .ZN(n14997) );
  AOI22_X1 U12701 ( .A1(n12898), .A2(n6655), .B1(n12560), .B2(n12896), .ZN(
        n10213) );
  OAI211_X1 U12702 ( .C1(n7523), .C2(n10211), .A(n14947), .B(n10210), .ZN(
        n10212) );
  OAI211_X1 U12703 ( .C1(n14966), .C2(n14997), .A(n10213), .B(n10212), .ZN(
        n14968) );
  INV_X1 U12704 ( .A(n14968), .ZN(n10221) );
  INV_X1 U12705 ( .A(n14966), .ZN(n10219) );
  INV_X1 U12706 ( .A(n14952), .ZN(n10214) );
  OR2_X1 U12707 ( .A1(n14955), .A2(n10214), .ZN(n12757) );
  INV_X1 U12708 ( .A(n12757), .ZN(n10850) );
  AOI22_X1 U12709 ( .A1(n12889), .A2(n10216), .B1(n12888), .B2(n10215), .ZN(
        n10217) );
  OAI21_X1 U12710 ( .B1(n9704), .B2(n14953), .A(n10217), .ZN(n10218) );
  AOI21_X1 U12711 ( .B1(n10219), .B2(n10850), .A(n10218), .ZN(n10220) );
  OAI21_X1 U12712 ( .B1(n10221), .B2(n14955), .A(n10220), .ZN(P3_U3230) );
  NOR2_X1 U12713 ( .A1(n10222), .A2(n12102), .ZN(n10224) );
  NAND2_X1 U12714 ( .A1(n10224), .A2(n10223), .ZN(n11757) );
  NAND2_X1 U12715 ( .A1(n11835), .A2(n11845), .ZN(n12035) );
  INV_X1 U12716 ( .A(n12035), .ZN(n10227) );
  AND2_X1 U12717 ( .A1(n14671), .A2(n10227), .ZN(n14655) );
  AOI21_X1 U12718 ( .B1(n14723), .B2(n14671), .A(n14655), .ZN(n14141) );
  AND2_X1 U12719 ( .A1(n14658), .A2(n12036), .ZN(n10228) );
  INV_X1 U12720 ( .A(n14662), .ZN(n14645) );
  AOI22_X1 U12721 ( .A1(n14646), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14645), .ZN(n10229) );
  OAI21_X1 U12722 ( .B1(n14175), .B2(n11848), .A(n10229), .ZN(n10232) );
  NOR2_X1 U12723 ( .A1(n10230), .A2(n14646), .ZN(n10231) );
  AOI211_X1 U12724 ( .C1(n10233), .C2(n14654), .A(n10232), .B(n10231), .ZN(
        n10234) );
  OAI21_X1 U12725 ( .B1(n14141), .B2(n10235), .A(n10234), .ZN(P1_U3291) );
  NOR2_X1 U12726 ( .A1(n14175), .A2(n10236), .ZN(n10239) );
  OAI22_X1 U12727 ( .A1(n14671), .A2(n10237), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14662), .ZN(n10238) );
  AOI211_X1 U12728 ( .C1(n10240), .C2(n14654), .A(n10239), .B(n10238), .ZN(
        n10243) );
  NAND2_X1 U12729 ( .A1(n10241), .A2(n14655), .ZN(n10242) );
  OAI211_X1 U12730 ( .C1(n10244), .C2(n14646), .A(n10243), .B(n10242), .ZN(
        P1_U3290) );
  INV_X1 U12731 ( .A(n14878), .ZN(n10436) );
  INV_X1 U12732 ( .A(n10245), .ZN(n10247) );
  NAND2_X1 U12733 ( .A1(n10247), .A2(n10246), .ZN(n10248) );
  XNOR2_X1 U12734 ( .A(n10567), .B(n11612), .ZN(n10250) );
  AND2_X1 U12735 ( .A1(n10911), .A2(n13208), .ZN(n10251) );
  NAND2_X1 U12736 ( .A1(n10250), .A2(n10251), .ZN(n10253) );
  NAND2_X1 U12737 ( .A1(n10253), .A2(n10252), .ZN(n10389) );
  XNOR2_X1 U12738 ( .A(n14878), .B(n11612), .ZN(n10254) );
  AND2_X1 U12739 ( .A1(n13492), .A2(n13207), .ZN(n10255) );
  NAND2_X1 U12740 ( .A1(n10254), .A2(n10255), .ZN(n10671) );
  INV_X1 U12741 ( .A(n10254), .ZN(n10257) );
  INV_X1 U12742 ( .A(n10255), .ZN(n10256) );
  NAND2_X1 U12743 ( .A1(n10257), .A2(n10256), .ZN(n10258) );
  AND2_X1 U12744 ( .A1(n10671), .A2(n10258), .ZN(n10259) );
  OAI211_X1 U12745 ( .C1(n10260), .C2(n10259), .A(n10672), .B(n13162), .ZN(
        n10264) );
  INV_X1 U12746 ( .A(n13206), .ZN(n10684) );
  OAI22_X1 U12747 ( .A1(n10427), .A2(n13139), .B1(n13138), .B2(n10684), .ZN(
        n10261) );
  AOI211_X1 U12748 ( .C1(n13151), .C2(n10434), .A(n10262), .B(n10261), .ZN(
        n10263) );
  OAI211_X1 U12749 ( .C1(n10436), .C2(n13154), .A(n10264), .B(n10263), .ZN(
        P2_U3185) );
  OR2_X1 U12750 ( .A1(n13210), .A2(n10336), .ZN(n10265) );
  INV_X1 U12751 ( .A(n10272), .ZN(n10267) );
  OR2_X1 U12752 ( .A1(n10268), .A2(n10267), .ZN(n10269) );
  AND2_X1 U12753 ( .A1(n10421), .A2(n10269), .ZN(n14872) );
  NAND2_X1 U12754 ( .A1(n10336), .A2(n10274), .ZN(n10270) );
  NAND2_X1 U12755 ( .A1(n10273), .A2(n10272), .ZN(n10426) );
  OAI21_X1 U12756 ( .B1(n10273), .B2(n10272), .A(n10426), .ZN(n10277) );
  OAI22_X1 U12757 ( .A1(n10274), .A2(n13445), .B1(n10427), .B2(n13447), .ZN(
        n10276) );
  NOR2_X1 U12758 ( .A1(n14872), .A2(n14849), .ZN(n10275) );
  AOI211_X1 U12759 ( .C1(n13488), .C2(n10277), .A(n10276), .B(n10275), .ZN(
        n14870) );
  MUX2_X1 U12760 ( .A(n10278), .B(n14870), .S(n13476), .Z(n10286) );
  NAND2_X1 U12761 ( .A1(n13495), .A2(n10279), .ZN(n10283) );
  AOI21_X1 U12762 ( .B1(n10280), .B2(n14868), .A(n13492), .ZN(n10281) );
  AND2_X1 U12763 ( .A1(n10281), .A2(n10532), .ZN(n14867) );
  NAND2_X1 U12764 ( .A1(n13507), .A2(n14867), .ZN(n10282) );
  OAI211_X1 U12765 ( .C1(n13498), .C2(n6997), .A(n10283), .B(n10282), .ZN(
        n10284) );
  INV_X1 U12766 ( .A(n10284), .ZN(n10285) );
  OAI211_X1 U12767 ( .C1(n14872), .C2(n13462), .A(n10286), .B(n10285), .ZN(
        P2_U3260) );
  INV_X1 U12768 ( .A(n10289), .ZN(n10290) );
  NAND2_X1 U12769 ( .A1(n10290), .A2(n10844), .ZN(n10291) );
  NAND2_X1 U12770 ( .A1(n10292), .A2(n10291), .ZN(n10295) );
  XNOR2_X1 U12771 ( .A(n10293), .B(n12194), .ZN(n10556) );
  XNOR2_X1 U12772 ( .A(n10556), .B(n10779), .ZN(n10294) );
  AOI21_X1 U12773 ( .B1(n10295), .B2(n10294), .A(n12311), .ZN(n10296) );
  NAND2_X1 U12774 ( .A1(n10296), .A2(n10559), .ZN(n10300) );
  OAI22_X1 U12775 ( .A1(n12288), .A2(n14983), .B1(n10844), .B2(n12291), .ZN(
        n10297) );
  AOI211_X1 U12776 ( .C1(n12294), .C2(n12558), .A(n10298), .B(n10297), .ZN(
        n10299) );
  OAI211_X1 U12777 ( .C1(n10840), .C2(n12307), .A(n10300), .B(n10299), .ZN(
        P3_U3179) );
  NAND2_X1 U12778 ( .A1(n10301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10302) );
  MUX2_X1 U12779 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10302), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10303) );
  AND2_X1 U12780 ( .A1(n10303), .A2(n10805), .ZN(n14033) );
  INV_X1 U12781 ( .A(n14033), .ZN(n14609) );
  INV_X1 U12782 ( .A(n11634), .ZN(n10305) );
  OAI222_X1 U12783 ( .A1(P1_U3086), .A2(n14609), .B1(n14382), .B2(n10305), 
        .C1(n10304), .C2(n14379), .ZN(P1_U3338) );
  OAI222_X1 U12784 ( .A1(n13636), .A2(n10306), .B1(n13637), .B2(n10305), .C1(
        n14823), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U12785 ( .A(n10307), .ZN(n10314) );
  MUX2_X1 U12786 ( .A(n10309), .B(n10308), .S(n12623), .Z(n10310) );
  NAND2_X1 U12787 ( .A1(n10310), .A2(n10491), .ZN(n10483) );
  INV_X1 U12788 ( .A(n10310), .ZN(n10311) );
  NAND2_X1 U12789 ( .A1(n10311), .A2(n14399), .ZN(n10312) );
  AND2_X1 U12790 ( .A1(n10483), .A2(n10312), .ZN(n10313) );
  OAI21_X1 U12791 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(n10484) );
  INV_X1 U12792 ( .A(n10484), .ZN(n10317) );
  NOR3_X1 U12793 ( .A1(n10315), .A2(n10314), .A3(n10313), .ZN(n10316) );
  OAI21_X1 U12794 ( .B1(n10317), .B2(n10316), .A(n12703), .ZN(n10320) );
  NOR2_X1 U12795 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10318), .ZN(n10945) );
  AOI21_X1 U12796 ( .B1(n14896), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10945), .ZN(
        n10319) );
  OAI211_X1 U12797 ( .C1(n14918), .C2(n14399), .A(n10320), .B(n10319), .ZN(
        n10330) );
  AND2_X2 U12798 ( .A1(n10322), .A2(n10321), .ZN(n10490) );
  AOI21_X1 U12799 ( .B1(n10309), .B2(n10323), .A(n10492), .ZN(n10328) );
  AOI21_X1 U12800 ( .B1(n10308), .B2(n10326), .A(n10473), .ZN(n10327) );
  OAI22_X1 U12801 ( .A1(n10328), .A2(n14934), .B1(n10327), .B2(n14926), .ZN(
        n10329) );
  OR2_X1 U12802 ( .A1(n10330), .A2(n10329), .ZN(P3_U3191) );
  INV_X1 U12803 ( .A(n10331), .ZN(n10332) );
  MUX2_X1 U12804 ( .A(n9353), .B(n10332), .S(n13476), .Z(n10338) );
  INV_X1 U12805 ( .A(n13507), .ZN(n13371) );
  OAI22_X1 U12806 ( .A1(n13371), .A2(n10334), .B1(n10333), .B2(n13473), .ZN(
        n10335) );
  AOI21_X1 U12807 ( .B1(n13483), .B2(n10336), .A(n10335), .ZN(n10337) );
  OAI211_X1 U12808 ( .C1(n10339), .C2(n13462), .A(n10338), .B(n10337), .ZN(
        P2_U3261) );
  INV_X1 U12809 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U12810 ( .A1(n12746), .A2(P3_U3897), .ZN(n10340) );
  OAI21_X1 U12811 ( .B1(P3_U3897), .B2(n15066), .A(n10340), .ZN(P3_U3518) );
  INV_X1 U12812 ( .A(n14849), .ZN(n13456) );
  OAI211_X2 U12813 ( .C1(n11500), .C2(n13456), .A(n13476), .B(n11612), .ZN(
        n13504) );
  NOR2_X1 U12814 ( .A1(n13371), .A2(n13492), .ZN(n13442) );
  OAI21_X1 U12815 ( .B1(n13442), .B2(n13483), .A(n10377), .ZN(n10344) );
  INV_X1 U12816 ( .A(n14850), .ZN(n14854) );
  AOI22_X1 U12817 ( .A1(n14854), .A2(n13488), .B1(n13437), .B2(n6748), .ZN(
        n14851) );
  INV_X1 U12818 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10341) );
  OAI22_X1 U12819 ( .A1(n13392), .A2(n14851), .B1(n10341), .B2(n13473), .ZN(
        n10342) );
  AOI21_X1 U12820 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13509), .A(n10342), .ZN(
        n10343) );
  OAI211_X1 U12821 ( .C1(n14850), .C2(n13504), .A(n10344), .B(n10343), .ZN(
        P2_U3265) );
  NAND2_X1 U12822 ( .A1(n10345), .A2(P2_U3947), .ZN(n10346) );
  OAI21_X1 U12823 ( .B1(n11622), .B2(P2_U3947), .A(n10346), .ZN(P2_U3560) );
  AOI21_X1 U12824 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10878), .A(n10347), 
        .ZN(n10350) );
  INV_X1 U12825 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10348) );
  MUX2_X1 U12826 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10348), .S(n11034), .Z(
        n10349) );
  NAND2_X1 U12827 ( .A1(n10350), .A2(n10349), .ZN(n10546) );
  OAI21_X1 U12828 ( .B1(n10350), .B2(n10349), .A(n10546), .ZN(n10358) );
  NAND2_X1 U12829 ( .A1(n14625), .A2(n11034), .ZN(n10351) );
  NAND2_X1 U12830 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14508)
         );
  OAI211_X1 U12831 ( .C1(n10352), .C2(n14633), .A(n10351), .B(n14508), .ZN(
        n10357) );
  XNOR2_X1 U12832 ( .A(n11034), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n10354) );
  NOR2_X1 U12833 ( .A1(n10355), .A2(n10354), .ZN(n10539) );
  AOI211_X1 U12834 ( .C1(n10355), .C2(n10354), .A(n14566), .B(n10539), .ZN(
        n10356) );
  AOI211_X1 U12835 ( .C1(n14617), .C2(n10358), .A(n10357), .B(n10356), .ZN(
        n10359) );
  INV_X1 U12836 ( .A(n10359), .ZN(P1_U3254) );
  NAND2_X1 U12837 ( .A1(n13946), .A2(n6487), .ZN(n10361) );
  NAND2_X1 U12838 ( .A1(n11862), .A2(n13800), .ZN(n10360) );
  NAND2_X1 U12839 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  XNOR2_X1 U12840 ( .A(n10362), .B(n13798), .ZN(n10440) );
  INV_X1 U12841 ( .A(n10363), .ZN(n10365) );
  NAND2_X1 U12842 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  AOI22_X1 U12843 ( .A1(n13946), .A2(n13764), .B1(n11862), .B2(n6487), .ZN(
        n10442) );
  XNOR2_X1 U12844 ( .A(n10444), .B(n10442), .ZN(n10441) );
  XOR2_X1 U12845 ( .A(n10440), .B(n10441), .Z(n10373) );
  INV_X1 U12846 ( .A(n10579), .ZN(n10371) );
  AND2_X1 U12847 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13995) );
  AOI21_X1 U12848 ( .B1(n10368), .B2(n14506), .A(n13995), .ZN(n10370) );
  NAND2_X1 U12849 ( .A1(n14502), .A2(n11862), .ZN(n10369) );
  OAI211_X1 U12850 ( .C1(n14511), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10372) );
  AOI21_X1 U12851 ( .B1(n10373), .B2(n14504), .A(n10372), .ZN(n10374) );
  INV_X1 U12852 ( .A(n10374), .ZN(P1_U3230) );
  INV_X1 U12853 ( .A(n10376), .ZN(n10375) );
  NAND2_X1 U12854 ( .A1(n13162), .A2(n10375), .ZN(n10379) );
  AOI21_X1 U12855 ( .B1(n13162), .B2(n10376), .A(n13185), .ZN(n10378) );
  MUX2_X1 U12856 ( .A(n10379), .B(n10378), .S(n10377), .Z(n10382) );
  OR2_X1 U12857 ( .A1(n10380), .A2(P2_U3088), .ZN(n13157) );
  NAND2_X1 U12858 ( .A1(n13157), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10381) );
  OAI211_X1 U12859 ( .C1(n9622), .C2(n13138), .A(n10382), .B(n10381), .ZN(
        P2_U3204) );
  INV_X1 U12860 ( .A(n10383), .ZN(n10385) );
  OAI222_X1 U12861 ( .A1(n10386), .A2(P3_U3151), .B1(n13057), .B2(n10385), 
        .C1(n10384), .C2(n13054), .ZN(P3_U3275) );
  NAND2_X1 U12862 ( .A1(n12562), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10387) );
  OAI21_X1 U12863 ( .B1(n12720), .B2(n12562), .A(n10387), .ZN(P3_U3520) );
  AOI211_X1 U12864 ( .C1(n10389), .C2(n10388), .A(n13187), .B(n6629), .ZN(
        n10394) );
  INV_X1 U12865 ( .A(n10567), .ZN(n10535) );
  OAI22_X1 U12866 ( .A1(n10535), .A2(n13154), .B1(n13138), .B2(n10597), .ZN(
        n10393) );
  NAND2_X1 U12867 ( .A1(n13151), .A2(n10533), .ZN(n10390) );
  OAI211_X1 U12868 ( .C1(n13139), .C2(n10527), .A(n10391), .B(n10390), .ZN(
        n10392) );
  OR3_X1 U12869 ( .A1(n10394), .A2(n10393), .A3(n10392), .ZN(P2_U3211) );
  INV_X1 U12870 ( .A(n13504), .ZN(n13387) );
  AOI22_X1 U12871 ( .A1(n13507), .A2(n10395), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13495), .ZN(n10396) );
  OAI21_X1 U12872 ( .B1(n10397), .B2(n13498), .A(n10396), .ZN(n10398) );
  AOI21_X1 U12873 ( .B1(n13387), .B2(n10399), .A(n10398), .ZN(n10402) );
  MUX2_X1 U12874 ( .A(n9349), .B(n10400), .S(n13476), .Z(n10401) );
  NAND2_X1 U12875 ( .A1(n10402), .A2(n10401), .ZN(P2_U3263) );
  OAI21_X1 U12876 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(n14864) );
  NAND2_X1 U12877 ( .A1(n10407), .A2(n10406), .ZN(n10408) );
  NAND2_X1 U12878 ( .A1(n10408), .A2(n10055), .ZN(n10409) );
  NOR2_X1 U12879 ( .A1(n10410), .A2(n10409), .ZN(n14857) );
  AOI22_X1 U12880 ( .A1(n13507), .A2(n14857), .B1(n13495), .B2(n10411), .ZN(
        n10412) );
  OAI21_X1 U12881 ( .B1(n14860), .B2(n13498), .A(n10412), .ZN(n10413) );
  AOI21_X1 U12882 ( .B1(n13387), .B2(n14864), .A(n10413), .ZN(n10419) );
  OAI21_X1 U12883 ( .B1(n10416), .B2(n10415), .A(n10414), .ZN(n10417) );
  AOI222_X1 U12884 ( .A1(n13488), .A2(n10417), .B1(n13210), .B2(n13437), .C1(
        n13212), .C2(n13435), .ZN(n14861) );
  MUX2_X1 U12885 ( .A(n9350), .B(n14861), .S(n13476), .Z(n10418) );
  NAND2_X1 U12886 ( .A1(n10419), .A2(n10418), .ZN(P2_U3262) );
  OR2_X1 U12887 ( .A1(n14868), .A2(n13209), .ZN(n10420) );
  INV_X1 U12888 ( .A(n10525), .ZN(n10521) );
  OR2_X1 U12889 ( .A1(n10567), .A2(n13208), .ZN(n10422) );
  OR2_X1 U12890 ( .A1(n10423), .A2(n10429), .ZN(n10424) );
  AND2_X1 U12891 ( .A1(n10590), .A2(n10424), .ZN(n14876) );
  NAND2_X1 U12892 ( .A1(n14868), .A2(n10527), .ZN(n10425) );
  NAND2_X1 U12893 ( .A1(n10426), .A2(n10425), .ZN(n10526) );
  NAND2_X1 U12894 ( .A1(n10567), .A2(n10427), .ZN(n10428) );
  XNOR2_X1 U12895 ( .A(n10596), .B(n7443), .ZN(n10430) );
  NAND2_X1 U12896 ( .A1(n10430), .A2(n13488), .ZN(n10432) );
  AOI22_X1 U12897 ( .A1(n13435), .A2(n13208), .B1(n13206), .B2(n13437), .ZN(
        n10431) );
  AND2_X1 U12898 ( .A1(n10432), .A2(n10431), .ZN(n14882) );
  MUX2_X1 U12899 ( .A(n15159), .B(n14882), .S(n13476), .Z(n10439) );
  OAI21_X1 U12900 ( .B1(n10531), .B2(n10436), .A(n10055), .ZN(n10433) );
  NOR2_X1 U12901 ( .A1(n10433), .A2(n10592), .ZN(n14880) );
  INV_X1 U12902 ( .A(n10434), .ZN(n10435) );
  OAI22_X1 U12903 ( .A1(n13498), .A2(n10436), .B1(n13473), .B2(n10435), .ZN(
        n10437) );
  AOI21_X1 U12904 ( .B1(n13507), .B2(n14880), .A(n10437), .ZN(n10438) );
  OAI211_X1 U12905 ( .C1(n14876), .C2(n13504), .A(n10439), .B(n10438), .ZN(
        P2_U3258) );
  INV_X1 U12906 ( .A(n10442), .ZN(n10443) );
  NAND2_X1 U12907 ( .A1(n10447), .A2(n12025), .ZN(n10450) );
  AOI22_X1 U12908 ( .A1(n11646), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11645), 
        .B2(n10448), .ZN(n10449) );
  OAI22_X1 U12909 ( .A1(n11865), .A2(n13682), .B1(n11866), .B2(n13690), .ZN(
        n10451) );
  XNOR2_X1 U12910 ( .A(n10451), .B(n13798), .ZN(n10454) );
  INV_X1 U12911 ( .A(n10452), .ZN(n13689) );
  OAI22_X1 U12912 ( .A1(n11865), .A2(n13690), .B1(n11866), .B2(n13689), .ZN(
        n10453) );
  OR2_X1 U12913 ( .A1(n10454), .A2(n10453), .ZN(n10658) );
  NAND2_X1 U12914 ( .A1(n10454), .A2(n10453), .ZN(n10660) );
  NAND2_X1 U12915 ( .A1(n10658), .A2(n10660), .ZN(n10455) );
  XNOR2_X1 U12916 ( .A(n10659), .B(n10455), .ZN(n10470) );
  INV_X1 U12917 ( .A(n10456), .ZN(n10515) );
  NAND2_X1 U12918 ( .A1(n13946), .A2(n13899), .ZN(n10464) );
  NAND2_X1 U12919 ( .A1(n11653), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12920 ( .A1(n6491), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10461) );
  NOR2_X1 U12921 ( .A1(n10457), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10458) );
  NOR2_X1 U12922 ( .A1(n10632), .A2(n10458), .ZN(n14644) );
  NAND2_X1 U12923 ( .A1(n11743), .A2(n14644), .ZN(n10460) );
  NAND2_X1 U12924 ( .A1(n11039), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U12925 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n13944) );
  NAND2_X1 U12926 ( .A1(n13944), .A2(n13898), .ZN(n10463) );
  NAND2_X1 U12927 ( .A1(n10464), .A2(n10463), .ZN(n10511) );
  INV_X1 U12928 ( .A(n10465), .ZN(n10466) );
  AOI21_X1 U12929 ( .B1(n10511), .B2(n14506), .A(n10466), .ZN(n10468) );
  INV_X1 U12930 ( .A(n11865), .ZN(n14690) );
  NAND2_X1 U12931 ( .A1(n14502), .A2(n14690), .ZN(n10467) );
  OAI211_X1 U12932 ( .C1(n14511), .C2(n10515), .A(n10468), .B(n10467), .ZN(
        n10469) );
  AOI21_X1 U12933 ( .B1(n10470), .B2(n14504), .A(n10469), .ZN(n10471) );
  INV_X1 U12934 ( .A(n10471), .ZN(P1_U3227) );
  NAND2_X1 U12935 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11186), .ZN(n10474) );
  OAI21_X1 U12936 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11186), .A(n10474), 
        .ZN(n10475) );
  AOI21_X1 U12937 ( .B1(n10476), .B2(n10475), .A(n11172), .ZN(n10499) );
  INV_X1 U12938 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n10477) );
  NAND2_X1 U12939 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n11083)
         );
  OAI21_X1 U12940 ( .B1(n14916), .B2(n10477), .A(n11083), .ZN(n10488) );
  MUX2_X1 U12941 ( .A(n11025), .B(n10478), .S(n12623), .Z(n10479) );
  NAND2_X1 U12942 ( .A1(n10479), .A2(n10489), .ZN(n11179) );
  INV_X1 U12943 ( .A(n10479), .ZN(n10480) );
  NAND2_X1 U12944 ( .A1(n10480), .A2(n11186), .ZN(n10481) );
  NAND2_X1 U12945 ( .A1(n11179), .A2(n10481), .ZN(n10482) );
  AOI21_X1 U12946 ( .B1(n10484), .B2(n10483), .A(n10482), .ZN(n11181) );
  INV_X1 U12947 ( .A(n11181), .ZN(n10486) );
  NAND3_X1 U12948 ( .A1(n10484), .A2(n10483), .A3(n10482), .ZN(n10485) );
  AOI21_X1 U12949 ( .B1(n10486), .B2(n10485), .A(n14928), .ZN(n10487) );
  AOI211_X1 U12950 ( .C1(n12669), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10498) );
  NAND2_X1 U12951 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11186), .ZN(n10494) );
  OAI21_X1 U12952 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11186), .A(n10494), 
        .ZN(n10495) );
  OR2_X1 U12953 ( .A1(n10496), .A2(n14934), .ZN(n10497) );
  OAI211_X1 U12954 ( .C1(n10499), .C2(n14926), .A(n10498), .B(n10497), .ZN(
        P3_U3192) );
  NAND2_X1 U12955 ( .A1(n13946), .A2(n11862), .ZN(n10500) );
  NAND2_X1 U12956 ( .A1(n10501), .A2(n10500), .ZN(n10503) );
  OR2_X1 U12957 ( .A1(n13946), .A2(n11862), .ZN(n10502) );
  NAND2_X1 U12958 ( .A1(n10503), .A2(n10502), .ZN(n10618) );
  INV_X1 U12959 ( .A(n11866), .ZN(n13945) );
  NAND2_X1 U12960 ( .A1(n11865), .A2(n13945), .ZN(n10504) );
  NAND2_X1 U12961 ( .A1(n14690), .A2(n11866), .ZN(n10637) );
  NAND2_X1 U12962 ( .A1(n10504), .A2(n10637), .ZN(n12066) );
  INV_X1 U12963 ( .A(n12066), .ZN(n10509) );
  XNOR2_X1 U12964 ( .A(n10618), .B(n10509), .ZN(n14694) );
  INV_X1 U12965 ( .A(n14655), .ZN(n10519) );
  OR2_X1 U12966 ( .A1(n13946), .A2(n10581), .ZN(n10506) );
  AND2_X1 U12967 ( .A1(n10581), .A2(n13946), .ZN(n10505) );
  NAND2_X1 U12968 ( .A1(n10508), .A2(n10509), .ZN(n10638) );
  OAI21_X1 U12969 ( .B1(n10509), .B2(n10508), .A(n10638), .ZN(n10512) );
  NOR2_X1 U12970 ( .A1(n14694), .A2(n14707), .ZN(n10510) );
  AOI211_X1 U12971 ( .C1(n14643), .C2(n10512), .A(n10511), .B(n10510), .ZN(
        n14693) );
  MUX2_X1 U12972 ( .A(n9217), .B(n14693), .S(n14671), .Z(n10518) );
  INV_X1 U12973 ( .A(n10513), .ZN(n10514) );
  INV_X1 U12974 ( .A(n10649), .ZN(n14652) );
  AOI211_X1 U12975 ( .C1(n14690), .C2(n10514), .A(n14683), .B(n14652), .ZN(
        n14689) );
  OAI22_X1 U12976 ( .A1(n14175), .A2(n11865), .B1(n10515), .B2(n14662), .ZN(
        n10516) );
  AOI21_X1 U12977 ( .B1(n14689), .B2(n14654), .A(n10516), .ZN(n10517) );
  OAI211_X1 U12978 ( .C1(n14694), .C2(n10519), .A(n10518), .B(n10517), .ZN(
        P1_U3288) );
  OAI21_X1 U12979 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(n10523) );
  INV_X1 U12980 ( .A(n10523), .ZN(n10570) );
  OAI21_X1 U12981 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(n10530) );
  OAI22_X1 U12982 ( .A1(n10527), .A2(n13445), .B1(n10597), .B2(n13447), .ZN(
        n10529) );
  NOR2_X1 U12983 ( .A1(n10570), .A2(n14849), .ZN(n10528) );
  AOI211_X1 U12984 ( .C1(n13488), .C2(n10530), .A(n10529), .B(n10528), .ZN(
        n10569) );
  MUX2_X1 U12985 ( .A(n9356), .B(n10569), .S(n13476), .Z(n10538) );
  AOI211_X1 U12986 ( .C1(n10567), .C2(n10532), .A(n13492), .B(n10531), .ZN(
        n10566) );
  INV_X1 U12987 ( .A(n10533), .ZN(n10534) );
  OAI22_X1 U12988 ( .A1(n13498), .A2(n10535), .B1(n13473), .B2(n10534), .ZN(
        n10536) );
  AOI21_X1 U12989 ( .B1(n10566), .B2(n13507), .A(n10536), .ZN(n10537) );
  OAI211_X1 U12990 ( .C1(n10570), .C2(n13462), .A(n10538), .B(n10537), .ZN(
        P2_U3259) );
  INV_X1 U12991 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10540) );
  MUX2_X1 U12992 ( .A(n10540), .B(P1_REG2_REG_12__SCAN_IN), .S(n14025), .Z(
        n10541) );
  INV_X1 U12993 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U12994 ( .A1(n10543), .A2(n10542), .ZN(n14013) );
  OAI21_X1 U12995 ( .B1(n10543), .B2(n10542), .A(n14013), .ZN(n10544) );
  INV_X1 U12996 ( .A(n14566), .ZN(n14620) );
  NAND2_X1 U12997 ( .A1(n10544), .A2(n14620), .ZN(n10555) );
  INV_X1 U12998 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U12999 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10545), .S(n14025), .Z(
        n10548) );
  OAI21_X1 U13000 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11034), .A(n10546), 
        .ZN(n10547) );
  NAND2_X1 U13001 ( .A1(n10547), .A2(n10548), .ZN(n14024) );
  OAI21_X1 U13002 ( .B1(n10548), .B2(n10547), .A(n14024), .ZN(n10553) );
  INV_X1 U13003 ( .A(n14625), .ZN(n14610) );
  NAND2_X1 U13004 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11476)
         );
  NAND2_X1 U13005 ( .A1(n10549), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10550) );
  OAI211_X1 U13006 ( .C1(n14610), .C2(n10551), .A(n11476), .B(n10550), .ZN(
        n10552) );
  AOI21_X1 U13007 ( .B1(n10553), .B2(n14617), .A(n10552), .ZN(n10554) );
  NAND2_X1 U13008 ( .A1(n10555), .A2(n10554), .ZN(P1_U3255) );
  INV_X1 U13009 ( .A(n10556), .ZN(n10557) );
  NAND2_X1 U13010 ( .A1(n12559), .A2(n10557), .ZN(n10558) );
  NAND2_X1 U13011 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  XNOR2_X1 U13012 ( .A(n10777), .B(n12153), .ZN(n10765) );
  OAI211_X1 U13013 ( .C1(n10560), .C2(n10765), .A(n10768), .B(n12280), .ZN(
        n10565) );
  OAI22_X1 U13014 ( .A1(n12288), .A2(n10561), .B1(n10779), .B2(n12291), .ZN(
        n10562) );
  AOI211_X1 U13015 ( .C1(n12294), .C2(n12557), .A(n10563), .B(n10562), .ZN(
        n10564) );
  OAI211_X1 U13016 ( .C1(n10784), .C2(n12307), .A(n10565), .B(n10564), .ZN(
        P3_U3153) );
  INV_X1 U13017 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10572) );
  AOI21_X1 U13018 ( .B1(n14877), .B2(n10567), .A(n10566), .ZN(n10568) );
  OAI211_X1 U13019 ( .C1(n10570), .C2(n14871), .A(n10569), .B(n10568), .ZN(
        n10573) );
  NAND2_X1 U13020 ( .A1(n10573), .A2(n14886), .ZN(n10571) );
  OAI21_X1 U13021 ( .B1(n14886), .B2(n10572), .A(n10571), .ZN(P2_U3448) );
  NAND2_X1 U13022 ( .A1(n10573), .A2(n14895), .ZN(n10574) );
  OAI21_X1 U13023 ( .B1(n14895), .B2(n10575), .A(n10574), .ZN(P2_U3505) );
  INV_X1 U13024 ( .A(SI_21_), .ZN(n10578) );
  INV_X1 U13025 ( .A(n10576), .ZN(n10577) );
  OAI222_X1 U13026 ( .A1(n12332), .A2(P3_U3151), .B1(n13054), .B2(n10578), 
        .C1(n13057), .C2(n10577), .ZN(P3_U3274) );
  AOI22_X1 U13027 ( .A1(n14646), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10579), 
        .B2(n14645), .ZN(n10580) );
  OAI21_X1 U13028 ( .B1(n14175), .B2(n10581), .A(n10580), .ZN(n10585) );
  NAND2_X1 U13029 ( .A1(n14671), .A2(n10582), .ZN(n14256) );
  NOR2_X1 U13030 ( .A1(n10583), .A2(n14256), .ZN(n10584) );
  AOI211_X1 U13031 ( .C1(n10586), .C2(n14654), .A(n10585), .B(n10584), .ZN(
        n10587) );
  OAI21_X1 U13032 ( .B1(n14646), .B2(n10588), .A(n10587), .ZN(P1_U3289) );
  OR2_X1 U13033 ( .A1(n14878), .A2(n13207), .ZN(n10589) );
  AOI21_X1 U13034 ( .B1(n7118), .B2(n10591), .A(n6630), .ZN(n10612) );
  INV_X1 U13035 ( .A(n6727), .ZN(n10610) );
  NAND2_X1 U13036 ( .A1(n10592), .A2(n10610), .ZN(n10694) );
  OAI211_X1 U13037 ( .C1(n10592), .C2(n10610), .A(n10055), .B(n10694), .ZN(
        n10608) );
  AOI22_X1 U13038 ( .A1(n13509), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10677), 
        .B2(n13495), .ZN(n10594) );
  OR2_X1 U13039 ( .A1(n13498), .A2(n10610), .ZN(n10593) );
  OAI211_X1 U13040 ( .C1(n10608), .C2(n13371), .A(n10594), .B(n10593), .ZN(
        n10606) );
  OR2_X1 U13041 ( .A1(n14878), .A2(n10597), .ZN(n10595) );
  NAND2_X1 U13042 ( .A1(n14878), .A2(n10597), .ZN(n10598) );
  INV_X1 U13043 ( .A(n13488), .ZN(n13451) );
  AOI21_X1 U13044 ( .B1(n10600), .B2(n6481), .A(n13451), .ZN(n10604) );
  NAND2_X1 U13045 ( .A1(n13435), .A2(n13207), .ZN(n10602) );
  NAND2_X1 U13046 ( .A1(n13205), .A2(n13437), .ZN(n10601) );
  AND2_X1 U13047 ( .A1(n10602), .A2(n10601), .ZN(n10680) );
  INV_X1 U13048 ( .A(n10680), .ZN(n10603) );
  AOI21_X1 U13049 ( .B1(n10604), .B2(n10687), .A(n10603), .ZN(n10609) );
  NOR2_X1 U13050 ( .A1(n10609), .A2(n13509), .ZN(n10605) );
  AOI211_X1 U13051 ( .C1(n10612), .C2(n13387), .A(n10606), .B(n10605), .ZN(
        n10607) );
  INV_X1 U13052 ( .A(n10607), .ZN(P2_U3257) );
  INV_X1 U13053 ( .A(n14875), .ZN(n14865) );
  OAI211_X1 U13054 ( .C1(n10610), .C2(n14859), .A(n10609), .B(n10608), .ZN(
        n10611) );
  AOI21_X1 U13055 ( .B1(n10612), .B2(n14865), .A(n10611), .ZN(n10617) );
  INV_X1 U13056 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10613) );
  OR2_X1 U13057 ( .A1(n14886), .A2(n10613), .ZN(n10614) );
  OAI21_X1 U13058 ( .B1(n10617), .B2(n14884), .A(n10614), .ZN(P2_U3454) );
  OR2_X1 U13059 ( .A1(n14895), .A2(n10615), .ZN(n10616) );
  OAI21_X1 U13060 ( .B1(n10617), .B2(n14893), .A(n10616), .ZN(P2_U3507) );
  NAND2_X1 U13061 ( .A1(n10618), .A2(n12066), .ZN(n10620) );
  NAND2_X1 U13062 ( .A1(n11865), .A2(n11866), .ZN(n10619) );
  NAND2_X1 U13063 ( .A1(n10621), .A2(n12025), .ZN(n10624) );
  AOI22_X1 U13064 ( .A1(n11646), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11645), 
        .B2(n10622), .ZN(n10623) );
  NAND2_X1 U13065 ( .A1(n10624), .A2(n10623), .ZN(n14648) );
  XNOR2_X1 U13066 ( .A(n14648), .B(n13944), .ZN(n14638) );
  INV_X1 U13067 ( .A(n14638), .ZN(n10625) );
  NAND2_X1 U13068 ( .A1(n14639), .A2(n10625), .ZN(n10627) );
  OR2_X1 U13069 ( .A1(n14648), .A2(n13944), .ZN(n10626) );
  NAND2_X1 U13070 ( .A1(n10627), .A2(n10626), .ZN(n10706) );
  NAND2_X1 U13071 ( .A1(n10628), .A2(n12025), .ZN(n10631) );
  AOI22_X1 U13072 ( .A1(n11646), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11645), 
        .B2(n10629), .ZN(n10630) );
  NAND2_X1 U13073 ( .A1(n10631), .A2(n10630), .ZN(n11875) );
  OAI21_X1 U13074 ( .B1(n10632), .B2(P1_REG3_REG_7__SCAN_IN), .A(n10641), .ZN(
        n10798) );
  OR2_X1 U13075 ( .A1(n11720), .A2(n10798), .ZN(n10636) );
  NAND2_X1 U13076 ( .A1(n6491), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13077 ( .A1(n12006), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10634) );
  NAND2_X1 U13078 ( .A1(n11039), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10633) );
  NAND4_X1 U13079 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n13943) );
  XNOR2_X1 U13080 ( .A(n11875), .B(n13943), .ZN(n12068) );
  XNOR2_X1 U13081 ( .A(n10706), .B(n12068), .ZN(n14706) );
  NAND2_X1 U13082 ( .A1(n10638), .A2(n10637), .ZN(n14636) );
  NAND2_X1 U13083 ( .A1(n14636), .A2(n14638), .ZN(n14635) );
  INV_X1 U13084 ( .A(n13944), .ZN(n10639) );
  NAND2_X1 U13085 ( .A1(n14648), .A2(n10639), .ZN(n10640) );
  NAND2_X1 U13086 ( .A1(n14635), .A2(n10640), .ZN(n10724) );
  XNOR2_X1 U13087 ( .A(n10724), .B(n12068), .ZN(n10648) );
  NAND2_X1 U13088 ( .A1(n12006), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U13089 ( .A1(n6491), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10645) );
  AND2_X1 U13090 ( .A1(n10641), .A2(n10976), .ZN(n10642) );
  NOR2_X1 U13091 ( .A1(n10717), .A2(n10642), .ZN(n10980) );
  NAND2_X1 U13092 ( .A1(n11743), .A2(n10980), .ZN(n10644) );
  NAND2_X1 U13093 ( .A1(n11039), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13094 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n13942) );
  AOI22_X1 U13095 ( .A1(n13899), .A2(n13944), .B1(n13942), .B2(n13898), .ZN(
        n10800) );
  INV_X1 U13096 ( .A(n10800), .ZN(n10647) );
  AOI21_X1 U13097 ( .B1(n10648), .B2(n14643), .A(n10647), .ZN(n14705) );
  MUX2_X1 U13098 ( .A(n9219), .B(n14705), .S(n14671), .Z(n10653) );
  OR2_X1 U13099 ( .A1(n10649), .A2(n14648), .ZN(n14650) );
  NOR2_X1 U13100 ( .A1(n14650), .A2(n11875), .ZN(n10757) );
  AOI211_X1 U13101 ( .C1(n11875), .C2(n14650), .A(n14683), .B(n10757), .ZN(
        n14710) );
  INV_X1 U13102 ( .A(n11875), .ZN(n10650) );
  OAI22_X1 U13103 ( .A1(n10650), .A2(n14175), .B1(n10798), .B2(n14662), .ZN(
        n10651) );
  AOI21_X1 U13104 ( .B1(n14710), .B2(n14654), .A(n10651), .ZN(n10652) );
  OAI211_X1 U13105 ( .C1(n14141), .C2(n14706), .A(n10653), .B(n10652), .ZN(
        P1_U3286) );
  NAND2_X1 U13106 ( .A1(n10654), .A2(n14953), .ZN(n10657) );
  AOI22_X1 U13107 ( .A1(n12889), .A2(n10655), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n12888), .ZN(n10656) );
  OAI211_X1 U13108 ( .C1(n8548), .C2(n14953), .A(n10657), .B(n10656), .ZN(
        P3_U3233) );
  INV_X1 U13109 ( .A(n14648), .ZN(n14699) );
  NAND2_X1 U13110 ( .A1(n14648), .A2(n13800), .ZN(n10662) );
  NAND2_X1 U13111 ( .A1(n13944), .A2(n6487), .ZN(n10661) );
  NAND2_X1 U13112 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  XNOR2_X1 U13113 ( .A(n10663), .B(n13798), .ZN(n10790) );
  AND2_X1 U13114 ( .A1(n13944), .A2(n13764), .ZN(n10664) );
  AOI21_X1 U13115 ( .B1(n14648), .B2(n6487), .A(n10664), .ZN(n10788) );
  XNOR2_X1 U13116 ( .A(n10790), .B(n10788), .ZN(n10665) );
  OAI211_X1 U13117 ( .C1(n10666), .C2(n10665), .A(n10792), .B(n14504), .ZN(
        n10670) );
  AOI22_X1 U13118 ( .A1(n13945), .A2(n13899), .B1(n13898), .B2(n13943), .ZN(
        n14637) );
  INV_X1 U13119 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10667) );
  OAI22_X1 U13120 ( .A1(n14637), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10667), .ZN(n10668) );
  AOI21_X1 U13121 ( .B1(n14644), .B2(n13904), .A(n10668), .ZN(n10669) );
  OAI211_X1 U13122 ( .C1(n14699), .C2(n13907), .A(n10670), .B(n10669), .ZN(
        P1_U3239) );
  XNOR2_X1 U13123 ( .A(n6727), .B(n11604), .ZN(n10857) );
  NAND2_X1 U13124 ( .A1(n13206), .A2(n13492), .ZN(n10856) );
  XNOR2_X1 U13125 ( .A(n10857), .B(n10856), .ZN(n10676) );
  INV_X1 U13126 ( .A(n10862), .ZN(n10674) );
  AOI21_X1 U13127 ( .B1(n10676), .B2(n10675), .A(n10674), .ZN(n10683) );
  INV_X1 U13128 ( .A(n13181), .ZN(n13149) );
  NAND2_X1 U13129 ( .A1(n13151), .A2(n10677), .ZN(n10678) );
  OAI211_X1 U13130 ( .C1(n13149), .C2(n10680), .A(n10679), .B(n10678), .ZN(
        n10681) );
  AOI21_X1 U13131 ( .B1(n6727), .B2(n13173), .A(n10681), .ZN(n10682) );
  OAI21_X1 U13132 ( .B1(n10683), .B2(n13187), .A(n10682), .ZN(P2_U3193) );
  INV_X1 U13133 ( .A(n10688), .ZN(n10809) );
  XNOR2_X1 U13134 ( .A(n10810), .B(n10809), .ZN(n10929) );
  OR2_X1 U13135 ( .A1(n6727), .A2(n10684), .ZN(n10686) );
  OAI211_X1 U13136 ( .C1(n10689), .C2(n10688), .A(n10815), .B(n13488), .ZN(
        n10693) );
  NAND2_X1 U13137 ( .A1(n13435), .A2(n13206), .ZN(n10691) );
  NAND2_X1 U13138 ( .A1(n13204), .A2(n13437), .ZN(n10690) );
  NAND2_X1 U13139 ( .A1(n10691), .A2(n10690), .ZN(n10853) );
  INV_X1 U13140 ( .A(n10853), .ZN(n10692) );
  NAND2_X1 U13141 ( .A1(n10693), .A2(n10692), .ZN(n10925) );
  INV_X1 U13142 ( .A(n10927), .ZN(n10698) );
  AOI21_X1 U13143 ( .B1(n10694), .B2(n10927), .A(n13492), .ZN(n10695) );
  AND2_X1 U13144 ( .A1(n10695), .A2(n10821), .ZN(n10926) );
  NAND2_X1 U13145 ( .A1(n10926), .A2(n13507), .ZN(n10697) );
  AOI22_X1 U13146 ( .A1(n13509), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10852), 
        .B2(n13495), .ZN(n10696) );
  OAI211_X1 U13147 ( .C1(n10698), .C2(n13498), .A(n10697), .B(n10696), .ZN(
        n10699) );
  AOI21_X1 U13148 ( .B1(n10925), .B2(n13476), .A(n10699), .ZN(n10700) );
  OAI21_X1 U13149 ( .B1(n13504), .B2(n10929), .A(n10700), .ZN(P2_U3256) );
  INV_X1 U13150 ( .A(n10701), .ZN(n10703) );
  INV_X1 U13151 ( .A(n13057), .ZN(n14413) );
  OAI22_X1 U13152 ( .A1(n12544), .A2(P3_U3151), .B1(SI_22_), .B2(n13054), .ZN(
        n10702) );
  AOI21_X1 U13153 ( .B1(n10703), .B2(n14413), .A(n10702), .ZN(P3_U3273) );
  INV_X1 U13154 ( .A(n11638), .ZN(n10807) );
  AOI22_X1 U13155 ( .A1(n15225), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n13633), .ZN(n10704) );
  OAI21_X1 U13156 ( .B1(n10807), .B2(n13637), .A(n10704), .ZN(P2_U3309) );
  INV_X1 U13157 ( .A(n12068), .ZN(n10705) );
  OR2_X1 U13158 ( .A1(n11875), .A2(n13943), .ZN(n10707) );
  NAND2_X1 U13159 ( .A1(n10708), .A2(n12025), .ZN(n10711) );
  AOI22_X1 U13160 ( .A1(n11646), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11645), 
        .B2(n10709), .ZN(n10710) );
  NAND2_X1 U13161 ( .A1(n10711), .A2(n10710), .ZN(n11883) );
  XNOR2_X1 U13162 ( .A(n11883), .B(n13942), .ZN(n12070) );
  INV_X1 U13163 ( .A(n12070), .ZN(n10756) );
  OR2_X1 U13164 ( .A1(n11883), .A2(n13942), .ZN(n10712) );
  NAND2_X1 U13165 ( .A1(n10713), .A2(n12025), .ZN(n10716) );
  AOI22_X1 U13166 ( .A1(n11646), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11645), 
        .B2(n10714), .ZN(n10715) );
  NAND2_X1 U13167 ( .A1(n10716), .A2(n10715), .ZN(n11893) );
  NAND2_X1 U13168 ( .A1(n6491), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13169 ( .A1(n12006), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10721) );
  OR2_X1 U13170 ( .A1(n10717), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10718) );
  AND2_X1 U13171 ( .A1(n10734), .A2(n10718), .ZN(n11222) );
  NAND2_X1 U13172 ( .A1(n11743), .A2(n11222), .ZN(n10720) );
  NAND2_X1 U13173 ( .A1(n11039), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13174 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n13941) );
  INV_X1 U13175 ( .A(n13941), .ZN(n10881) );
  XNOR2_X1 U13176 ( .A(n11893), .B(n10881), .ZN(n12072) );
  XNOR2_X1 U13177 ( .A(n10874), .B(n12072), .ZN(n14724) );
  INV_X1 U13178 ( .A(n14724), .ZN(n10749) );
  INV_X1 U13179 ( .A(n13943), .ZN(n10725) );
  OR2_X1 U13180 ( .A1(n11875), .A2(n10725), .ZN(n10723) );
  NAND2_X1 U13181 ( .A1(n10724), .A2(n10723), .ZN(n10727) );
  NAND2_X1 U13182 ( .A1(n11875), .A2(n10725), .ZN(n10726) );
  INV_X1 U13183 ( .A(n13942), .ZN(n10728) );
  OR2_X1 U13184 ( .A1(n11883), .A2(n10728), .ZN(n10729) );
  NAND2_X1 U13185 ( .A1(n10730), .A2(n12072), .ZN(n10731) );
  NAND2_X1 U13186 ( .A1(n10882), .A2(n10731), .ZN(n10732) );
  NAND2_X1 U13187 ( .A1(n10732), .A2(n14643), .ZN(n10743) );
  NAND2_X1 U13188 ( .A1(n13942), .A2(n13899), .ZN(n10741) );
  NAND2_X1 U13189 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  NAND2_X1 U13190 ( .A1(n10891), .A2(n10735), .ZN(n14487) );
  OR2_X1 U13191 ( .A1(n11720), .A2(n14487), .ZN(n10739) );
  NAND2_X1 U13192 ( .A1(n12006), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13193 ( .A1(n11039), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13194 ( .A1(n6491), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10736) );
  NAND4_X1 U13195 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n13940) );
  NAND2_X1 U13196 ( .A1(n13940), .A2(n13898), .ZN(n10740) );
  NAND2_X1 U13197 ( .A1(n10741), .A2(n10740), .ZN(n11223) );
  INV_X1 U13198 ( .A(n11223), .ZN(n10742) );
  NAND2_X1 U13199 ( .A1(n10743), .A2(n10742), .ZN(n14731) );
  INV_X1 U13200 ( .A(n11883), .ZN(n10761) );
  AND2_X2 U13201 ( .A1(n10757), .A2(n10761), .ZN(n10887) );
  XNOR2_X1 U13202 ( .A(n10887), .B(n11893), .ZN(n10744) );
  INV_X1 U13203 ( .A(n14683), .ZN(n14651) );
  NAND2_X1 U13204 ( .A1(n10744), .A2(n14651), .ZN(n14727) );
  INV_X1 U13205 ( .A(n14654), .ZN(n14234) );
  AOI22_X1 U13206 ( .A1(n14646), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11222), 
        .B2(n14645), .ZN(n10746) );
  NAND2_X1 U13207 ( .A1(n11893), .A2(n14647), .ZN(n10745) );
  OAI211_X1 U13208 ( .C1(n14727), .C2(n14234), .A(n10746), .B(n10745), .ZN(
        n10747) );
  AOI21_X1 U13209 ( .B1(n14731), .B2(n14671), .A(n10747), .ZN(n10748) );
  OAI21_X1 U13210 ( .B1(n14141), .B2(n10749), .A(n10748), .ZN(P1_U3284) );
  XNOR2_X1 U13211 ( .A(n10750), .B(n12070), .ZN(n10751) );
  NAND2_X1 U13212 ( .A1(n10751), .A2(n14643), .ZN(n10754) );
  NAND2_X1 U13213 ( .A1(n13943), .A2(n13899), .ZN(n10753) );
  NAND2_X1 U13214 ( .A1(n13941), .A2(n13898), .ZN(n10752) );
  AND2_X1 U13215 ( .A1(n10753), .A2(n10752), .ZN(n10977) );
  NAND2_X1 U13216 ( .A1(n10754), .A2(n10977), .ZN(n14719) );
  INV_X1 U13217 ( .A(n14719), .ZN(n10764) );
  XNOR2_X1 U13218 ( .A(n10755), .B(n10756), .ZN(n14715) );
  INV_X1 U13219 ( .A(n14256), .ZN(n14668) );
  OAI21_X1 U13220 ( .B1(n10757), .B2(n10761), .A(n14651), .ZN(n10758) );
  NOR2_X1 U13221 ( .A1(n10758), .A2(n10887), .ZN(n14717) );
  NAND2_X1 U13222 ( .A1(n14717), .A2(n14654), .ZN(n10760) );
  AOI22_X1 U13223 ( .A1(n14646), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n10980), 
        .B2(n14645), .ZN(n10759) );
  OAI211_X1 U13224 ( .C1(n10761), .C2(n14175), .A(n10760), .B(n10759), .ZN(
        n10762) );
  AOI21_X1 U13225 ( .B1(n14715), .B2(n14668), .A(n10762), .ZN(n10763) );
  OAI21_X1 U13226 ( .B1(n10764), .B2(n14646), .A(n10763), .ZN(P1_U3285) );
  INV_X1 U13227 ( .A(n10765), .ZN(n10766) );
  NAND2_X1 U13228 ( .A1(n10766), .A2(n12558), .ZN(n10767) );
  XNOR2_X1 U13229 ( .A(n12153), .B(n15000), .ZN(n10938) );
  XNOR2_X1 U13230 ( .A(n10938), .B(n10986), .ZN(n10769) );
  NAND2_X1 U13231 ( .A1(n10770), .A2(n10769), .ZN(n10940) );
  OAI211_X1 U13232 ( .C1(n10770), .C2(n10769), .A(n10940), .B(n12280), .ZN(
        n10774) );
  OAI22_X1 U13233 ( .A1(n12288), .A2(n10961), .B1(n10959), .B2(n12291), .ZN(
        n10771) );
  AOI211_X1 U13234 ( .C1(n12294), .C2(n12556), .A(n10772), .B(n10771), .ZN(
        n10773) );
  OAI211_X1 U13235 ( .C1(n12307), .C2(n10960), .A(n10774), .B(n10773), .ZN(
        P3_U3161) );
  XNOR2_X1 U13236 ( .A(n10775), .B(n10777), .ZN(n14991) );
  OAI211_X1 U13237 ( .C1(n10778), .C2(n10777), .A(n10776), .B(n14947), .ZN(
        n10782) );
  OAI22_X1 U13238 ( .A1(n10779), .A2(n14943), .B1(n10986), .B2(n14944), .ZN(
        n10780) );
  INV_X1 U13239 ( .A(n10780), .ZN(n10781) );
  AND2_X1 U13240 ( .A1(n10782), .A2(n10781), .ZN(n14990) );
  MUX2_X1 U13241 ( .A(n14990), .B(n10783), .S(n14955), .Z(n10787) );
  INV_X1 U13242 ( .A(n10784), .ZN(n10785) );
  AOI22_X1 U13243 ( .A1(n12889), .A2(n14988), .B1(n12888), .B2(n10785), .ZN(
        n10786) );
  OAI211_X1 U13244 ( .C1(n12892), .C2(n14991), .A(n10787), .B(n10786), .ZN(
        P3_U3226) );
  INV_X1 U13245 ( .A(n14480), .ZN(n13779) );
  NAND2_X1 U13246 ( .A1(n11875), .A2(n14691), .ZN(n14709) );
  INV_X1 U13247 ( .A(n10788), .ZN(n10789) );
  NAND2_X1 U13248 ( .A1(n10790), .A2(n10789), .ZN(n10791) );
  NAND2_X1 U13249 ( .A1(n11875), .A2(n13800), .ZN(n10794) );
  NAND2_X1 U13250 ( .A1(n13943), .A2(n6487), .ZN(n10793) );
  NAND2_X1 U13251 ( .A1(n10794), .A2(n10793), .ZN(n10795) );
  XNOR2_X1 U13252 ( .A(n10795), .B(n13798), .ZN(n10971) );
  AOI21_X1 U13253 ( .B1(n11875), .B2(n6487), .A(n6587), .ZN(n10969) );
  XNOR2_X1 U13254 ( .A(n10971), .B(n10969), .ZN(n10796) );
  OAI211_X1 U13255 ( .C1(n10797), .C2(n10796), .A(n10973), .B(n14504), .ZN(
        n10804) );
  INV_X1 U13256 ( .A(n10798), .ZN(n10802) );
  INV_X1 U13257 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10799) );
  OAI22_X1 U13258 ( .A1(n10800), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10799), .ZN(n10801) );
  AOI21_X1 U13259 ( .B1(n10802), .B2(n13904), .A(n10801), .ZN(n10803) );
  OAI211_X1 U13260 ( .C1(n13779), .C2(n14709), .A(n10804), .B(n10803), .ZN(
        P1_U3213) );
  NAND2_X1 U13261 ( .A1(n10805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10806) );
  XNOR2_X1 U13262 ( .A(n10806), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14624) );
  INV_X1 U13263 ( .A(n14624), .ZN(n10808) );
  OAI222_X1 U13264 ( .A1(P1_U3086), .A2(n10808), .B1(n14382), .B2(n10807), 
        .C1(n7013), .C2(n14379), .ZN(P1_U3337) );
  NAND2_X1 U13265 ( .A1(n10810), .A2(n10809), .ZN(n10812) );
  NAND2_X1 U13266 ( .A1(n10927), .A2(n13205), .ZN(n10811) );
  XNOR2_X1 U13267 ( .A(n11057), .B(n11056), .ZN(n11015) );
  OR2_X1 U13268 ( .A1(n10927), .A2(n10813), .ZN(n10814) );
  NAND2_X1 U13269 ( .A1(n10815), .A2(n10814), .ZN(n10817) );
  INV_X1 U13270 ( .A(n11056), .ZN(n10816) );
  OAI211_X1 U13271 ( .C1(n10817), .C2(n10816), .A(n11064), .B(n13488), .ZN(
        n10820) );
  NAND2_X1 U13272 ( .A1(n13435), .A2(n13205), .ZN(n10819) );
  NAND2_X1 U13273 ( .A1(n13203), .A2(n13437), .ZN(n10818) );
  AND2_X1 U13274 ( .A1(n10819), .A2(n10818), .ZN(n10916) );
  NAND2_X1 U13275 ( .A1(n10820), .A2(n10916), .ZN(n11012) );
  INV_X1 U13276 ( .A(n11062), .ZN(n10921) );
  AOI211_X1 U13277 ( .C1(n11062), .C2(n10821), .A(n13492), .B(n11070), .ZN(
        n11013) );
  NAND2_X1 U13278 ( .A1(n11013), .A2(n13507), .ZN(n10823) );
  AOI22_X1 U13279 ( .A1(n13509), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10918), 
        .B2(n13495), .ZN(n10822) );
  OAI211_X1 U13280 ( .C1(n10921), .C2(n13498), .A(n10823), .B(n10822), .ZN(
        n10824) );
  AOI21_X1 U13281 ( .B1(n11012), .B2(n13476), .A(n10824), .ZN(n10825) );
  OAI21_X1 U13282 ( .B1(n13504), .B2(n11015), .A(n10825), .ZN(P2_U3255) );
  AND2_X1 U13283 ( .A1(n10826), .A2(n15001), .ZN(n14957) );
  XNOR2_X1 U13284 ( .A(n10827), .B(n10828), .ZN(n10829) );
  NAND2_X1 U13285 ( .A1(n10829), .A2(n14947), .ZN(n10832) );
  AOI22_X1 U13286 ( .A1(n12898), .A2(n10830), .B1(n6655), .B2(n12896), .ZN(
        n10831) );
  NAND2_X1 U13287 ( .A1(n10832), .A2(n10831), .ZN(n14956) );
  AOI21_X1 U13288 ( .B1(n14957), .B2(n14938), .A(n14956), .ZN(n10833) );
  MUX2_X1 U13289 ( .A(n10834), .B(n10833), .S(n14953), .Z(n10836) );
  XNOR2_X1 U13290 ( .A(n12501), .B(n12333), .ZN(n14958) );
  INV_X1 U13291 ( .A(n12892), .ZN(n12905) );
  AOI22_X1 U13292 ( .A1(n14958), .A2(n12905), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n12888), .ZN(n10835) );
  NAND2_X1 U13293 ( .A1(n10836), .A2(n10835), .ZN(P3_U3232) );
  OR2_X1 U13294 ( .A1(n10837), .A2(n12503), .ZN(n10838) );
  NAND2_X1 U13295 ( .A1(n10839), .A2(n10838), .ZN(n14986) );
  OAI22_X1 U13296 ( .A1(n12903), .A2(n14983), .B1(n10840), .B2(n14940), .ZN(
        n10849) );
  OAI211_X1 U13297 ( .C1(n10843), .C2(n10842), .A(n10841), .B(n14947), .ZN(
        n10847) );
  OAI22_X1 U13298 ( .A1(n10844), .A2(n14943), .B1(n10959), .B2(n14944), .ZN(
        n10845) );
  AOI21_X1 U13299 ( .B1(n14986), .B2(n14993), .A(n10845), .ZN(n10846) );
  NAND2_X1 U13300 ( .A1(n10847), .A2(n10846), .ZN(n14984) );
  MUX2_X1 U13301 ( .A(n14984), .B(P3_REG2_REG_6__SCAN_IN), .S(n14955), .Z(
        n10848) );
  AOI211_X1 U13302 ( .C1(n10850), .C2(n14986), .A(n10849), .B(n10848), .ZN(
        n10851) );
  INV_X1 U13303 ( .A(n10851), .ZN(P3_U3227) );
  INV_X1 U13304 ( .A(n10852), .ZN(n10855) );
  AOI22_X1 U13305 ( .A1(n13181), .A2(n10853), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10854) );
  OAI21_X1 U13306 ( .B1(n10855), .B2(n13183), .A(n10854), .ZN(n10865) );
  NAND2_X1 U13307 ( .A1(n10857), .A2(n10856), .ZN(n10860) );
  XNOR2_X1 U13308 ( .A(n10927), .B(n11612), .ZN(n10906) );
  NAND2_X1 U13309 ( .A1(n13205), .A2(n13492), .ZN(n10907) );
  XNOR2_X1 U13310 ( .A(n10906), .B(n10907), .ZN(n10859) );
  INV_X1 U13311 ( .A(n10859), .ZN(n10861) );
  NAND3_X1 U13312 ( .A1(n10862), .A2(n10861), .A3(n10860), .ZN(n10863) );
  AOI21_X1 U13313 ( .B1(n10910), .B2(n10863), .A(n13187), .ZN(n10864) );
  AOI211_X1 U13314 ( .C1(n10927), .C2(n13173), .A(n10865), .B(n10864), .ZN(
        n10866) );
  INV_X1 U13315 ( .A(n10866), .ZN(P2_U3203) );
  OAI21_X1 U13316 ( .B1(n6634), .B2(n8620), .A(n10867), .ZN(n10868) );
  AOI222_X1 U13317 ( .A1(n14947), .A2(n10868), .B1(n12559), .B2(n12896), .C1(
        n12560), .C2(n12898), .ZN(n14978) );
  MUX2_X1 U13318 ( .A(n10869), .B(n14978), .S(n14953), .Z(n10873) );
  INV_X1 U13319 ( .A(n10870), .ZN(n10871) );
  AOI22_X1 U13320 ( .A1(n12889), .A2(n14976), .B1(n12888), .B2(n10871), .ZN(
        n10872) );
  OAI211_X1 U13321 ( .C1(n12892), .C2(n14979), .A(n10873), .B(n10872), .ZN(
        P3_U3228) );
  NAND2_X1 U13322 ( .A1(n10874), .A2(n12072), .ZN(n10876) );
  OR2_X1 U13323 ( .A1(n11893), .A2(n13941), .ZN(n10875) );
  NAND2_X1 U13324 ( .A1(n10876), .A2(n10875), .ZN(n11050) );
  NAND2_X1 U13325 ( .A1(n10877), .A2(n12025), .ZN(n10880) );
  AOI22_X1 U13326 ( .A1(n11646), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11645), 
        .B2(n10878), .ZN(n10879) );
  INV_X1 U13327 ( .A(n13940), .ZN(n11030) );
  XNOR2_X1 U13328 ( .A(n14471), .B(n11030), .ZN(n12073) );
  XNOR2_X1 U13329 ( .A(n11050), .B(n12073), .ZN(n14734) );
  INV_X1 U13330 ( .A(n14734), .ZN(n10904) );
  OR2_X1 U13331 ( .A1(n10883), .A2(n12073), .ZN(n11032) );
  NAND2_X1 U13332 ( .A1(n10883), .A2(n12073), .ZN(n10884) );
  NAND3_X1 U13333 ( .A1(n11032), .A2(n14643), .A3(n10884), .ZN(n10885) );
  NAND2_X1 U13334 ( .A1(n13941), .A2(n13899), .ZN(n14483) );
  NAND2_X1 U13335 ( .A1(n10885), .A2(n14483), .ZN(n14739) );
  NAND2_X1 U13336 ( .A1(n14739), .A2(n14671), .ZN(n10903) );
  INV_X1 U13337 ( .A(n11893), .ZN(n10886) );
  NAND2_X1 U13338 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  OR2_X2 U13339 ( .A1(n10888), .A2(n14471), .ZN(n11047) );
  NAND2_X1 U13340 ( .A1(n10888), .A2(n14471), .ZN(n10889) );
  NAND3_X1 U13341 ( .A1(n11047), .A2(n14651), .A3(n10889), .ZN(n10897) );
  AND2_X1 U13342 ( .A1(n10891), .A2(n10890), .ZN(n10892) );
  OR2_X1 U13343 ( .A1(n11037), .A2(n10892), .ZN(n14510) );
  OR2_X1 U13344 ( .A1(n11720), .A2(n14510), .ZN(n10896) );
  NAND2_X1 U13345 ( .A1(n12006), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10895) );
  NAND2_X1 U13346 ( .A1(n11039), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13347 ( .A1(n6491), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U13348 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n13939) );
  NAND2_X1 U13349 ( .A1(n13939), .A2(n13898), .ZN(n14482) );
  NAND2_X1 U13350 ( .A1(n10897), .A2(n14482), .ZN(n14736) );
  INV_X1 U13351 ( .A(n14471), .ZN(n10898) );
  NOR2_X1 U13352 ( .A1(n10898), .A2(n14175), .ZN(n10901) );
  INV_X1 U13353 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10899) );
  OAI22_X1 U13354 ( .A1(n14671), .A2(n10899), .B1(n14487), .B2(n14662), .ZN(
        n10900) );
  AOI211_X1 U13355 ( .C1(n14736), .C2(n14654), .A(n10901), .B(n10900), .ZN(
        n10902) );
  OAI211_X1 U13356 ( .C1(n10904), .C2(n14256), .A(n10903), .B(n10902), .ZN(
        P1_U3283) );
  INV_X1 U13357 ( .A(n11644), .ZN(n10951) );
  OAI222_X1 U13358 ( .A1(n13636), .A2(n10905), .B1(n13637), .B2(n10951), .C1(
        n6754), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U13359 ( .A(n10906), .ZN(n10908) );
  NAND2_X1 U13360 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  XNOR2_X1 U13361 ( .A(n11062), .B(n11604), .ZN(n10998) );
  NAND2_X1 U13362 ( .A1(n13204), .A2(n13492), .ZN(n10999) );
  XNOR2_X1 U13363 ( .A(n10998), .B(n10999), .ZN(n10913) );
  AOI21_X1 U13364 ( .B1(n10912), .B2(n10913), .A(n13187), .ZN(n10914) );
  NAND2_X1 U13365 ( .A1(n10914), .A2(n11003), .ZN(n10920) );
  OAI21_X1 U13366 ( .B1(n13149), .B2(n10916), .A(n10915), .ZN(n10917) );
  AOI21_X1 U13367 ( .B1(n10918), .B2(n13151), .A(n10917), .ZN(n10919) );
  OAI211_X1 U13368 ( .C1(n10921), .C2(n13154), .A(n10920), .B(n10919), .ZN(
        P2_U3189) );
  OAI222_X1 U13369 ( .A1(n12030), .A2(P1_U3086), .B1(n14382), .B2(n11659), 
        .C1(n11660), .C2(n14379), .ZN(P1_U3335) );
  OAI222_X1 U13370 ( .A1(n12037), .A2(P1_U3086), .B1(n14382), .B2(n11672), 
        .C1(n15204), .C2(n14379), .ZN(P1_U3334) );
  OAI222_X1 U13371 ( .A1(n13636), .A2(n10923), .B1(P2_U3088), .B2(n10922), 
        .C1(n13637), .C2(n11659), .ZN(P2_U3307) );
  OAI222_X1 U13372 ( .A1(n13636), .A2(n15043), .B1(P2_U3088), .B2(n10924), 
        .C1(n13637), .C2(n11672), .ZN(P2_U3306) );
  INV_X1 U13373 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10931) );
  AOI211_X1 U13374 ( .C1(n14877), .C2(n10927), .A(n10926), .B(n10925), .ZN(
        n10928) );
  OAI21_X1 U13375 ( .B1(n14875), .B2(n10929), .A(n10928), .ZN(n10932) );
  NAND2_X1 U13376 ( .A1(n10932), .A2(n14886), .ZN(n10930) );
  OAI21_X1 U13377 ( .B1(n14886), .B2(n10931), .A(n10930), .ZN(P2_U3457) );
  NAND2_X1 U13378 ( .A1(n10932), .A2(n14895), .ZN(n10933) );
  OAI21_X1 U13379 ( .B1(n14895), .B2(n10934), .A(n10933), .ZN(P2_U3508) );
  INV_X1 U13380 ( .A(SI_23_), .ZN(n10937) );
  NAND2_X1 U13381 ( .A1(n10935), .A2(n14413), .ZN(n10936) );
  OAI211_X1 U13382 ( .C1(n10937), .C2(n13054), .A(n10936), .B(n12547), .ZN(
        P3_U3272) );
  XNOR2_X1 U13383 ( .A(n12153), .B(n15005), .ZN(n11079) );
  XNOR2_X1 U13384 ( .A(n11079), .B(n11085), .ZN(n10943) );
  NAND2_X1 U13385 ( .A1(n12557), .A2(n10938), .ZN(n10939) );
  INV_X1 U13386 ( .A(n11081), .ZN(n10941) );
  AOI21_X1 U13387 ( .B1(n10943), .B2(n10942), .A(n10941), .ZN(n10949) );
  OAI22_X1 U13388 ( .A1(n12288), .A2(n15005), .B1(n10986), .B2(n12291), .ZN(
        n10944) );
  AOI211_X1 U13389 ( .C1(n12294), .C2(n12555), .A(n10945), .B(n10944), .ZN(
        n10948) );
  NAND2_X1 U13390 ( .A1(n12257), .A2(n10946), .ZN(n10947) );
  OAI211_X1 U13391 ( .C1(n10949), .C2(n12311), .A(n10948), .B(n10947), .ZN(
        P3_U3171) );
  OAI222_X1 U13392 ( .A1(P1_U3086), .A2(n14044), .B1(n14382), .B2(n10951), 
        .C1(n10950), .C2(n14379), .ZN(P1_U3336) );
  OAI222_X1 U13393 ( .A1(n13636), .A2(n10953), .B1(P2_U3088), .B2(n8263), .C1(
        n13637), .C2(n10952), .ZN(P2_U3305) );
  XOR2_X1 U13394 ( .A(n10954), .B(n12505), .Z(n14995) );
  INV_X1 U13395 ( .A(n10955), .ZN(n10956) );
  AOI21_X1 U13396 ( .B1(n12505), .B2(n10957), .A(n10956), .ZN(n10958) );
  OAI222_X1 U13397 ( .A1(n14944), .A2(n11085), .B1(n14943), .B2(n10959), .C1(
        n12861), .C2(n10958), .ZN(n14998) );
  NAND2_X1 U13398 ( .A1(n14998), .A2(n14953), .ZN(n10964) );
  OAI22_X1 U13399 ( .A1(n12903), .A2(n10961), .B1(n10960), .B2(n14940), .ZN(
        n10962) );
  AOI21_X1 U13400 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14955), .A(n10962), .ZN(
        n10963) );
  OAI211_X1 U13401 ( .C1(n12892), .C2(n14995), .A(n10964), .B(n10963), .ZN(
        P3_U3225) );
  NAND2_X1 U13402 ( .A1(n11883), .A2(n13800), .ZN(n10966) );
  NAND2_X1 U13403 ( .A1(n13942), .A2(n6487), .ZN(n10965) );
  NAND2_X1 U13404 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  XNOR2_X1 U13405 ( .A(n10967), .B(n13752), .ZN(n11216) );
  AND2_X1 U13406 ( .A1(n13942), .A2(n13764), .ZN(n10968) );
  AOI21_X1 U13407 ( .B1(n11883), .B2(n6487), .A(n10968), .ZN(n11215) );
  XNOR2_X1 U13408 ( .A(n11216), .B(n11215), .ZN(n10975) );
  INV_X1 U13409 ( .A(n10969), .ZN(n10970) );
  NAND2_X1 U13410 ( .A1(n10971), .A2(n10970), .ZN(n10972) );
  AOI21_X1 U13411 ( .B1(n10975), .B2(n10974), .A(n6631), .ZN(n10982) );
  OAI22_X1 U13412 ( .A1(n10977), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10976), .ZN(n10979) );
  NAND2_X1 U13413 ( .A1(n11883), .A2(n14691), .ZN(n14716) );
  NOR2_X1 U13414 ( .A1(n14716), .A2(n13779), .ZN(n10978) );
  AOI211_X1 U13415 ( .C1(n10980), .C2(n13904), .A(n10979), .B(n10978), .ZN(
        n10981) );
  OAI21_X1 U13416 ( .B1(n10982), .B2(n14475), .A(n10981), .ZN(P1_U3221) );
  XNOR2_X1 U13417 ( .A(n10983), .B(n12368), .ZN(n15003) );
  OAI211_X1 U13418 ( .C1(n10985), .C2(n12368), .A(n10984), .B(n14947), .ZN(
        n10989) );
  OAI22_X1 U13419 ( .A1(n10986), .A2(n14943), .B1(n11274), .B2(n14944), .ZN(
        n10987) );
  INV_X1 U13420 ( .A(n10987), .ZN(n10988) );
  OAI211_X1 U13421 ( .C1(n14997), .C2(n15003), .A(n10989), .B(n10988), .ZN(
        n15006) );
  NAND2_X1 U13422 ( .A1(n15006), .A2(n14953), .ZN(n10993) );
  OAI22_X1 U13423 ( .A1(n12903), .A2(n15005), .B1(n10990), .B2(n14940), .ZN(
        n10991) );
  AOI21_X1 U13424 ( .B1(n14955), .B2(P3_REG2_REG_9__SCAN_IN), .A(n10991), .ZN(
        n10992) );
  OAI211_X1 U13425 ( .C1(n15003), .C2(n12757), .A(n10993), .B(n10992), .ZN(
        P3_U3224) );
  XNOR2_X1 U13426 ( .A(n11291), .B(n11604), .ZN(n10994) );
  NAND2_X1 U13427 ( .A1(n13203), .A2(n13492), .ZN(n10995) );
  NAND2_X1 U13428 ( .A1(n10994), .A2(n10995), .ZN(n11234) );
  INV_X1 U13429 ( .A(n10994), .ZN(n10997) );
  INV_X1 U13430 ( .A(n10995), .ZN(n10996) );
  NAND2_X1 U13431 ( .A1(n10997), .A2(n10996), .ZN(n11236) );
  NAND2_X1 U13432 ( .A1(n11234), .A2(n11236), .ZN(n11004) );
  INV_X1 U13433 ( .A(n10998), .ZN(n11001) );
  INV_X1 U13434 ( .A(n10999), .ZN(n11000) );
  NAND2_X1 U13435 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  XOR2_X1 U13436 ( .A(n11004), .B(n11235), .Z(n11011) );
  INV_X1 U13437 ( .A(n11073), .ZN(n11008) );
  NAND2_X1 U13438 ( .A1(n13435), .A2(n13204), .ZN(n11006) );
  NAND2_X1 U13439 ( .A1(n13202), .A2(n13437), .ZN(n11005) );
  NAND2_X1 U13440 ( .A1(n11006), .A2(n11005), .ZN(n11067) );
  AOI22_X1 U13441 ( .A1(n13181), .A2(n11067), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11007) );
  OAI21_X1 U13442 ( .B1(n11008), .B2(n13183), .A(n11007), .ZN(n11009) );
  AOI21_X1 U13443 ( .B1(n11291), .B2(n13173), .A(n11009), .ZN(n11010) );
  OAI21_X1 U13444 ( .B1(n11011), .B2(n13187), .A(n11010), .ZN(P2_U3208) );
  INV_X1 U13445 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11017) );
  AOI211_X1 U13446 ( .C1(n14877), .C2(n11062), .A(n11013), .B(n11012), .ZN(
        n11014) );
  OAI21_X1 U13447 ( .B1(n14875), .B2(n11015), .A(n11014), .ZN(n11018) );
  NAND2_X1 U13448 ( .A1(n11018), .A2(n14886), .ZN(n11016) );
  OAI21_X1 U13449 ( .B1(n14886), .B2(n11017), .A(n11016), .ZN(P2_U3460) );
  NAND2_X1 U13450 ( .A1(n11018), .A2(n14895), .ZN(n11019) );
  OAI21_X1 U13451 ( .B1(n14895), .B2(n13215), .A(n11019), .ZN(P2_U3509) );
  OAI211_X1 U13452 ( .C1(n11021), .C2(n12511), .A(n11020), .B(n14947), .ZN(
        n11023) );
  AOI22_X1 U13453 ( .A1(n12898), .A2(n12556), .B1(n12554), .B2(n12896), .ZN(
        n11022) );
  NAND2_X1 U13454 ( .A1(n11023), .A2(n11022), .ZN(n11248) );
  INV_X1 U13455 ( .A(n11248), .ZN(n11029) );
  XNOR2_X1 U13456 ( .A(n11024), .B(n12511), .ZN(n11249) );
  NOR2_X1 U13457 ( .A1(n14953), .A2(n11025), .ZN(n11027) );
  OAI22_X1 U13458 ( .A1(n12903), .A2(n11254), .B1(n11086), .B2(n14940), .ZN(
        n11026) );
  AOI211_X1 U13459 ( .C1(n11249), .C2(n12905), .A(n11027), .B(n11026), .ZN(
        n11028) );
  OAI21_X1 U13460 ( .B1(n11029), .B2(n14955), .A(n11028), .ZN(P3_U3223) );
  OR2_X1 U13461 ( .A1(n14471), .A2(n11030), .ZN(n11031) );
  NAND2_X1 U13462 ( .A1(n11033), .A2(n12025), .ZN(n11036) );
  AOI22_X1 U13463 ( .A1(n11646), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11645), 
        .B2(n11034), .ZN(n11035) );
  INV_X1 U13464 ( .A(n13939), .ZN(n11119) );
  XNOR2_X1 U13465 ( .A(n14503), .B(n11119), .ZN(n12074) );
  XNOR2_X1 U13466 ( .A(n11118), .B(n12074), .ZN(n11046) );
  NAND2_X1 U13467 ( .A1(n13940), .A2(n13899), .ZN(n11045) );
  NAND2_X1 U13468 ( .A1(n6491), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U13469 ( .A1(n12006), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11042) );
  OR2_X1 U13470 ( .A1(n11037), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11038) );
  AND2_X1 U13471 ( .A1(n11150), .A2(n11038), .ZN(n11479) );
  NAND2_X1 U13472 ( .A1(n11743), .A2(n11479), .ZN(n11041) );
  NAND2_X1 U13473 ( .A1(n11039), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11040) );
  NAND4_X1 U13474 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n13938) );
  NAND2_X1 U13475 ( .A1(n13938), .A2(n13898), .ZN(n11044) );
  NAND2_X1 U13476 ( .A1(n11045), .A2(n11044), .ZN(n14507) );
  AOI21_X1 U13477 ( .B1(n11046), .B2(n14643), .A(n14507), .ZN(n11135) );
  AOI211_X1 U13478 ( .C1(n14503), .C2(n11047), .A(n14683), .B(n11127), .ZN(
        n11133) );
  INV_X1 U13479 ( .A(n14510), .ZN(n11048) );
  AOI22_X1 U13480 ( .A1(n14646), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11048), 
        .B2(n14645), .ZN(n11049) );
  OAI21_X1 U13481 ( .B1(n7200), .B2(n14175), .A(n11049), .ZN(n11054) );
  NAND2_X1 U13482 ( .A1(n11050), .A2(n12073), .ZN(n11052) );
  OR2_X1 U13483 ( .A1(n14471), .A2(n13940), .ZN(n11051) );
  NAND2_X1 U13484 ( .A1(n11052), .A2(n11051), .ZN(n11112) );
  XOR2_X1 U13485 ( .A(n11112), .B(n12074), .Z(n11136) );
  NOR2_X1 U13486 ( .A1(n11136), .A2(n14256), .ZN(n11053) );
  AOI211_X1 U13487 ( .C1(n11133), .C2(n14654), .A(n11054), .B(n11053), .ZN(
        n11055) );
  OAI21_X1 U13488 ( .B1(n14646), .B2(n11135), .A(n11055), .ZN(P1_U3282) );
  NAND2_X1 U13489 ( .A1(n11057), .A2(n11056), .ZN(n11059) );
  NAND2_X1 U13490 ( .A1(n11062), .A2(n13204), .ZN(n11058) );
  XNOR2_X1 U13491 ( .A(n11093), .B(n11066), .ZN(n11293) );
  OR2_X1 U13492 ( .A1(n11062), .A2(n11061), .ZN(n11063) );
  AOI21_X1 U13493 ( .B1(n11066), .B2(n11065), .A(n6611), .ZN(n11069) );
  INV_X1 U13494 ( .A(n11067), .ZN(n11068) );
  OAI21_X1 U13495 ( .B1(n11069), .B2(n13451), .A(n11068), .ZN(n11289) );
  INV_X1 U13496 ( .A(n11291), .ZN(n11076) );
  INV_X1 U13497 ( .A(n11070), .ZN(n11072) );
  NAND2_X1 U13498 ( .A1(n11070), .A2(n11076), .ZN(n11102) );
  INV_X1 U13499 ( .A(n11102), .ZN(n11071) );
  AOI211_X1 U13500 ( .C1(n11291), .C2(n11072), .A(n13492), .B(n11071), .ZN(
        n11290) );
  NAND2_X1 U13501 ( .A1(n11290), .A2(n13507), .ZN(n11075) );
  AOI22_X1 U13502 ( .A1(n13509), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11073), 
        .B2(n13495), .ZN(n11074) );
  OAI211_X1 U13503 ( .C1(n11076), .C2(n13498), .A(n11075), .B(n11074), .ZN(
        n11077) );
  AOI21_X1 U13504 ( .B1(n11289), .B2(n13476), .A(n11077), .ZN(n11078) );
  OAI21_X1 U13505 ( .B1(n11293), .B2(n13504), .A(n11078), .ZN(P2_U3254) );
  NAND2_X1 U13506 ( .A1(n11079), .A2(n11085), .ZN(n11080) );
  XNOR2_X1 U13507 ( .A(n11089), .B(n12153), .ZN(n11325) );
  XNOR2_X1 U13508 ( .A(n11325), .B(n11274), .ZN(n11082) );
  OAI211_X1 U13509 ( .C1(n6635), .C2(n11082), .A(n11327), .B(n12280), .ZN(
        n11091) );
  NAND2_X1 U13510 ( .A1(n12554), .A2(n12294), .ZN(n11084) );
  OAI211_X1 U13511 ( .C1(n11085), .C2(n12291), .A(n11084), .B(n11083), .ZN(
        n11088) );
  NOR2_X1 U13512 ( .A1(n12307), .A2(n11086), .ZN(n11087) );
  AOI211_X1 U13513 ( .C1(n11089), .C2(n9993), .A(n11088), .B(n11087), .ZN(
        n11090) );
  NAND2_X1 U13514 ( .A1(n11091), .A2(n11090), .ZN(P3_U3157) );
  AND2_X1 U13515 ( .A1(n11291), .A2(n13203), .ZN(n11092) );
  OR2_X1 U13516 ( .A1(n11291), .A2(n13203), .ZN(n11094) );
  XNOR2_X1 U13517 ( .A(n11199), .B(n11198), .ZN(n11260) );
  INV_X1 U13518 ( .A(n11260), .ZN(n11108) );
  AND2_X1 U13519 ( .A1(n11291), .A2(n11095), .ZN(n11096) );
  OAI21_X1 U13520 ( .B1(n6611), .B2(n11096), .A(n11198), .ZN(n11098) );
  NOR2_X1 U13521 ( .A1(n11198), .A2(n11096), .ZN(n11097) );
  NAND3_X1 U13522 ( .A1(n11098), .A2(n13488), .A3(n11204), .ZN(n11101) );
  NAND2_X1 U13523 ( .A1(n13435), .A2(n13203), .ZN(n11100) );
  NAND2_X1 U13524 ( .A1(n13201), .A2(n13437), .ZN(n11099) );
  AND2_X1 U13525 ( .A1(n11100), .A2(n11099), .ZN(n11242) );
  NAND2_X1 U13526 ( .A1(n11101), .A2(n11242), .ZN(n11258) );
  AOI21_X1 U13527 ( .B1(n11255), .B2(n11102), .A(n13492), .ZN(n11103) );
  NAND2_X1 U13528 ( .A1(n11103), .A2(n11210), .ZN(n11256) );
  AOI22_X1 U13529 ( .A1(n13392), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11244), 
        .B2(n13495), .ZN(n11105) );
  NAND2_X1 U13530 ( .A1(n11255), .A2(n13483), .ZN(n11104) );
  OAI211_X1 U13531 ( .C1(n11256), .C2(n13371), .A(n11105), .B(n11104), .ZN(
        n11106) );
  AOI21_X1 U13532 ( .B1(n11258), .B2(n13476), .A(n11106), .ZN(n11107) );
  OAI21_X1 U13533 ( .B1(n11108), .B2(n13504), .A(n11107), .ZN(P2_U3253) );
  NAND2_X1 U13534 ( .A1(n13633), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11109) );
  OAI211_X1 U13535 ( .C1(n11693), .C2(n13637), .A(n11110), .B(n11109), .ZN(
        P2_U3304) );
  NAND2_X1 U13536 ( .A1(n14369), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11111) );
  OAI211_X1 U13537 ( .C1(n11693), .C2(n14382), .A(n12105), .B(n11111), .ZN(
        P1_U3332) );
  NAND2_X1 U13538 ( .A1(n14503), .A2(n13939), .ZN(n11113) );
  NAND2_X1 U13539 ( .A1(n11114), .A2(n12025), .ZN(n11116) );
  AOI22_X1 U13540 ( .A1(n11646), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11645), 
        .B2(n14025), .ZN(n11115) );
  INV_X1 U13541 ( .A(n13938), .ZN(n11143) );
  XNOR2_X1 U13542 ( .A(n14424), .B(n11143), .ZN(n12076) );
  XNOR2_X1 U13543 ( .A(n11165), .B(n12076), .ZN(n14426) );
  NAND2_X1 U13544 ( .A1(n14503), .A2(n11119), .ZN(n11117) );
  OR2_X1 U13545 ( .A1(n14503), .A2(n11119), .ZN(n11120) );
  INV_X1 U13546 ( .A(n12076), .ZN(n11141) );
  XNOR2_X1 U13547 ( .A(n11142), .B(n11141), .ZN(n11126) );
  XNOR2_X1 U13548 ( .A(n11150), .B(n11149), .ZN(n14496) );
  OR2_X1 U13549 ( .A1(n11720), .A2(n14496), .ZN(n11125) );
  NAND2_X1 U13550 ( .A1(n12006), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U13551 ( .A1(n11039), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U13552 ( .A1(n6491), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11122) );
  NAND4_X1 U13553 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n13937) );
  AOI22_X1 U13554 ( .A1(n13899), .A2(n13939), .B1(n13937), .B2(n13898), .ZN(
        n11477) );
  OAI21_X1 U13555 ( .B1(n11126), .B2(n14676), .A(n11477), .ZN(n14428) );
  NAND2_X1 U13556 ( .A1(n14428), .A2(n14671), .ZN(n11132) );
  INV_X1 U13557 ( .A(n11127), .ZN(n11128) );
  INV_X1 U13558 ( .A(n14424), .ZN(n11482) );
  AOI211_X1 U13559 ( .C1(n14424), .C2(n11128), .A(n14683), .B(n11160), .ZN(
        n14423) );
  AOI22_X1 U13560 ( .A1(n14646), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11479), 
        .B2(n14645), .ZN(n11129) );
  OAI21_X1 U13561 ( .B1(n11482), .B2(n14175), .A(n11129), .ZN(n11130) );
  AOI21_X1 U13562 ( .B1(n14423), .B2(n14654), .A(n11130), .ZN(n11131) );
  OAI211_X1 U13563 ( .C1(n14426), .C2(n14256), .A(n11132), .B(n11131), .ZN(
        P1_U3281) );
  AOI21_X1 U13564 ( .B1(n14691), .B2(n14503), .A(n11133), .ZN(n11134) );
  OAI211_X1 U13565 ( .C1(n14677), .C2(n11136), .A(n11135), .B(n11134), .ZN(
        n11138) );
  NAND2_X1 U13566 ( .A1(n11138), .A2(n14753), .ZN(n11137) );
  OAI21_X1 U13567 ( .B1(n14753), .B2(n10348), .A(n11137), .ZN(P1_U3539) );
  INV_X1 U13568 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U13569 ( .A1(n11138), .A2(n14742), .ZN(n11139) );
  OAI21_X1 U13570 ( .B1(n14742), .B2(n11140), .A(n11139), .ZN(P1_U3492) );
  OR2_X1 U13571 ( .A1(n14424), .A2(n11143), .ZN(n11144) );
  NAND2_X1 U13572 ( .A1(n11145), .A2(n12025), .ZN(n11147) );
  AOI22_X1 U13573 ( .A1(n11646), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11645), 
        .B2(n14557), .ZN(n11146) );
  XNOR2_X1 U13574 ( .A(n14492), .B(n13937), .ZN(n12077) );
  INV_X1 U13575 ( .A(n12077), .ZN(n11168) );
  XNOR2_X1 U13576 ( .A(n11349), .B(n11168), .ZN(n11159) );
  NAND2_X1 U13577 ( .A1(n11039), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11157) );
  OAI21_X1 U13578 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n11151) );
  NAND2_X1 U13579 ( .A1(n11151), .A2(n11352), .ZN(n14470) );
  OR2_X1 U13580 ( .A1(n11720), .A2(n14470), .ZN(n11156) );
  INV_X1 U13581 ( .A(n11152), .ZN(n12009) );
  INV_X1 U13582 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11363) );
  OR2_X1 U13583 ( .A1(n12009), .A2(n11363), .ZN(n11155) );
  INV_X1 U13584 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11153) );
  OR2_X1 U13585 ( .A1(n7529), .A2(n11153), .ZN(n11154) );
  NAND2_X1 U13586 ( .A1(n13938), .A2(n13899), .ZN(n11158) );
  OAI21_X1 U13587 ( .B1(n13661), .B2(n13848), .A(n11158), .ZN(n14491) );
  AOI21_X1 U13588 ( .B1(n11159), .B2(n14643), .A(n14491), .ZN(n11282) );
  INV_X1 U13589 ( .A(n11160), .ZN(n11161) );
  INV_X1 U13590 ( .A(n14492), .ZN(n11913) );
  AOI211_X1 U13591 ( .C1(n14492), .C2(n11161), .A(n14683), .B(n7197), .ZN(
        n11280) );
  NOR2_X1 U13592 ( .A1(n11913), .A2(n14175), .ZN(n11164) );
  INV_X1 U13593 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11162) );
  OAI22_X1 U13594 ( .A1(n14671), .A2(n11162), .B1(n14496), .B2(n14662), .ZN(
        n11163) );
  AOI211_X1 U13595 ( .C1(n11280), .C2(n14654), .A(n11164), .B(n11163), .ZN(
        n11171) );
  OR2_X1 U13596 ( .A1(n14424), .A2(n13938), .ZN(n11166) );
  NAND2_X1 U13597 ( .A1(n11167), .A2(n11166), .ZN(n11169) );
  OAI21_X1 U13598 ( .B1(n11169), .B2(n11168), .A(n11345), .ZN(n11279) );
  NAND2_X1 U13599 ( .A1(n11279), .A2(n14668), .ZN(n11170) );
  OAI211_X1 U13600 ( .C1(n11282), .C2(n14646), .A(n11171), .B(n11170), .ZN(
        P1_U3280) );
  NOR2_X1 U13601 ( .A1(n11188), .A2(n11173), .ZN(n11174) );
  MUX2_X1 U13602 ( .A(n11175), .B(P3_REG1_REG_12__SCAN_IN), .S(n12582), .Z(
        n11177) );
  INV_X1 U13603 ( .A(n12566), .ZN(n11176) );
  AOI21_X1 U13604 ( .B1(n11178), .B2(n11177), .A(n11176), .ZN(n11197) );
  INV_X1 U13605 ( .A(n11179), .ZN(n11180) );
  NOR2_X1 U13606 ( .A1(n11181), .A2(n11180), .ZN(n14903) );
  MUX2_X1 U13607 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12623), .Z(n11182) );
  XNOR2_X1 U13608 ( .A(n11182), .B(n14900), .ZN(n14902) );
  NOR2_X1 U13609 ( .A1(n11182), .A2(n14900), .ZN(n11184) );
  MUX2_X1 U13610 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12623), .Z(n12581) );
  XNOR2_X1 U13611 ( .A(n12581), .B(n12582), .ZN(n11183) );
  NOR3_X1 U13612 ( .A1(n14901), .A2(n11184), .A3(n11183), .ZN(n14920) );
  NOR2_X1 U13613 ( .A1(n14920), .A2(n14928), .ZN(n11195) );
  OAI21_X1 U13614 ( .B1(n14901), .B2(n11184), .A(n11183), .ZN(n11194) );
  INV_X1 U13615 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11185) );
  NOR2_X1 U13616 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11185), .ZN(n11373) );
  AOI21_X1 U13617 ( .B1(n14896), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11373), 
        .ZN(n11192) );
  NOR2_X1 U13618 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  MUX2_X1 U13619 ( .A(n11302), .B(P3_REG2_REG_12__SCAN_IN), .S(n12582), .Z(
        n12570) );
  XNOR2_X1 U13620 ( .A(n12571), .B(n12570), .ZN(n11190) );
  NAND2_X1 U13621 ( .A1(n12592), .A2(n11190), .ZN(n11191) );
  OAI211_X1 U13622 ( .C1(n14918), .C2(n12582), .A(n11192), .B(n11191), .ZN(
        n11193) );
  AOI21_X1 U13623 ( .B1(n11195), .B2(n11194), .A(n11193), .ZN(n11196) );
  OAI21_X1 U13624 ( .B1(n11197), .B2(n14926), .A(n11196), .ZN(P3_U3194) );
  OR2_X1 U13625 ( .A1(n11255), .A2(n13202), .ZN(n11200) );
  NAND2_X1 U13626 ( .A1(n11201), .A2(n11200), .ZN(n11307) );
  INV_X1 U13627 ( .A(n11202), .ZN(n11205) );
  XNOR2_X1 U13628 ( .A(n11307), .B(n11205), .ZN(n13605) );
  NAND2_X1 U13629 ( .A1(n11204), .A2(n11203), .ZN(n11206) );
  OAI211_X1 U13630 ( .C1(n11206), .C2(n11205), .A(n11311), .B(n13488), .ZN(
        n11209) );
  NAND2_X1 U13631 ( .A1(n13435), .A2(n13202), .ZN(n11208) );
  NAND2_X1 U13632 ( .A1(n13200), .A2(n13437), .ZN(n11207) );
  AND2_X1 U13633 ( .A1(n11208), .A2(n11207), .ZN(n11266) );
  NAND2_X1 U13634 ( .A1(n11209), .A2(n11266), .ZN(n13601) );
  AOI211_X1 U13635 ( .C1(n13603), .C2(n11210), .A(n13492), .B(n7008), .ZN(
        n13602) );
  NAND2_X1 U13636 ( .A1(n13602), .A2(n13507), .ZN(n11212) );
  AOI22_X1 U13637 ( .A1(n13392), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11268), 
        .B2(n13495), .ZN(n11211) );
  OAI211_X1 U13638 ( .C1(n7009), .C2(n13498), .A(n11212), .B(n11211), .ZN(
        n11213) );
  AOI21_X1 U13639 ( .B1(n13601), .B2(n13476), .A(n11213), .ZN(n11214) );
  OAI21_X1 U13640 ( .B1(n13504), .B2(n13605), .A(n11214), .ZN(P2_U3252) );
  NAND2_X1 U13641 ( .A1(n11893), .A2(n6487), .ZN(n11218) );
  NAND2_X1 U13642 ( .A1(n13941), .A2(n13764), .ZN(n11217) );
  NAND2_X1 U13643 ( .A1(n11218), .A2(n11217), .ZN(n11449) );
  NAND2_X1 U13644 ( .A1(n11893), .A2(n13800), .ZN(n11220) );
  NAND2_X1 U13645 ( .A1(n13941), .A2(n6487), .ZN(n11219) );
  NAND2_X1 U13646 ( .A1(n11220), .A2(n11219), .ZN(n11221) );
  XNOR2_X1 U13647 ( .A(n11221), .B(n13752), .ZN(n11447) );
  XOR2_X1 U13648 ( .A(n11448), .B(n11447), .Z(n11228) );
  AND2_X1 U13649 ( .A1(n11893), .A2(n14691), .ZN(n14725) );
  INV_X1 U13650 ( .A(n11222), .ZN(n11225) );
  AOI22_X1 U13651 ( .A1(n11223), .A2(n14506), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11224) );
  OAI21_X1 U13652 ( .B1(n14511), .B2(n11225), .A(n11224), .ZN(n11226) );
  AOI21_X1 U13653 ( .B1(n14725), .B2(n14480), .A(n11226), .ZN(n11227) );
  OAI21_X1 U13654 ( .B1(n11228), .B2(n14475), .A(n11227), .ZN(P1_U3231) );
  XNOR2_X1 U13655 ( .A(n11255), .B(n11604), .ZN(n11229) );
  NAND2_X1 U13656 ( .A1(n13202), .A2(n13492), .ZN(n11230) );
  NAND2_X1 U13657 ( .A1(n11229), .A2(n11230), .ZN(n11264) );
  INV_X1 U13658 ( .A(n11229), .ZN(n11232) );
  INV_X1 U13659 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U13660 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  NAND2_X1 U13661 ( .A1(n11264), .A2(n11233), .ZN(n11241) );
  INV_X1 U13662 ( .A(n11241), .ZN(n11239) );
  INV_X1 U13663 ( .A(n11265), .ZN(n11240) );
  AOI21_X1 U13664 ( .B1(n11241), .B2(n11238), .A(n11240), .ZN(n11247) );
  OAI22_X1 U13665 ( .A1(n13149), .A2(n11242), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13240), .ZN(n11243) );
  AOI21_X1 U13666 ( .B1(n11244), .B2(n13151), .A(n11243), .ZN(n11246) );
  NAND2_X1 U13667 ( .A1(n11255), .A2(n13185), .ZN(n11245) );
  OAI211_X1 U13668 ( .C1(n11247), .C2(n13187), .A(n11246), .B(n11245), .ZN(
        P2_U3196) );
  INV_X1 U13669 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11250) );
  AOI21_X1 U13670 ( .B1(n14959), .B2(n11249), .A(n11248), .ZN(n11252) );
  MUX2_X1 U13671 ( .A(n11250), .B(n11252), .S(n15010), .Z(n11251) );
  OAI21_X1 U13672 ( .B1(n13039), .B2(n11254), .A(n11251), .ZN(P3_U3420) );
  MUX2_X1 U13673 ( .A(n10478), .B(n11252), .S(n15025), .Z(n11253) );
  OAI21_X1 U13674 ( .B1(n12961), .B2(n11254), .A(n11253), .ZN(P3_U3469) );
  INV_X1 U13675 ( .A(n11255), .ZN(n11257) );
  OAI21_X1 U13676 ( .B1(n11257), .B2(n14859), .A(n11256), .ZN(n11259) );
  AOI211_X1 U13677 ( .C1(n14865), .C2(n11260), .A(n11259), .B(n11258), .ZN(
        n11263) );
  NAND2_X1 U13678 ( .A1(n14893), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11261) );
  OAI21_X1 U13679 ( .B1(n11263), .B2(n14893), .A(n11261), .ZN(P2_U3511) );
  NAND2_X1 U13680 ( .A1(n14884), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11262) );
  OAI21_X1 U13681 ( .B1(n11263), .B2(n14884), .A(n11262), .ZN(P2_U3466) );
  XNOR2_X1 U13682 ( .A(n13603), .B(n11604), .ZN(n11397) );
  NAND2_X1 U13683 ( .A1(n13201), .A2(n13492), .ZN(n11396) );
  XNOR2_X1 U13684 ( .A(n11397), .B(n11396), .ZN(n11399) );
  XNOR2_X1 U13685 ( .A(n11400), .B(n11399), .ZN(n11271) );
  AND2_X1 U13686 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14777) );
  NOR2_X1 U13687 ( .A1(n13149), .A2(n11266), .ZN(n11267) );
  AOI211_X1 U13688 ( .C1(n13151), .C2(n11268), .A(n14777), .B(n11267), .ZN(
        n11270) );
  NAND2_X1 U13689 ( .A1(n13603), .A2(n13185), .ZN(n11269) );
  OAI211_X1 U13690 ( .C1(n11271), .C2(n13187), .A(n11270), .B(n11269), .ZN(
        P2_U3206) );
  INV_X1 U13691 ( .A(n12382), .ZN(n12516) );
  XNOR2_X1 U13692 ( .A(n11272), .B(n12516), .ZN(n14450) );
  XNOR2_X1 U13693 ( .A(n11273), .B(n12516), .ZN(n11275) );
  OAI222_X1 U13694 ( .A1(n14944), .A2(n12264), .B1(n11275), .B2(n12861), .C1(
        n14943), .C2(n11274), .ZN(n14452) );
  NAND2_X1 U13695 ( .A1(n14452), .A2(n14953), .ZN(n11278) );
  OAI22_X1 U13696 ( .A1(n14953), .A2(n8692), .B1(n11332), .B2(n14940), .ZN(
        n11276) );
  AOI21_X1 U13697 ( .B1(n12379), .B2(n12889), .A(n11276), .ZN(n11277) );
  OAI211_X1 U13698 ( .C1(n12892), .C2(n14450), .A(n11278), .B(n11277), .ZN(
        P3_U3222) );
  INV_X1 U13699 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11285) );
  INV_X1 U13700 ( .A(n11279), .ZN(n11283) );
  AOI21_X1 U13701 ( .B1(n14691), .B2(n14492), .A(n11280), .ZN(n11281) );
  OAI211_X1 U13702 ( .C1(n14677), .C2(n11283), .A(n11282), .B(n11281), .ZN(
        n11286) );
  NAND2_X1 U13703 ( .A1(n11286), .A2(n14742), .ZN(n11284) );
  OAI21_X1 U13704 ( .B1(n14742), .B2(n11285), .A(n11284), .ZN(P1_U3498) );
  INV_X1 U13705 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U13706 ( .A1(n11286), .A2(n14753), .ZN(n11287) );
  OAI21_X1 U13707 ( .B1(n14753), .B2(n11288), .A(n11287), .ZN(P1_U3541) );
  INV_X1 U13708 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11295) );
  AOI211_X1 U13709 ( .C1(n14877), .C2(n11291), .A(n11290), .B(n11289), .ZN(
        n11292) );
  OAI21_X1 U13710 ( .B1(n14875), .B2(n11293), .A(n11292), .ZN(n11296) );
  NAND2_X1 U13711 ( .A1(n11296), .A2(n14886), .ZN(n11294) );
  OAI21_X1 U13712 ( .B1(n14886), .B2(n11295), .A(n11294), .ZN(P2_U3463) );
  INV_X1 U13713 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U13714 ( .A1(n11296), .A2(n14895), .ZN(n11297) );
  OAI21_X1 U13715 ( .B1(n14895), .B2(n13217), .A(n11297), .ZN(P2_U3510) );
  XNOR2_X1 U13716 ( .A(n11298), .B(n11300), .ZN(n14445) );
  XNOR2_X1 U13717 ( .A(n11299), .B(n11300), .ZN(n11301) );
  OAI222_X1 U13718 ( .A1(n14944), .A2(n12171), .B1(n11301), .B2(n12861), .C1(
        n14943), .C2(n12380), .ZN(n14447) );
  NAND2_X1 U13719 ( .A1(n14447), .A2(n14953), .ZN(n11305) );
  OAI22_X1 U13720 ( .A1(n14953), .A2(n11302), .B1(n11371), .B2(n14940), .ZN(
        n11303) );
  AOI21_X1 U13721 ( .B1(n12889), .B2(n11377), .A(n11303), .ZN(n11304) );
  OAI211_X1 U13722 ( .C1(n12892), .C2(n14445), .A(n11305), .B(n11304), .ZN(
        P3_U3221) );
  NOR2_X1 U13723 ( .A1(n13603), .A2(n13201), .ZN(n11306) );
  NAND2_X1 U13724 ( .A1(n13603), .A2(n13201), .ZN(n11308) );
  XNOR2_X1 U13725 ( .A(n11413), .B(n11312), .ZN(n13600) );
  OR2_X1 U13726 ( .A1(n13603), .A2(n11309), .ZN(n11310) );
  XOR2_X1 U13727 ( .A(n11312), .B(n11415), .Z(n11315) );
  NAND2_X1 U13728 ( .A1(n13435), .A2(n13201), .ZN(n11314) );
  NAND2_X1 U13729 ( .A1(n13199), .A2(n13437), .ZN(n11313) );
  AND2_X1 U13730 ( .A1(n11314), .A2(n11313), .ZN(n11405) );
  OAI21_X1 U13731 ( .B1(n11315), .B2(n13451), .A(n11405), .ZN(n13596) );
  INV_X1 U13732 ( .A(n11417), .ZN(n11316) );
  AOI211_X1 U13733 ( .C1(n13598), .C2(n11317), .A(n13492), .B(n11316), .ZN(
        n13597) );
  NAND2_X1 U13734 ( .A1(n13597), .A2(n13507), .ZN(n11319) );
  AOI22_X1 U13735 ( .A1(n13509), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11407), 
        .B2(n13495), .ZN(n11318) );
  OAI211_X1 U13736 ( .C1(n7011), .C2(n13498), .A(n11319), .B(n11318), .ZN(
        n11320) );
  AOI21_X1 U13737 ( .B1(n13596), .B2(n13476), .A(n11320), .ZN(n11321) );
  OAI21_X1 U13738 ( .B1(n13600), .B2(n13504), .A(n11321), .ZN(P2_U3251) );
  OAI222_X1 U13739 ( .A1(n11322), .A2(P1_U3086), .B1(n14382), .B2(n11703), 
        .C1(n11704), .C2(n14379), .ZN(P1_U3331) );
  OAI222_X1 U13740 ( .A1(n11324), .A2(P2_U3088), .B1(n13637), .B2(n11703), 
        .C1(n11323), .C2(n13636), .ZN(P2_U3303) );
  NAND2_X1 U13741 ( .A1(n12555), .A2(n11325), .ZN(n11326) );
  XNOR2_X1 U13742 ( .A(n14448), .B(n12194), .ZN(n11328) );
  NAND2_X1 U13743 ( .A1(n11329), .A2(n11328), .ZN(n11369) );
  NAND2_X1 U13744 ( .A1(n11368), .A2(n11369), .ZN(n11330) );
  XNOR2_X1 U13745 ( .A(n11330), .B(n12554), .ZN(n11339) );
  NOR2_X1 U13746 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11331), .ZN(n14910) );
  AOI21_X1 U13747 ( .B1(n12553), .B2(n12294), .A(n14910), .ZN(n11337) );
  INV_X1 U13748 ( .A(n11332), .ZN(n11333) );
  NAND2_X1 U13749 ( .A1(n12257), .A2(n11333), .ZN(n11336) );
  NAND2_X1 U13750 ( .A1(n9993), .A2(n12379), .ZN(n11335) );
  INV_X1 U13751 ( .A(n12291), .ZN(n12305) );
  NAND2_X1 U13752 ( .A1(n12555), .A2(n12305), .ZN(n11334) );
  NAND4_X1 U13753 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11338) );
  AOI21_X1 U13754 ( .B1(n11339), .B2(n12280), .A(n11338), .ZN(n11340) );
  INV_X1 U13755 ( .A(n11340), .ZN(P3_U3176) );
  INV_X1 U13756 ( .A(n11341), .ZN(n11342) );
  OAI222_X1 U13757 ( .A1(n11343), .A2(P3_U3151), .B1(n13054), .B2(n6970), .C1(
        n13057), .C2(n11342), .ZN(P3_U3271) );
  OR2_X1 U13758 ( .A1(n14492), .A2(n13937), .ZN(n11344) );
  NAND2_X1 U13759 ( .A1(n11346), .A2(n12025), .ZN(n11348) );
  AOI22_X1 U13760 ( .A1(n14564), .A2(n11645), .B1(n11646), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11347) );
  OR2_X1 U13761 ( .A1(n14518), .A2(n13661), .ZN(n11916) );
  NAND2_X1 U13762 ( .A1(n14518), .A2(n13661), .ZN(n11924) );
  XNOR2_X1 U13763 ( .A(n11423), .B(n12079), .ZN(n14521) );
  INV_X1 U13764 ( .A(n13937), .ZN(n11914) );
  XNOR2_X1 U13765 ( .A(n11429), .B(n6755), .ZN(n11359) );
  NAND2_X1 U13766 ( .A1(n6491), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U13767 ( .A1(n12006), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U13768 ( .A1(n11039), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11355) );
  INV_X1 U13769 ( .A(n11350), .ZN(n11433) );
  NAND2_X1 U13770 ( .A1(n11352), .A2(n11351), .ZN(n11353) );
  NAND2_X1 U13771 ( .A1(n11433), .A2(n11353), .ZN(n13916) );
  OR2_X1 U13772 ( .A1(n11720), .A2(n13916), .ZN(n11354) );
  NAND2_X1 U13773 ( .A1(n13937), .A2(n13899), .ZN(n11358) );
  OAI21_X1 U13774 ( .B1(n13674), .B2(n13848), .A(n11358), .ZN(n14468) );
  AOI21_X1 U13775 ( .B1(n11359), .B2(n14643), .A(n14468), .ZN(n14524) );
  OAI21_X1 U13776 ( .B1(n14470), .B2(n14662), .A(n14524), .ZN(n11360) );
  NAND2_X1 U13777 ( .A1(n11360), .A2(n14671), .ZN(n11367) );
  AOI21_X1 U13778 ( .B1(n14518), .B2(n11361), .A(n14683), .ZN(n11362) );
  AND2_X1 U13779 ( .A1(n11362), .A2(n11440), .ZN(n14520) );
  INV_X1 U13780 ( .A(n14518), .ZN(n11364) );
  OAI22_X1 U13781 ( .A1(n11364), .A2(n14175), .B1(n14671), .B2(n11363), .ZN(
        n11365) );
  AOI21_X1 U13782 ( .B1(n14654), .B2(n14520), .A(n11365), .ZN(n11366) );
  OAI211_X1 U13783 ( .C1(n14521), .C2(n14256), .A(n11367), .B(n11366), .ZN(
        P1_U3279) );
  XNOR2_X1 U13784 ( .A(n11377), .B(n12194), .ZN(n12117) );
  XNOR2_X1 U13785 ( .A(n12553), .B(n12117), .ZN(n11370) );
  XNOR2_X1 U13786 ( .A(n12116), .B(n11370), .ZN(n11379) );
  INV_X1 U13787 ( .A(n11371), .ZN(n11372) );
  NAND2_X1 U13788 ( .A1(n12257), .A2(n11372), .ZN(n11375) );
  AOI21_X1 U13789 ( .B1(n12294), .B2(n12899), .A(n11373), .ZN(n11374) );
  OAI211_X1 U13790 ( .C1(n12380), .C2(n12291), .A(n11375), .B(n11374), .ZN(
        n11376) );
  AOI21_X1 U13791 ( .B1(n11377), .B2(n9993), .A(n11376), .ZN(n11378) );
  OAI21_X1 U13792 ( .B1(n11379), .B2(n12311), .A(n11378), .ZN(P3_U3164) );
  XNOR2_X1 U13793 ( .A(n11380), .B(n12395), .ZN(n14441) );
  XNOR2_X1 U13794 ( .A(n11381), .B(n12395), .ZN(n11382) );
  OAI222_X1 U13795 ( .A1(n14944), .A2(n12124), .B1(n11382), .B2(n12861), .C1(
        n14943), .C2(n12264), .ZN(n14443) );
  NAND2_X1 U13796 ( .A1(n14443), .A2(n14953), .ZN(n11386) );
  INV_X1 U13797 ( .A(n14440), .ZN(n12269) );
  OAI22_X1 U13798 ( .A1(n14953), .A2(n11383), .B1(n12267), .B2(n14940), .ZN(
        n11384) );
  AOI21_X1 U13799 ( .B1(n12269), .B2(n12889), .A(n11384), .ZN(n11385) );
  OAI211_X1 U13800 ( .C1(n12892), .C2(n14441), .A(n11386), .B(n11385), .ZN(
        P3_U3220) );
  INV_X1 U13801 ( .A(n11387), .ZN(n11389) );
  OAI222_X1 U13802 ( .A1(n13054), .A2(n11390), .B1(n13057), .B2(n11389), .C1(
        n11388), .C2(P3_U3151), .ZN(P3_U3270) );
  XNOR2_X1 U13803 ( .A(n13598), .B(n11604), .ZN(n11391) );
  NAND2_X1 U13804 ( .A1(n13200), .A2(n13492), .ZN(n11392) );
  NAND2_X1 U13805 ( .A1(n11391), .A2(n11392), .ZN(n11535) );
  INV_X1 U13806 ( .A(n11391), .ZN(n11394) );
  INV_X1 U13807 ( .A(n11392), .ZN(n11393) );
  NAND2_X1 U13808 ( .A1(n11394), .A2(n11393), .ZN(n11395) );
  NAND2_X1 U13809 ( .A1(n11535), .A2(n11395), .ZN(n11403) );
  INV_X1 U13810 ( .A(n11536), .ZN(n11401) );
  AOI21_X1 U13811 ( .B1(n11403), .B2(n11402), .A(n11401), .ZN(n11410) );
  OAI22_X1 U13812 ( .A1(n13149), .A2(n11405), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11404), .ZN(n11406) );
  AOI21_X1 U13813 ( .B1(n11407), .B2(n13151), .A(n11406), .ZN(n11409) );
  NAND2_X1 U13814 ( .A1(n13598), .A2(n13185), .ZN(n11408) );
  OAI211_X1 U13815 ( .C1(n11410), .C2(n13187), .A(n11409), .B(n11408), .ZN(
        P2_U3187) );
  INV_X1 U13816 ( .A(n11411), .ZN(n11412) );
  XNOR2_X1 U13817 ( .A(n11484), .B(n11492), .ZN(n13595) );
  INV_X1 U13818 ( .A(n13200), .ZN(n11539) );
  XNOR2_X1 U13819 ( .A(n11493), .B(n11492), .ZN(n11416) );
  OAI222_X1 U13820 ( .A1(n13447), .A2(n13117), .B1(n13445), .B2(n11539), .C1(
        n11416), .C2(n13451), .ZN(n13591) );
  AOI211_X1 U13821 ( .C1(n13593), .C2(n11417), .A(n13492), .B(n11487), .ZN(
        n13592) );
  INV_X1 U13822 ( .A(n13592), .ZN(n11419) );
  INV_X1 U13823 ( .A(n11418), .ZN(n11538) );
  OAI22_X1 U13824 ( .A1(n11419), .A2(n11500), .B1(n13473), .B2(n11538), .ZN(
        n11420) );
  OAI21_X1 U13825 ( .B1(n13591), .B2(n11420), .A(n13476), .ZN(n11422) );
  AOI22_X1 U13826 ( .A1(n13593), .A2(n13483), .B1(n13392), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n11421) );
  OAI211_X1 U13827 ( .C1(n13595), .C2(n13504), .A(n11422), .B(n11421), .ZN(
        P2_U3250) );
  INV_X1 U13828 ( .A(n13661), .ZN(n13936) );
  NAND2_X1 U13829 ( .A1(n14518), .A2(n13936), .ZN(n11424) );
  NAND2_X1 U13830 ( .A1(n11425), .A2(n12025), .ZN(n11427) );
  INV_X1 U13831 ( .A(n14026), .ZN(n14583) );
  AOI22_X1 U13832 ( .A1(n11646), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11645), 
        .B2(n14583), .ZN(n11426) );
  NAND2_X1 U13833 ( .A1(n14345), .A2(n13674), .ZN(n11925) );
  XNOR2_X1 U13834 ( .A(n11522), .B(n11523), .ZN(n14347) );
  INV_X1 U13835 ( .A(n11916), .ZN(n11428) );
  OAI211_X1 U13836 ( .C1(n6619), .C2(n12080), .A(n11512), .B(n14643), .ZN(
        n11439) );
  NAND2_X1 U13837 ( .A1(n6491), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U13838 ( .A1(n12006), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11437) );
  INV_X1 U13839 ( .A(n11431), .ZN(n11516) );
  INV_X1 U13840 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U13841 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  AND2_X1 U13842 ( .A1(n11516), .A2(n11434), .ZN(n13835) );
  NAND2_X1 U13843 ( .A1(n11743), .A2(n13835), .ZN(n11436) );
  NAND2_X1 U13844 ( .A1(n11039), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11435) );
  NAND4_X1 U13845 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n13934) );
  AOI22_X1 U13846 ( .A1(n13936), .A2(n13899), .B1(n13898), .B2(n13934), .ZN(
        n13917) );
  NAND2_X1 U13847 ( .A1(n11439), .A2(n13917), .ZN(n14343) );
  NAND2_X1 U13848 ( .A1(n14343), .A2(n14671), .ZN(n11446) );
  AOI21_X1 U13849 ( .B1(n14345), .B2(n11440), .A(n14683), .ZN(n11441) );
  AND2_X1 U13850 ( .A1(n11441), .A2(n11527), .ZN(n14344) );
  NAND2_X1 U13851 ( .A1(n14345), .A2(n14647), .ZN(n11443) );
  NAND2_X1 U13852 ( .A1(n14646), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11442) );
  OAI211_X1 U13853 ( .C1(n14662), .C2(n13916), .A(n11443), .B(n11442), .ZN(
        n11444) );
  AOI21_X1 U13854 ( .B1(n14344), .B2(n14654), .A(n11444), .ZN(n11445) );
  OAI211_X1 U13855 ( .C1(n14347), .C2(n14256), .A(n11446), .B(n11445), .ZN(
        P1_U3278) );
  INV_X1 U13856 ( .A(n11449), .ZN(n11450) );
  NAND2_X1 U13857 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  NAND2_X1 U13858 ( .A1(n14471), .A2(n13800), .ZN(n11454) );
  NAND2_X1 U13859 ( .A1(n13940), .A2(n6487), .ZN(n11453) );
  NAND2_X1 U13860 ( .A1(n11454), .A2(n11453), .ZN(n11455) );
  XNOR2_X1 U13861 ( .A(n11455), .B(n13752), .ZN(n11460) );
  AND2_X1 U13862 ( .A1(n13940), .A2(n13764), .ZN(n11456) );
  AOI21_X1 U13863 ( .B1(n14471), .B2(n9526), .A(n11456), .ZN(n11461) );
  XNOR2_X1 U13864 ( .A(n11460), .B(n11461), .ZN(n14477) );
  NAND2_X1 U13865 ( .A1(n14503), .A2(n13800), .ZN(n11458) );
  NAND2_X1 U13866 ( .A1(n13939), .A2(n6487), .ZN(n11457) );
  NAND2_X1 U13867 ( .A1(n11458), .A2(n11457), .ZN(n11459) );
  XNOR2_X1 U13868 ( .A(n11459), .B(n13798), .ZN(n11465) );
  AOI21_X1 U13869 ( .B1(n14503), .B2(n6487), .A(n6625), .ZN(n11466) );
  XNOR2_X1 U13870 ( .A(n11465), .B(n11466), .ZN(n14500) );
  INV_X1 U13871 ( .A(n11460), .ZN(n11463) );
  INV_X1 U13872 ( .A(n11461), .ZN(n11462) );
  NAND2_X1 U13873 ( .A1(n11463), .A2(n11462), .ZN(n14497) );
  AND2_X1 U13874 ( .A1(n14500), .A2(n14497), .ZN(n11464) );
  INV_X1 U13875 ( .A(n11465), .ZN(n11467) );
  NAND2_X1 U13876 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  NAND2_X1 U13877 ( .A1(n14424), .A2(n13800), .ZN(n11470) );
  NAND2_X1 U13878 ( .A1(n13938), .A2(n6487), .ZN(n11469) );
  NAND2_X1 U13879 ( .A1(n11470), .A2(n11469), .ZN(n11471) );
  XNOR2_X1 U13880 ( .A(n11471), .B(n13752), .ZN(n13648) );
  AND2_X1 U13881 ( .A1(n13938), .A2(n13764), .ZN(n11472) );
  AOI21_X1 U13882 ( .B1(n14424), .B2(n9526), .A(n11472), .ZN(n13649) );
  XNOR2_X1 U13883 ( .A(n13648), .B(n13649), .ZN(n11473) );
  AOI21_X1 U13884 ( .B1(n11474), .B2(n11473), .A(n14475), .ZN(n11475) );
  NAND2_X1 U13885 ( .A1(n11475), .A2(n13653), .ZN(n11481) );
  OAI21_X1 U13886 ( .B1(n11477), .B2(n14481), .A(n11476), .ZN(n11478) );
  AOI21_X1 U13887 ( .B1(n11479), .B2(n13904), .A(n11478), .ZN(n11480) );
  OAI211_X1 U13888 ( .C1(n11482), .C2(n13907), .A(n11481), .B(n11480), .ZN(
        P1_U3224) );
  NAND2_X1 U13889 ( .A1(n11484), .A2(n11483), .ZN(n11486) );
  OR2_X1 U13890 ( .A1(n13593), .A2(n13199), .ZN(n11485) );
  NAND2_X1 U13891 ( .A1(n11486), .A2(n11485), .ZN(n11812) );
  XNOR2_X1 U13892 ( .A(n11812), .B(n11811), .ZN(n13590) );
  INV_X1 U13893 ( .A(n11487), .ZN(n11490) );
  INV_X1 U13894 ( .A(n13587), .ZN(n11488) );
  NAND2_X1 U13895 ( .A1(n11488), .A2(n11487), .ZN(n13493) );
  INV_X1 U13896 ( .A(n13493), .ZN(n11489) );
  AOI211_X1 U13897 ( .C1(n13587), .C2(n11490), .A(n13492), .B(n11489), .ZN(
        n13585) );
  INV_X1 U13898 ( .A(n13585), .ZN(n11501) );
  INV_X1 U13899 ( .A(n13110), .ZN(n11491) );
  OAI22_X1 U13900 ( .A1(n13169), .A2(n13447), .B1(n11494), .B2(n13445), .ZN(
        n13586) );
  AOI21_X1 U13901 ( .B1(n13495), .B2(n11491), .A(n13586), .ZN(n11499) );
  NAND2_X1 U13902 ( .A1(n11493), .A2(n11492), .ZN(n11496) );
  OR2_X1 U13903 ( .A1(n13593), .A2(n11494), .ZN(n11495) );
  XNOR2_X1 U13904 ( .A(n11785), .B(n11497), .ZN(n11498) );
  NAND2_X1 U13905 ( .A1(n11498), .A2(n13488), .ZN(n13588) );
  OAI211_X1 U13906 ( .C1(n11501), .C2(n11500), .A(n11499), .B(n13588), .ZN(
        n11502) );
  NAND2_X1 U13907 ( .A1(n11502), .A2(n13476), .ZN(n11504) );
  AOI22_X1 U13908 ( .A1(n13587), .A2(n13483), .B1(n13392), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n11503) );
  OAI211_X1 U13909 ( .C1(n13590), .C2(n13504), .A(n11504), .B(n11503), .ZN(
        P2_U3249) );
  INV_X1 U13910 ( .A(n11714), .ZN(n11507) );
  OAI222_X1 U13911 ( .A1(n13636), .A2(n15202), .B1(n13637), .B2(n11507), .C1(
        n11505), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U13912 ( .A(n11506), .ZN(n11508) );
  OAI222_X1 U13913 ( .A1(P1_U3086), .A2(n11508), .B1(n14382), .B2(n11507), 
        .C1(n11715), .C2(n14379), .ZN(P1_U3330) );
  NAND2_X1 U13914 ( .A1(n11509), .A2(n12025), .ZN(n11511) );
  INV_X1 U13915 ( .A(n14596), .ZN(n14030) );
  AOI22_X1 U13916 ( .A1(n11646), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11645), 
        .B2(n14030), .ZN(n11510) );
  INV_X1 U13917 ( .A(n13934), .ZN(n13847) );
  XNOR2_X1 U13918 ( .A(n13839), .B(n13847), .ZN(n12083) );
  XOR2_X1 U13919 ( .A(n12083), .B(n11759), .Z(n11521) );
  INV_X1 U13920 ( .A(n13674), .ZN(n13935) );
  INV_X1 U13921 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U13922 ( .A1(n6491), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U13923 ( .A1(n12006), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11513) );
  AND2_X1 U13924 ( .A1(n11514), .A2(n11513), .ZN(n11520) );
  INV_X1 U13925 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U13926 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U13927 ( .A1(n11518), .A2(n11517), .ZN(n14249) );
  OR2_X1 U13928 ( .A1(n14249), .A2(n11720), .ZN(n11519) );
  OAI211_X1 U13929 ( .C1(n11656), .C2(n14032), .A(n11520), .B(n11519), .ZN(
        n13933) );
  AOI22_X1 U13930 ( .A1(n13935), .A2(n13899), .B1(n13898), .B2(n13933), .ZN(
        n13837) );
  OAI21_X1 U13931 ( .B1(n11521), .B2(n14676), .A(n13837), .ZN(n14514) );
  INV_X1 U13932 ( .A(n14514), .ZN(n11534) );
  INV_X1 U13933 ( .A(n12080), .ZN(n11523) );
  OR2_X1 U13934 ( .A1(n14345), .A2(n13935), .ZN(n11524) );
  OAI21_X1 U13935 ( .B1(n6742), .B2(n12083), .A(n11633), .ZN(n14516) );
  INV_X1 U13936 ( .A(n13839), .ZN(n14513) );
  INV_X1 U13937 ( .A(n11527), .ZN(n11529) );
  INV_X1 U13938 ( .A(n14245), .ZN(n11528) );
  OAI211_X1 U13939 ( .C1(n14513), .C2(n11529), .A(n11528), .B(n14651), .ZN(
        n14512) );
  AOI22_X1 U13940 ( .A1(n14646), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13835), 
        .B2(n14645), .ZN(n11531) );
  NAND2_X1 U13941 ( .A1(n13839), .A2(n14647), .ZN(n11530) );
  OAI211_X1 U13942 ( .C1(n14512), .C2(n14234), .A(n11531), .B(n11530), .ZN(
        n11532) );
  AOI21_X1 U13943 ( .B1(n14516), .B2(n14668), .A(n11532), .ZN(n11533) );
  OAI21_X1 U13944 ( .B1(n11534), .B2(n14646), .A(n11533), .ZN(P1_U3277) );
  XOR2_X1 U13945 ( .A(n11612), .B(n13593), .Z(n11569) );
  NAND2_X1 U13946 ( .A1(n13199), .A2(n13492), .ZN(n11570) );
  XNOR2_X1 U13947 ( .A(n11571), .B(n11570), .ZN(n11543) );
  OAI22_X1 U13948 ( .A1(n13183), .A2(n11538), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11537), .ZN(n11541) );
  OAI22_X1 U13949 ( .A1(n11539), .A2(n13139), .B1(n13138), .B2(n13117), .ZN(
        n11540) );
  AOI211_X1 U13950 ( .C1(n13593), .C2(n13185), .A(n11541), .B(n11540), .ZN(
        n11542) );
  OAI21_X1 U13951 ( .B1(n11543), .B2(n13187), .A(n11542), .ZN(P2_U3213) );
  NOR2_X1 U13952 ( .A1(n11544), .A2(n14660), .ZN(n11545) );
  OR2_X1 U13953 ( .A1(n11546), .A2(n11545), .ZN(n14684) );
  XNOR2_X1 U13954 ( .A(n14684), .B(n11547), .ZN(n11548) );
  MUX2_X1 U13955 ( .A(n11548), .B(n12063), .S(n11844), .Z(n11554) );
  NAND2_X1 U13956 ( .A1(n12063), .A2(n11549), .ZN(n11550) );
  NAND2_X1 U13957 ( .A1(n11551), .A2(n11550), .ZN(n14687) );
  AOI21_X1 U13958 ( .B1(n14687), .B2(n14723), .A(n11552), .ZN(n11553) );
  OAI21_X1 U13959 ( .B1(n11554), .B2(n14676), .A(n11553), .ZN(n14685) );
  MUX2_X1 U13960 ( .A(n14685), .B(P1_REG2_REG_1__SCAN_IN), .S(n14646), .Z(
        n11561) );
  NAND2_X1 U13961 ( .A1(n14687), .A2(n14655), .ZN(n11559) );
  AOI22_X1 U13962 ( .A1(n14647), .A2(n11555), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14645), .ZN(n11558) );
  INV_X1 U13963 ( .A(n14684), .ZN(n11556) );
  NAND3_X1 U13964 ( .A1(n14654), .A2(n11556), .A3(n14651), .ZN(n11557) );
  NAND3_X1 U13965 ( .A1(n11559), .A2(n11558), .A3(n11557), .ZN(n11560) );
  OR2_X1 U13966 ( .A1(n11561), .A2(n11560), .ZN(P1_U3292) );
  OAI222_X1 U13967 ( .A1(n14382), .A2(n12012), .B1(n11562), .B2(P1_U3086), 
        .C1(n12472), .C2(n14379), .ZN(P1_U3325) );
  INV_X1 U13968 ( .A(n11737), .ZN(n14377) );
  OAI222_X1 U13969 ( .A1(n13636), .A2(n11563), .B1(n13637), .B2(n14377), .C1(
        P2_U3088), .C2(n6719), .ZN(P2_U3300) );
  INV_X1 U13970 ( .A(n11564), .ZN(n11565) );
  OAI222_X1 U13971 ( .A1(n13637), .A2(n12012), .B1(P2_U3088), .B2(n11566), 
        .C1(n7022), .C2(n13636), .ZN(P2_U3297) );
  XNOR2_X1 U13972 ( .A(n13587), .B(n11604), .ZN(n11573) );
  NAND2_X1 U13973 ( .A1(n13198), .A2(n13492), .ZN(n11572) );
  NAND2_X1 U13974 ( .A1(n11573), .A2(n11572), .ZN(n11574) );
  OAI21_X1 U13975 ( .B1(n11573), .B2(n11572), .A(n11574), .ZN(n13108) );
  INV_X1 U13976 ( .A(n11574), .ZN(n11575) );
  XNOR2_X1 U13977 ( .A(n13581), .B(n11604), .ZN(n11577) );
  NAND2_X1 U13978 ( .A1(n13197), .A2(n13492), .ZN(n11576) );
  NAND2_X1 U13979 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  OAI21_X1 U13980 ( .B1(n11577), .B2(n11576), .A(n11578), .ZN(n13115) );
  INV_X1 U13981 ( .A(n11578), .ZN(n11579) );
  XNOR2_X1 U13982 ( .A(n13576), .B(n11612), .ZN(n11582) );
  NAND2_X1 U13983 ( .A1(n13196), .A2(n13492), .ZN(n11580) );
  XNOR2_X1 U13984 ( .A(n11582), .B(n11580), .ZN(n13167) );
  INV_X1 U13985 ( .A(n11580), .ZN(n11581) );
  XNOR2_X1 U13986 ( .A(n13571), .B(n11612), .ZN(n11585) );
  AND2_X1 U13987 ( .A1(n13436), .A2(n13492), .ZN(n11584) );
  NOR2_X1 U13988 ( .A1(n11585), .A2(n11584), .ZN(n13072) );
  NAND2_X1 U13989 ( .A1(n11585), .A2(n11584), .ZN(n13073) );
  XNOR2_X1 U13990 ( .A(n13565), .B(n11604), .ZN(n11587) );
  NAND2_X1 U13991 ( .A1(n13195), .A2(n13492), .ZN(n11586) );
  NAND2_X1 U13992 ( .A1(n11587), .A2(n11586), .ZN(n13131) );
  NOR2_X1 U13993 ( .A1(n11587), .A2(n11586), .ZN(n13133) );
  NAND2_X1 U13994 ( .A1(n13438), .A2(n13492), .ZN(n11589) );
  XNOR2_X1 U13995 ( .A(n13561), .B(n11612), .ZN(n11588) );
  XOR2_X1 U13996 ( .A(n11589), .B(n11588), .Z(n13089) );
  INV_X1 U13997 ( .A(n11588), .ZN(n11590) );
  INV_X1 U13998 ( .A(n11591), .ZN(n11594) );
  XNOR2_X1 U13999 ( .A(n13557), .B(n11612), .ZN(n11592) );
  XNOR2_X1 U14000 ( .A(n11594), .B(n11592), .ZN(n13146) );
  NAND2_X1 U14001 ( .A1(n13375), .A2(n13492), .ZN(n13145) );
  NAND2_X1 U14002 ( .A1(n13146), .A2(n13145), .ZN(n13144) );
  INV_X1 U14003 ( .A(n11592), .ZN(n11593) );
  NAND2_X1 U14004 ( .A1(n13144), .A2(n11595), .ZN(n11596) );
  XNOR2_X1 U14005 ( .A(n13549), .B(n11612), .ZN(n11597) );
  NAND2_X1 U14006 ( .A1(n13194), .A2(n13492), .ZN(n13066) );
  XNOR2_X1 U14007 ( .A(n13369), .B(n11612), .ZN(n11600) );
  NAND2_X1 U14008 ( .A1(n13377), .A2(n13492), .ZN(n11598) );
  XNOR2_X1 U14009 ( .A(n11600), .B(n11598), .ZN(n13124) );
  INV_X1 U14010 ( .A(n11598), .ZN(n11599) );
  AND2_X1 U14011 ( .A1(n11600), .A2(n11599), .ZN(n11601) );
  XNOR2_X1 U14012 ( .A(n13537), .B(n11612), .ZN(n11602) );
  NOR2_X1 U14013 ( .A1(n13180), .A2(n10055), .ZN(n11603) );
  XNOR2_X1 U14014 ( .A(n11602), .B(n11603), .ZN(n13097) );
  XNOR2_X1 U14015 ( .A(n13532), .B(n11604), .ZN(n11606) );
  NAND2_X1 U14016 ( .A1(n13192), .A2(n13492), .ZN(n11605) );
  NAND2_X1 U14017 ( .A1(n11606), .A2(n11605), .ZN(n11607) );
  OAI21_X1 U14018 ( .B1(n11606), .B2(n11605), .A(n11607), .ZN(n13178) );
  NAND2_X1 U14019 ( .A1(n13191), .A2(n13492), .ZN(n11609) );
  XNOR2_X1 U14020 ( .A(n13526), .B(n11612), .ZN(n11608) );
  XOR2_X1 U14021 ( .A(n11609), .B(n11608), .Z(n13061) );
  INV_X1 U14022 ( .A(n11608), .ZN(n11610) );
  NAND2_X1 U14023 ( .A1(n13190), .A2(n13492), .ZN(n11611) );
  XOR2_X1 U14024 ( .A(n11612), .B(n11611), .Z(n11613) );
  XNOR2_X1 U14025 ( .A(n13520), .B(n11613), .ZN(n11614) );
  XNOR2_X1 U14026 ( .A(n11615), .B(n11614), .ZN(n11616) );
  NAND2_X1 U14027 ( .A1(n11616), .A2(n13162), .ZN(n11621) );
  OAI22_X1 U14028 ( .A1(n13312), .A2(n13183), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11617), .ZN(n11619) );
  INV_X1 U14029 ( .A(n13191), .ZN(n13306) );
  OAI22_X1 U14030 ( .A1(n13306), .A2(n13139), .B1(n13305), .B2(n13138), .ZN(
        n11618) );
  AOI211_X1 U14031 ( .C1(n13520), .C2(n13173), .A(n11619), .B(n11618), .ZN(
        n11620) );
  NAND2_X1 U14032 ( .A1(n11621), .A2(n11620), .ZN(P2_U3192) );
  NAND2_X1 U14033 ( .A1(n13629), .A2(n12025), .ZN(n11624) );
  OR2_X1 U14034 ( .A1(n12013), .A2(n11622), .ZN(n11623) );
  INV_X1 U14035 ( .A(n13804), .ZN(n11625) );
  NAND2_X1 U14036 ( .A1(n6491), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U14037 ( .A1(n12006), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11628) );
  INV_X1 U14038 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13807) );
  XNOR2_X1 U14039 ( .A(n11742), .B(n13807), .ZN(n14074) );
  NAND2_X1 U14040 ( .A1(n11743), .A2(n14074), .ZN(n11627) );
  NAND2_X1 U14041 ( .A1(n11039), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11626) );
  NAND4_X1 U14042 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n13923) );
  OR2_X1 U14043 ( .A1(n12013), .A2(n14374), .ZN(n11630) );
  OR2_X1 U14044 ( .A1(n13839), .A2(n13934), .ZN(n11632) );
  NAND2_X1 U14045 ( .A1(n11634), .A2(n12025), .ZN(n11636) );
  AOI22_X1 U14046 ( .A1(n11646), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11645), 
        .B2(n14033), .ZN(n11635) );
  INV_X1 U14047 ( .A(n13933), .ZN(n13681) );
  AND2_X1 U14048 ( .A1(n14246), .A2(n13681), .ZN(n11637) );
  NAND2_X1 U14049 ( .A1(n11638), .A2(n12025), .ZN(n11640) );
  AOI22_X1 U14050 ( .A1(n11646), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11645), 
        .B2(n14624), .ZN(n11639) );
  NAND2_X2 U14051 ( .A1(n11640), .A2(n11639), .ZN(n14232) );
  OR2_X1 U14052 ( .A1(n14232), .A2(n13691), .ZN(n11641) );
  NAND2_X1 U14053 ( .A1(n14232), .A2(n13691), .ZN(n11642) );
  INV_X1 U14054 ( .A(n14209), .ZN(n11658) );
  NAND2_X1 U14055 ( .A1(n11644), .A2(n12025), .ZN(n11648) );
  AOI22_X1 U14056 ( .A1(n11646), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11835), 
        .B2(n11645), .ZN(n11647) );
  INV_X1 U14057 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14038) );
  INV_X1 U14058 ( .A(n11663), .ZN(n11652) );
  NAND2_X1 U14059 ( .A1(n11650), .A2(n11649), .ZN(n11651) );
  NAND2_X1 U14060 ( .A1(n11652), .A2(n11651), .ZN(n14214) );
  OR2_X1 U14061 ( .A1(n14214), .A2(n11720), .ZN(n11655) );
  AOI22_X1 U14062 ( .A1(n6491), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n12006), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n11654) );
  OAI211_X1 U14063 ( .C1(n11656), .C2(n14038), .A(n11655), .B(n11654), .ZN(
        n13932) );
  XNOR2_X1 U14064 ( .A(n14327), .B(n13932), .ZN(n14216) );
  OR2_X1 U14065 ( .A1(n12013), .A2(n11660), .ZN(n11661) );
  NAND2_X2 U14066 ( .A1(n11662), .A2(n11661), .ZN(n14319) );
  NOR2_X1 U14067 ( .A1(n11663), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11664) );
  OR2_X1 U14068 ( .A1(n11675), .A2(n11664), .ZN(n13868) );
  OR2_X1 U14069 ( .A1(n13868), .A2(n11720), .ZN(n11670) );
  INV_X1 U14070 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U14071 ( .A1(n12006), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14072 ( .A1(n11039), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11665) );
  OAI211_X1 U14073 ( .C1(n11667), .C2(n12009), .A(n11666), .B(n11665), .ZN(
        n11668) );
  INV_X1 U14074 ( .A(n11668), .ZN(n11669) );
  NAND2_X1 U14075 ( .A1(n11670), .A2(n11669), .ZN(n13931) );
  INV_X1 U14076 ( .A(n13931), .ZN(n13792) );
  XNOR2_X1 U14077 ( .A(n14319), .B(n13792), .ZN(n14204) );
  NAND2_X1 U14078 ( .A1(n14319), .A2(n13931), .ZN(n11671) );
  OR2_X1 U14079 ( .A1(n11672), .A2(n6686), .ZN(n11674) );
  OR2_X1 U14080 ( .A1(n12023), .A2(n15204), .ZN(n11673) );
  OR2_X1 U14081 ( .A1(n11675), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14082 ( .A1(n11676), .A2(n11687), .ZN(n14189) );
  OR2_X1 U14083 ( .A1(n14189), .A2(n11720), .ZN(n11681) );
  INV_X1 U14084 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U14085 ( .A1(n11039), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U14086 ( .A1(n12006), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11677) );
  OAI211_X1 U14087 ( .C1(n12009), .C2(n14188), .A(n11678), .B(n11677), .ZN(
        n11679) );
  INV_X1 U14088 ( .A(n11679), .ZN(n11680) );
  NAND2_X1 U14089 ( .A1(n11681), .A2(n11680), .ZN(n13930) );
  XNOR2_X1 U14090 ( .A(n14314), .B(n13930), .ZN(n14181) );
  OR2_X1 U14091 ( .A1(n11683), .A2(n9517), .ZN(n11684) );
  XNOR2_X1 U14092 ( .A(n11684), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14384) );
  NAND2_X1 U14093 ( .A1(n6491), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14094 ( .A1(n12006), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11690) );
  INV_X1 U14095 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13880) );
  AOI21_X1 U14096 ( .B1(n13880), .B2(n11687), .A(n11686), .ZN(n14171) );
  NAND2_X1 U14097 ( .A1(n11743), .A2(n14171), .ZN(n11689) );
  NAND2_X1 U14098 ( .A1(n11039), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11688) );
  NAND4_X1 U14099 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n13929) );
  INV_X1 U14100 ( .A(n13929), .ZN(n11767) );
  XNOR2_X1 U14101 ( .A(n14174), .B(n11767), .ZN(n14162) );
  INV_X1 U14102 ( .A(n14162), .ZN(n14167) );
  OR2_X1 U14103 ( .A1(n14308), .A2(n13929), .ZN(n11692) );
  NAND2_X1 U14104 ( .A1(n14166), .A2(n11692), .ZN(n14149) );
  OR2_X1 U14105 ( .A1(n11693), .A2(n6686), .ZN(n11696) );
  OR2_X1 U14106 ( .A1(n12013), .A2(n11694), .ZN(n11695) );
  NAND2_X1 U14107 ( .A1(n6491), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U14108 ( .A1(n12006), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11700) );
  INV_X1 U14109 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13784) );
  AOI21_X1 U14110 ( .B1(n13784), .B2(n11697), .A(n11708), .ZN(n14153) );
  NAND2_X1 U14111 ( .A1(n11743), .A2(n14153), .ZN(n11699) );
  NAND2_X1 U14112 ( .A1(n11039), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U14113 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n13928) );
  INV_X1 U14114 ( .A(n13928), .ZN(n11769) );
  XNOR2_X1 U14115 ( .A(n14156), .B(n11769), .ZN(n14145) );
  INV_X1 U14116 ( .A(n14145), .ZN(n14150) );
  NAND2_X1 U14117 ( .A1(n14156), .A2(n13928), .ZN(n11702) );
  OR2_X1 U14118 ( .A1(n11703), .A2(n6686), .ZN(n11706) );
  OR2_X1 U14119 ( .A1(n12023), .A2(n11704), .ZN(n11705) );
  OAI21_X1 U14120 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11708), .A(n11707), 
        .ZN(n14134) );
  OR2_X1 U14121 ( .A1(n11720), .A2(n14134), .ZN(n11712) );
  NAND2_X1 U14122 ( .A1(n6491), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U14123 ( .A1(n12006), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14124 ( .A1(n11039), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14125 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n13927) );
  INV_X1 U14126 ( .A(n13927), .ZN(n11770) );
  XNOR2_X1 U14127 ( .A(n14295), .B(n11770), .ZN(n14127) );
  INV_X1 U14128 ( .A(n14127), .ZN(n14137) );
  OR2_X1 U14129 ( .A1(n14295), .A2(n13927), .ZN(n11713) );
  NAND2_X1 U14130 ( .A1(n11714), .A2(n12025), .ZN(n11717) );
  OR2_X1 U14131 ( .A1(n12013), .A2(n11715), .ZN(n11716) );
  INV_X1 U14132 ( .A(n11718), .ZN(n11728) );
  OAI21_X1 U14133 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11719), .A(n11728), 
        .ZN(n14121) );
  OR2_X1 U14134 ( .A1(n11720), .A2(n14121), .ZN(n11724) );
  NAND2_X1 U14135 ( .A1(n6491), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11723) );
  NAND2_X1 U14136 ( .A1(n12006), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U14137 ( .A1(n11039), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11721) );
  NAND4_X1 U14138 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n13926) );
  INV_X1 U14139 ( .A(n13926), .ZN(n11772) );
  XNOR2_X1 U14140 ( .A(n14290), .B(n11772), .ZN(n14113) );
  NAND2_X1 U14141 ( .A1(n14290), .A2(n13926), .ZN(n11725) );
  NAND2_X1 U14142 ( .A1(n13635), .A2(n12025), .ZN(n11727) );
  OR2_X1 U14143 ( .A1(n12013), .A2(n14380), .ZN(n11726) );
  NAND2_X1 U14144 ( .A1(n6491), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11734) );
  NAND2_X1 U14145 ( .A1(n12006), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11733) );
  INV_X1 U14146 ( .A(n11740), .ZN(n11730) );
  INV_X1 U14147 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13902) );
  NAND2_X1 U14148 ( .A1(n11728), .A2(n13902), .ZN(n11729) );
  NAND2_X1 U14149 ( .A1(n11743), .A2(n14099), .ZN(n11732) );
  NAND2_X1 U14150 ( .A1(n11039), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11731) );
  NAND4_X1 U14151 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n13925) );
  INV_X1 U14152 ( .A(n13925), .ZN(n11774) );
  XNOR2_X1 U14153 ( .A(n14283), .B(n11774), .ZN(n14100) );
  NAND2_X1 U14154 ( .A1(n14098), .A2(n14100), .ZN(n11736) );
  NAND2_X1 U14155 ( .A1(n14283), .A2(n13925), .ZN(n11735) );
  NAND2_X1 U14156 ( .A1(n11737), .A2(n12025), .ZN(n11739) );
  OR2_X1 U14157 ( .A1(n12013), .A2(n7036), .ZN(n11738) );
  NAND2_X1 U14158 ( .A1(n12006), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14159 ( .A1(n6491), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11746) );
  NOR2_X1 U14160 ( .A1(n11740), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11741) );
  NOR2_X1 U14161 ( .A1(n11742), .A2(n11741), .ZN(n14092) );
  NAND2_X1 U14162 ( .A1(n11743), .A2(n14092), .ZN(n11745) );
  NAND2_X1 U14163 ( .A1(n11039), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11744) );
  NAND4_X1 U14164 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n13924) );
  INV_X1 U14165 ( .A(n13924), .ZN(n11776) );
  OR2_X1 U14166 ( .A1(n14093), .A2(n13924), .ZN(n11748) );
  OR2_X2 U14167 ( .A1(n14210), .A2(n14319), .ZN(n14199) );
  NAND2_X1 U14168 ( .A1(n14174), .A2(n14187), .ZN(n14151) );
  NOR2_X2 U14169 ( .A1(n14266), .A2(n14072), .ZN(n14060) );
  AOI211_X1 U14170 ( .C1(n14266), .C2(n14072), .A(n14683), .B(n14060), .ZN(
        n14264) );
  AOI21_X1 U14171 ( .B1(n11750), .B2(P1_B_REG_SCAN_IN), .A(n13848), .ZN(n14055) );
  INV_X1 U14172 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14061) );
  NAND2_X1 U14173 ( .A1(n9188), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14174 ( .A1(n12006), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11751) );
  OAI211_X1 U14175 ( .C1(n12009), .C2(n14061), .A(n11752), .B(n11751), .ZN(
        n13922) );
  NAND2_X1 U14176 ( .A1(n14055), .A2(n13922), .ZN(n14263) );
  NAND2_X1 U14177 ( .A1(n14266), .A2(n14647), .ZN(n11756) );
  INV_X1 U14178 ( .A(n11753), .ZN(n11754) );
  AOI22_X1 U14179 ( .A1(n14646), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n14645), 
        .B2(n11754), .ZN(n11755) );
  OAI211_X1 U14180 ( .C1(n11757), .C2(n14263), .A(n11756), .B(n11755), .ZN(
        n11758) );
  AOI21_X1 U14181 ( .B1(n14264), .B2(n14654), .A(n11758), .ZN(n11784) );
  NAND2_X1 U14182 ( .A1(n14340), .A2(n13681), .ZN(n11760) );
  NAND2_X1 U14183 ( .A1(n11761), .A2(n11760), .ZN(n12082) );
  NAND2_X1 U14184 ( .A1(n14240), .A2(n14241), .ZN(n14239) );
  NAND2_X1 U14185 ( .A1(n14232), .A2(n13849), .ZN(n11950) );
  INV_X1 U14186 ( .A(n13932), .ZN(n11762) );
  NAND2_X1 U14187 ( .A1(n14327), .A2(n11762), .ZN(n11763) );
  OR2_X1 U14188 ( .A1(n13792), .A2(n14319), .ZN(n11764) );
  INV_X1 U14189 ( .A(n13930), .ZN(n11765) );
  OR2_X1 U14190 ( .A1(n14314), .A2(n11765), .ZN(n14160) );
  AND2_X1 U14191 ( .A1(n14162), .A2(n14160), .ZN(n11766) );
  NAND2_X1 U14192 ( .A1(n14308), .A2(n11767), .ZN(n11768) );
  OR2_X1 U14193 ( .A1(n14295), .A2(n11770), .ZN(n11771) );
  OR2_X2 U14194 ( .A1(n14112), .A2(n14113), .ZN(n14114) );
  NAND2_X1 U14195 ( .A1(n14290), .A2(n11772), .ZN(n11773) );
  AND2_X1 U14196 ( .A1(n14283), .A2(n11774), .ZN(n11775) );
  INV_X1 U14197 ( .A(n14270), .ZN(n11777) );
  NAND2_X1 U14198 ( .A1(n11777), .A2(n13923), .ZN(n11779) );
  INV_X1 U14199 ( .A(n13923), .ZN(n11778) );
  XNOR2_X1 U14200 ( .A(n11780), .B(n12089), .ZN(n11781) );
  NAND2_X1 U14201 ( .A1(n13923), .A2(n13899), .ZN(n14262) );
  AOI21_X1 U14202 ( .B1(n14267), .B2(n14262), .A(n14646), .ZN(n11782) );
  INV_X1 U14203 ( .A(n11782), .ZN(n11783) );
  OAI211_X1 U14204 ( .C1(n14269), .C2(n14256), .A(n11784), .B(n11783), .ZN(
        P1_U3356) );
  INV_X1 U14205 ( .A(n13520), .ZN(n11797) );
  NAND2_X1 U14206 ( .A1(n11785), .A2(n11811), .ZN(n11787) );
  OR2_X1 U14207 ( .A1(n13587), .A2(n13117), .ZN(n11786) );
  NAND2_X1 U14208 ( .A1(n13581), .A2(n13169), .ZN(n11788) );
  AND2_X1 U14209 ( .A1(n13576), .A2(n13446), .ZN(n11790) );
  OR2_X1 U14210 ( .A1(n13576), .A2(n13446), .ZN(n11791) );
  INV_X1 U14211 ( .A(n13432), .ZN(n11792) );
  NAND2_X1 U14212 ( .A1(n13565), .A2(n13448), .ZN(n11794) );
  OR2_X1 U14213 ( .A1(n13561), .A2(n13137), .ZN(n11795) );
  NAND2_X1 U14214 ( .A1(n13561), .A2(n13137), .ZN(n11796) );
  INV_X1 U14215 ( .A(n13353), .ZN(n13344) );
  INV_X1 U14216 ( .A(n13192), .ZN(n13100) );
  INV_X1 U14217 ( .A(n13526), .ZN(n11821) );
  NAND2_X1 U14218 ( .A1(n13190), .A2(n13435), .ZN(n11803) );
  INV_X1 U14219 ( .A(n6719), .ZN(n11801) );
  AOI21_X1 U14220 ( .B1(n11801), .B2(P2_B_REG_SCAN_IN), .A(n13447), .ZN(n13293) );
  NAND2_X1 U14221 ( .A1(n13293), .A2(n13189), .ZN(n11802) );
  OR2_X2 U14222 ( .A1(n13493), .A2(n13581), .ZN(n13490) );
  NAND2_X1 U14223 ( .A1(n13549), .A2(n13399), .ZN(n13374) );
  NOR2_X2 U14224 ( .A1(n13369), .A2(n13374), .ZN(n13365) );
  NAND2_X1 U14225 ( .A1(n13352), .A2(n13365), .ZN(n13349) );
  AOI211_X1 U14226 ( .C1(n13515), .C2(n13309), .A(n13492), .B(n13297), .ZN(
        n13514) );
  INV_X1 U14227 ( .A(n11806), .ZN(n11807) );
  AOI22_X1 U14228 ( .A1(n11807), .A2(n13495), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13509), .ZN(n11808) );
  OAI21_X1 U14229 ( .B1(n11809), .B2(n13498), .A(n11808), .ZN(n11825) );
  NAND2_X1 U14230 ( .A1(n13587), .A2(n13198), .ZN(n11810) );
  NAND2_X1 U14231 ( .A1(n13581), .A2(n13197), .ZN(n11813) );
  OR2_X1 U14232 ( .A1(n13576), .A2(n13196), .ZN(n11815) );
  NOR2_X1 U14233 ( .A1(n13571), .A2(n13436), .ZN(n11816) );
  INV_X1 U14234 ( .A(n13411), .ZN(n13413) );
  INV_X1 U14235 ( .A(n13393), .ZN(n13405) );
  NOR2_X1 U14236 ( .A1(n13537), .A2(n13193), .ZN(n11817) );
  NAND2_X1 U14237 ( .A1(n13532), .A2(n13192), .ZN(n11819) );
  OAI21_X1 U14238 ( .B1(n13517), .B2(n13509), .A(n11826), .ZN(P2_U3236) );
  OAI21_X1 U14239 ( .B1(n11829), .B2(n11828), .A(n11827), .ZN(n11830) );
  NAND2_X1 U14240 ( .A1(n11830), .A2(n14504), .ZN(n11834) );
  AOI22_X1 U14241 ( .A1(n11832), .A2(n14506), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n11831), .ZN(n11833) );
  OAI211_X1 U14242 ( .C1(n11848), .C2(n13907), .A(n11834), .B(n11833), .ZN(
        P1_U3237) );
  NAND2_X1 U14243 ( .A1(n11837), .A2(n11836), .ZN(n12018) );
  MUX2_X1 U14244 ( .A(n12037), .B(n12036), .S(n12018), .Z(n11846) );
  NAND2_X1 U14245 ( .A1(n13949), .A2(n11846), .ZN(n11838) );
  NAND2_X1 U14246 ( .A1(n11840), .A2(n11953), .ZN(n11841) );
  NOR2_X1 U14247 ( .A1(n13949), .A2(n12026), .ZN(n11842) );
  NAND2_X1 U14248 ( .A1(n11842), .A2(n11849), .ZN(n11843) );
  NAND2_X1 U14249 ( .A1(n11844), .A2(n14660), .ZN(n12060) );
  AND2_X1 U14250 ( .A1(n12060), .A2(n11845), .ZN(n11853) );
  AND2_X1 U14251 ( .A1(n11847), .A2(n12026), .ZN(n11851) );
  NAND2_X1 U14252 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  OAI211_X1 U14253 ( .C1(n11853), .C2(n11852), .A(n11851), .B(n11850), .ZN(
        n11855) );
  AOI21_X1 U14254 ( .B1(n11856), .B2(n11855), .A(n11854), .ZN(n11861) );
  AND2_X1 U14255 ( .A1(n13947), .A2(n11953), .ZN(n11859) );
  NOR2_X1 U14256 ( .A1(n13947), .A2(n11953), .ZN(n11858) );
  MUX2_X1 U14257 ( .A(n11859), .B(n11858), .S(n11857), .Z(n11860) );
  MUX2_X1 U14258 ( .A(n13946), .B(n11862), .S(n12026), .Z(n11863) );
  MUX2_X1 U14259 ( .A(n13946), .B(n11862), .S(n11953), .Z(n11864) );
  MUX2_X1 U14260 ( .A(n11866), .B(n11865), .S(n11953), .Z(n11870) );
  INV_X1 U14261 ( .A(n11870), .ZN(n11867) );
  MUX2_X1 U14262 ( .A(n13945), .B(n14690), .S(n12026), .Z(n11868) );
  NAND2_X1 U14263 ( .A1(n11869), .A2(n11868), .ZN(n11872) );
  MUX2_X1 U14264 ( .A(n13944), .B(n14648), .S(n12026), .Z(n11873) );
  MUX2_X1 U14265 ( .A(n13944), .B(n14648), .S(n11953), .Z(n11874) );
  MUX2_X1 U14266 ( .A(n13943), .B(n11875), .S(n11953), .Z(n11879) );
  MUX2_X1 U14267 ( .A(n13943), .B(n11875), .S(n11998), .Z(n11876) );
  NAND2_X1 U14268 ( .A1(n11877), .A2(n11876), .ZN(n11890) );
  INV_X1 U14269 ( .A(n11878), .ZN(n11881) );
  INV_X1 U14270 ( .A(n11879), .ZN(n11880) );
  NAND2_X1 U14271 ( .A1(n11881), .A2(n11880), .ZN(n11887) );
  NAND2_X1 U14272 ( .A1(n11890), .A2(n11887), .ZN(n11882) );
  MUX2_X1 U14273 ( .A(n13942), .B(n11883), .S(n12026), .Z(n11886) );
  NAND2_X1 U14274 ( .A1(n11882), .A2(n11886), .ZN(n11885) );
  MUX2_X1 U14275 ( .A(n13942), .B(n11883), .S(n11953), .Z(n11884) );
  NAND2_X1 U14276 ( .A1(n11885), .A2(n11884), .ZN(n11892) );
  INV_X1 U14277 ( .A(n11886), .ZN(n11888) );
  AND2_X1 U14278 ( .A1(n11888), .A2(n11887), .ZN(n11889) );
  NAND2_X1 U14279 ( .A1(n11890), .A2(n11889), .ZN(n11891) );
  NAND2_X1 U14280 ( .A1(n11892), .A2(n11891), .ZN(n11896) );
  INV_X1 U14281 ( .A(n12026), .ZN(n11999) );
  MUX2_X1 U14282 ( .A(n13941), .B(n11893), .S(n11999), .Z(n11897) );
  NAND2_X1 U14283 ( .A1(n11896), .A2(n11897), .ZN(n11895) );
  MUX2_X1 U14284 ( .A(n13941), .B(n11893), .S(n12026), .Z(n11894) );
  NAND2_X1 U14285 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  INV_X1 U14286 ( .A(n11896), .ZN(n11899) );
  INV_X1 U14287 ( .A(n11897), .ZN(n11898) );
  NAND2_X1 U14288 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  MUX2_X1 U14289 ( .A(n13940), .B(n14471), .S(n11998), .Z(n11904) );
  MUX2_X1 U14290 ( .A(n13940), .B(n14471), .S(n11999), .Z(n11902) );
  INV_X1 U14291 ( .A(n11904), .ZN(n11905) );
  MUX2_X1 U14292 ( .A(n13939), .B(n14503), .S(n11999), .Z(n11908) );
  MUX2_X1 U14293 ( .A(n13939), .B(n14503), .S(n11998), .Z(n11906) );
  NAND2_X1 U14294 ( .A1(n11907), .A2(n11906), .ZN(n11910) );
  MUX2_X1 U14295 ( .A(n13938), .B(n14424), .S(n11998), .Z(n11912) );
  MUX2_X1 U14296 ( .A(n13938), .B(n14424), .S(n11999), .Z(n11911) );
  MUX2_X1 U14297 ( .A(n13937), .B(n14492), .S(n11999), .Z(n11917) );
  MUX2_X1 U14298 ( .A(n11914), .B(n11913), .S(n11998), .Z(n11915) );
  OAI21_X1 U14299 ( .B1(n11918), .B2(n11917), .A(n11915), .ZN(n11920) );
  AOI21_X1 U14300 ( .B1(n11934), .B2(n11916), .A(n11999), .ZN(n11921) );
  AOI21_X1 U14301 ( .B1(n11918), .B2(n11917), .A(n11921), .ZN(n11919) );
  NAND2_X1 U14302 ( .A1(n11920), .A2(n11919), .ZN(n11923) );
  NAND2_X1 U14303 ( .A1(n11925), .A2(n11924), .ZN(n11926) );
  NAND2_X1 U14304 ( .A1(n11944), .A2(n13933), .ZN(n11927) );
  NAND2_X1 U14305 ( .A1(n13847), .A2(n11999), .ZN(n11929) );
  AOI21_X1 U14306 ( .B1(n11927), .B2(n11929), .A(n14246), .ZN(n11933) );
  NAND2_X1 U14307 ( .A1(n11944), .A2(n13681), .ZN(n11928) );
  OR2_X1 U14308 ( .A1(n13839), .A2(n11953), .ZN(n11940) );
  AOI21_X1 U14309 ( .B1(n11928), .B2(n11940), .A(n14340), .ZN(n11932) );
  NAND2_X1 U14310 ( .A1(n13933), .A2(n11998), .ZN(n11941) );
  OR2_X1 U14311 ( .A1(n13839), .A2(n11941), .ZN(n11931) );
  INV_X1 U14312 ( .A(n11929), .ZN(n11937) );
  NAND2_X1 U14313 ( .A1(n11937), .A2(n13681), .ZN(n11930) );
  NAND2_X1 U14314 ( .A1(n11931), .A2(n11930), .ZN(n11938) );
  AOI22_X1 U14315 ( .A1(n11939), .A2(n14340), .B1(n11944), .B2(n11938), .ZN(
        n11948) );
  INV_X1 U14316 ( .A(n11940), .ZN(n11943) );
  INV_X1 U14317 ( .A(n11941), .ZN(n11942) );
  AOI21_X1 U14318 ( .B1(n11944), .B2(n11943), .A(n11942), .ZN(n11945) );
  INV_X1 U14319 ( .A(n11945), .ZN(n11946) );
  MUX2_X1 U14320 ( .A(n11950), .B(n11949), .S(n11998), .Z(n11951) );
  NAND2_X1 U14321 ( .A1(n11952), .A2(n14216), .ZN(n11957) );
  NAND2_X1 U14322 ( .A1(n14327), .A2(n11999), .ZN(n11955) );
  OR2_X1 U14323 ( .A1(n14327), .A2(n11953), .ZN(n11954) );
  MUX2_X1 U14324 ( .A(n11955), .B(n11954), .S(n13932), .Z(n11956) );
  MUX2_X1 U14325 ( .A(n13931), .B(n14319), .S(n11999), .Z(n11959) );
  MUX2_X1 U14326 ( .A(n13931), .B(n14319), .S(n11998), .Z(n11958) );
  MUX2_X1 U14327 ( .A(n13930), .B(n14314), .S(n11998), .Z(n11963) );
  MUX2_X1 U14328 ( .A(n13930), .B(n14314), .S(n11999), .Z(n11961) );
  NAND2_X1 U14329 ( .A1(n11962), .A2(n11961), .ZN(n11971) );
  NAND2_X1 U14330 ( .A1(n11971), .A2(n11969), .ZN(n11964) );
  MUX2_X1 U14331 ( .A(n13929), .B(n14308), .S(n11999), .Z(n11967) );
  NAND2_X1 U14332 ( .A1(n11964), .A2(n11967), .ZN(n11966) );
  MUX2_X1 U14333 ( .A(n13929), .B(n14308), .S(n11998), .Z(n11965) );
  NAND2_X1 U14334 ( .A1(n11966), .A2(n11965), .ZN(n11973) );
  INV_X1 U14335 ( .A(n11967), .ZN(n11968) );
  AND2_X1 U14336 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U14337 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  MUX2_X1 U14338 ( .A(n13928), .B(n14156), .S(n11998), .Z(n11977) );
  NAND2_X1 U14339 ( .A1(n11976), .A2(n11977), .ZN(n11975) );
  MUX2_X1 U14340 ( .A(n13928), .B(n14156), .S(n11999), .Z(n11974) );
  MUX2_X1 U14341 ( .A(n13927), .B(n14295), .S(n11999), .Z(n11980) );
  MUX2_X1 U14342 ( .A(n13927), .B(n14295), .S(n11998), .Z(n11979) );
  MUX2_X1 U14343 ( .A(n13926), .B(n14290), .S(n11998), .Z(n11983) );
  MUX2_X1 U14344 ( .A(n13926), .B(n14290), .S(n11999), .Z(n11981) );
  INV_X1 U14345 ( .A(n11983), .ZN(n11984) );
  MUX2_X1 U14346 ( .A(n13925), .B(n14283), .S(n11999), .Z(n11988) );
  MUX2_X1 U14347 ( .A(n13925), .B(n14283), .S(n11998), .Z(n11985) );
  NAND2_X1 U14348 ( .A1(n11986), .A2(n11985), .ZN(n11992) );
  INV_X1 U14349 ( .A(n11987), .ZN(n11990) );
  INV_X1 U14350 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U14351 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  MUX2_X1 U14352 ( .A(n13924), .B(n14093), .S(n11998), .Z(n11995) );
  MUX2_X1 U14353 ( .A(n13924), .B(n14093), .S(n11999), .Z(n11993) );
  MUX2_X1 U14354 ( .A(n13923), .B(n14270), .S(n11999), .Z(n11997) );
  MUX2_X1 U14355 ( .A(n13923), .B(n14270), .S(n11998), .Z(n11996) );
  MUX2_X1 U14356 ( .A(n13804), .B(n14266), .S(n11998), .Z(n12001) );
  NAND2_X1 U14357 ( .A1(n12000), .A2(n12001), .ZN(n12005) );
  MUX2_X1 U14358 ( .A(n13804), .B(n14266), .S(n11999), .Z(n12004) );
  INV_X1 U14359 ( .A(n12000), .ZN(n12003) );
  INV_X1 U14360 ( .A(n12001), .ZN(n12002) );
  INV_X1 U14361 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U14362 ( .A1(n9188), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U14363 ( .A1(n12006), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12007) );
  OAI211_X1 U14364 ( .C1(n12009), .C2(n14053), .A(n12008), .B(n12007), .ZN(
        n14054) );
  OAI21_X1 U14365 ( .B1(n14054), .B2(n12010), .A(n13922), .ZN(n12016) );
  OR2_X1 U14366 ( .A1(n12012), .A2(n6686), .ZN(n12015) );
  OR2_X1 U14367 ( .A1(n12013), .A2(n12472), .ZN(n12014) );
  MUX2_X1 U14368 ( .A(n12016), .B(n14261), .S(n11999), .Z(n12039) );
  NAND2_X1 U14369 ( .A1(n14064), .A2(n11998), .ZN(n12022) );
  NAND2_X1 U14370 ( .A1(n14054), .A2(n11999), .ZN(n12017) );
  OAI21_X1 U14371 ( .B1(n12019), .B2(n12018), .A(n12017), .ZN(n12020) );
  NAND2_X1 U14372 ( .A1(n12020), .A2(n13922), .ZN(n12021) );
  NAND2_X1 U14373 ( .A1(n12022), .A2(n12021), .ZN(n12040) );
  AND2_X1 U14374 ( .A1(n12039), .A2(n12040), .ZN(n12046) );
  INV_X1 U14375 ( .A(n14054), .ZN(n12027) );
  INV_X1 U14376 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12473) );
  NOR2_X1 U14377 ( .A1(n12013), .A2(n12473), .ZN(n12024) );
  MUX2_X1 U14378 ( .A(n12027), .B(n14258), .S(n12026), .Z(n12029) );
  NAND2_X1 U14379 ( .A1(n14258), .A2(n12027), .ZN(n12028) );
  NAND2_X1 U14380 ( .A1(n12029), .A2(n12028), .ZN(n12053) );
  NAND2_X1 U14381 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  NAND2_X1 U14382 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  NAND2_X1 U14383 ( .A1(n12035), .A2(n12034), .ZN(n12038) );
  NAND2_X1 U14384 ( .A1(n12037), .A2(n12036), .ZN(n12094) );
  AND2_X1 U14385 ( .A1(n12038), .A2(n12094), .ZN(n12050) );
  NAND2_X1 U14386 ( .A1(n12053), .A2(n12050), .ZN(n12047) );
  NOR3_X1 U14387 ( .A1(n12045), .A2(n12046), .A3(n12047), .ZN(n12101) );
  INV_X1 U14388 ( .A(n14258), .ZN(n14057) );
  XNOR2_X1 U14389 ( .A(n14057), .B(n14054), .ZN(n12091) );
  INV_X1 U14390 ( .A(n12038), .ZN(n12054) );
  NAND2_X1 U14391 ( .A1(n12091), .A2(n12054), .ZN(n12057) );
  INV_X1 U14392 ( .A(n12057), .ZN(n12044) );
  INV_X1 U14393 ( .A(n12039), .ZN(n12042) );
  INV_X1 U14394 ( .A(n12040), .ZN(n12041) );
  INV_X1 U14395 ( .A(n12048), .ZN(n12043) );
  NAND3_X1 U14396 ( .A1(n12045), .A2(n12044), .A3(n12043), .ZN(n12099) );
  INV_X1 U14397 ( .A(n12046), .ZN(n12058) );
  INV_X1 U14398 ( .A(n12047), .ZN(n12049) );
  NAND2_X1 U14399 ( .A1(n12049), .A2(n12048), .ZN(n12056) );
  INV_X1 U14400 ( .A(n12050), .ZN(n12051) );
  OAI21_X1 U14401 ( .B1(n12091), .B2(n12051), .A(n12053), .ZN(n12052) );
  OAI21_X1 U14402 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n12055) );
  OAI211_X1 U14403 ( .C1(n12058), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12059) );
  XNOR2_X1 U14404 ( .A(n14064), .B(n13922), .ZN(n12092) );
  NAND2_X1 U14405 ( .A1(n12061), .A2(n12060), .ZN(n14666) );
  INV_X1 U14406 ( .A(n14666), .ZN(n14675) );
  NAND4_X1 U14407 ( .A1(n14675), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n12067) );
  NOR3_X1 U14408 ( .A1(n12067), .A2(n12066), .A3(n12065), .ZN(n12069) );
  NAND4_X1 U14409 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n14638), .ZN(
        n12071) );
  OR4_X1 U14410 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12075) );
  NOR2_X1 U14411 ( .A1(n12076), .A2(n12075), .ZN(n12078) );
  NAND4_X1 U14412 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12081) );
  OR4_X1 U14413 ( .A1(n6837), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12084) );
  NOR2_X1 U14414 ( .A1(n14204), .A2(n12084), .ZN(n12085) );
  NAND4_X1 U14415 ( .A1(n14162), .A2(n12085), .A3(n14216), .A4(n14181), .ZN(
        n12086) );
  OR4_X1 U14416 ( .A1(n14113), .A2(n14127), .A3(n14145), .A4(n12086), .ZN(
        n12087) );
  NOR2_X1 U14417 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  NAND4_X1 U14418 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n14070), .ZN(
        n12093) );
  XNOR2_X1 U14419 ( .A(n12093), .B(n11835), .ZN(n12096) );
  INV_X1 U14420 ( .A(n12094), .ZN(n12095) );
  NAND3_X1 U14421 ( .A1(n12099), .A2(n12098), .A3(n12097), .ZN(n12100) );
  NOR2_X1 U14422 ( .A1(n12101), .A2(n12100), .ZN(n12106) );
  NOR3_X1 U14423 ( .A1(n12102), .A2(n14378), .A3(n13846), .ZN(n12104) );
  OAI21_X1 U14424 ( .B1(n14385), .B2(n12105), .A(P1_B_REG_SCAN_IN), .ZN(n12103) );
  OAI22_X1 U14425 ( .A1(n12106), .A2(n12105), .B1(n12104), .B2(n12103), .ZN(
        P1_U3242) );
  INV_X1 U14426 ( .A(n12107), .ZN(n12109) );
  OAI222_X1 U14427 ( .A1(n13054), .A2(n12110), .B1(n13057), .B2(n12109), .C1(
        P3_U3151), .C2(n12108), .ZN(P3_U3266) );
  AOI22_X1 U14428 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n7022), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n12472), .ZN(n12470) );
  XNOR2_X1 U14429 ( .A(n12471), .B(n12470), .ZN(n12466) );
  INV_X1 U14430 ( .A(n12466), .ZN(n12113) );
  XNOR2_X1 U14431 ( .A(n12739), .B(n12194), .ZN(n12191) );
  XNOR2_X1 U14432 ( .A(n12191), .B(n12746), .ZN(n12192) );
  NAND2_X1 U14433 ( .A1(n12117), .A2(n12264), .ZN(n12115) );
  NAND2_X1 U14434 ( .A1(n12116), .A2(n12115), .ZN(n12120) );
  INV_X1 U14435 ( .A(n12117), .ZN(n12118) );
  NAND2_X1 U14436 ( .A1(n12553), .A2(n12118), .ZN(n12119) );
  NAND2_X1 U14437 ( .A1(n12120), .A2(n12119), .ZN(n12263) );
  XNOR2_X1 U14438 ( .A(n14440), .B(n12194), .ZN(n12121) );
  XNOR2_X1 U14439 ( .A(n12121), .B(n12171), .ZN(n12262) );
  NAND2_X1 U14440 ( .A1(n12263), .A2(n12262), .ZN(n12123) );
  NAND2_X1 U14441 ( .A1(n12121), .A2(n12899), .ZN(n12122) );
  XNOR2_X1 U14442 ( .A(n13038), .B(n12194), .ZN(n12125) );
  XNOR2_X1 U14443 ( .A(n12125), .B(n12124), .ZN(n12167) );
  NAND2_X1 U14444 ( .A1(n12168), .A2(n12167), .ZN(n12127) );
  NAND2_X1 U14445 ( .A1(n12125), .A2(n12885), .ZN(n12126) );
  XNOR2_X1 U14446 ( .A(n13027), .B(n12153), .ZN(n12300) );
  AND2_X1 U14447 ( .A1(n12300), .A2(n12897), .ZN(n12128) );
  INV_X1 U14448 ( .A(n12300), .ZN(n12129) );
  NAND2_X1 U14449 ( .A1(n12129), .A2(n12299), .ZN(n12130) );
  XNOR2_X1 U14450 ( .A(n13021), .B(n12194), .ZN(n12131) );
  XNOR2_X1 U14451 ( .A(n12131), .B(n12884), .ZN(n12223) );
  INV_X1 U14452 ( .A(n12131), .ZN(n12132) );
  NAND2_X1 U14453 ( .A1(n12132), .A2(n12884), .ZN(n12133) );
  XNOR2_X1 U14454 ( .A(n13015), .B(n12194), .ZN(n12134) );
  XNOR2_X1 U14455 ( .A(n12134), .B(n12873), .ZN(n12232) );
  NAND2_X1 U14456 ( .A1(n12233), .A2(n12232), .ZN(n12231) );
  INV_X1 U14457 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U14458 ( .A1(n12135), .A2(n12873), .ZN(n12136) );
  XNOR2_X1 U14459 ( .A(n12944), .B(n12194), .ZN(n12137) );
  XNOR2_X1 U14460 ( .A(n12137), .B(n12834), .ZN(n12282) );
  INV_X1 U14461 ( .A(n12137), .ZN(n12138) );
  NAND2_X1 U14462 ( .A1(n12138), .A2(n12834), .ZN(n12139) );
  XNOR2_X1 U14463 ( .A(n12522), .B(n12194), .ZN(n12140) );
  XNOR2_X1 U14464 ( .A(n12140), .B(n12552), .ZN(n12185) );
  INV_X1 U14465 ( .A(n12140), .ZN(n12141) );
  NAND2_X1 U14466 ( .A1(n12141), .A2(n12851), .ZN(n12142) );
  XNOR2_X1 U14467 ( .A(n12937), .B(n12194), .ZN(n12143) );
  XNOR2_X1 U14468 ( .A(n12143), .B(n12811), .ZN(n12251) );
  INV_X1 U14469 ( .A(n12143), .ZN(n12144) );
  NAND2_X1 U14470 ( .A1(n12144), .A2(n12835), .ZN(n12145) );
  XNOR2_X1 U14471 ( .A(n12933), .B(n12194), .ZN(n12146) );
  XNOR2_X1 U14472 ( .A(n12146), .B(n12800), .ZN(n12205) );
  NAND2_X1 U14473 ( .A1(n12146), .A2(n12824), .ZN(n12147) );
  XNOR2_X1 U14474 ( .A(n12991), .B(n12153), .ZN(n12148) );
  INV_X1 U14475 ( .A(n12148), .ZN(n12149) );
  AND2_X1 U14476 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  XNOR2_X1 U14477 ( .A(n12152), .B(n12153), .ZN(n12243) );
  XNOR2_X1 U14478 ( .A(n12154), .B(n12153), .ZN(n12155) );
  OAI22_X1 U14479 ( .A1(n12243), .A2(n12791), .B1(n12447), .B2(n12155), .ZN(
        n12159) );
  OAI21_X1 U14480 ( .B1(n12240), .B2(n12801), .A(n12764), .ZN(n12157) );
  NOR3_X1 U14481 ( .A1(n12240), .A2(n12801), .A3(n12764), .ZN(n12156) );
  AOI21_X1 U14482 ( .B1(n12243), .B2(n12157), .A(n12156), .ZN(n12158) );
  XNOR2_X1 U14483 ( .A(n12975), .B(n12194), .ZN(n12160) );
  XNOR2_X1 U14484 ( .A(n12160), .B(n12778), .ZN(n12215) );
  XNOR2_X1 U14485 ( .A(n12753), .B(n12194), .ZN(n12161) );
  XNOR2_X1 U14486 ( .A(n12161), .B(n12218), .ZN(n12290) );
  XOR2_X1 U14487 ( .A(n12192), .B(n12193), .Z(n12166) );
  OAI22_X1 U14488 ( .A1(n12218), .A2(n12291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15182), .ZN(n12162) );
  AOI21_X1 U14489 ( .B1(n12294), .B2(n12732), .A(n12162), .ZN(n12163) );
  OAI21_X1 U14490 ( .B1(n12736), .B2(n12307), .A(n12163), .ZN(n12164) );
  AOI21_X1 U14491 ( .B1(n12739), .B2(n9993), .A(n12164), .ZN(n12165) );
  OAI21_X1 U14492 ( .B1(n12166), .B2(n12311), .A(n12165), .ZN(P3_U3154) );
  XNOR2_X1 U14493 ( .A(n12168), .B(n12167), .ZN(n12176) );
  NOR2_X1 U14494 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12169), .ZN(n12578) );
  AOI21_X1 U14495 ( .B1(n12897), .B2(n12294), .A(n12578), .ZN(n12170) );
  OAI21_X1 U14496 ( .B1(n12171), .B2(n12291), .A(n12170), .ZN(n12173) );
  NOR2_X1 U14497 ( .A1(n13038), .A2(n12288), .ZN(n12172) );
  AOI211_X1 U14498 ( .C1(n12174), .C2(n12257), .A(n12173), .B(n12172), .ZN(
        n12175) );
  OAI21_X1 U14499 ( .B1(n12176), .B2(n12311), .A(n12175), .ZN(P3_U3155) );
  XNOR2_X1 U14500 ( .A(n12241), .B(n12240), .ZN(n12242) );
  XNOR2_X1 U14501 ( .A(n12242), .B(n12447), .ZN(n12181) );
  NOR2_X1 U14502 ( .A1(n12307), .A2(n12792), .ZN(n12179) );
  AOI22_X1 U14503 ( .A1(n12294), .A2(n12764), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12177) );
  OAI21_X1 U14504 ( .B1(n12812), .B2(n12291), .A(n12177), .ZN(n12178) );
  AOI211_X1 U14505 ( .C1(n12926), .C2(n9993), .A(n12179), .B(n12178), .ZN(
        n12180) );
  OAI21_X1 U14506 ( .B1(n12181), .B2(n12311), .A(n12180), .ZN(P3_U3156) );
  INV_X1 U14507 ( .A(n12182), .ZN(n12183) );
  AOI21_X1 U14508 ( .B1(n12185), .B2(n12184), .A(n12183), .ZN(n12190) );
  NAND2_X1 U14509 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12701)
         );
  OAI21_X1 U14510 ( .B1(n12811), .B2(n12303), .A(n12701), .ZN(n12186) );
  AOI21_X1 U14511 ( .B1(n12305), .B2(n12834), .A(n12186), .ZN(n12187) );
  OAI21_X1 U14512 ( .B1(n12838), .B2(n12307), .A(n12187), .ZN(n12188) );
  AOI21_X1 U14513 ( .B1(n13005), .B2(n9993), .A(n12188), .ZN(n12189) );
  OAI21_X1 U14514 ( .B1(n12190), .B2(n12311), .A(n12189), .ZN(P3_U3159) );
  XNOR2_X1 U14515 ( .A(n12530), .B(n12194), .ZN(n12195) );
  NOR2_X1 U14516 ( .A1(n12720), .A2(n12303), .ZN(n12199) );
  OAI22_X1 U14517 ( .A1(n12197), .A2(n12291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12196), .ZN(n12198) );
  AOI211_X1 U14518 ( .C1(n12724), .C2(n12257), .A(n12199), .B(n12198), .ZN(
        n12202) );
  NAND2_X1 U14519 ( .A1(n12200), .A2(n9993), .ZN(n12201) );
  OAI211_X1 U14520 ( .C1(n12203), .C2(n12311), .A(n12202), .B(n12201), .ZN(
        P3_U3160) );
  OAI21_X1 U14521 ( .B1(n12206), .B2(n12205), .A(n12204), .ZN(n12207) );
  NAND2_X1 U14522 ( .A1(n12207), .A2(n12280), .ZN(n12212) );
  INV_X1 U14523 ( .A(n12813), .ZN(n12210) );
  AOI22_X1 U14524 ( .A1(n12294), .A2(n12551), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12208) );
  OAI21_X1 U14525 ( .B1(n12811), .B2(n12291), .A(n12208), .ZN(n12209) );
  AOI21_X1 U14526 ( .B1(n12210), .B2(n12257), .A(n12209), .ZN(n12211) );
  OAI211_X1 U14527 ( .C1(n12213), .C2(n12288), .A(n12212), .B(n12211), .ZN(
        P3_U3163) );
  XOR2_X1 U14528 ( .A(n12215), .B(n12214), .Z(n12221) );
  AOI22_X1 U14529 ( .A1(n12305), .A2(n12764), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12217) );
  NAND2_X1 U14530 ( .A1(n12257), .A2(n12768), .ZN(n12216) );
  OAI211_X1 U14531 ( .C1(n12218), .C2(n12303), .A(n12217), .B(n12216), .ZN(
        n12219) );
  AOI21_X1 U14532 ( .B1(n12975), .B2(n9993), .A(n12219), .ZN(n12220) );
  OAI21_X1 U14533 ( .B1(n12221), .B2(n12311), .A(n12220), .ZN(P3_U3165) );
  OAI211_X1 U14534 ( .C1(n12224), .C2(n12223), .A(n12222), .B(n12280), .ZN(
        n12229) );
  INV_X1 U14535 ( .A(n12225), .ZN(n12876) );
  NAND2_X1 U14536 ( .A1(n12897), .A2(n12305), .ZN(n12226) );
  NAND2_X1 U14537 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12635)
         );
  OAI211_X1 U14538 ( .C1(n12850), .C2(n12303), .A(n12226), .B(n12635), .ZN(
        n12227) );
  AOI21_X1 U14539 ( .B1(n12876), .B2(n12257), .A(n12227), .ZN(n12228) );
  OAI211_X1 U14540 ( .C1(n12230), .C2(n12288), .A(n12229), .B(n12228), .ZN(
        P3_U3166) );
  INV_X1 U14541 ( .A(n13015), .ZN(n12239) );
  OAI211_X1 U14542 ( .C1(n12233), .C2(n12232), .A(n12231), .B(n12280), .ZN(
        n12238) );
  INV_X1 U14543 ( .A(n12234), .ZN(n12867) );
  NAND2_X1 U14544 ( .A1(n12305), .A2(n12884), .ZN(n12235) );
  NAND2_X1 U14545 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12648)
         );
  OAI211_X1 U14546 ( .C1(n12858), .C2(n12303), .A(n12235), .B(n12648), .ZN(
        n12236) );
  AOI21_X1 U14547 ( .B1(n12867), .B2(n12257), .A(n12236), .ZN(n12237) );
  OAI211_X1 U14548 ( .C1(n12239), .C2(n12288), .A(n12238), .B(n12237), .ZN(
        P3_U3168) );
  OAI22_X1 U14549 ( .A1(n12242), .A2(n12801), .B1(n12241), .B2(n12240), .ZN(
        n12245) );
  XNOR2_X1 U14550 ( .A(n12243), .B(n12791), .ZN(n12244) );
  XNOR2_X1 U14551 ( .A(n12245), .B(n12244), .ZN(n12250) );
  NOR2_X1 U14552 ( .A1(n12307), .A2(n12780), .ZN(n12248) );
  AOI22_X1 U14553 ( .A1(n12778), .A2(n12294), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12246) );
  OAI21_X1 U14554 ( .B1(n12447), .B2(n12291), .A(n12246), .ZN(n12247) );
  AOI211_X1 U14555 ( .C1(n12981), .C2(n9993), .A(n12248), .B(n12247), .ZN(
        n12249) );
  OAI21_X1 U14556 ( .B1(n12250), .B2(n12311), .A(n12249), .ZN(P3_U3169) );
  AOI21_X1 U14557 ( .B1(n12252), .B2(n12251), .A(n12311), .ZN(n12254) );
  NAND2_X1 U14558 ( .A1(n12254), .A2(n12253), .ZN(n12260) );
  INV_X1 U14559 ( .A(n12826), .ZN(n12258) );
  AOI22_X1 U14560 ( .A1(n12294), .A2(n12800), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12255) );
  OAI21_X1 U14561 ( .B1(n12851), .B2(n12291), .A(n12255), .ZN(n12256) );
  AOI21_X1 U14562 ( .B1(n12258), .B2(n12257), .A(n12256), .ZN(n12259) );
  OAI211_X1 U14563 ( .C1(n12261), .C2(n12288), .A(n12260), .B(n12259), .ZN(
        P3_U3173) );
  XNOR2_X1 U14564 ( .A(n12263), .B(n12262), .ZN(n12271) );
  AND2_X1 U14565 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14932) );
  NOR2_X1 U14566 ( .A1(n12264), .A2(n12291), .ZN(n12265) );
  AOI211_X1 U14567 ( .C1(n12294), .C2(n12885), .A(n14932), .B(n12265), .ZN(
        n12266) );
  OAI21_X1 U14568 ( .B1(n12267), .B2(n12307), .A(n12266), .ZN(n12268) );
  AOI21_X1 U14569 ( .B1(n12269), .B2(n9993), .A(n12268), .ZN(n12270) );
  OAI21_X1 U14570 ( .B1(n12271), .B2(n12311), .A(n12270), .ZN(P3_U3174) );
  XNOR2_X1 U14571 ( .A(n12272), .B(n12551), .ZN(n12279) );
  OAI22_X1 U14572 ( .A1(n12447), .A2(n12303), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12273), .ZN(n12274) );
  AOI21_X1 U14573 ( .B1(n12305), .B2(n12800), .A(n12274), .ZN(n12275) );
  OAI21_X1 U14574 ( .B1(n12276), .B2(n12307), .A(n12275), .ZN(n12277) );
  AOI21_X1 U14575 ( .B1(n12991), .B2(n9993), .A(n12277), .ZN(n12278) );
  OAI21_X1 U14576 ( .B1(n12279), .B2(n12311), .A(n12278), .ZN(P3_U3175) );
  INV_X1 U14577 ( .A(n12944), .ZN(n12289) );
  OAI211_X1 U14578 ( .C1(n12283), .C2(n12282), .A(n12281), .B(n12280), .ZN(
        n12287) );
  NAND2_X1 U14579 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12668)
         );
  OAI21_X1 U14580 ( .B1(n12851), .B2(n12303), .A(n12668), .ZN(n12285) );
  NOR2_X1 U14581 ( .A1(n12307), .A2(n12853), .ZN(n12284) );
  AOI211_X1 U14582 ( .C1(n12305), .C2(n12873), .A(n12285), .B(n12284), .ZN(
        n12286) );
  OAI211_X1 U14583 ( .C1(n12289), .C2(n12288), .A(n12287), .B(n12286), .ZN(
        P3_U3178) );
  OAI22_X1 U14584 ( .A1(n12292), .A2(n12291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15029), .ZN(n12293) );
  AOI21_X1 U14585 ( .B1(n12294), .B2(n12746), .A(n12293), .ZN(n12295) );
  OAI21_X1 U14586 ( .B1(n12307), .B2(n12750), .A(n12295), .ZN(n12296) );
  AOI21_X1 U14587 ( .B1(n12753), .B2(n9993), .A(n12296), .ZN(n12297) );
  OAI21_X1 U14588 ( .B1(n12298), .B2(n12311), .A(n12297), .ZN(P3_U3180) );
  XNOR2_X1 U14589 ( .A(n12300), .B(n12299), .ZN(n12301) );
  XNOR2_X1 U14590 ( .A(n12302), .B(n12301), .ZN(n12312) );
  NAND2_X1 U14591 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12598)
         );
  OAI21_X1 U14592 ( .B1(n12406), .B2(n12303), .A(n12598), .ZN(n12304) );
  AOI21_X1 U14593 ( .B1(n12305), .B2(n12885), .A(n12304), .ZN(n12306) );
  OAI21_X1 U14594 ( .B1(n12308), .B2(n12307), .A(n12306), .ZN(n12309) );
  AOI21_X1 U14595 ( .B1(n13027), .B2(n9993), .A(n12309), .ZN(n12310) );
  OAI21_X1 U14596 ( .B1(n12312), .B2(n12311), .A(n12310), .ZN(P3_U3181) );
  NAND2_X1 U14597 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  NAND2_X1 U14598 ( .A1(n12317), .A2(n12315), .ZN(n12316) );
  INV_X1 U14599 ( .A(n12533), .ZN(n12458) );
  INV_X1 U14600 ( .A(n12317), .ZN(n12456) );
  NAND2_X1 U14601 ( .A1(n6509), .A2(n12453), .ZN(n12528) );
  INV_X1 U14602 ( .A(n12772), .ZN(n12318) );
  NAND2_X1 U14603 ( .A1(n12321), .A2(n12318), .ZN(n12320) );
  NAND2_X1 U14604 ( .A1(n12320), .A2(n12319), .ZN(n12323) );
  INV_X1 U14605 ( .A(n12321), .ZN(n12322) );
  MUX2_X1 U14606 ( .A(n12323), .B(n12322), .S(n12446), .Z(n12328) );
  MUX2_X1 U14607 ( .A(n12325), .B(n12324), .S(n12463), .Z(n12326) );
  OAI21_X1 U14608 ( .B1(n12328), .B2(n12327), .A(n12326), .ZN(n12452) );
  MUX2_X1 U14609 ( .A(n12439), .B(n12438), .S(n12463), .Z(n12445) );
  NAND3_X1 U14610 ( .A1(n12338), .A2(n12330), .A3(n12544), .ZN(n12335) );
  NAND2_X1 U14611 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND2_X1 U14612 ( .A1(n12331), .A2(n12463), .ZN(n12334) );
  AOI22_X1 U14613 ( .A1(n12335), .A2(n12334), .B1(n12333), .B2(n12332), .ZN(
        n12336) );
  MUX2_X1 U14614 ( .A(n12446), .B(n12336), .S(n8979), .Z(n12342) );
  OAI21_X1 U14615 ( .B1(n12446), .B2(n12338), .A(n12337), .ZN(n12341) );
  NAND2_X1 U14616 ( .A1(n6655), .A2(n14937), .ZN(n12339) );
  AND2_X1 U14617 ( .A1(n12347), .A2(n12339), .ZN(n12340) );
  OAI22_X1 U14618 ( .A1(n12342), .A2(n12341), .B1(n12340), .B2(n12463), .ZN(
        n12346) );
  AOI21_X1 U14619 ( .B1(n12345), .B2(n12343), .A(n12446), .ZN(n12344) );
  AOI21_X1 U14620 ( .B1(n12346), .B2(n12345), .A(n12344), .ZN(n12349) );
  NOR2_X1 U14621 ( .A1(n12347), .A2(n12446), .ZN(n12348) );
  OAI21_X1 U14622 ( .B1(n12349), .B2(n12348), .A(n12514), .ZN(n12354) );
  NAND2_X1 U14623 ( .A1(n12560), .A2(n12463), .ZN(n12352) );
  NAND2_X1 U14624 ( .A1(n12350), .A2(n12446), .ZN(n12351) );
  MUX2_X1 U14625 ( .A(n12352), .B(n12351), .S(n6914), .Z(n12353) );
  AOI21_X1 U14626 ( .B1(n12354), .B2(n12353), .A(n8620), .ZN(n12363) );
  NAND2_X1 U14627 ( .A1(n12359), .A2(n12355), .ZN(n12358) );
  NAND2_X1 U14628 ( .A1(n12360), .A2(n12356), .ZN(n12357) );
  MUX2_X1 U14629 ( .A(n12358), .B(n12357), .S(n12446), .Z(n12362) );
  MUX2_X1 U14630 ( .A(n12360), .B(n12359), .S(n12446), .Z(n12361) );
  OAI211_X1 U14631 ( .C1(n12363), .C2(n12362), .A(n12507), .B(n12361), .ZN(
        n12367) );
  MUX2_X1 U14632 ( .A(n12365), .B(n12364), .S(n12446), .Z(n12366) );
  NAND3_X1 U14633 ( .A1(n12367), .A2(n12505), .A3(n12366), .ZN(n12372) );
  INV_X1 U14634 ( .A(n12368), .ZN(n12508) );
  MUX2_X1 U14635 ( .A(n12370), .B(n12369), .S(n12463), .Z(n12371) );
  NAND3_X1 U14636 ( .A1(n12372), .A2(n12508), .A3(n12371), .ZN(n12374) );
  NOR2_X1 U14637 ( .A1(n12516), .A2(n12511), .ZN(n12373) );
  NAND2_X1 U14638 ( .A1(n12374), .A2(n12373), .ZN(n12389) );
  NAND2_X1 U14639 ( .A1(n12390), .A2(n12376), .ZN(n12377) );
  AOI21_X1 U14640 ( .B1(n7073), .B2(n12382), .A(n12377), .ZN(n12378) );
  OAI21_X1 U14641 ( .B1(n12389), .B2(n12556), .A(n12378), .ZN(n12387) );
  OAI21_X1 U14642 ( .B1(n12380), .B2(n12379), .A(n12391), .ZN(n12381) );
  AOI21_X1 U14643 ( .B1(n12383), .B2(n12382), .A(n12381), .ZN(n12384) );
  OAI21_X1 U14644 ( .B1(n12389), .B2(n12385), .A(n12384), .ZN(n12386) );
  MUX2_X1 U14645 ( .A(n12387), .B(n12386), .S(n12446), .Z(n12394) );
  NOR2_X1 U14646 ( .A1(n12389), .A2(n12388), .ZN(n12393) );
  MUX2_X1 U14647 ( .A(n12391), .B(n12390), .S(n12446), .Z(n12392) );
  OAI21_X1 U14648 ( .B1(n12394), .B2(n12393), .A(n12392), .ZN(n12396) );
  INV_X1 U14649 ( .A(n12395), .ZN(n12519) );
  NAND2_X1 U14650 ( .A1(n12396), .A2(n12519), .ZN(n12400) );
  INV_X1 U14651 ( .A(n12900), .ZN(n12894) );
  MUX2_X1 U14652 ( .A(n12398), .B(n12397), .S(n12463), .Z(n12399) );
  NAND3_X1 U14653 ( .A1(n12400), .A2(n12894), .A3(n12399), .ZN(n12404) );
  MUX2_X1 U14654 ( .A(n12402), .B(n12401), .S(n12446), .Z(n12403) );
  NAND3_X1 U14655 ( .A1(n12404), .A2(n7327), .A3(n12403), .ZN(n12410) );
  OAI21_X1 U14656 ( .B1(n13021), .B2(n12406), .A(n12405), .ZN(n12407) );
  NAND2_X1 U14657 ( .A1(n12407), .A2(n12463), .ZN(n12409) );
  INV_X1 U14658 ( .A(n12412), .ZN(n12408) );
  AOI21_X1 U14659 ( .B1(n12410), .B2(n12409), .A(n12408), .ZN(n12415) );
  AOI21_X1 U14660 ( .B1(n12412), .B2(n12411), .A(n12463), .ZN(n12414) );
  NAND2_X1 U14661 ( .A1(n12884), .A2(n12446), .ZN(n12413) );
  OAI22_X1 U14662 ( .A1(n12415), .A2(n12414), .B1(n13021), .B2(n12413), .ZN(
        n12422) );
  INV_X1 U14663 ( .A(n12416), .ZN(n12421) );
  INV_X1 U14664 ( .A(n12417), .ZN(n12418) );
  AOI21_X1 U14665 ( .B1(n12423), .B2(n12418), .A(n12463), .ZN(n12419) );
  NAND2_X1 U14666 ( .A1(n12420), .A2(n12419), .ZN(n12425) );
  AOI22_X1 U14667 ( .A1(n12422), .A2(n12863), .B1(n12421), .B2(n12425), .ZN(
        n12427) );
  NAND3_X1 U14668 ( .A1(n12429), .A2(n12463), .A3(n12423), .ZN(n12424) );
  NAND2_X1 U14669 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  OAI21_X1 U14670 ( .B1(n12427), .B2(n12842), .A(n12426), .ZN(n12431) );
  MUX2_X1 U14671 ( .A(n12429), .B(n12428), .S(n12463), .Z(n12430) );
  NAND3_X1 U14672 ( .A1(n12431), .A2(n7318), .A3(n12430), .ZN(n12437) );
  NAND2_X1 U14673 ( .A1(n12937), .A2(n12811), .ZN(n12432) );
  MUX2_X1 U14674 ( .A(n12433), .B(n12432), .S(n12463), .Z(n12436) );
  AND2_X1 U14675 ( .A1(n12435), .A2(n12434), .ZN(n12525) );
  NAND3_X1 U14676 ( .A1(n12437), .A2(n12436), .A3(n12808), .ZN(n12443) );
  NAND2_X1 U14677 ( .A1(n12800), .A2(n12463), .ZN(n12440) );
  OR2_X1 U14678 ( .A1(n12933), .A2(n12440), .ZN(n12442) );
  NAND3_X1 U14679 ( .A1(n12933), .A2(n12824), .A3(n12446), .ZN(n12441) );
  NAND4_X1 U14680 ( .A1(n12443), .A2(n12799), .A3(n12442), .A4(n12441), .ZN(
        n12444) );
  NAND3_X1 U14681 ( .A1(n12445), .A2(n12784), .A3(n12444), .ZN(n12449) );
  NAND3_X1 U14682 ( .A1(n12926), .A2(n12447), .A3(n12446), .ZN(n12448) );
  NAND2_X1 U14683 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  NAND3_X1 U14684 ( .A1(n12758), .A2(n12775), .A3(n12450), .ZN(n12451) );
  NAND3_X1 U14685 ( .A1(n12744), .A2(n12452), .A3(n12451), .ZN(n12455) );
  MUX2_X1 U14686 ( .A(n12453), .B(n6509), .S(n12463), .Z(n12454) );
  NAND3_X1 U14687 ( .A1(n12456), .A2(n12455), .A3(n12454), .ZN(n12457) );
  NAND2_X1 U14688 ( .A1(n12458), .A2(n12457), .ZN(n12459) );
  NOR2_X2 U14689 ( .A1(n6521), .A2(n12459), .ZN(n12462) );
  INV_X1 U14690 ( .A(n12462), .ZN(n12460) );
  NAND2_X1 U14691 ( .A1(n12460), .A2(n12491), .ZN(n12465) );
  INV_X1 U14692 ( .A(n12461), .ZN(n12492) );
  NOR2_X1 U14693 ( .A1(n12462), .A2(n12492), .ZN(n12464) );
  NAND2_X1 U14694 ( .A1(n12466), .A2(n12477), .ZN(n12468) );
  NAND2_X1 U14695 ( .A1(n6483), .A2(SI_30_), .ZN(n12467) );
  INV_X1 U14696 ( .A(n12550), .ZN(n12469) );
  NAND2_X1 U14697 ( .A1(n14438), .A2(n12469), .ZN(n12531) );
  AOI22_X1 U14698 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n12474), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n12473), .ZN(n12475) );
  XNOR2_X1 U14699 ( .A(n12476), .B(n12475), .ZN(n13043) );
  NAND2_X1 U14700 ( .A1(n6483), .A2(SI_31_), .ZN(n12479) );
  NAND2_X1 U14701 ( .A1(n6497), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12485) );
  INV_X1 U14702 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12480) );
  OR2_X1 U14703 ( .A1(n6694), .A2(n12480), .ZN(n12484) );
  INV_X1 U14704 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12482) );
  OR2_X1 U14705 ( .A1(n6484), .A2(n12482), .ZN(n12483) );
  NAND2_X1 U14706 ( .A1(n12488), .A2(n12709), .ZN(n12497) );
  INV_X1 U14707 ( .A(n14438), .ZN(n12715) );
  NAND2_X1 U14708 ( .A1(n12715), .A2(n12550), .ZN(n12499) );
  NAND2_X1 U14709 ( .A1(n12497), .A2(n12499), .ZN(n12534) );
  INV_X1 U14710 ( .A(n12488), .ZN(n12712) );
  INV_X1 U14711 ( .A(n12491), .ZN(n12496) );
  INV_X1 U14712 ( .A(n12709), .ZN(n12549) );
  NAND2_X1 U14713 ( .A1(n12549), .A2(n12550), .ZN(n12493) );
  OAI211_X1 U14714 ( .C1(n12712), .C2(n12499), .A(n12498), .B(n12497), .ZN(
        n12500) );
  INV_X1 U14715 ( .A(n12871), .ZN(n12521) );
  NAND4_X1 U14716 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12510) );
  NAND4_X1 U14717 ( .A1(n12508), .A2(n12507), .A3(n12506), .A4(n12505), .ZN(
        n12509) );
  NOR2_X1 U14718 ( .A1(n12510), .A2(n12509), .ZN(n12515) );
  NOR2_X1 U14719 ( .A1(n12511), .A2(n14942), .ZN(n12512) );
  NAND4_X1 U14720 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12517) );
  NOR2_X1 U14721 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  NAND3_X1 U14722 ( .A1(n12894), .A2(n12519), .A3(n12518), .ZN(n12520) );
  NOR3_X1 U14723 ( .A1(n12521), .A2(n12879), .A3(n12520), .ZN(n12523) );
  XNOR2_X1 U14724 ( .A(n12522), .B(n12851), .ZN(n12833) );
  NAND4_X1 U14725 ( .A1(n12863), .A2(n7070), .A3(n12523), .A4(n12833), .ZN(
        n12524) );
  NOR4_X1 U14726 ( .A1(n12525), .A2(n12788), .A3(n12821), .A4(n12524), .ZN(
        n12526) );
  NAND4_X1 U14727 ( .A1(n12799), .A2(n12758), .A3(n12775), .A4(n12526), .ZN(
        n12527) );
  NOR2_X1 U14728 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  NAND4_X1 U14729 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n6924), .ZN(
        n12532) );
  NOR4_X1 U14730 ( .A1(n12535), .A2(n12534), .A3(n12533), .A4(n12532), .ZN(
        n12536) );
  XNOR2_X1 U14731 ( .A(n12536), .B(n12690), .ZN(n12537) );
  NOR2_X1 U14732 ( .A1(n12543), .A2(n12542), .ZN(n12546) );
  OAI21_X1 U14733 ( .B1(n12547), .B2(n12544), .A(P3_B_REG_SCAN_IN), .ZN(n12545) );
  OAI22_X1 U14734 ( .A1(n12548), .A2(n12547), .B1(n12546), .B2(n12545), .ZN(
        P3_U3296) );
  MUX2_X1 U14735 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12549), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14736 ( .A(n12550), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12562), .Z(
        P3_U3521) );
  MUX2_X1 U14737 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12732), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14738 ( .A(n12763), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12562), .Z(
        P3_U3517) );
  MUX2_X1 U14739 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12778), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14740 ( .A(n12764), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12562), .Z(
        P3_U3515) );
  MUX2_X1 U14741 ( .A(n12801), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12562), .Z(
        P3_U3514) );
  MUX2_X1 U14742 ( .A(n12551), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12562), .Z(
        P3_U3513) );
  MUX2_X1 U14743 ( .A(n12800), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12562), .Z(
        P3_U3512) );
  MUX2_X1 U14744 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12835), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14745 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12552), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14746 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12834), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14747 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12873), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14748 ( .A(n12884), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12562), .Z(
        P3_U3507) );
  MUX2_X1 U14749 ( .A(n12885), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12562), .Z(
        P3_U3505) );
  MUX2_X1 U14750 ( .A(n12899), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12562), .Z(
        P3_U3504) );
  MUX2_X1 U14751 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12553), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14752 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12554), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14753 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12555), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14754 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14755 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14756 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12558), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14757 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12559), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14758 ( .A(n12560), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12562), .Z(
        P3_U3495) );
  MUX2_X1 U14759 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12561), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14760 ( .A(n6655), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12562), .Z(
        P3_U3493) );
  MUX2_X1 U14761 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12564), .S(P3_U3897), .Z(
        P3_U3492) );
  INV_X1 U14762 ( .A(n14917), .ZN(n12575) );
  NAND2_X1 U14763 ( .A1(n12582), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12565) );
  AND2_X2 U14764 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  NOR2_X1 U14765 ( .A1(n12575), .A2(n12567), .ZN(n12568) );
  AND2_X1 U14766 ( .A1(n12580), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12600) );
  NOR2_X1 U14767 ( .A1(n12580), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12569) );
  OR2_X1 U14768 ( .A1(n12600), .A2(n12569), .ZN(n12586) );
  AOI21_X1 U14769 ( .B1(n6615), .B2(n12586), .A(n12596), .ZN(n12595) );
  NAND2_X1 U14770 ( .A1(n12582), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12572) );
  NOR2_X1 U14771 ( .A1(n12575), .A2(n12574), .ZN(n12576) );
  NAND2_X1 U14772 ( .A1(n12580), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12611) );
  OR2_X1 U14773 ( .A1(n12580), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12577) );
  NAND2_X1 U14774 ( .A1(n12611), .A2(n12577), .ZN(n12609) );
  XNOR2_X1 U14775 ( .A(n12610), .B(n12609), .ZN(n12593) );
  AOI21_X1 U14776 ( .B1(n14896), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12578), 
        .ZN(n12579) );
  OAI21_X1 U14777 ( .B1(n14918), .B2(n12580), .A(n12579), .ZN(n12591) );
  INV_X1 U14778 ( .A(n12581), .ZN(n12584) );
  INV_X1 U14779 ( .A(n12582), .ZN(n12583) );
  NOR2_X1 U14780 ( .A1(n12584), .A2(n12583), .ZN(n14919) );
  MUX2_X1 U14781 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12623), .Z(n12585) );
  XNOR2_X1 U14782 ( .A(n12585), .B(n14917), .ZN(n14923) );
  NOR2_X1 U14783 ( .A1(n12585), .A2(n14917), .ZN(n12587) );
  OR2_X1 U14784 ( .A1(n14921), .A2(n12587), .ZN(n12589) );
  MUX2_X1 U14785 ( .A(n12609), .B(n12586), .S(n12623), .Z(n12588) );
  NOR3_X1 U14786 ( .A1(n14921), .A2(n12587), .A3(n12588), .ZN(n12603) );
  AOI211_X1 U14787 ( .C1(n12589), .C2(n12588), .A(n14928), .B(n12603), .ZN(
        n12590) );
  AOI211_X1 U14788 ( .C1(n12593), .C2(n12592), .A(n12591), .B(n12590), .ZN(
        n12594) );
  OAI21_X1 U14789 ( .B1(n12595), .B2(n14926), .A(n12594), .ZN(P3_U3196) );
  INV_X1 U14790 ( .A(n12628), .ZN(n14411) );
  AOI21_X1 U14791 ( .B1(n12952), .B2(n12597), .A(n12629), .ZN(n12616) );
  OAI21_X1 U14792 ( .B1(n14916), .B2(n12599), .A(n12598), .ZN(n12608) );
  INV_X1 U14793 ( .A(n12611), .ZN(n12601) );
  MUX2_X1 U14794 ( .A(n12601), .B(n12600), .S(n12623), .Z(n12602) );
  NOR2_X1 U14795 ( .A1(n12603), .A2(n12602), .ZN(n12622) );
  XNOR2_X1 U14796 ( .A(n12622), .B(n12628), .ZN(n12605) );
  MUX2_X1 U14797 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12623), .Z(n12604) );
  NOR2_X1 U14798 ( .A1(n12605), .A2(n12604), .ZN(n12621) );
  AOI21_X1 U14799 ( .B1(n12605), .B2(n12604), .A(n12621), .ZN(n12606) );
  NOR2_X1 U14800 ( .A1(n12606), .A2(n14928), .ZN(n12607) );
  AOI211_X1 U14801 ( .C1(n12669), .C2(n12628), .A(n12608), .B(n12607), .ZN(
        n12615) );
  AOI21_X1 U14802 ( .B1(n12886), .B2(n12612), .A(n12618), .ZN(n12613) );
  OR2_X1 U14803 ( .A1(n12613), .A2(n14934), .ZN(n12614) );
  OAI211_X1 U14804 ( .C1(n12616), .C2(n14926), .A(n12615), .B(n12614), .ZN(
        P3_U3197) );
  AND2_X1 U14805 ( .A1(n14411), .A2(n12617), .ZN(n12619) );
  INV_X1 U14806 ( .A(n12634), .ZN(n14416) );
  AOI22_X1 U14807 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12634), .B1(n14416), 
        .B2(n12875), .ZN(n12620) );
  AOI21_X1 U14808 ( .B1(n6551), .B2(n12620), .A(n12645), .ZN(n12642) );
  MUX2_X1 U14809 ( .A(n12875), .B(n12949), .S(n12623), .Z(n12624) );
  NOR2_X1 U14810 ( .A1(n12624), .A2(n12634), .ZN(n12651) );
  INV_X1 U14811 ( .A(n12651), .ZN(n12625) );
  NAND2_X1 U14812 ( .A1(n12624), .A2(n12634), .ZN(n12650) );
  NAND2_X1 U14813 ( .A1(n12625), .A2(n12650), .ZN(n12626) );
  XNOR2_X1 U14814 ( .A(n12652), .B(n12626), .ZN(n12640) );
  NOR2_X1 U14815 ( .A1(n12628), .A2(n12627), .ZN(n12630) );
  AOI22_X1 U14816 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12634), .B1(n14416), 
        .B2(n12949), .ZN(n12631) );
  AOI21_X1 U14817 ( .B1(n12632), .B2(n12631), .A(n12643), .ZN(n12633) );
  NOR2_X1 U14818 ( .A1(n12633), .A2(n14926), .ZN(n12639) );
  NAND2_X1 U14819 ( .A1(n12669), .A2(n12634), .ZN(n12636) );
  OAI211_X1 U14820 ( .C1(n12637), .C2(n14916), .A(n12636), .B(n12635), .ZN(
        n12638) );
  AOI211_X1 U14821 ( .C1(n12640), .C2(n12703), .A(n12639), .B(n12638), .ZN(
        n12641) );
  OAI21_X1 U14822 ( .B1(n12642), .B2(n14934), .A(n12641), .ZN(P3_U3198) );
  AOI21_X1 U14823 ( .B1(n15058), .B2(n12644), .A(n12670), .ZN(n12658) );
  AOI21_X1 U14824 ( .B1(n12866), .B2(n12646), .A(n12663), .ZN(n12649) );
  NAND2_X1 U14825 ( .A1(n14896), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12647) );
  OAI211_X1 U14826 ( .C1(n14934), .C2(n12649), .A(n12648), .B(n12647), .ZN(
        n12656) );
  MUX2_X1 U14827 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12623), .Z(n12660) );
  XNOR2_X1 U14828 ( .A(n12660), .B(n12664), .ZN(n12654) );
  NOR2_X1 U14829 ( .A1(n12653), .A2(n12654), .ZN(n12659) );
  AOI211_X1 U14830 ( .C1(n12654), .C2(n12653), .A(n14928), .B(n12659), .ZN(
        n12655) );
  AOI211_X1 U14831 ( .C1(n12669), .C2(n12671), .A(n12656), .B(n12655), .ZN(
        n12657) );
  OAI21_X1 U14832 ( .B1(n12658), .B2(n14926), .A(n12657), .ZN(P3_U3199) );
  MUX2_X1 U14833 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12623), .Z(n12662) );
  AOI21_X1 U14834 ( .B1(n12660), .B2(n12664), .A(n12659), .ZN(n12689) );
  XNOR2_X1 U14835 ( .A(n12689), .B(n12688), .ZN(n12661) );
  NOR2_X1 U14836 ( .A1(n12661), .A2(n12662), .ZN(n12687) );
  AOI21_X1 U14837 ( .B1(n12662), .B2(n12661), .A(n12687), .ZN(n12681) );
  NAND2_X1 U14838 ( .A1(n12673), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12695) );
  OAI21_X1 U14839 ( .B1(n12673), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12695), 
        .ZN(n12665) );
  NAND2_X1 U14840 ( .A1(n14896), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12667) );
  OR2_X1 U14841 ( .A1(n12672), .A2(n12671), .ZN(n12676) );
  NAND2_X1 U14842 ( .A1(n12673), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U14843 ( .A1(n12688), .A2(n12945), .ZN(n12674) );
  NAND2_X1 U14844 ( .A1(n12682), .A2(n12674), .ZN(n12675) );
  AND3_X1 U14845 ( .A1(n12677), .A2(n12676), .A3(n12675), .ZN(n12679) );
  OAI21_X1 U14846 ( .B1(n12684), .B2(n12679), .A(n12678), .ZN(n12680) );
  INV_X1 U14847 ( .A(n12682), .ZN(n12683) );
  NOR2_X1 U14848 ( .A1(n12684), .A2(n12683), .ZN(n12686) );
  XNOR2_X1 U14849 ( .A(n12690), .B(n12940), .ZN(n12691) );
  INV_X1 U14850 ( .A(n12691), .ZN(n12685) );
  XNOR2_X1 U14851 ( .A(n12686), .B(n12685), .ZN(n12705) );
  AOI21_X1 U14852 ( .B1(n12689), .B2(n12688), .A(n12687), .ZN(n12693) );
  XNOR2_X1 U14853 ( .A(n12690), .B(n12837), .ZN(n12698) );
  MUX2_X1 U14854 ( .A(n12698), .B(n12691), .S(n12623), .Z(n12692) );
  XNOR2_X1 U14855 ( .A(n12693), .B(n12692), .ZN(n12704) );
  NOR2_X1 U14856 ( .A1(n14918), .A2(n12694), .ZN(n12702) );
  INV_X1 U14857 ( .A(n12695), .ZN(n12696) );
  INV_X1 U14858 ( .A(n12698), .ZN(n12699) );
  NAND2_X1 U14859 ( .A1(n14896), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U14860 ( .A1(n12706), .A2(n12888), .ZN(n12710) );
  INV_X1 U14861 ( .A(n12707), .ZN(n12708) );
  OR2_X1 U14862 ( .A1(n12709), .A2(n12708), .ZN(n14436) );
  AOI21_X1 U14863 ( .B1(n12710), .B2(n14436), .A(n14955), .ZN(n12713) );
  AOI21_X1 U14864 ( .B1(n14955), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12713), 
        .ZN(n12711) );
  OAI21_X1 U14865 ( .B1(n12712), .B2(n12903), .A(n12711), .ZN(P3_U3202) );
  AOI21_X1 U14866 ( .B1(n14955), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12713), 
        .ZN(n12714) );
  OAI21_X1 U14867 ( .B1(n12715), .B2(n12903), .A(n12714), .ZN(P3_U3203) );
  OAI211_X1 U14868 ( .C1(n12717), .C2(n12723), .A(n12716), .B(n14947), .ZN(
        n12719) );
  NAND2_X1 U14869 ( .A1(n12746), .A2(n12898), .ZN(n12718) );
  OAI211_X1 U14870 ( .C1(n12720), .C2(n14944), .A(n12719), .B(n12718), .ZN(
        n12908) );
  INV_X1 U14871 ( .A(n12908), .ZN(n12728) );
  NAND2_X1 U14872 ( .A1(n12729), .A2(n12721), .ZN(n12722) );
  XOR2_X1 U14873 ( .A(n12723), .B(n12722), .Z(n12909) );
  AOI22_X1 U14874 ( .A1(n14955), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n12888), 
        .B2(n12724), .ZN(n12725) );
  OAI21_X1 U14875 ( .B1(n12965), .B2(n12903), .A(n12725), .ZN(n12726) );
  AOI21_X1 U14876 ( .B1(n12909), .B2(n12905), .A(n12726), .ZN(n12727) );
  OAI21_X1 U14877 ( .B1(n12728), .B2(n14955), .A(n12727), .ZN(P3_U3205) );
  INV_X1 U14878 ( .A(n12913), .ZN(n12742) );
  AOI22_X1 U14879 ( .A1(n12732), .A2(n12896), .B1(n12898), .B2(n12763), .ZN(
        n12734) );
  OAI211_X1 U14880 ( .C1(n12735), .C2(n12861), .A(n12734), .B(n12733), .ZN(
        n12912) );
  NAND2_X1 U14881 ( .A1(n12912), .A2(n14953), .ZN(n12741) );
  INV_X1 U14882 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12737) );
  OAI22_X1 U14883 ( .A1(n14953), .A2(n12737), .B1(n12736), .B2(n14940), .ZN(
        n12738) );
  AOI21_X1 U14884 ( .B1(n12739), .B2(n12889), .A(n12738), .ZN(n12740) );
  OAI211_X1 U14885 ( .C1(n12742), .C2(n12757), .A(n12741), .B(n12740), .ZN(
        P3_U3206) );
  XNOR2_X1 U14886 ( .A(n12743), .B(n12744), .ZN(n12916) );
  INV_X1 U14887 ( .A(n12916), .ZN(n12756) );
  XNOR2_X1 U14888 ( .A(n12745), .B(n12744), .ZN(n12749) );
  AOI22_X1 U14889 ( .A1(n12778), .A2(n12898), .B1(n12896), .B2(n12746), .ZN(
        n12748) );
  NAND2_X1 U14890 ( .A1(n12916), .A2(n14993), .ZN(n12747) );
  OAI211_X1 U14891 ( .C1(n12749), .C2(n12861), .A(n12748), .B(n12747), .ZN(
        n12915) );
  NAND2_X1 U14892 ( .A1(n12915), .A2(n14953), .ZN(n12755) );
  OAI22_X1 U14893 ( .A1(n14953), .A2(n12751), .B1(n12750), .B2(n14940), .ZN(
        n12752) );
  AOI21_X1 U14894 ( .B1(n12753), .B2(n12889), .A(n12752), .ZN(n12754) );
  OAI211_X1 U14895 ( .C1(n12757), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        P3_U3207) );
  XNOR2_X1 U14896 ( .A(n6584), .B(n12758), .ZN(n12978) );
  NAND2_X1 U14897 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  NAND2_X1 U14898 ( .A1(n12760), .A2(n14947), .ZN(n12762) );
  OR2_X1 U14899 ( .A1(n12762), .A2(n12761), .ZN(n12766) );
  AOI22_X1 U14900 ( .A1(n12898), .A2(n12764), .B1(n12763), .B2(n12896), .ZN(
        n12765) );
  MUX2_X1 U14901 ( .A(n12974), .B(n12767), .S(n14955), .Z(n12770) );
  AOI22_X1 U14902 ( .A1(n12975), .A2(n12889), .B1(n12888), .B2(n12768), .ZN(
        n12769) );
  OAI211_X1 U14903 ( .C1(n12978), .C2(n12892), .A(n12770), .B(n12769), .ZN(
        P3_U3208) );
  INV_X1 U14904 ( .A(n12771), .ZN(n12774) );
  AOI21_X1 U14905 ( .B1(n12787), .B2(n12772), .A(n12775), .ZN(n12773) );
  NOR2_X1 U14906 ( .A1(n12774), .A2(n12773), .ZN(n12984) );
  XNOR2_X1 U14907 ( .A(n12776), .B(n12775), .ZN(n12777) );
  AOI222_X1 U14908 ( .A1(n12801), .A2(n12898), .B1(n12778), .B2(n12896), .C1(
        n14947), .C2(n12777), .ZN(n12979) );
  MUX2_X1 U14909 ( .A(n12779), .B(n12979), .S(n14953), .Z(n12783) );
  INV_X1 U14910 ( .A(n12780), .ZN(n12781) );
  AOI22_X1 U14911 ( .A1(n12981), .A2(n12889), .B1(n12888), .B2(n12781), .ZN(
        n12782) );
  OAI211_X1 U14912 ( .C1(n12984), .C2(n12892), .A(n12783), .B(n12782), .ZN(
        P3_U3209) );
  OR2_X1 U14913 ( .A1(n12785), .A2(n12784), .ZN(n12786) );
  NAND2_X1 U14914 ( .A1(n12787), .A2(n12786), .ZN(n12988) );
  XNOR2_X1 U14915 ( .A(n12789), .B(n12788), .ZN(n12790) );
  OAI222_X1 U14916 ( .A1(n14944), .A2(n12791), .B1(n12790), .B2(n12861), .C1(
        n14943), .C2(n12812), .ZN(n12925) );
  NAND2_X1 U14917 ( .A1(n12925), .A2(n14953), .ZN(n12796) );
  OAI22_X1 U14918 ( .A1(n14953), .A2(n12793), .B1(n12792), .B2(n14940), .ZN(
        n12794) );
  AOI21_X1 U14919 ( .B1(n12926), .B2(n12889), .A(n12794), .ZN(n12795) );
  OAI211_X1 U14920 ( .C1(n12988), .C2(n12892), .A(n12796), .B(n12795), .ZN(
        P3_U3210) );
  XNOR2_X1 U14921 ( .A(n12797), .B(n12799), .ZN(n12994) );
  XOR2_X1 U14922 ( .A(n12798), .B(n12799), .Z(n12802) );
  AOI222_X1 U14923 ( .A1(n14947), .A2(n12802), .B1(n12801), .B2(n12896), .C1(
        n12800), .C2(n12898), .ZN(n12989) );
  MUX2_X1 U14924 ( .A(n12803), .B(n12989), .S(n14953), .Z(n12806) );
  AOI22_X1 U14925 ( .A1(n12991), .A2(n12889), .B1(n12888), .B2(n12804), .ZN(
        n12805) );
  OAI211_X1 U14926 ( .C1(n12994), .C2(n12892), .A(n12806), .B(n12805), .ZN(
        P3_U3211) );
  XNOR2_X1 U14927 ( .A(n12807), .B(n12808), .ZN(n12998) );
  XNOR2_X1 U14928 ( .A(n12809), .B(n12808), .ZN(n12810) );
  OAI222_X1 U14929 ( .A1(n14944), .A2(n12812), .B1(n14943), .B2(n12811), .C1(
        n12861), .C2(n12810), .ZN(n12932) );
  NAND2_X1 U14930 ( .A1(n12932), .A2(n14953), .ZN(n12817) );
  OAI22_X1 U14931 ( .A1(n14953), .A2(n12814), .B1(n12813), .B2(n14940), .ZN(
        n12815) );
  AOI21_X1 U14932 ( .B1(n12933), .B2(n12889), .A(n12815), .ZN(n12816) );
  OAI211_X1 U14933 ( .C1(n12998), .C2(n12892), .A(n12817), .B(n12816), .ZN(
        P3_U3212) );
  NAND2_X1 U14934 ( .A1(n12818), .A2(n12821), .ZN(n12819) );
  NAND2_X1 U14935 ( .A1(n12820), .A2(n12819), .ZN(n13002) );
  XNOR2_X1 U14936 ( .A(n12822), .B(n12821), .ZN(n12823) );
  OAI222_X1 U14937 ( .A1(n14944), .A2(n12824), .B1(n14943), .B2(n12851), .C1(
        n12861), .C2(n12823), .ZN(n12936) );
  NAND2_X1 U14938 ( .A1(n12936), .A2(n14953), .ZN(n12829) );
  NAND2_X1 U14939 ( .A1(n14955), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n12825) );
  OAI21_X1 U14940 ( .B1(n12826), .B2(n14940), .A(n12825), .ZN(n12827) );
  AOI21_X1 U14941 ( .B1(n12937), .B2(n12889), .A(n12827), .ZN(n12828) );
  OAI211_X1 U14942 ( .C1(n13002), .C2(n12892), .A(n12829), .B(n12828), .ZN(
        P3_U3213) );
  NAND2_X1 U14943 ( .A1(n12845), .A2(n12830), .ZN(n12831) );
  XNOR2_X1 U14944 ( .A(n12831), .B(n12833), .ZN(n13008) );
  XOR2_X1 U14945 ( .A(n12833), .B(n12832), .Z(n12836) );
  AOI222_X1 U14946 ( .A1(n14947), .A2(n12836), .B1(n12835), .B2(n12896), .C1(
        n12834), .C2(n12898), .ZN(n13003) );
  MUX2_X1 U14947 ( .A(n12837), .B(n13003), .S(n14953), .Z(n12841) );
  INV_X1 U14948 ( .A(n12838), .ZN(n12839) );
  AOI22_X1 U14949 ( .A1(n13005), .A2(n12889), .B1(n12888), .B2(n12839), .ZN(
        n12840) );
  OAI211_X1 U14950 ( .C1(n13008), .C2(n12892), .A(n12841), .B(n12840), .ZN(
        P3_U3214) );
  NAND2_X1 U14951 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  NAND2_X1 U14952 ( .A1(n12845), .A2(n12844), .ZN(n13012) );
  INV_X1 U14953 ( .A(n12846), .ZN(n12847) );
  AOI21_X1 U14954 ( .B1(n7070), .B2(n12848), .A(n12847), .ZN(n12849) );
  OAI222_X1 U14955 ( .A1(n14944), .A2(n12851), .B1(n14943), .B2(n12850), .C1(
        n12861), .C2(n12849), .ZN(n12943) );
  NAND2_X1 U14956 ( .A1(n12943), .A2(n14953), .ZN(n12856) );
  NAND2_X1 U14957 ( .A1(n14955), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U14958 ( .B1(n12853), .B2(n14940), .A(n12852), .ZN(n12854) );
  AOI21_X1 U14959 ( .B1(n12944), .B2(n12889), .A(n12854), .ZN(n12855) );
  OAI211_X1 U14960 ( .C1(n13012), .C2(n12892), .A(n12856), .B(n12855), .ZN(
        P3_U3215) );
  XOR2_X1 U14961 ( .A(n12863), .B(n12857), .Z(n13018) );
  NOR2_X1 U14962 ( .A1(n12858), .A2(n14944), .ZN(n12865) );
  INV_X1 U14963 ( .A(n12859), .ZN(n12860) );
  AOI211_X1 U14964 ( .C1(n12863), .C2(n12862), .A(n12861), .B(n12860), .ZN(
        n12864) );
  AOI211_X1 U14965 ( .C1(n12898), .C2(n12884), .A(n12865), .B(n12864), .ZN(
        n13013) );
  MUX2_X1 U14966 ( .A(n12866), .B(n13013), .S(n14953), .Z(n12869) );
  AOI22_X1 U14967 ( .A1(n13015), .A2(n12889), .B1(n12888), .B2(n12867), .ZN(
        n12868) );
  OAI211_X1 U14968 ( .C1(n13018), .C2(n12892), .A(n12869), .B(n12868), .ZN(
        P3_U3216) );
  XOR2_X1 U14969 ( .A(n12870), .B(n12871), .Z(n13024) );
  XNOR2_X1 U14970 ( .A(n12872), .B(n12871), .ZN(n12874) );
  AOI222_X1 U14971 ( .A1(n14947), .A2(n12874), .B1(n12873), .B2(n12896), .C1(
        n12897), .C2(n12898), .ZN(n13019) );
  MUX2_X1 U14972 ( .A(n12875), .B(n13019), .S(n14953), .Z(n12878) );
  AOI22_X1 U14973 ( .A1(n13021), .A2(n12889), .B1(n12888), .B2(n12876), .ZN(
        n12877) );
  OAI211_X1 U14974 ( .C1(n13024), .C2(n12892), .A(n12878), .B(n12877), .ZN(
        P3_U3217) );
  XNOR2_X1 U14975 ( .A(n12880), .B(n12879), .ZN(n13030) );
  XNOR2_X1 U14976 ( .A(n12882), .B(n7327), .ZN(n12883) );
  AOI222_X1 U14977 ( .A1(n12885), .A2(n12898), .B1(n12884), .B2(n12896), .C1(
        n14947), .C2(n12883), .ZN(n13025) );
  MUX2_X1 U14978 ( .A(n12886), .B(n13025), .S(n14953), .Z(n12891) );
  AOI22_X1 U14979 ( .A1(n13027), .A2(n12889), .B1(n12888), .B2(n12887), .ZN(
        n12890) );
  OAI211_X1 U14980 ( .C1(n13030), .C2(n12892), .A(n12891), .B(n12890), .ZN(
        P3_U3218) );
  XNOR2_X1 U14981 ( .A(n12893), .B(n12894), .ZN(n12895) );
  AOI222_X1 U14982 ( .A1(n12899), .A2(n12898), .B1(n12897), .B2(n12896), .C1(
        n14947), .C2(n12895), .ZN(n13031) );
  MUX2_X1 U14983 ( .A(n8745), .B(n13031), .S(n14953), .Z(n12907) );
  XNOR2_X1 U14984 ( .A(n12901), .B(n12900), .ZN(n13035) );
  OAI22_X1 U14985 ( .A1(n13038), .A2(n12903), .B1(n12902), .B2(n14940), .ZN(
        n12904) );
  AOI21_X1 U14986 ( .B1(n13035), .B2(n12905), .A(n12904), .ZN(n12906) );
  NAND2_X1 U14987 ( .A1(n12907), .A2(n12906), .ZN(P3_U3219) );
  AOI21_X1 U14988 ( .B1(n12909), .B2(n14959), .A(n12908), .ZN(n12962) );
  MUX2_X1 U14989 ( .A(n12910), .B(n12962), .S(n15025), .Z(n12911) );
  INV_X1 U14990 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12914) );
  AOI21_X1 U14991 ( .B1(n15009), .B2(n12916), .A(n12915), .ZN(n12969) );
  MUX2_X1 U14992 ( .A(n12917), .B(n12969), .S(n15025), .Z(n12918) );
  OAI21_X1 U14993 ( .B1(n12972), .B2(n12961), .A(n12918), .ZN(P3_U3485) );
  MUX2_X1 U14994 ( .A(n12919), .B(n12974), .S(n15025), .Z(n12921) );
  INV_X1 U14995 ( .A(n12961), .ZN(n12953) );
  NAND2_X1 U14996 ( .A1(n12975), .A2(n12953), .ZN(n12920) );
  OAI211_X1 U14997 ( .C1(n12957), .C2(n12978), .A(n12921), .B(n12920), .ZN(
        P3_U3484) );
  MUX2_X1 U14998 ( .A(n12922), .B(n12979), .S(n15025), .Z(n12924) );
  NAND2_X1 U14999 ( .A1(n12981), .A2(n12953), .ZN(n12923) );
  OAI211_X1 U15000 ( .C1(n12984), .C2(n12957), .A(n12924), .B(n12923), .ZN(
        P3_U3483) );
  AOI21_X1 U15001 ( .B1(n15001), .B2(n12926), .A(n12925), .ZN(n12985) );
  MUX2_X1 U15002 ( .A(n12927), .B(n12985), .S(n15025), .Z(n12928) );
  OAI21_X1 U15003 ( .B1(n12957), .B2(n12988), .A(n12928), .ZN(P3_U3482) );
  MUX2_X1 U15004 ( .A(n12929), .B(n12989), .S(n15025), .Z(n12931) );
  NAND2_X1 U15005 ( .A1(n12991), .A2(n12953), .ZN(n12930) );
  OAI211_X1 U15006 ( .C1(n12994), .C2(n12957), .A(n12931), .B(n12930), .ZN(
        P3_U3481) );
  AOI21_X1 U15007 ( .B1(n15001), .B2(n12933), .A(n12932), .ZN(n12995) );
  MUX2_X1 U15008 ( .A(n12934), .B(n12995), .S(n15025), .Z(n12935) );
  OAI21_X1 U15009 ( .B1(n12957), .B2(n12998), .A(n12935), .ZN(P3_U3480) );
  AOI21_X1 U15010 ( .B1(n15001), .B2(n12937), .A(n12936), .ZN(n12999) );
  MUX2_X1 U15011 ( .A(n12938), .B(n12999), .S(n15025), .Z(n12939) );
  OAI21_X1 U15012 ( .B1(n12957), .B2(n13002), .A(n12939), .ZN(P3_U3479) );
  MUX2_X1 U15013 ( .A(n12940), .B(n13003), .S(n15025), .Z(n12942) );
  NAND2_X1 U15014 ( .A1(n13005), .A2(n12953), .ZN(n12941) );
  OAI211_X1 U15015 ( .C1(n13008), .C2(n12957), .A(n12942), .B(n12941), .ZN(
        P3_U3478) );
  AOI21_X1 U15016 ( .B1(n15001), .B2(n12944), .A(n12943), .ZN(n13009) );
  MUX2_X1 U15017 ( .A(n12945), .B(n13009), .S(n15025), .Z(n12946) );
  OAI21_X1 U15018 ( .B1(n12957), .B2(n13012), .A(n12946), .ZN(P3_U3477) );
  MUX2_X1 U15019 ( .A(n15058), .B(n13013), .S(n15025), .Z(n12948) );
  NAND2_X1 U15020 ( .A1(n13015), .A2(n12953), .ZN(n12947) );
  OAI211_X1 U15021 ( .C1(n12957), .C2(n13018), .A(n12948), .B(n12947), .ZN(
        P3_U3476) );
  MUX2_X1 U15022 ( .A(n12949), .B(n13019), .S(n15025), .Z(n12951) );
  NAND2_X1 U15023 ( .A1(n13021), .A2(n12953), .ZN(n12950) );
  OAI211_X1 U15024 ( .C1(n13024), .C2(n12957), .A(n12951), .B(n12950), .ZN(
        P3_U3475) );
  MUX2_X1 U15025 ( .A(n12952), .B(n13025), .S(n15025), .Z(n12955) );
  NAND2_X1 U15026 ( .A1(n13027), .A2(n12953), .ZN(n12954) );
  OAI211_X1 U15027 ( .C1(n12957), .C2(n13030), .A(n12955), .B(n12954), .ZN(
        P3_U3474) );
  MUX2_X1 U15028 ( .A(n12956), .B(n13031), .S(n15025), .Z(n12960) );
  INV_X1 U15029 ( .A(n12957), .ZN(n12958) );
  NAND2_X1 U15030 ( .A1(n13035), .A2(n12958), .ZN(n12959) );
  OAI211_X1 U15031 ( .C1(n12961), .C2(n13038), .A(n12960), .B(n12959), .ZN(
        P3_U3473) );
  MUX2_X1 U15032 ( .A(n12963), .B(n12962), .S(n15010), .Z(n12964) );
  OAI21_X1 U15033 ( .B1(n12965), .B2(n13039), .A(n12964), .ZN(P3_U3455) );
  INV_X1 U15034 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12967) );
  INV_X1 U15035 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12970) );
  MUX2_X1 U15036 ( .A(n12970), .B(n12969), .S(n15010), .Z(n12971) );
  OAI21_X1 U15037 ( .B1(n12972), .B2(n13039), .A(n12971), .ZN(P3_U3453) );
  INV_X1 U15038 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12973) );
  MUX2_X1 U15039 ( .A(n12974), .B(n12973), .S(n15012), .Z(n12977) );
  INV_X1 U15040 ( .A(n13039), .ZN(n13026) );
  NAND2_X1 U15041 ( .A1(n12975), .A2(n13026), .ZN(n12976) );
  OAI211_X1 U15042 ( .C1(n12978), .C2(n13033), .A(n12977), .B(n12976), .ZN(
        P3_U3452) );
  INV_X1 U15043 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12980) );
  MUX2_X1 U15044 ( .A(n12980), .B(n12979), .S(n15010), .Z(n12983) );
  NAND2_X1 U15045 ( .A1(n12981), .A2(n13026), .ZN(n12982) );
  OAI211_X1 U15046 ( .C1(n12984), .C2(n13033), .A(n12983), .B(n12982), .ZN(
        P3_U3451) );
  INV_X1 U15047 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12986) );
  MUX2_X1 U15048 ( .A(n12986), .B(n12985), .S(n15010), .Z(n12987) );
  OAI21_X1 U15049 ( .B1(n12988), .B2(n13033), .A(n12987), .ZN(P3_U3450) );
  INV_X1 U15050 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12990) );
  MUX2_X1 U15051 ( .A(n12990), .B(n12989), .S(n15010), .Z(n12993) );
  NAND2_X1 U15052 ( .A1(n12991), .A2(n13026), .ZN(n12992) );
  OAI211_X1 U15053 ( .C1(n12994), .C2(n13033), .A(n12993), .B(n12992), .ZN(
        P3_U3449) );
  INV_X1 U15054 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12996) );
  MUX2_X1 U15055 ( .A(n12996), .B(n12995), .S(n15010), .Z(n12997) );
  OAI21_X1 U15056 ( .B1(n12998), .B2(n13033), .A(n12997), .ZN(P3_U3448) );
  INV_X1 U15057 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13000) );
  MUX2_X1 U15058 ( .A(n13000), .B(n12999), .S(n15010), .Z(n13001) );
  OAI21_X1 U15059 ( .B1(n13002), .B2(n13033), .A(n13001), .ZN(P3_U3447) );
  INV_X1 U15060 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13004) );
  MUX2_X1 U15061 ( .A(n13004), .B(n13003), .S(n15010), .Z(n13007) );
  NAND2_X1 U15062 ( .A1(n13005), .A2(n13026), .ZN(n13006) );
  OAI211_X1 U15063 ( .C1(n13008), .C2(n13033), .A(n13007), .B(n13006), .ZN(
        P3_U3446) );
  INV_X1 U15064 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13010) );
  MUX2_X1 U15065 ( .A(n13010), .B(n13009), .S(n15010), .Z(n13011) );
  OAI21_X1 U15066 ( .B1(n13012), .B2(n13033), .A(n13011), .ZN(P3_U3444) );
  INV_X1 U15067 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13014) );
  MUX2_X1 U15068 ( .A(n13014), .B(n13013), .S(n15010), .Z(n13017) );
  NAND2_X1 U15069 ( .A1(n13015), .A2(n13026), .ZN(n13016) );
  OAI211_X1 U15070 ( .C1(n13018), .C2(n13033), .A(n13017), .B(n13016), .ZN(
        P3_U3441) );
  INV_X1 U15071 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13020) );
  MUX2_X1 U15072 ( .A(n13020), .B(n13019), .S(n15010), .Z(n13023) );
  NAND2_X1 U15073 ( .A1(n13021), .A2(n13026), .ZN(n13022) );
  OAI211_X1 U15074 ( .C1(n13024), .C2(n13033), .A(n13023), .B(n13022), .ZN(
        P3_U3438) );
  INV_X1 U15075 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n15186) );
  MUX2_X1 U15076 ( .A(n15186), .B(n13025), .S(n15010), .Z(n13029) );
  NAND2_X1 U15077 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  OAI211_X1 U15078 ( .C1(n13030), .C2(n13033), .A(n13029), .B(n13028), .ZN(
        P3_U3435) );
  INV_X1 U15079 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13032) );
  MUX2_X1 U15080 ( .A(n13032), .B(n13031), .S(n15010), .Z(n13037) );
  INV_X1 U15081 ( .A(n13033), .ZN(n13034) );
  NAND2_X1 U15082 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  OAI211_X1 U15083 ( .C1(n13039), .C2(n13038), .A(n13037), .B(n13036), .ZN(
        P3_U3432) );
  MUX2_X1 U15084 ( .A(P3_D_REG_1__SCAN_IN), .B(n13040), .S(n13041), .Z(
        P3_U3377) );
  MUX2_X1 U15085 ( .A(P3_D_REG_0__SCAN_IN), .B(n13042), .S(n13041), .Z(
        P3_U3376) );
  INV_X1 U15086 ( .A(n13043), .ZN(n13048) );
  INV_X1 U15087 ( .A(n13054), .ZN(n14412) );
  NOR4_X1 U15088 ( .A1(n13045), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n13044), .ZN(n13046) );
  AOI21_X1 U15089 ( .B1(SI_31_), .B2(n14412), .A(n13046), .ZN(n13047) );
  OAI21_X1 U15090 ( .B1(n13048), .B2(n13057), .A(n13047), .ZN(P3_U3264) );
  INV_X1 U15091 ( .A(n13049), .ZN(n13051) );
  OAI222_X1 U15092 ( .A1(n13054), .A2(n15031), .B1(n13057), .B2(n13051), .C1(
        n12623), .C2(P3_U3151), .ZN(P3_U3268) );
  INV_X1 U15093 ( .A(n13052), .ZN(n13058) );
  INV_X1 U15094 ( .A(n13053), .ZN(n13056) );
  OAI222_X1 U15095 ( .A1(P3_U3151), .A2(n13058), .B1(n13057), .B2(n13056), 
        .C1(n13055), .C2(n13054), .ZN(P3_U3269) );
  MUX2_X1 U15096 ( .A(n13059), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15097 ( .A(n13060), .B(n13061), .ZN(n13065) );
  AOI22_X1 U15098 ( .A1(n13190), .A2(n13437), .B1(n13435), .B2(n13192), .ZN(
        n13317) );
  AOI22_X1 U15099 ( .A1(n13324), .A2(n13151), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13062) );
  OAI21_X1 U15100 ( .B1(n13317), .B2(n13149), .A(n13062), .ZN(n13063) );
  AOI21_X1 U15101 ( .B1(n13526), .B2(n13185), .A(n13063), .ZN(n13064) );
  OAI21_X1 U15102 ( .B1(n13065), .B2(n13187), .A(n13064), .ZN(P2_U3186) );
  OAI22_X1 U15103 ( .A1(n13183), .A2(n13378), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13067), .ZN(n13069) );
  OAI22_X1 U15104 ( .A1(n13091), .A2(n13139), .B1(n13138), .B2(n13099), .ZN(
        n13068) );
  AOI211_X1 U15105 ( .C1(n13388), .C2(n13173), .A(n13069), .B(n13068), .ZN(
        n13070) );
  OAI21_X1 U15106 ( .B1(n13071), .B2(n13187), .A(n13070), .ZN(P2_U3188) );
  INV_X1 U15107 ( .A(n13072), .ZN(n13074) );
  NAND2_X1 U15108 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  XNOR2_X1 U15109 ( .A(n13076), .B(n13075), .ZN(n13080) );
  NAND2_X1 U15110 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13290)
         );
  OAI21_X1 U15111 ( .B1(n13183), .B2(n13458), .A(n13290), .ZN(n13078) );
  OAI22_X1 U15112 ( .A1(n13448), .A2(n13138), .B1(n13139), .B2(n13446), .ZN(
        n13077) );
  AOI211_X1 U15113 ( .C1(n13571), .C2(n13173), .A(n13078), .B(n13077), .ZN(
        n13079) );
  OAI21_X1 U15114 ( .B1(n13080), .B2(n13187), .A(n13079), .ZN(P2_U3191) );
  INV_X1 U15115 ( .A(n13138), .ZN(n13155) );
  AOI22_X1 U15116 ( .A1(n13173), .A2(n13081), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13157), .ZN(n13087) );
  OAI21_X1 U15117 ( .B1(n13084), .B2(n13083), .A(n13082), .ZN(n13085) );
  NAND2_X1 U15118 ( .A1(n13162), .A2(n13085), .ZN(n13086) );
  NAND3_X1 U15119 ( .A1(n13088), .A2(n13087), .A3(n13086), .ZN(P2_U3194) );
  XNOR2_X1 U15120 ( .A(n13090), .B(n13089), .ZN(n13095) );
  OAI22_X1 U15121 ( .A1(n13091), .A2(n13447), .B1(n13448), .B2(n13445), .ZN(
        n13415) );
  AOI22_X1 U15122 ( .A1(n13181), .A2(n13415), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13092) );
  OAI21_X1 U15123 ( .B1(n13417), .B2(n13183), .A(n13092), .ZN(n13093) );
  AOI21_X1 U15124 ( .B1(n13561), .B2(n13185), .A(n13093), .ZN(n13094) );
  OAI21_X1 U15125 ( .B1(n13095), .B2(n13187), .A(n13094), .ZN(P2_U3195) );
  XNOR2_X1 U15126 ( .A(n13098), .B(n13097), .ZN(n13105) );
  INV_X1 U15127 ( .A(n13350), .ZN(n13102) );
  OAI22_X1 U15128 ( .A1(n13100), .A2(n13447), .B1(n13099), .B2(n13445), .ZN(
        n13346) );
  AOI22_X1 U15129 ( .A1(n13346), .A2(n13181), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13101) );
  OAI21_X1 U15130 ( .B1(n13102), .B2(n13183), .A(n13101), .ZN(n13103) );
  AOI21_X1 U15131 ( .B1(n13537), .B2(n13185), .A(n13103), .ZN(n13104) );
  OAI21_X1 U15132 ( .B1(n13105), .B2(n13187), .A(n13104), .ZN(P2_U3197) );
  AOI21_X1 U15133 ( .B1(n13108), .B2(n13107), .A(n13106), .ZN(n13113) );
  AOI22_X1 U15134 ( .A1(n13181), .A2(n13586), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13109) );
  OAI21_X1 U15135 ( .B1(n13110), .B2(n13183), .A(n13109), .ZN(n13111) );
  AOI21_X1 U15136 ( .B1(n13587), .B2(n13173), .A(n13111), .ZN(n13112) );
  OAI21_X1 U15137 ( .B1(n13113), .B2(n13187), .A(n13112), .ZN(P2_U3198) );
  AOI21_X1 U15138 ( .B1(n13116), .B2(n13115), .A(n13114), .ZN(n13122) );
  OAI22_X1 U15139 ( .A1(n13446), .A2(n13447), .B1(n13117), .B2(n13445), .ZN(
        n13487) );
  NOR2_X1 U15140 ( .A1(n13118), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14826) );
  AOI21_X1 U15141 ( .B1(n13181), .B2(n13487), .A(n14826), .ZN(n13119) );
  OAI21_X1 U15142 ( .B1(n13494), .B2(n13183), .A(n13119), .ZN(n13120) );
  AOI21_X1 U15143 ( .B1(n13581), .B2(n13185), .A(n13120), .ZN(n13121) );
  OAI21_X1 U15144 ( .B1(n13122), .B2(n13187), .A(n13121), .ZN(P2_U3200) );
  XNOR2_X1 U15145 ( .A(n13125), .B(n13124), .ZN(n13130) );
  OAI22_X1 U15146 ( .A1(n13180), .A2(n13447), .B1(n13126), .B2(n13445), .ZN(
        n13359) );
  AOI22_X1 U15147 ( .A1(n13359), .A2(n13181), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13127) );
  OAI21_X1 U15148 ( .B1(n13366), .B2(n13183), .A(n13127), .ZN(n13128) );
  AOI21_X1 U15149 ( .B1(n13369), .B2(n13185), .A(n13128), .ZN(n13129) );
  OAI21_X1 U15150 ( .B1(n13130), .B2(n13187), .A(n13129), .ZN(P2_U3201) );
  INV_X1 U15151 ( .A(n13131), .ZN(n13132) );
  NOR2_X1 U15152 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  XNOR2_X1 U15153 ( .A(n13135), .B(n13134), .ZN(n13143) );
  OAI22_X1 U15154 ( .A1(n13183), .A2(n13428), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13136), .ZN(n13141) );
  OAI22_X1 U15155 ( .A1(n13170), .A2(n13139), .B1(n13138), .B2(n13137), .ZN(
        n13140) );
  AOI211_X1 U15156 ( .C1(n13565), .C2(n13185), .A(n13141), .B(n13140), .ZN(
        n13142) );
  OAI21_X1 U15157 ( .B1(n13143), .B2(n13187), .A(n13142), .ZN(P2_U3205) );
  OAI21_X1 U15158 ( .B1(n13146), .B2(n13145), .A(n13144), .ZN(n13147) );
  NAND2_X1 U15159 ( .A1(n13147), .A2(n13162), .ZN(n13153) );
  AOI22_X1 U15160 ( .A1(n13194), .A2(n13437), .B1(n13435), .B2(n13438), .ZN(
        n13395) );
  OAI22_X1 U15161 ( .A1(n13395), .A2(n13149), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13148), .ZN(n13150) );
  AOI21_X1 U15162 ( .B1(n13400), .B2(n13151), .A(n13150), .ZN(n13152) );
  OAI211_X1 U15163 ( .C1(n13403), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        P2_U3207) );
  AOI22_X1 U15164 ( .A1(n13156), .A2(n6748), .B1(n13155), .B2(n13211), .ZN(
        n13166) );
  AOI22_X1 U15165 ( .A1(n13185), .A2(n13158), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13157), .ZN(n13165) );
  OAI21_X1 U15166 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13163) );
  NAND2_X1 U15167 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  NAND3_X1 U15168 ( .A1(n13166), .A2(n13165), .A3(n13164), .ZN(P2_U3209) );
  XNOR2_X1 U15169 ( .A(n13168), .B(n13167), .ZN(n13175) );
  OAI22_X1 U15170 ( .A1(n13170), .A2(n13447), .B1(n13169), .B2(n13445), .ZN(
        n13469) );
  AOI22_X1 U15171 ( .A1(n13181), .A2(n13469), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13171) );
  OAI21_X1 U15172 ( .B1(n13474), .B2(n13183), .A(n13171), .ZN(n13172) );
  AOI21_X1 U15173 ( .B1(n13576), .B2(n13173), .A(n13172), .ZN(n13174) );
  OAI21_X1 U15174 ( .B1(n13175), .B2(n13187), .A(n13174), .ZN(P2_U3210) );
  INV_X1 U15175 ( .A(n13176), .ZN(n13177) );
  AOI21_X1 U15176 ( .B1(n13179), .B2(n13178), .A(n13177), .ZN(n13188) );
  OAI22_X1 U15177 ( .A1(n13306), .A2(n13447), .B1(n13180), .B2(n13445), .ZN(
        n13331) );
  AOI22_X1 U15178 ( .A1(n13331), .A2(n13181), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13182) );
  OAI21_X1 U15179 ( .B1(n13336), .B2(n13183), .A(n13182), .ZN(n13184) );
  AOI21_X1 U15180 ( .B1(n13532), .B2(n13185), .A(n13184), .ZN(n13186) );
  OAI21_X1 U15181 ( .B1(n13188), .B2(n13187), .A(n13186), .ZN(P2_U3212) );
  INV_X2 U15182 ( .A(P2_U3947), .ZN(n13214) );
  MUX2_X1 U15183 ( .A(n13292), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13214), .Z(
        P2_U3562) );
  MUX2_X1 U15184 ( .A(n13189), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13214), .Z(
        P2_U3561) );
  MUX2_X1 U15185 ( .A(n13190), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13214), .Z(
        P2_U3559) );
  MUX2_X1 U15186 ( .A(n13191), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13214), .Z(
        P2_U3558) );
  MUX2_X1 U15187 ( .A(n13192), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13214), .Z(
        P2_U3557) );
  MUX2_X1 U15188 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13193), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15189 ( .A(n13377), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13214), .Z(
        P2_U3555) );
  MUX2_X1 U15190 ( .A(n13194), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13214), .Z(
        P2_U3554) );
  MUX2_X1 U15191 ( .A(n13375), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13214), .Z(
        P2_U3553) );
  MUX2_X1 U15192 ( .A(n13438), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13214), .Z(
        P2_U3552) );
  MUX2_X1 U15193 ( .A(n13195), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13214), .Z(
        P2_U3551) );
  MUX2_X1 U15194 ( .A(n13436), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13214), .Z(
        P2_U3550) );
  MUX2_X1 U15195 ( .A(n13196), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13214), .Z(
        P2_U3549) );
  MUX2_X1 U15196 ( .A(n13197), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13214), .Z(
        P2_U3548) );
  MUX2_X1 U15197 ( .A(n13198), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13214), .Z(
        P2_U3547) );
  MUX2_X1 U15198 ( .A(n13199), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13214), .Z(
        P2_U3546) );
  MUX2_X1 U15199 ( .A(n13200), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13214), .Z(
        P2_U3545) );
  MUX2_X1 U15200 ( .A(n13201), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13214), .Z(
        P2_U3544) );
  MUX2_X1 U15201 ( .A(n13202), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13214), .Z(
        P2_U3543) );
  MUX2_X1 U15202 ( .A(n13203), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13214), .Z(
        P2_U3542) );
  MUX2_X1 U15203 ( .A(n13204), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13214), .Z(
        P2_U3541) );
  MUX2_X1 U15204 ( .A(n13205), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13214), .Z(
        P2_U3540) );
  MUX2_X1 U15205 ( .A(n13206), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13214), .Z(
        P2_U3539) );
  MUX2_X1 U15206 ( .A(n13207), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13214), .Z(
        P2_U3538) );
  MUX2_X1 U15207 ( .A(n13208), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13214), .Z(
        P2_U3537) );
  MUX2_X1 U15208 ( .A(n13209), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13214), .Z(
        P2_U3536) );
  MUX2_X1 U15209 ( .A(n13210), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13214), .Z(
        P2_U3535) );
  MUX2_X1 U15210 ( .A(n13211), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13214), .Z(
        P2_U3534) );
  MUX2_X1 U15211 ( .A(n13212), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13214), .Z(
        P2_U3533) );
  MUX2_X1 U15212 ( .A(n6748), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13214), .Z(
        P2_U3532) );
  NOR2_X1 U15213 ( .A1(n13216), .A2(n13215), .ZN(n13221) );
  INV_X1 U15214 ( .A(n13221), .ZN(n13219) );
  MUX2_X1 U15215 ( .A(n13217), .B(P2_REG1_REG_11__SCAN_IN), .S(n13234), .Z(
        n13218) );
  NAND2_X1 U15216 ( .A1(n13219), .A2(n13218), .ZN(n13222) );
  MUX2_X1 U15217 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13217), .S(n13234), .Z(
        n13220) );
  OAI211_X1 U15218 ( .C1(n13223), .C2(n13222), .A(n13237), .B(n15223), .ZN(
        n13232) );
  OAI22_X1 U15219 ( .A1(n14774), .A2(n14531), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7875), .ZN(n13224) );
  AOI21_X1 U15220 ( .B1(n13234), .B2(n15226), .A(n13224), .ZN(n13231) );
  AOI21_X1 U15221 ( .B1(n13226), .B2(P2_REG2_REG_10__SCAN_IN), .A(n13225), 
        .ZN(n13228) );
  INV_X1 U15222 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13242) );
  MUX2_X1 U15223 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13242), .S(n13234), .Z(
        n13227) );
  NAND2_X1 U15224 ( .A1(n13228), .A2(n13227), .ZN(n13247) );
  OAI21_X1 U15225 ( .B1(n13228), .B2(n13227), .A(n13247), .ZN(n13229) );
  NAND2_X1 U15226 ( .A1(n13229), .A2(n14833), .ZN(n13230) );
  NAND3_X1 U15227 ( .A1(n13232), .A2(n13231), .A3(n13230), .ZN(P2_U3225) );
  INV_X1 U15228 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13233) );
  XNOR2_X1 U15229 ( .A(n13270), .B(n13233), .ZN(n13235) );
  NAND2_X1 U15230 ( .A1(n13234), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n13236) );
  NAND3_X1 U15231 ( .A1(n13237), .A2(n13235), .A3(n13236), .ZN(n13269) );
  INV_X1 U15232 ( .A(n13269), .ZN(n13239) );
  AOI21_X1 U15233 ( .B1(n13237), .B2(n13236), .A(n13235), .ZN(n13238) );
  OAI21_X1 U15234 ( .B1(n13239), .B2(n13238), .A(n15223), .ZN(n13252) );
  NOR2_X1 U15235 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13240), .ZN(n13241) );
  AOI21_X1 U15236 ( .B1(n15233), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n13241), 
        .ZN(n13251) );
  NAND2_X1 U15237 ( .A1(n13243), .A2(n13242), .ZN(n13245) );
  INV_X1 U15238 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13244) );
  MUX2_X1 U15239 ( .A(n13244), .B(P2_REG2_REG_12__SCAN_IN), .S(n13270), .Z(
        n13246) );
  AOI21_X1 U15240 ( .B1(n13247), .B2(n13245), .A(n13246), .ZN(n13253) );
  AND3_X1 U15241 ( .A1(n13247), .A2(n13246), .A3(n13245), .ZN(n13248) );
  OAI21_X1 U15242 ( .B1(n13253), .B2(n13248), .A(n14833), .ZN(n13250) );
  NAND2_X1 U15243 ( .A1(n15226), .A2(n13270), .ZN(n13249) );
  NAND4_X1 U15244 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n13249), .ZN(
        P2_U3226) );
  INV_X1 U15245 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13265) );
  INV_X1 U15246 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13258) );
  AOI21_X1 U15247 ( .B1(n13244), .B2(n13254), .A(n13253), .ZN(n14786) );
  NAND2_X1 U15248 ( .A1(n14778), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13255) );
  OAI21_X1 U15249 ( .B1(n14778), .B2(P2_REG2_REG_13__SCAN_IN), .A(n13255), 
        .ZN(n13256) );
  INV_X1 U15250 ( .A(n13256), .ZN(n14785) );
  NAND2_X1 U15251 ( .A1(n14786), .A2(n14785), .ZN(n14784) );
  OAI21_X1 U15252 ( .B1(n13258), .B2(n13257), .A(n14784), .ZN(n13259) );
  NAND2_X1 U15253 ( .A1(n14790), .A2(n13259), .ZN(n13260) );
  XNOR2_X1 U15254 ( .A(n13259), .B(n13272), .ZN(n14792) );
  NAND2_X1 U15255 ( .A1(n14792), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U15256 ( .A1(n13260), .A2(n14791), .ZN(n13261) );
  NAND2_X1 U15257 ( .A1(n14800), .A2(n13261), .ZN(n13262) );
  XNOR2_X1 U15258 ( .A(n13273), .B(n13261), .ZN(n14802) );
  NAND2_X1 U15259 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14802), .ZN(n14801) );
  NAND2_X1 U15260 ( .A1(n13262), .A2(n14801), .ZN(n14813) );
  XNOR2_X1 U15261 ( .A(n13276), .B(n13263), .ZN(n14814) );
  AOI22_X1 U15262 ( .A1(n14813), .A2(n14814), .B1(n13276), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U15263 ( .A1(n14823), .A2(n13265), .ZN(n13264) );
  OAI21_X1 U15264 ( .B1(n14823), .B2(n13265), .A(n13264), .ZN(n14830) );
  OAI21_X1 U15265 ( .B1(n14823), .B2(n13265), .A(n14834), .ZN(n13266) );
  NOR2_X1 U15266 ( .A1(n15225), .A2(n13266), .ZN(n13267) );
  XNOR2_X1 U15267 ( .A(n15225), .B(n13266), .ZN(n15221) );
  NOR2_X1 U15268 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15221), .ZN(n15220) );
  NOR2_X1 U15269 ( .A1(n13267), .A2(n15220), .ZN(n13268) );
  XOR2_X1 U15270 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13268), .Z(n13287) );
  INV_X1 U15271 ( .A(n13287), .ZN(n13285) );
  INV_X1 U15272 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13279) );
  OAI21_X1 U15273 ( .B1(n13270), .B2(P2_REG1_REG_12__SCAN_IN), .A(n13269), 
        .ZN(n14781) );
  XNOR2_X1 U15274 ( .A(n14778), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14782) );
  NOR2_X1 U15275 ( .A1(n14781), .A2(n14782), .ZN(n14779) );
  XNOR2_X1 U15276 ( .A(n14790), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14794) );
  INV_X1 U15277 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13271) );
  OAI22_X1 U15278 ( .A1(n14793), .A2(n14794), .B1(n13272), .B2(n13271), .ZN(
        n13274) );
  NAND2_X1 U15279 ( .A1(n14800), .A2(n13274), .ZN(n13275) );
  NAND2_X1 U15280 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14804), .ZN(n14803) );
  NAND2_X1 U15281 ( .A1(n13275), .A2(n14803), .ZN(n14817) );
  INV_X1 U15282 ( .A(n14817), .ZN(n13278) );
  XNOR2_X1 U15283 ( .A(n13276), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14816) );
  XNOR2_X1 U15284 ( .A(n14823), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U15285 ( .A1(n14829), .A2(n14828), .ZN(n14827) );
  OAI21_X1 U15286 ( .B1(n14823), .B2(n13279), .A(n14827), .ZN(n13280) );
  XOR2_X1 U15287 ( .A(n13280), .B(n15225), .Z(n15224) );
  NAND2_X1 U15288 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n15224), .ZN(n15222) );
  NAND2_X1 U15289 ( .A1(n15225), .A2(n13280), .ZN(n13281) );
  NAND2_X1 U15290 ( .A1(n15222), .A2(n13281), .ZN(n13283) );
  INV_X1 U15291 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13282) );
  XNOR2_X1 U15292 ( .A(n13283), .B(n13282), .ZN(n13286) );
  NOR2_X1 U15293 ( .A1(n13286), .A2(n14780), .ZN(n13284) );
  AOI211_X1 U15294 ( .C1(n13285), .C2(n14833), .A(n15226), .B(n13284), .ZN(
        n13289) );
  AOI22_X1 U15295 ( .A1(n13287), .A2(n14833), .B1(n15223), .B2(n13286), .ZN(
        n13288) );
  MUX2_X1 U15296 ( .A(n13289), .B(n13288), .S(n6754), .Z(n13291) );
  OAI211_X1 U15297 ( .C1(n7532), .C2(n14774), .A(n13291), .B(n13290), .ZN(
        P2_U3233) );
  NAND2_X1 U15298 ( .A1(n13513), .A2(n13297), .ZN(n13296) );
  NAND2_X1 U15299 ( .A1(n13293), .A2(n13292), .ZN(n13511) );
  NOR2_X1 U15300 ( .A1(n13509), .A2(n13511), .ZN(n13299) );
  NOR2_X1 U15301 ( .A1(n6992), .A2(n13498), .ZN(n13294) );
  AOI211_X1 U15302 ( .C1(n13392), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13299), 
        .B(n13294), .ZN(n13295) );
  OAI21_X1 U15303 ( .B1(n13510), .B2(n13371), .A(n13295), .ZN(P2_U3234) );
  OAI211_X1 U15304 ( .C1(n13513), .C2(n13297), .A(n10055), .B(n13296), .ZN(
        n13512) );
  NOR2_X1 U15305 ( .A1(n13513), .A2(n13498), .ZN(n13298) );
  AOI211_X1 U15306 ( .C1(n13392), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13299), 
        .B(n13298), .ZN(n13300) );
  OAI21_X1 U15307 ( .B1(n13371), .B2(n13512), .A(n13300), .ZN(P2_U3235) );
  OAI21_X1 U15308 ( .B1(n13302), .B2(n13304), .A(n13301), .ZN(n13523) );
  AOI22_X1 U15309 ( .A1(n13520), .A2(n13483), .B1(n13392), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13315) );
  OAI22_X1 U15310 ( .A1(n13306), .A2(n13445), .B1(n13305), .B2(n13447), .ZN(
        n13307) );
  AOI21_X1 U15311 ( .B1(n13520), .B2(n13322), .A(n13492), .ZN(n13310) );
  NAND2_X1 U15312 ( .A1(n13519), .A2(n6754), .ZN(n13311) );
  NAND2_X1 U15313 ( .A1(n13313), .A2(n13476), .ZN(n13314) );
  OAI211_X1 U15314 ( .C1(n13523), .C2(n13504), .A(n13315), .B(n13314), .ZN(
        P2_U3237) );
  XNOR2_X1 U15315 ( .A(n13316), .B(n13320), .ZN(n13319) );
  INV_X1 U15316 ( .A(n13317), .ZN(n13318) );
  AOI21_X1 U15317 ( .B1(n13319), .B2(n13488), .A(n13318), .ZN(n13529) );
  OR2_X1 U15318 ( .A1(n13321), .A2(n13320), .ZN(n13525) );
  NAND3_X1 U15319 ( .A1(n13525), .A2(n13524), .A3(n13387), .ZN(n13329) );
  AOI21_X1 U15320 ( .B1(n13526), .B2(n13338), .A(n13492), .ZN(n13323) );
  NAND2_X1 U15321 ( .A1(n13323), .A2(n13322), .ZN(n13528) );
  AOI22_X1 U15322 ( .A1(n13324), .A2(n13495), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13509), .ZN(n13326) );
  NAND2_X1 U15323 ( .A1(n13526), .A2(n13483), .ZN(n13325) );
  OAI211_X1 U15324 ( .C1(n13528), .C2(n13371), .A(n13326), .B(n13325), .ZN(
        n13327) );
  INV_X1 U15325 ( .A(n13327), .ZN(n13328) );
  OAI211_X1 U15326 ( .C1(n13392), .C2(n13529), .A(n13329), .B(n13328), .ZN(
        P2_U3238) );
  XNOR2_X1 U15327 ( .A(n13330), .B(n13334), .ZN(n13332) );
  AOI21_X1 U15328 ( .B1(n13332), .B2(n13488), .A(n13331), .ZN(n13534) );
  XOR2_X1 U15329 ( .A(n13333), .B(n13334), .Z(n13535) );
  INV_X1 U15330 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13335) );
  OAI22_X1 U15331 ( .A1(n13336), .A2(n13473), .B1(n13335), .B2(n13476), .ZN(
        n13337) );
  AOI21_X1 U15332 ( .B1(n13532), .B2(n13483), .A(n13337), .ZN(n13341) );
  AOI21_X1 U15333 ( .B1(n13532), .B2(n13349), .A(n13492), .ZN(n13339) );
  AND2_X1 U15334 ( .A1(n13339), .A2(n13338), .ZN(n13531) );
  NAND2_X1 U15335 ( .A1(n13531), .A2(n13507), .ZN(n13340) );
  OAI211_X1 U15336 ( .C1(n13535), .C2(n13504), .A(n13341), .B(n13340), .ZN(
        n13342) );
  INV_X1 U15337 ( .A(n13342), .ZN(n13343) );
  OAI21_X1 U15338 ( .B1(n13392), .B2(n13534), .A(n13343), .ZN(P2_U3239) );
  XNOR2_X1 U15339 ( .A(n13345), .B(n13344), .ZN(n13347) );
  AOI21_X1 U15340 ( .B1(n13347), .B2(n13488), .A(n13346), .ZN(n13539) );
  OR2_X1 U15341 ( .A1(n13352), .A2(n13365), .ZN(n13348) );
  AND3_X1 U15342 ( .A1(n13349), .A2(n13348), .A3(n10055), .ZN(n13536) );
  AOI22_X1 U15343 ( .A1(n13350), .A2(n13495), .B1(n13509), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n13351) );
  OAI21_X1 U15344 ( .B1(n13352), .B2(n13498), .A(n13351), .ZN(n13356) );
  XNOR2_X1 U15345 ( .A(n13354), .B(n13353), .ZN(n13540) );
  NOR2_X1 U15346 ( .A1(n13540), .A2(n13504), .ZN(n13355) );
  AOI211_X1 U15347 ( .C1(n13536), .C2(n13507), .A(n13356), .B(n13355), .ZN(
        n13357) );
  OAI21_X1 U15348 ( .B1(n13392), .B2(n13539), .A(n13357), .ZN(P2_U3240) );
  XNOR2_X1 U15349 ( .A(n13358), .B(n13363), .ZN(n13360) );
  AOI21_X1 U15350 ( .B1(n13360), .B2(n13488), .A(n13359), .ZN(n13542) );
  AOI21_X1 U15351 ( .B1(n13363), .B2(n13362), .A(n13361), .ZN(n13545) );
  AND2_X1 U15352 ( .A1(n13369), .A2(n13374), .ZN(n13364) );
  OR3_X1 U15353 ( .A1(n13365), .A2(n13364), .A3(n13492), .ZN(n13541) );
  INV_X1 U15354 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13367) );
  OAI22_X1 U15355 ( .A1(n13476), .A2(n13367), .B1(n13366), .B2(n13473), .ZN(
        n13368) );
  AOI21_X1 U15356 ( .B1(n13369), .B2(n13483), .A(n13368), .ZN(n13370) );
  OAI21_X1 U15357 ( .B1(n13541), .B2(n13371), .A(n13370), .ZN(n13372) );
  AOI21_X1 U15358 ( .B1(n13545), .B2(n13387), .A(n13372), .ZN(n13373) );
  OAI21_X1 U15359 ( .B1(n13392), .B2(n13542), .A(n13373), .ZN(P2_U3241) );
  OAI211_X1 U15360 ( .C1(n13549), .C2(n13399), .A(n10055), .B(n13374), .ZN(
        n13548) );
  INV_X1 U15361 ( .A(n13548), .ZN(n13383) );
  AND2_X1 U15362 ( .A1(n13375), .A2(n13435), .ZN(n13376) );
  AOI21_X1 U15363 ( .B1(n13377), .B2(n13437), .A(n13376), .ZN(n13547) );
  OAI21_X1 U15364 ( .B1(n13378), .B2(n13473), .A(n13547), .ZN(n13382) );
  NAND2_X1 U15365 ( .A1(n13379), .A2(n13385), .ZN(n13380) );
  AOI21_X1 U15366 ( .B1(n13381), .B2(n13380), .A(n13451), .ZN(n13551) );
  AOI211_X1 U15367 ( .C1(n13383), .C2(n6754), .A(n13382), .B(n13551), .ZN(
        n13391) );
  OAI21_X1 U15368 ( .B1(n13386), .B2(n13385), .A(n13384), .ZN(n13552) );
  NAND2_X1 U15369 ( .A1(n13552), .A2(n13387), .ZN(n13390) );
  AOI22_X1 U15370 ( .A1(n13388), .A2(n13483), .B1(n13392), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13389) );
  OAI211_X1 U15371 ( .C1(n13392), .C2(n13391), .A(n13390), .B(n13389), .ZN(
        P2_U3242) );
  XNOR2_X1 U15372 ( .A(n13394), .B(n13393), .ZN(n13396) );
  OAI21_X1 U15373 ( .B1(n13396), .B2(n13451), .A(n13395), .ZN(n13555) );
  NAND2_X1 U15374 ( .A1(n13421), .A2(n13557), .ZN(n13397) );
  NAND2_X1 U15375 ( .A1(n13397), .A2(n10055), .ZN(n13398) );
  NOR2_X1 U15376 ( .A1(n13399), .A2(n13398), .ZN(n13556) );
  NAND2_X1 U15377 ( .A1(n13556), .A2(n13507), .ZN(n13402) );
  AOI22_X1 U15378 ( .A1(n13509), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13400), 
        .B2(n13495), .ZN(n13401) );
  OAI211_X1 U15379 ( .C1(n13403), .C2(n13498), .A(n13402), .B(n13401), .ZN(
        n13409) );
  NAND2_X1 U15380 ( .A1(n13406), .A2(n13405), .ZN(n13554) );
  INV_X1 U15381 ( .A(n13554), .ZN(n13407) );
  NOR3_X1 U15382 ( .A1(n13404), .A2(n13407), .A3(n13504), .ZN(n13408) );
  AOI211_X1 U15383 ( .C1(n13476), .C2(n13555), .A(n13409), .B(n13408), .ZN(
        n13410) );
  INV_X1 U15384 ( .A(n13410), .ZN(P2_U3243) );
  XNOR2_X1 U15385 ( .A(n6649), .B(n13411), .ZN(n13564) );
  XNOR2_X1 U15386 ( .A(n13414), .B(n13413), .ZN(n13416) );
  AOI21_X1 U15387 ( .B1(n13416), .B2(n13488), .A(n13415), .ZN(n13563) );
  INV_X1 U15388 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13418) );
  OAI22_X1 U15389 ( .A1(n13476), .A2(n13418), .B1(n13417), .B2(n13473), .ZN(
        n13419) );
  AOI21_X1 U15390 ( .B1(n13561), .B2(n13483), .A(n13419), .ZN(n13423) );
  AOI21_X1 U15391 ( .B1(n13427), .B2(n13561), .A(n13492), .ZN(n13420) );
  AND2_X1 U15392 ( .A1(n13421), .A2(n13420), .ZN(n13560) );
  NAND2_X1 U15393 ( .A1(n13560), .A2(n13507), .ZN(n13422) );
  OAI211_X1 U15394 ( .C1(n13563), .C2(n13509), .A(n13423), .B(n13422), .ZN(
        n13424) );
  INV_X1 U15395 ( .A(n13424), .ZN(n13425) );
  OAI21_X1 U15396 ( .B1(n13564), .B2(n13504), .A(n13425), .ZN(P2_U3244) );
  XNOR2_X1 U15397 ( .A(n13426), .B(n13432), .ZN(n13569) );
  AOI21_X1 U15398 ( .B1(n13565), .B2(n13457), .A(n6489), .ZN(n13566) );
  INV_X1 U15399 ( .A(n13428), .ZN(n13429) );
  AOI22_X1 U15400 ( .A1(n13509), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13429), 
        .B2(n13495), .ZN(n13430) );
  OAI21_X1 U15401 ( .B1(n7004), .B2(n13498), .A(n13430), .ZN(n13441) );
  NAND3_X1 U15402 ( .A1(n13453), .A2(n13432), .A3(n13431), .ZN(n13433) );
  NAND2_X1 U15403 ( .A1(n13434), .A2(n13433), .ZN(n13439) );
  AOI222_X1 U15404 ( .A1(n13488), .A2(n13439), .B1(n13438), .B2(n13437), .C1(
        n13436), .C2(n13435), .ZN(n13568) );
  NOR2_X1 U15405 ( .A1(n13568), .A2(n13509), .ZN(n13440) );
  AOI211_X1 U15406 ( .C1(n13566), .C2(n13442), .A(n13441), .B(n13440), .ZN(
        n13443) );
  OAI21_X1 U15407 ( .B1(n13569), .B2(n13504), .A(n13443), .ZN(P2_U3245) );
  XNOR2_X1 U15408 ( .A(n13444), .B(n13449), .ZN(n13461) );
  OAI22_X1 U15409 ( .A1(n13448), .A2(n13447), .B1(n13446), .B2(n13445), .ZN(
        n13455) );
  NAND2_X1 U15410 ( .A1(n13450), .A2(n13449), .ZN(n13452) );
  AOI21_X1 U15411 ( .B1(n13453), .B2(n13452), .A(n13451), .ZN(n13454) );
  AOI211_X1 U15412 ( .C1(n13461), .C2(n13456), .A(n13455), .B(n13454), .ZN(
        n13573) );
  AOI211_X1 U15413 ( .C1(n13571), .C2(n13466), .A(n13492), .B(n7005), .ZN(
        n13570) );
  INV_X1 U15414 ( .A(n13458), .ZN(n13459) );
  AOI22_X1 U15415 ( .A1(n13509), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13459), 
        .B2(n13495), .ZN(n13460) );
  OAI21_X1 U15416 ( .B1(n7006), .B2(n13498), .A(n13460), .ZN(n13464) );
  INV_X1 U15417 ( .A(n13461), .ZN(n13574) );
  NOR2_X1 U15418 ( .A1(n13574), .A2(n13462), .ZN(n13463) );
  AOI211_X1 U15419 ( .C1(n13570), .C2(n13507), .A(n13464), .B(n13463), .ZN(
        n13465) );
  OAI21_X1 U15420 ( .B1(n13509), .B2(n13573), .A(n13465), .ZN(P2_U3246) );
  INV_X1 U15421 ( .A(n13466), .ZN(n13467) );
  AOI211_X1 U15422 ( .C1(n13576), .C2(n13490), .A(n13492), .B(n13467), .ZN(
        n13575) );
  XNOR2_X1 U15423 ( .A(n13480), .B(n13468), .ZN(n13470) );
  AOI21_X1 U15424 ( .B1(n13470), .B2(n13488), .A(n13469), .ZN(n13578) );
  INV_X1 U15425 ( .A(n13578), .ZN(n13471) );
  AOI21_X1 U15426 ( .B1(n13575), .B2(n6754), .A(n13471), .ZN(n13485) );
  INV_X1 U15427 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13475) );
  OAI22_X1 U15428 ( .A1(n13476), .A2(n13475), .B1(n13474), .B2(n13473), .ZN(
        n13482) );
  INV_X1 U15429 ( .A(n13477), .ZN(n13478) );
  AOI21_X1 U15430 ( .B1(n13480), .B2(n13479), .A(n13478), .ZN(n13579) );
  NOR2_X1 U15431 ( .A1(n13579), .A2(n13504), .ZN(n13481) );
  AOI211_X1 U15432 ( .C1(n13483), .C2(n13576), .A(n13482), .B(n13481), .ZN(
        n13484) );
  OAI21_X1 U15433 ( .B1(n13509), .B2(n13485), .A(n13484), .ZN(P2_U3247) );
  XNOR2_X1 U15434 ( .A(n13486), .B(n13500), .ZN(n13489) );
  AOI21_X1 U15435 ( .B1(n13489), .B2(n13488), .A(n13487), .ZN(n13583) );
  INV_X1 U15436 ( .A(n13490), .ZN(n13491) );
  AOI211_X1 U15437 ( .C1(n13581), .C2(n13493), .A(n13492), .B(n13491), .ZN(
        n13580) );
  INV_X1 U15438 ( .A(n13581), .ZN(n13499) );
  INV_X1 U15439 ( .A(n13494), .ZN(n13496) );
  AOI22_X1 U15440 ( .A1(n13509), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13496), 
        .B2(n13495), .ZN(n13497) );
  OAI21_X1 U15441 ( .B1(n13499), .B2(n13498), .A(n13497), .ZN(n13506) );
  OR2_X1 U15442 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  NAND2_X1 U15443 ( .A1(n13503), .A2(n13502), .ZN(n13584) );
  NOR2_X1 U15444 ( .A1(n13584), .A2(n13504), .ZN(n13505) );
  AOI211_X1 U15445 ( .C1(n13580), .C2(n13507), .A(n13506), .B(n13505), .ZN(
        n13508) );
  OAI21_X1 U15446 ( .B1(n13509), .B2(n13583), .A(n13508), .ZN(P2_U3248) );
  OAI211_X1 U15447 ( .C1(n13513), .C2(n14859), .A(n13512), .B(n13511), .ZN(
        n13607) );
  MUX2_X1 U15448 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13607), .S(n14895), .Z(
        P2_U3529) );
  AOI21_X1 U15449 ( .B1(n14877), .B2(n13515), .A(n13514), .ZN(n13516) );
  MUX2_X1 U15450 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13608), .S(n14895), .Z(
        P2_U3528) );
  AOI21_X1 U15451 ( .B1(n14877), .B2(n13520), .A(n13519), .ZN(n13521) );
  OAI211_X1 U15452 ( .C1(n13523), .C2(n14875), .A(n13522), .B(n13521), .ZN(
        n13609) );
  MUX2_X1 U15453 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13609), .S(n14895), .Z(
        P2_U3527) );
  NAND3_X1 U15454 ( .A1(n13525), .A2(n13524), .A3(n14865), .ZN(n13530) );
  NAND2_X1 U15455 ( .A1(n13526), .A2(n14877), .ZN(n13527) );
  NAND4_X1 U15456 ( .A1(n13530), .A2(n13529), .A3(n13528), .A4(n13527), .ZN(
        n13610) );
  MUX2_X1 U15457 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13610), .S(n14895), .Z(
        P2_U3526) );
  AOI21_X1 U15458 ( .B1(n14877), .B2(n13532), .A(n13531), .ZN(n13533) );
  OAI211_X1 U15459 ( .C1(n13535), .C2(n14875), .A(n13534), .B(n13533), .ZN(
        n13611) );
  MUX2_X1 U15460 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13611), .S(n14895), .Z(
        P2_U3525) );
  AOI21_X1 U15461 ( .B1(n14877), .B2(n13537), .A(n13536), .ZN(n13538) );
  OAI211_X1 U15462 ( .C1(n13540), .C2(n14875), .A(n13539), .B(n13538), .ZN(
        n13612) );
  MUX2_X1 U15463 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13612), .S(n14895), .Z(
        P2_U3524) );
  OAI211_X1 U15464 ( .C1(n13543), .C2(n14859), .A(n13542), .B(n13541), .ZN(
        n13544) );
  AOI21_X1 U15465 ( .B1(n13545), .B2(n14865), .A(n13544), .ZN(n13546) );
  INV_X1 U15466 ( .A(n13546), .ZN(n13613) );
  MUX2_X1 U15467 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13613), .S(n14895), .Z(
        P2_U3523) );
  OAI211_X1 U15468 ( .C1(n13549), .C2(n14859), .A(n13548), .B(n13547), .ZN(
        n13550) );
  AOI211_X1 U15469 ( .C1(n13552), .C2(n14865), .A(n13551), .B(n13550), .ZN(
        n13553) );
  INV_X1 U15470 ( .A(n13553), .ZN(n13614) );
  MUX2_X1 U15471 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13614), .S(n14895), .Z(
        P2_U3522) );
  NAND2_X1 U15472 ( .A1(n13554), .A2(n14865), .ZN(n13559) );
  AOI211_X1 U15473 ( .C1(n14877), .C2(n13557), .A(n13556), .B(n13555), .ZN(
        n13558) );
  OAI21_X1 U15474 ( .B1(n13404), .B2(n13559), .A(n13558), .ZN(n13615) );
  MUX2_X1 U15475 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13615), .S(n14895), .Z(
        P2_U3521) );
  AOI21_X1 U15476 ( .B1(n14877), .B2(n13561), .A(n13560), .ZN(n13562) );
  OAI211_X1 U15477 ( .C1(n13564), .C2(n14875), .A(n13563), .B(n13562), .ZN(
        n13616) );
  MUX2_X1 U15478 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13616), .S(n14895), .Z(
        P2_U3520) );
  AOI22_X1 U15479 ( .A1(n13566), .A2(n10055), .B1(n14877), .B2(n13565), .ZN(
        n13567) );
  OAI211_X1 U15480 ( .C1(n14875), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        n13617) );
  MUX2_X1 U15481 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13617), .S(n14895), .Z(
        P2_U3519) );
  AOI21_X1 U15482 ( .B1(n14877), .B2(n13571), .A(n13570), .ZN(n13572) );
  OAI211_X1 U15483 ( .C1(n13574), .C2(n14871), .A(n13573), .B(n13572), .ZN(
        n13618) );
  MUX2_X1 U15484 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13618), .S(n14895), .Z(
        P2_U3518) );
  AOI21_X1 U15485 ( .B1(n14877), .B2(n13576), .A(n13575), .ZN(n13577) );
  OAI211_X1 U15486 ( .C1(n13579), .C2(n14875), .A(n13578), .B(n13577), .ZN(
        n13619) );
  MUX2_X1 U15487 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13619), .S(n14895), .Z(
        P2_U3517) );
  AOI21_X1 U15488 ( .B1(n14877), .B2(n13581), .A(n13580), .ZN(n13582) );
  OAI211_X1 U15489 ( .C1(n13584), .C2(n14875), .A(n13583), .B(n13582), .ZN(
        n13620) );
  MUX2_X1 U15490 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13620), .S(n14895), .Z(
        P2_U3516) );
  AOI211_X1 U15491 ( .C1(n14877), .C2(n13587), .A(n13586), .B(n13585), .ZN(
        n13589) );
  OAI211_X1 U15492 ( .C1(n14875), .C2(n13590), .A(n13589), .B(n13588), .ZN(
        n13621) );
  MUX2_X1 U15493 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13621), .S(n14895), .Z(
        P2_U3515) );
  AOI211_X1 U15494 ( .C1(n14877), .C2(n13593), .A(n13592), .B(n13591), .ZN(
        n13594) );
  OAI21_X1 U15495 ( .B1(n14875), .B2(n13595), .A(n13594), .ZN(n13622) );
  MUX2_X1 U15496 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13622), .S(n14895), .Z(
        P2_U3514) );
  AOI211_X1 U15497 ( .C1(n14877), .C2(n13598), .A(n13597), .B(n13596), .ZN(
        n13599) );
  OAI21_X1 U15498 ( .B1(n14875), .B2(n13600), .A(n13599), .ZN(n13623) );
  MUX2_X1 U15499 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13623), .S(n14895), .Z(
        P2_U3513) );
  AOI211_X1 U15500 ( .C1(n14877), .C2(n13603), .A(n13602), .B(n13601), .ZN(
        n13604) );
  OAI21_X1 U15501 ( .B1(n14875), .B2(n13605), .A(n13604), .ZN(n13624) );
  MUX2_X1 U15502 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13624), .S(n14895), .Z(
        P2_U3512) );
  MUX2_X1 U15503 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13606), .S(n14886), .Z(
        P2_U3498) );
  MUX2_X1 U15504 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13607), .S(n14886), .Z(
        P2_U3497) );
  MUX2_X1 U15505 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13608), .S(n14886), .Z(
        P2_U3496) );
  MUX2_X1 U15506 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13609), .S(n14886), .Z(
        P2_U3495) );
  MUX2_X1 U15507 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13610), .S(n14886), .Z(
        P2_U3494) );
  MUX2_X1 U15508 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13611), .S(n14886), .Z(
        P2_U3493) );
  MUX2_X1 U15509 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13612), .S(n14886), .Z(
        P2_U3492) );
  MUX2_X1 U15510 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13613), .S(n14886), .Z(
        P2_U3491) );
  MUX2_X1 U15511 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13614), .S(n14886), .Z(
        P2_U3490) );
  MUX2_X1 U15512 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13615), .S(n14886), .Z(
        P2_U3489) );
  MUX2_X1 U15513 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13616), .S(n14886), .Z(
        P2_U3488) );
  MUX2_X1 U15514 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13617), .S(n14886), .Z(
        P2_U3487) );
  MUX2_X1 U15515 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13618), .S(n14886), .Z(
        P2_U3486) );
  MUX2_X1 U15516 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13619), .S(n14886), .Z(
        P2_U3484) );
  MUX2_X1 U15517 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13620), .S(n14886), .Z(
        P2_U3481) );
  MUX2_X1 U15518 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13621), .S(n14886), .Z(
        P2_U3478) );
  MUX2_X1 U15519 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13622), .S(n14886), .Z(
        P2_U3475) );
  MUX2_X1 U15520 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13623), .S(n14886), .Z(
        P2_U3472) );
  MUX2_X1 U15521 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13624), .S(n14886), .Z(
        P2_U3469) );
  INV_X1 U15522 ( .A(n13625), .ZN(n14371) );
  NOR4_X1 U15523 ( .A1(n13626), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7709), .A4(
        P2_U3088), .ZN(n13627) );
  AOI21_X1 U15524 ( .B1(n13633), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13627), 
        .ZN(n13628) );
  OAI21_X1 U15525 ( .B1(n14371), .B2(n13637), .A(n13628), .ZN(P2_U3296) );
  INV_X1 U15526 ( .A(n13629), .ZN(n14372) );
  OAI222_X1 U15527 ( .A1(P2_U3088), .A2(n13630), .B1(n13637), .B2(n14372), 
        .C1(n13636), .C2(n8237), .ZN(P2_U3298) );
  INV_X1 U15528 ( .A(n13631), .ZN(n14375) );
  AOI21_X1 U15529 ( .B1(n13633), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13632), 
        .ZN(n13634) );
  OAI21_X1 U15530 ( .B1(n14375), .B2(n13637), .A(n13634), .ZN(P2_U3299) );
  INV_X1 U15531 ( .A(n13635), .ZN(n14381) );
  OAI222_X1 U15532 ( .A1(n13638), .A2(P2_U3088), .B1(n13637), .B2(n14381), 
        .C1(n7043), .C2(n13636), .ZN(P2_U3301) );
  INV_X1 U15533 ( .A(n13639), .ZN(n13640) );
  MUX2_X1 U15534 ( .A(n13640), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15535 ( .A1(n14093), .A2(n14691), .ZN(n14279) );
  NAND2_X1 U15536 ( .A1(n14093), .A2(n13800), .ZN(n13642) );
  NAND2_X1 U15537 ( .A1(n13924), .A2(n6487), .ZN(n13641) );
  NAND2_X1 U15538 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  XNOR2_X1 U15539 ( .A(n13643), .B(n13798), .ZN(n13647) );
  NAND2_X1 U15540 ( .A1(n14093), .A2(n6487), .ZN(n13645) );
  NAND2_X1 U15541 ( .A1(n13924), .A2(n13764), .ZN(n13644) );
  NAND2_X1 U15542 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  NOR2_X1 U15543 ( .A1(n13647), .A2(n13646), .ZN(n13796) );
  AOI21_X1 U15544 ( .B1(n13647), .B2(n13646), .A(n13796), .ZN(n13772) );
  INV_X1 U15545 ( .A(n13648), .ZN(n13651) );
  INV_X1 U15546 ( .A(n13649), .ZN(n13650) );
  NAND2_X1 U15547 ( .A1(n13651), .A2(n13650), .ZN(n13652) );
  NAND2_X1 U15548 ( .A1(n14492), .A2(n13800), .ZN(n13655) );
  NAND2_X1 U15549 ( .A1(n13937), .A2(n6487), .ZN(n13654) );
  NAND2_X1 U15550 ( .A1(n13655), .A2(n13654), .ZN(n13656) );
  XNOR2_X1 U15551 ( .A(n13656), .B(n13798), .ZN(n13665) );
  AND2_X1 U15552 ( .A1(n13937), .A2(n13764), .ZN(n13657) );
  AOI21_X1 U15553 ( .B1(n14492), .B2(n6487), .A(n13657), .ZN(n13663) );
  XNOR2_X1 U15554 ( .A(n13665), .B(n13663), .ZN(n14490) );
  NAND2_X1 U15555 ( .A1(n14489), .A2(n14490), .ZN(n14488) );
  NAND2_X1 U15556 ( .A1(n14518), .A2(n13800), .ZN(n13659) );
  NAND2_X1 U15557 ( .A1(n13936), .A2(n6487), .ZN(n13658) );
  NAND2_X1 U15558 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  XNOR2_X1 U15559 ( .A(n13660), .B(n13798), .ZN(n13667) );
  NOR2_X1 U15560 ( .A1(n13661), .A2(n13689), .ZN(n13662) );
  AOI21_X1 U15561 ( .B1(n14518), .B2(n6487), .A(n13662), .ZN(n13668) );
  XNOR2_X1 U15562 ( .A(n13667), .B(n13668), .ZN(n14465) );
  INV_X1 U15563 ( .A(n13663), .ZN(n13664) );
  NAND2_X1 U15564 ( .A1(n13665), .A2(n13664), .ZN(n14463) );
  AND2_X1 U15565 ( .A1(n14465), .A2(n14463), .ZN(n13666) );
  NAND2_X1 U15566 ( .A1(n14488), .A2(n13666), .ZN(n14464) );
  INV_X1 U15567 ( .A(n13667), .ZN(n13669) );
  NAND2_X1 U15568 ( .A1(n13669), .A2(n13668), .ZN(n13670) );
  NAND2_X1 U15569 ( .A1(n14464), .A2(n13670), .ZN(n13677) );
  NAND2_X1 U15570 ( .A1(n14345), .A2(n13800), .ZN(n13672) );
  NAND2_X1 U15571 ( .A1(n13935), .A2(n6487), .ZN(n13671) );
  NAND2_X1 U15572 ( .A1(n13672), .A2(n13671), .ZN(n13673) );
  XNOR2_X1 U15573 ( .A(n13673), .B(n13752), .ZN(n13676) );
  NAND2_X1 U15574 ( .A1(n13677), .A2(n13676), .ZN(n13914) );
  OAI22_X1 U15575 ( .A1(n6744), .A2(n13690), .B1(n13674), .B2(n13689), .ZN(
        n13912) );
  NAND2_X1 U15576 ( .A1(n13914), .A2(n13912), .ZN(n13909) );
  AOI22_X1 U15577 ( .A1(n13839), .A2(n13800), .B1(n6487), .B2(n13934), .ZN(
        n13678) );
  XNOR2_X1 U15578 ( .A(n13678), .B(n13798), .ZN(n13680) );
  AOI22_X1 U15579 ( .A1(n13839), .A2(n9526), .B1(n13764), .B2(n13934), .ZN(
        n13679) );
  XNOR2_X1 U15580 ( .A(n13680), .B(n13679), .ZN(n13834) );
  OAI22_X1 U15581 ( .A1(n14246), .A2(n13682), .B1(n13681), .B2(n13690), .ZN(
        n13683) );
  XNOR2_X1 U15582 ( .A(n13683), .B(n13752), .ZN(n13843) );
  OR2_X1 U15583 ( .A1(n14246), .A2(n13690), .ZN(n13685) );
  NAND2_X1 U15584 ( .A1(n13933), .A2(n13764), .ZN(n13684) );
  AND2_X1 U15585 ( .A1(n13685), .A2(n13684), .ZN(n13686) );
  NAND2_X1 U15586 ( .A1(n13843), .A2(n13686), .ZN(n13688) );
  INV_X1 U15587 ( .A(n13843), .ZN(n13687) );
  INV_X1 U15588 ( .A(n13686), .ZN(n13842) );
  INV_X1 U15589 ( .A(n14232), .ZN(n14334) );
  OAI22_X1 U15590 ( .A1(n14334), .A2(n13690), .B1(n13849), .B2(n13689), .ZN(
        n13700) );
  NAND2_X1 U15591 ( .A1(n14232), .A2(n13800), .ZN(n13693) );
  NAND2_X1 U15592 ( .A1(n13691), .A2(n6487), .ZN(n13692) );
  NAND2_X1 U15593 ( .A1(n13693), .A2(n13692), .ZN(n13694) );
  XNOR2_X1 U15594 ( .A(n13694), .B(n13798), .ZN(n13699) );
  XOR2_X1 U15595 ( .A(n13700), .B(n13699), .Z(n13887) );
  NAND2_X1 U15596 ( .A1(n14327), .A2(n13800), .ZN(n13696) );
  NAND2_X1 U15597 ( .A1(n13932), .A2(n6487), .ZN(n13695) );
  NAND2_X1 U15598 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  XNOR2_X1 U15599 ( .A(n13697), .B(n13798), .ZN(n13703) );
  AND2_X1 U15600 ( .A1(n13932), .A2(n13764), .ZN(n13698) );
  AOI21_X1 U15601 ( .B1(n14327), .B2(n9526), .A(n13698), .ZN(n13704) );
  XNOR2_X1 U15602 ( .A(n13703), .B(n13704), .ZN(n13790) );
  INV_X1 U15603 ( .A(n13699), .ZN(n13702) );
  INV_X1 U15604 ( .A(n13700), .ZN(n13701) );
  NAND2_X1 U15605 ( .A1(n13702), .A2(n13701), .ZN(n13788) );
  AND2_X1 U15606 ( .A1(n13931), .A2(n13764), .ZN(n13707) );
  AOI21_X1 U15607 ( .B1(n14319), .B2(n6487), .A(n13707), .ZN(n13710) );
  AOI22_X1 U15608 ( .A1(n14319), .A2(n13800), .B1(n6487), .B2(n13931), .ZN(
        n13708) );
  XNOR2_X1 U15609 ( .A(n13708), .B(n13798), .ZN(n13709) );
  XOR2_X1 U15610 ( .A(n13710), .B(n13709), .Z(n13865) );
  INV_X1 U15611 ( .A(n13709), .ZN(n13712) );
  INV_X1 U15612 ( .A(n13710), .ZN(n13711) );
  NAND2_X1 U15613 ( .A1(n14314), .A2(n13800), .ZN(n13714) );
  NAND2_X1 U15614 ( .A1(n13930), .A2(n6487), .ZN(n13713) );
  NAND2_X1 U15615 ( .A1(n13714), .A2(n13713), .ZN(n13715) );
  XNOR2_X1 U15616 ( .A(n13715), .B(n13798), .ZN(n13719) );
  NAND2_X1 U15617 ( .A1(n14314), .A2(n6487), .ZN(n13717) );
  NAND2_X1 U15618 ( .A1(n13930), .A2(n13764), .ZN(n13716) );
  NAND2_X1 U15619 ( .A1(n13717), .A2(n13716), .ZN(n13718) );
  NOR2_X1 U15620 ( .A1(n13719), .A2(n13718), .ZN(n13720) );
  AOI21_X1 U15621 ( .B1(n13719), .B2(n13718), .A(n13720), .ZN(n13812) );
  INV_X1 U15622 ( .A(n13720), .ZN(n13874) );
  NAND2_X1 U15623 ( .A1(n14308), .A2(n13800), .ZN(n13722) );
  NAND2_X1 U15624 ( .A1(n13929), .A2(n6487), .ZN(n13721) );
  NAND2_X1 U15625 ( .A1(n13722), .A2(n13721), .ZN(n13723) );
  XNOR2_X1 U15626 ( .A(n13723), .B(n13752), .ZN(n13725) );
  AND2_X1 U15627 ( .A1(n13929), .A2(n13764), .ZN(n13724) );
  AOI21_X1 U15628 ( .B1(n14308), .B2(n6487), .A(n13724), .ZN(n13726) );
  NAND2_X1 U15629 ( .A1(n13725), .A2(n13726), .ZN(n13730) );
  INV_X1 U15630 ( .A(n13725), .ZN(n13728) );
  INV_X1 U15631 ( .A(n13726), .ZN(n13727) );
  NAND2_X1 U15632 ( .A1(n13728), .A2(n13727), .ZN(n13729) );
  NAND2_X1 U15633 ( .A1(n13730), .A2(n13729), .ZN(n13873) );
  INV_X1 U15634 ( .A(n13730), .ZN(n13781) );
  NAND2_X1 U15635 ( .A1(n14156), .A2(n13800), .ZN(n13732) );
  NAND2_X1 U15636 ( .A1(n13928), .A2(n6487), .ZN(n13731) );
  NAND2_X1 U15637 ( .A1(n13732), .A2(n13731), .ZN(n13733) );
  XNOR2_X1 U15638 ( .A(n13733), .B(n13752), .ZN(n13735) );
  AND2_X1 U15639 ( .A1(n13928), .A2(n13764), .ZN(n13734) );
  AOI21_X1 U15640 ( .B1(n14156), .B2(n6487), .A(n13734), .ZN(n13736) );
  NAND2_X1 U15641 ( .A1(n13735), .A2(n13736), .ZN(n13858) );
  INV_X1 U15642 ( .A(n13735), .ZN(n13738) );
  INV_X1 U15643 ( .A(n13736), .ZN(n13737) );
  NAND2_X1 U15644 ( .A1(n13738), .A2(n13737), .ZN(n13739) );
  AND2_X1 U15645 ( .A1(n13858), .A2(n13739), .ZN(n13780) );
  NAND2_X1 U15646 ( .A1(n14295), .A2(n13800), .ZN(n13741) );
  NAND2_X1 U15647 ( .A1(n13927), .A2(n6487), .ZN(n13740) );
  NAND2_X1 U15648 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  XNOR2_X1 U15649 ( .A(n13742), .B(n13752), .ZN(n13744) );
  AND2_X1 U15650 ( .A1(n13927), .A2(n13764), .ZN(n13743) );
  AOI21_X1 U15651 ( .B1(n14295), .B2(n6487), .A(n13743), .ZN(n13745) );
  NAND2_X1 U15652 ( .A1(n13744), .A2(n13745), .ZN(n13749) );
  INV_X1 U15653 ( .A(n13744), .ZN(n13747) );
  INV_X1 U15654 ( .A(n13745), .ZN(n13746) );
  NAND2_X1 U15655 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U15656 ( .A1(n13749), .A2(n13748), .ZN(n13857) );
  INV_X1 U15657 ( .A(n13749), .ZN(n13827) );
  NAND2_X1 U15658 ( .A1(n14290), .A2(n13800), .ZN(n13751) );
  NAND2_X1 U15659 ( .A1(n13926), .A2(n6487), .ZN(n13750) );
  NAND2_X1 U15660 ( .A1(n13751), .A2(n13750), .ZN(n13753) );
  XNOR2_X1 U15661 ( .A(n13753), .B(n13752), .ZN(n13755) );
  AND2_X1 U15662 ( .A1(n13926), .A2(n13764), .ZN(n13754) );
  AOI21_X1 U15663 ( .B1(n14290), .B2(n6487), .A(n13754), .ZN(n13756) );
  NAND2_X1 U15664 ( .A1(n13755), .A2(n13756), .ZN(n13760) );
  INV_X1 U15665 ( .A(n13755), .ZN(n13758) );
  INV_X1 U15666 ( .A(n13756), .ZN(n13757) );
  NAND2_X1 U15667 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  AND2_X1 U15668 ( .A1(n13760), .A2(n13759), .ZN(n13826) );
  NAND2_X1 U15669 ( .A1(n14283), .A2(n13800), .ZN(n13762) );
  NAND2_X1 U15670 ( .A1(n13925), .A2(n6487), .ZN(n13761) );
  NAND2_X1 U15671 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  XNOR2_X1 U15672 ( .A(n13763), .B(n13798), .ZN(n13768) );
  NAND2_X1 U15673 ( .A1(n14283), .A2(n6487), .ZN(n13766) );
  NAND2_X1 U15674 ( .A1(n13925), .A2(n13764), .ZN(n13765) );
  NAND2_X1 U15675 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  NOR2_X1 U15676 ( .A1(n13768), .A2(n13767), .ZN(n13769) );
  AOI21_X1 U15677 ( .B1(n13768), .B2(n13767), .A(n13769), .ZN(n13896) );
  NAND2_X1 U15678 ( .A1(n13895), .A2(n13896), .ZN(n13894) );
  INV_X1 U15679 ( .A(n13769), .ZN(n13770) );
  OAI21_X1 U15680 ( .B1(n13772), .B2(n13771), .A(n13797), .ZN(n13773) );
  NAND2_X1 U15681 ( .A1(n13923), .A2(n13898), .ZN(n13775) );
  NAND2_X1 U15682 ( .A1(n13925), .A2(n13899), .ZN(n13774) );
  AND2_X1 U15683 ( .A1(n13775), .A2(n13774), .ZN(n14086) );
  INV_X1 U15684 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13776) );
  OAI22_X1 U15685 ( .A1(n14086), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13776), .ZN(n13777) );
  AOI21_X1 U15686 ( .B1(n13904), .B2(n14092), .A(n13777), .ZN(n13778) );
  INV_X1 U15687 ( .A(n14156), .ZN(n14301) );
  INV_X1 U15688 ( .A(n13859), .ZN(n13783) );
  NOR3_X1 U15689 ( .A1(n13877), .A2(n13781), .A3(n13780), .ZN(n13782) );
  OAI21_X1 U15690 ( .B1(n13783), .B2(n13782), .A(n14504), .ZN(n13787) );
  AOI22_X1 U15691 ( .A1(n13899), .A2(n13929), .B1(n13927), .B2(n13898), .ZN(
        n14299) );
  OAI22_X1 U15692 ( .A1(n14299), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13784), .ZN(n13785) );
  AOI21_X1 U15693 ( .B1(n14153), .B2(n13904), .A(n13785), .ZN(n13786) );
  OAI211_X1 U15694 ( .C1(n14301), .C2(n13907), .A(n13787), .B(n13786), .ZN(
        P1_U3216) );
  AND2_X1 U15695 ( .A1(n13885), .A2(n13788), .ZN(n13791) );
  OAI211_X1 U15696 ( .C1(n13791), .C2(n13790), .A(n14504), .B(n13789), .ZN(
        n13795) );
  OAI22_X1 U15697 ( .A1(n13792), .A2(n13848), .B1(n13849), .B2(n13846), .ZN(
        n14217) );
  NAND2_X1 U15698 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14047)
         );
  OAI21_X1 U15699 ( .B1(n14511), .B2(n14214), .A(n14047), .ZN(n13793) );
  AOI21_X1 U15700 ( .B1(n14217), .B2(n14506), .A(n13793), .ZN(n13794) );
  OAI211_X1 U15701 ( .C1(n7201), .C2(n13907), .A(n13795), .B(n13794), .ZN(
        P1_U3219) );
  XNOR2_X1 U15702 ( .A(n13799), .B(n13798), .ZN(n13802) );
  AOI22_X1 U15703 ( .A1(n14270), .A2(n13800), .B1(n6487), .B2(n13923), .ZN(
        n13801) );
  XNOR2_X1 U15704 ( .A(n13802), .B(n13801), .ZN(n13803) );
  NAND2_X1 U15705 ( .A1(n13804), .A2(n13898), .ZN(n13806) );
  NAND2_X1 U15706 ( .A1(n13924), .A2(n13899), .ZN(n13805) );
  AND2_X1 U15707 ( .A1(n13806), .A2(n13805), .ZN(n14067) );
  OAI22_X1 U15708 ( .A1(n14067), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13807), .ZN(n13808) );
  AOI21_X1 U15709 ( .B1(n13904), .B2(n14074), .A(n13808), .ZN(n13810) );
  NAND2_X1 U15710 ( .A1(n14270), .A2(n14502), .ZN(n13809) );
  OAI211_X1 U15711 ( .C1(n13811), .C2(n14475), .A(n13810), .B(n13809), .ZN(
        P1_U3220) );
  INV_X1 U15712 ( .A(n14314), .ZN(n13821) );
  OAI21_X1 U15713 ( .B1(n13813), .B2(n13812), .A(n13875), .ZN(n13814) );
  NAND2_X1 U15714 ( .A1(n13814), .A2(n14504), .ZN(n13820) );
  NAND2_X1 U15715 ( .A1(n13931), .A2(n13899), .ZN(n13816) );
  NAND2_X1 U15716 ( .A1(n13929), .A2(n13898), .ZN(n13815) );
  NAND2_X1 U15717 ( .A1(n13816), .A2(n13815), .ZN(n14182) );
  INV_X1 U15718 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13817) );
  OAI22_X1 U15719 ( .A1(n14189), .A2(n14511), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13817), .ZN(n13818) );
  AOI21_X1 U15720 ( .B1(n14182), .B2(n14506), .A(n13818), .ZN(n13819) );
  OAI211_X1 U15721 ( .C1(n13821), .C2(n13907), .A(n13820), .B(n13819), .ZN(
        P1_U3223) );
  NAND2_X1 U15722 ( .A1(n13927), .A2(n13899), .ZN(n13823) );
  NAND2_X1 U15723 ( .A1(n13925), .A2(n13898), .ZN(n13822) );
  NAND2_X1 U15724 ( .A1(n13823), .A2(n13822), .ZN(n14289) );
  AOI22_X1 U15725 ( .A1(n14289), .A2(n14506), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13824) );
  OAI21_X1 U15726 ( .B1(n14511), .B2(n14121), .A(n13824), .ZN(n13831) );
  OR3_X1 U15727 ( .A1(n13825), .A2(n13827), .A3(n13826), .ZN(n13828) );
  AOI21_X1 U15728 ( .B1(n13829), .B2(n13828), .A(n14475), .ZN(n13830) );
  AOI211_X1 U15729 ( .C1(n14502), .C2(n14290), .A(n13831), .B(n13830), .ZN(
        n13832) );
  INV_X1 U15730 ( .A(n13832), .ZN(P1_U3225) );
  AOI21_X1 U15731 ( .B1(n13834), .B2(n13908), .A(n13833), .ZN(n13841) );
  NAND2_X1 U15732 ( .A1(n13904), .A2(n13835), .ZN(n13836) );
  NAND2_X1 U15733 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14598)
         );
  OAI211_X1 U15734 ( .C1(n13837), .C2(n14481), .A(n13836), .B(n14598), .ZN(
        n13838) );
  AOI21_X1 U15735 ( .B1(n13839), .B2(n14502), .A(n13838), .ZN(n13840) );
  OAI21_X1 U15736 ( .B1(n13841), .B2(n14475), .A(n13840), .ZN(P1_U3226) );
  XNOR2_X1 U15737 ( .A(n13843), .B(n13842), .ZN(n13844) );
  XNOR2_X1 U15738 ( .A(n13845), .B(n13844), .ZN(n13853) );
  OAI22_X1 U15739 ( .A1(n13849), .A2(n13848), .B1(n13847), .B2(n13846), .ZN(
        n14242) );
  NAND2_X1 U15740 ( .A1(n14242), .A2(n14506), .ZN(n13850) );
  NAND2_X1 U15741 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14612)
         );
  OAI211_X1 U15742 ( .C1(n14511), .C2(n14249), .A(n13850), .B(n14612), .ZN(
        n13851) );
  AOI21_X1 U15743 ( .B1(n14340), .B2(n14502), .A(n13851), .ZN(n13852) );
  OAI21_X1 U15744 ( .B1(n13853), .B2(n14475), .A(n13852), .ZN(P1_U3228) );
  NAND2_X1 U15745 ( .A1(n13928), .A2(n13899), .ZN(n13855) );
  NAND2_X1 U15746 ( .A1(n13926), .A2(n13898), .ZN(n13854) );
  NAND2_X1 U15747 ( .A1(n13855), .A2(n13854), .ZN(n14129) );
  AOI22_X1 U15748 ( .A1(n14129), .A2(n14506), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13856) );
  OAI21_X1 U15749 ( .B1(n14511), .B2(n14134), .A(n13856), .ZN(n13863) );
  INV_X1 U15750 ( .A(n13825), .ZN(n13861) );
  NAND3_X1 U15751 ( .A1(n13859), .A2(n13858), .A3(n13857), .ZN(n13860) );
  AOI21_X1 U15752 ( .B1(n13861), .B2(n13860), .A(n14475), .ZN(n13862) );
  AOI211_X1 U15753 ( .C1(n14502), .C2(n14295), .A(n13863), .B(n13862), .ZN(
        n13864) );
  INV_X1 U15754 ( .A(n13864), .ZN(P1_U3229) );
  XNOR2_X1 U15755 ( .A(n13866), .B(n13865), .ZN(n13872) );
  AND2_X1 U15756 ( .A1(n13932), .A2(n13899), .ZN(n13867) );
  AOI21_X1 U15757 ( .B1(n13930), .B2(n13898), .A(n13867), .ZN(n14317) );
  INV_X1 U15758 ( .A(n13868), .ZN(n14197) );
  AOI22_X1 U15759 ( .A1(n13904), .A2(n14197), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13869) );
  OAI21_X1 U15760 ( .B1(n14317), .B2(n14481), .A(n13869), .ZN(n13870) );
  AOI21_X1 U15761 ( .B1(n14319), .B2(n14502), .A(n13870), .ZN(n13871) );
  OAI21_X1 U15762 ( .B1(n13872), .B2(n14475), .A(n13871), .ZN(P1_U3233) );
  AND3_X1 U15763 ( .A1(n13875), .A2(n13874), .A3(n13873), .ZN(n13876) );
  OAI21_X1 U15764 ( .B1(n13877), .B2(n13876), .A(n14504), .ZN(n13884) );
  NAND2_X1 U15765 ( .A1(n13930), .A2(n13899), .ZN(n13879) );
  NAND2_X1 U15766 ( .A1(n13928), .A2(n13898), .ZN(n13878) );
  NAND2_X1 U15767 ( .A1(n13879), .A2(n13878), .ZN(n14164) );
  INV_X1 U15768 ( .A(n14171), .ZN(n13881) );
  OAI22_X1 U15769 ( .A1(n14511), .A2(n13881), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13880), .ZN(n13882) );
  AOI21_X1 U15770 ( .B1(n14164), .B2(n14506), .A(n13882), .ZN(n13883) );
  OAI211_X1 U15771 ( .C1(n13907), .C2(n14174), .A(n13884), .B(n13883), .ZN(
        P1_U3235) );
  OAI21_X1 U15772 ( .B1(n13887), .B2(n13886), .A(n13885), .ZN(n13888) );
  NAND2_X1 U15773 ( .A1(n13888), .A2(n14504), .ZN(n13893) );
  INV_X1 U15774 ( .A(n13889), .ZN(n14229) );
  AND2_X1 U15775 ( .A1(n13933), .A2(n13899), .ZN(n13890) );
  AOI21_X1 U15776 ( .B1(n13932), .B2(n13898), .A(n13890), .ZN(n14227) );
  NAND2_X1 U15777 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14631)
         );
  OAI21_X1 U15778 ( .B1(n14227), .B2(n14481), .A(n14631), .ZN(n13891) );
  AOI21_X1 U15779 ( .B1(n14229), .B2(n13904), .A(n13891), .ZN(n13892) );
  OAI211_X1 U15780 ( .C1(n14334), .C2(n13907), .A(n13893), .B(n13892), .ZN(
        P1_U3238) );
  OAI21_X1 U15781 ( .B1(n13896), .B2(n13895), .A(n13894), .ZN(n13897) );
  NAND2_X1 U15782 ( .A1(n13897), .A2(n14504), .ZN(n13906) );
  NAND2_X1 U15783 ( .A1(n13924), .A2(n13898), .ZN(n13901) );
  NAND2_X1 U15784 ( .A1(n13926), .A2(n13899), .ZN(n13900) );
  AND2_X1 U15785 ( .A1(n13901), .A2(n13900), .ZN(n14280) );
  OAI22_X1 U15786 ( .A1(n14280), .A2(n14481), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13902), .ZN(n13903) );
  AOI21_X1 U15787 ( .B1(n13904), .B2(n14099), .A(n13903), .ZN(n13905) );
  OAI211_X1 U15788 ( .C1(n7204), .C2(n13907), .A(n13906), .B(n13905), .ZN(
        P1_U3240) );
  INV_X1 U15789 ( .A(n13908), .ZN(n13915) );
  INV_X1 U15790 ( .A(n13909), .ZN(n13911) );
  NAND2_X1 U15791 ( .A1(n13911), .A2(n13910), .ZN(n13913) );
  AOI22_X1 U15792 ( .A1(n13915), .A2(n13914), .B1(n13913), .B2(n13912), .ZN(
        n13921) );
  NOR2_X1 U15793 ( .A1(n14511), .A2(n13916), .ZN(n13919) );
  NAND2_X1 U15794 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14585)
         );
  OAI21_X1 U15795 ( .B1(n13917), .B2(n14481), .A(n14585), .ZN(n13918) );
  AOI211_X1 U15796 ( .C1(n14345), .C2(n14502), .A(n13919), .B(n13918), .ZN(
        n13920) );
  OAI21_X1 U15797 ( .B1(n13921), .B2(n14475), .A(n13920), .ZN(P1_U3241) );
  MUX2_X1 U15798 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14054), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15799 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13922), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15800 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13923), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15801 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13924), .S(n13948), .Z(
        P1_U3587) );
  MUX2_X1 U15802 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13925), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15803 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13926), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15804 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13927), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15805 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13928), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15806 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13929), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15807 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13930), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15808 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13931), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15809 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13932), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15810 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13933), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15811 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13934), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15812 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13935), .S(n13948), .Z(
        P1_U3575) );
  MUX2_X1 U15813 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13936), .S(n13948), .Z(
        P1_U3574) );
  MUX2_X1 U15814 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13937), .S(n13948), .Z(
        P1_U3573) );
  MUX2_X1 U15815 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13938), .S(n13948), .Z(
        P1_U3572) );
  MUX2_X1 U15816 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13939), .S(n13948), .Z(
        P1_U3571) );
  MUX2_X1 U15817 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13940), .S(n13948), .Z(
        P1_U3570) );
  MUX2_X1 U15818 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13941), .S(n13948), .Z(
        P1_U3569) );
  MUX2_X1 U15819 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13942), .S(n13948), .Z(
        P1_U3568) );
  MUX2_X1 U15820 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13943), .S(n13948), .Z(
        P1_U3567) );
  MUX2_X1 U15821 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13944), .S(n13948), .Z(
        P1_U3566) );
  MUX2_X1 U15822 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13945), .S(n13948), .Z(
        P1_U3565) );
  MUX2_X1 U15823 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13946), .S(n13948), .Z(
        P1_U3564) );
  MUX2_X1 U15824 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13947), .S(n13948), .Z(
        P1_U3563) );
  MUX2_X1 U15825 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13949), .S(n13948), .Z(
        P1_U3562) );
  MUX2_X1 U15826 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6678), .S(P1_U4016), .Z(
        P1_U3561) );
  INV_X1 U15827 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13951) );
  OAI22_X1 U15828 ( .A1(n14633), .A2(n7095), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13951), .ZN(n13952) );
  AOI21_X1 U15829 ( .B1(n13953), .B2(n14625), .A(n13952), .ZN(n13961) );
  OAI211_X1 U15830 ( .C1(n13956), .C2(n13955), .A(n14617), .B(n13954), .ZN(
        n13960) );
  OAI211_X1 U15831 ( .C1(n13958), .C2(n13963), .A(n14620), .B(n13957), .ZN(
        n13959) );
  NAND3_X1 U15832 ( .A1(n13961), .A2(n13960), .A3(n13959), .ZN(P1_U3244) );
  MUX2_X1 U15833 ( .A(n13963), .B(n13962), .S(n14378), .Z(n13965) );
  NAND2_X1 U15834 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  OAI211_X1 U15835 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13967), .A(n13966), .B(
        n13948), .ZN(n14011) );
  INV_X1 U15836 ( .A(n13968), .ZN(n13971) );
  INV_X1 U15837 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13969) );
  OAI22_X1 U15838 ( .A1(n14633), .A2(n7092), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13969), .ZN(n13970) );
  AOI21_X1 U15839 ( .B1(n13971), .B2(n14625), .A(n13970), .ZN(n13980) );
  OAI211_X1 U15840 ( .C1(n13974), .C2(n13973), .A(n14620), .B(n13972), .ZN(
        n13979) );
  OAI211_X1 U15841 ( .C1(n13977), .C2(n13976), .A(n14617), .B(n13975), .ZN(
        n13978) );
  NAND4_X1 U15842 ( .A1(n14011), .A2(n13980), .A3(n13979), .A4(n13978), .ZN(
        P1_U3245) );
  INV_X1 U15843 ( .A(n13981), .ZN(n13985) );
  NAND2_X1 U15844 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13982) );
  OAI21_X1 U15845 ( .B1(n14633), .B2(n13983), .A(n13982), .ZN(n13984) );
  AOI21_X1 U15846 ( .B1(n13985), .B2(n14625), .A(n13984), .ZN(n13994) );
  OAI211_X1 U15847 ( .C1(n13988), .C2(n13987), .A(n14620), .B(n13986), .ZN(
        n13993) );
  OAI211_X1 U15848 ( .C1(n13991), .C2(n13990), .A(n14617), .B(n13989), .ZN(
        n13992) );
  NAND3_X1 U15849 ( .A1(n13994), .A2(n13993), .A3(n13992), .ZN(P1_U3246) );
  INV_X1 U15850 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n13997) );
  INV_X1 U15851 ( .A(n13995), .ZN(n13996) );
  OAI21_X1 U15852 ( .B1(n14633), .B2(n13997), .A(n13996), .ZN(n13998) );
  AOI21_X1 U15853 ( .B1(n13999), .B2(n14625), .A(n13998), .ZN(n14010) );
  INV_X1 U15854 ( .A(n14000), .ZN(n14001) );
  OAI211_X1 U15855 ( .C1(n14003), .C2(n14002), .A(n14617), .B(n14001), .ZN(
        n14009) );
  INV_X1 U15856 ( .A(n14004), .ZN(n14005) );
  OAI211_X1 U15857 ( .C1(n14007), .C2(n14006), .A(n14620), .B(n14005), .ZN(
        n14008) );
  NAND4_X1 U15858 ( .A1(n14011), .A2(n14010), .A3(n14009), .A4(n14008), .ZN(
        P1_U3247) );
  MUX2_X1 U15859 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n11162), .S(n14557), .Z(
        n14012) );
  INV_X1 U15860 ( .A(n14012), .ZN(n14553) );
  OAI21_X1 U15861 ( .B1(n14025), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14013), 
        .ZN(n14554) );
  NAND2_X1 U15862 ( .A1(n14564), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n14014) );
  OAI21_X1 U15863 ( .B1(n14564), .B2(P1_REG2_REG_14__SCAN_IN), .A(n14014), 
        .ZN(n14568) );
  NOR2_X1 U15864 ( .A1(n14569), .A2(n14568), .ZN(n14567) );
  NAND2_X1 U15865 ( .A1(n14015), .A2(n14026), .ZN(n14016) );
  INV_X1 U15866 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U15867 ( .A1(n14578), .A2(n14577), .ZN(n14576) );
  AND2_X2 U15868 ( .A1(n14016), .A2(n14576), .ZN(n14590) );
  XNOR2_X1 U15869 ( .A(n14596), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U15870 ( .A1(n14590), .A2(n14589), .ZN(n14588) );
  NAND2_X1 U15871 ( .A1(n14030), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U15872 ( .A1(n14588), .A2(n14017), .ZN(n14603) );
  INV_X1 U15873 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U15874 ( .A1(n14033), .A2(n14250), .ZN(n14018) );
  OAI21_X1 U15875 ( .B1(n14033), .B2(n14250), .A(n14018), .ZN(n14602) );
  NAND2_X1 U15876 ( .A1(n14603), .A2(n14602), .ZN(n14601) );
  NAND2_X1 U15877 ( .A1(n14033), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U15878 ( .A1(n14601), .A2(n14019), .ZN(n14020) );
  AND2_X1 U15879 ( .A1(n14020), .A2(n14624), .ZN(n14022) );
  NOR2_X1 U15880 ( .A1(n14020), .A2(n14624), .ZN(n14021) );
  INV_X1 U15881 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15192) );
  NAND2_X1 U15882 ( .A1(n14043), .A2(n14620), .ZN(n14041) );
  INV_X1 U15883 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14023) );
  MUX2_X1 U15884 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14023), .S(n14564), .Z(
        n14563) );
  OAI21_X1 U15885 ( .B1(n14025), .B2(P1_REG1_REG_12__SCAN_IN), .A(n14024), 
        .ZN(n14551) );
  MUX2_X1 U15886 ( .A(n11288), .B(P1_REG1_REG_13__SCAN_IN), .S(n14557), .Z(
        n14550) );
  NOR2_X1 U15887 ( .A1(n14551), .A2(n14550), .ZN(n14549) );
  AOI21_X1 U15888 ( .B1(n14557), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14549), 
        .ZN(n14562) );
  NAND2_X1 U15889 ( .A1(n14563), .A2(n14562), .ZN(n14561) );
  OAI21_X1 U15890 ( .B1(n14564), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14561), 
        .ZN(n14027) );
  NAND2_X1 U15891 ( .A1(n14026), .A2(n14027), .ZN(n14028) );
  XNOR2_X1 U15892 ( .A(n14583), .B(n14027), .ZN(n14581) );
  INV_X1 U15893 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U15894 ( .A1(n14581), .A2(n14580), .ZN(n14579) );
  NAND2_X1 U15895 ( .A1(n14596), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14029) );
  OAI21_X1 U15896 ( .B1(n14596), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14029), 
        .ZN(n14592) );
  NAND2_X1 U15897 ( .A1(n14593), .A2(n14592), .ZN(n14591) );
  NAND2_X1 U15898 ( .A1(n14030), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U15899 ( .A1(n14591), .A2(n14031), .ZN(n14606) );
  XNOR2_X1 U15900 ( .A(n14033), .B(n14032), .ZN(n14605) );
  NAND2_X1 U15901 ( .A1(n14606), .A2(n14605), .ZN(n14604) );
  NAND2_X1 U15902 ( .A1(n14033), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U15903 ( .A1(n14604), .A2(n14034), .ZN(n14035) );
  AND2_X1 U15904 ( .A1(n14035), .A2(n14624), .ZN(n14037) );
  NOR2_X1 U15905 ( .A1(n14035), .A2(n14624), .ZN(n14036) );
  OR2_X1 U15906 ( .A1(n14037), .A2(n14036), .ZN(n14616) );
  INV_X1 U15907 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14615) );
  NOR2_X1 U15908 ( .A1(n14616), .A2(n14615), .ZN(n14629) );
  NOR2_X1 U15909 ( .A1(n14629), .A2(n14037), .ZN(n14039) );
  XNOR2_X1 U15910 ( .A(n14039), .B(n14038), .ZN(n14042) );
  AOI21_X1 U15911 ( .B1(n14042), .B2(n14617), .A(n14625), .ZN(n14040) );
  NAND2_X1 U15912 ( .A1(n14041), .A2(n14040), .ZN(n14046) );
  OAI22_X1 U15913 ( .A1(n14043), .A2(n14566), .B1(n14042), .B2(n14548), .ZN(
        n14045) );
  MUX2_X1 U15914 ( .A(n14046), .B(n14045), .S(n14044), .Z(n14050) );
  OAI21_X1 U15915 ( .B1(n14633), .B2(n14048), .A(n14047), .ZN(n14049) );
  NOR2_X1 U15916 ( .A1(n14050), .A2(n14049), .ZN(n14051) );
  INV_X1 U15917 ( .A(n14051), .ZN(P1_U3262) );
  NAND2_X1 U15918 ( .A1(n14261), .A2(n14060), .ZN(n14059) );
  XNOR2_X1 U15919 ( .A(n14059), .B(n14258), .ZN(n14052) );
  NAND2_X1 U15920 ( .A1(n14052), .A2(n14651), .ZN(n14257) );
  NOR2_X1 U15921 ( .A1(n14671), .A2(n14053), .ZN(n14056) );
  NAND2_X1 U15922 ( .A1(n14055), .A2(n14054), .ZN(n14259) );
  NOR2_X1 U15923 ( .A1(n14646), .A2(n14259), .ZN(n14062) );
  AOI211_X1 U15924 ( .C1(n14057), .C2(n14647), .A(n14056), .B(n14062), .ZN(
        n14058) );
  OAI21_X1 U15925 ( .B1(n14257), .B2(n14234), .A(n14058), .ZN(P1_U3263) );
  OAI211_X1 U15926 ( .C1(n14261), .C2(n14060), .A(n14651), .B(n14059), .ZN(
        n14260) );
  NOR2_X1 U15927 ( .A1(n14671), .A2(n14061), .ZN(n14063) );
  AOI211_X1 U15928 ( .C1(n14064), .C2(n14647), .A(n14063), .B(n14062), .ZN(
        n14065) );
  OAI21_X1 U15929 ( .B1(n14260), .B2(n14234), .A(n14065), .ZN(P1_U3264) );
  XNOR2_X1 U15930 ( .A(n14066), .B(n14070), .ZN(n14069) );
  INV_X1 U15931 ( .A(n14067), .ZN(n14068) );
  INV_X1 U15932 ( .A(n14275), .ZN(n14080) );
  AOI21_X1 U15933 ( .B1(n14270), .B2(n14090), .A(n14683), .ZN(n14073) );
  NAND2_X1 U15934 ( .A1(n14073), .A2(n14072), .ZN(n14272) );
  INV_X1 U15935 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14076) );
  INV_X1 U15936 ( .A(n14074), .ZN(n14075) );
  OAI22_X1 U15937 ( .A1(n14671), .A2(n14076), .B1(n14075), .B2(n14662), .ZN(
        n14077) );
  AOI21_X1 U15938 ( .B1(n14270), .B2(n14647), .A(n14077), .ZN(n14078) );
  OAI21_X1 U15939 ( .B1(n14272), .B2(n14234), .A(n14078), .ZN(n14079) );
  AOI21_X1 U15940 ( .B1(n14080), .B2(n14668), .A(n14079), .ZN(n14081) );
  OAI21_X1 U15941 ( .B1(n14274), .B2(n14646), .A(n14081), .ZN(P1_U3265) );
  INV_X1 U15942 ( .A(n14082), .ZN(n14084) );
  OAI21_X1 U15943 ( .B1(n14087), .B2(n14676), .A(n14086), .ZN(n14088) );
  INV_X1 U15944 ( .A(n14093), .ZN(n14091) );
  INV_X1 U15945 ( .A(n14089), .ZN(n14105) );
  OAI211_X1 U15946 ( .C1(n14091), .C2(n14105), .A(n14651), .B(n14090), .ZN(
        n14277) );
  AOI22_X1 U15947 ( .A1(n14646), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14092), 
        .B2(n14645), .ZN(n14095) );
  NAND2_X1 U15948 ( .A1(n14093), .A2(n14647), .ZN(n14094) );
  OAI211_X1 U15949 ( .C1(n14277), .C2(n14234), .A(n14095), .B(n14094), .ZN(
        n14096) );
  AOI21_X1 U15950 ( .B1(n14276), .B2(n14655), .A(n14096), .ZN(n14097) );
  OAI21_X1 U15951 ( .B1(n6552), .B2(n14646), .A(n14097), .ZN(P1_U3266) );
  XNOR2_X1 U15952 ( .A(n14098), .B(n14100), .ZN(n14286) );
  INV_X1 U15953 ( .A(n14099), .ZN(n14103) );
  XOR2_X1 U15954 ( .A(n14101), .B(n14100), .Z(n14102) );
  NAND2_X1 U15955 ( .A1(n14102), .A2(n14643), .ZN(n14285) );
  OAI211_X1 U15956 ( .C1(n14662), .C2(n14103), .A(n14285), .B(n14280), .ZN(
        n14104) );
  NAND2_X1 U15957 ( .A1(n14104), .A2(n14671), .ZN(n14109) );
  AOI211_X1 U15958 ( .C1(n14283), .C2(n14117), .A(n14683), .B(n14105), .ZN(
        n14281) );
  INV_X1 U15959 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14106) );
  OAI22_X1 U15960 ( .A1(n7204), .A2(n14175), .B1(n14106), .B2(n14671), .ZN(
        n14107) );
  AOI21_X1 U15961 ( .B1(n14281), .B2(n14654), .A(n14107), .ZN(n14108) );
  OAI211_X1 U15962 ( .C1(n14286), .C2(n14256), .A(n14109), .B(n14108), .ZN(
        P1_U3267) );
  OAI21_X1 U15963 ( .B1(n14111), .B2(n14113), .A(n14110), .ZN(n14293) );
  INV_X1 U15964 ( .A(n14112), .ZN(n14116) );
  INV_X1 U15965 ( .A(n14113), .ZN(n14115) );
  OAI21_X1 U15966 ( .B1(n14116), .B2(n14115), .A(n14114), .ZN(n14287) );
  AND2_X1 U15967 ( .A1(n14671), .A2(n14643), .ZN(n14667) );
  AOI21_X1 U15968 ( .B1(n14290), .B2(n14132), .A(n14683), .ZN(n14118) );
  AND2_X1 U15969 ( .A1(n14118), .A2(n14117), .ZN(n14288) );
  NAND2_X1 U15970 ( .A1(n14288), .A2(n14654), .ZN(n14124) );
  NAND2_X1 U15971 ( .A1(n14646), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U15972 ( .A1(n14289), .A2(n14671), .ZN(n14119) );
  OAI211_X1 U15973 ( .C1(n14662), .C2(n14121), .A(n14120), .B(n14119), .ZN(
        n14122) );
  AOI21_X1 U15974 ( .B1(n14290), .B2(n14647), .A(n14122), .ZN(n14123) );
  NAND2_X1 U15975 ( .A1(n14124), .A2(n14123), .ZN(n14125) );
  AOI21_X1 U15976 ( .B1(n14287), .B2(n14667), .A(n14125), .ZN(n14126) );
  OAI21_X1 U15977 ( .B1(n14256), .B2(n14293), .A(n14126), .ZN(P1_U3268) );
  AOI21_X1 U15978 ( .B1(n14128), .B2(n14127), .A(n14676), .ZN(n14131) );
  AOI21_X1 U15979 ( .B1(n14131), .B2(n14130), .A(n14129), .ZN(n14297) );
  INV_X1 U15980 ( .A(n14132), .ZN(n14133) );
  AOI211_X1 U15981 ( .C1(n14295), .C2(n14152), .A(n14683), .B(n14133), .ZN(
        n14294) );
  INV_X1 U15982 ( .A(n14134), .ZN(n14135) );
  AOI22_X1 U15983 ( .A1(n14646), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14135), 
        .B2(n14645), .ZN(n14136) );
  OAI21_X1 U15984 ( .B1(n7206), .B2(n14175), .A(n14136), .ZN(n14143) );
  NAND2_X1 U15985 ( .A1(n14138), .A2(n14137), .ZN(n14139) );
  AND2_X1 U15986 ( .A1(n14140), .A2(n14139), .ZN(n14298) );
  NOR2_X1 U15987 ( .A1(n14298), .A2(n14141), .ZN(n14142) );
  AOI211_X1 U15988 ( .C1(n14294), .C2(n14654), .A(n14143), .B(n14142), .ZN(
        n14144) );
  OAI21_X1 U15989 ( .B1(n14646), .B2(n14297), .A(n14144), .ZN(P1_U3269) );
  XNOR2_X1 U15990 ( .A(n14146), .B(n14145), .ZN(n14305) );
  INV_X1 U15991 ( .A(n14667), .ZN(n14208) );
  INV_X1 U15992 ( .A(n14147), .ZN(n14148) );
  AOI21_X1 U15993 ( .B1(n14150), .B2(n14149), .A(n14148), .ZN(n14303) );
  INV_X1 U15994 ( .A(n14151), .ZN(n14169) );
  OAI211_X1 U15995 ( .C1(n14169), .C2(n14301), .A(n14651), .B(n14152), .ZN(
        n14300) );
  AOI22_X1 U15996 ( .A1(n14646), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14153), 
        .B2(n14645), .ZN(n14154) );
  OAI21_X1 U15997 ( .B1(n14299), .B2(n14646), .A(n14154), .ZN(n14155) );
  AOI21_X1 U15998 ( .B1(n14156), .B2(n14647), .A(n14155), .ZN(n14157) );
  OAI21_X1 U15999 ( .B1(n14300), .B2(n14234), .A(n14157), .ZN(n14158) );
  AOI21_X1 U16000 ( .B1(n14303), .B2(n14668), .A(n14158), .ZN(n14159) );
  OAI21_X1 U16001 ( .B1(n14305), .B2(n14208), .A(n14159), .ZN(P1_U3270) );
  AND2_X1 U16002 ( .A1(n14179), .A2(n14160), .ZN(n14163) );
  OAI21_X1 U16003 ( .B1(n14163), .B2(n14162), .A(n14161), .ZN(n14165) );
  AOI21_X1 U16004 ( .B1(n14165), .B2(n14643), .A(n14164), .ZN(n14310) );
  OAI21_X1 U16005 ( .B1(n14168), .B2(n14167), .A(n14166), .ZN(n14306) );
  INV_X1 U16006 ( .A(n14187), .ZN(n14170) );
  AOI211_X1 U16007 ( .C1(n14308), .C2(n14170), .A(n14683), .B(n14169), .ZN(
        n14307) );
  NAND2_X1 U16008 ( .A1(n14307), .A2(n14654), .ZN(n14173) );
  AOI22_X1 U16009 ( .A1(n14646), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14171), 
        .B2(n14645), .ZN(n14172) );
  OAI211_X1 U16010 ( .C1(n14175), .C2(n14174), .A(n14173), .B(n14172), .ZN(
        n14176) );
  AOI21_X1 U16011 ( .B1(n14668), .B2(n14306), .A(n14176), .ZN(n14177) );
  OAI21_X1 U16012 ( .B1(n14310), .B2(n14646), .A(n14177), .ZN(P1_U3271) );
  XOR2_X1 U16013 ( .A(n14181), .B(n14178), .Z(n14316) );
  OAI211_X1 U16014 ( .C1(n14181), .C2(n14180), .A(n14179), .B(n14643), .ZN(
        n14184) );
  INV_X1 U16015 ( .A(n14182), .ZN(n14183) );
  NAND2_X1 U16016 ( .A1(n14184), .A2(n14183), .ZN(n14312) );
  NAND2_X1 U16017 ( .A1(n14199), .A2(n14314), .ZN(n14185) );
  NAND2_X1 U16018 ( .A1(n14185), .A2(n14651), .ZN(n14186) );
  NOR2_X1 U16019 ( .A1(n14187), .A2(n14186), .ZN(n14313) );
  NAND2_X1 U16020 ( .A1(n14313), .A2(n14654), .ZN(n14192) );
  OAI22_X1 U16021 ( .A1(n14189), .A2(n14662), .B1(n14188), .B2(n14671), .ZN(
        n14190) );
  AOI21_X1 U16022 ( .B1(n14314), .B2(n14647), .A(n14190), .ZN(n14191) );
  NAND2_X1 U16023 ( .A1(n14192), .A2(n14191), .ZN(n14193) );
  AOI21_X1 U16024 ( .B1(n14312), .B2(n14671), .A(n14193), .ZN(n14194) );
  OAI21_X1 U16025 ( .B1(n14316), .B2(n14256), .A(n14194), .ZN(P1_U3272) );
  OAI21_X1 U16026 ( .B1(n14196), .B2(n7130), .A(n14195), .ZN(n14325) );
  AOI22_X1 U16027 ( .A1(n14197), .A2(n14645), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n14646), .ZN(n14198) );
  OAI21_X1 U16028 ( .B1(n14317), .B2(n14646), .A(n14198), .ZN(n14202) );
  AOI21_X1 U16029 ( .B1(n14210), .B2(n14319), .A(n14683), .ZN(n14200) );
  NAND2_X1 U16030 ( .A1(n14200), .A2(n14199), .ZN(n14320) );
  NOR2_X1 U16031 ( .A1(n14320), .A2(n14234), .ZN(n14201) );
  AOI211_X1 U16032 ( .C1(n14647), .C2(n14319), .A(n14202), .B(n14201), .ZN(
        n14207) );
  OAI21_X1 U16033 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n14322) );
  OR2_X1 U16034 ( .A1(n14322), .A2(n14256), .ZN(n14206) );
  OAI211_X1 U16035 ( .C1(n14325), .C2(n14208), .A(n14207), .B(n14206), .ZN(
        P1_U3273) );
  XNOR2_X1 U16036 ( .A(n14209), .B(n11657), .ZN(n14330) );
  AOI21_X1 U16037 ( .B1(n14327), .B2(n14230), .A(n14683), .ZN(n14211) );
  AND2_X1 U16038 ( .A1(n14211), .A2(n14210), .ZN(n14326) );
  NAND2_X1 U16039 ( .A1(n14327), .A2(n14647), .ZN(n14213) );
  NAND2_X1 U16040 ( .A1(n14646), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14212) );
  OAI211_X1 U16041 ( .C1(n14662), .C2(n14214), .A(n14213), .B(n14212), .ZN(
        n14220) );
  OAI21_X1 U16042 ( .B1(n6616), .B2(n14216), .A(n14215), .ZN(n14218) );
  AOI21_X1 U16043 ( .B1(n14218), .B2(n14643), .A(n14217), .ZN(n14329) );
  NOR2_X1 U16044 ( .A1(n14329), .A2(n14646), .ZN(n14219) );
  AOI211_X1 U16045 ( .C1(n14326), .C2(n14654), .A(n14220), .B(n14219), .ZN(
        n14221) );
  OAI21_X1 U16046 ( .B1(n14330), .B2(n14256), .A(n14221), .ZN(P1_U3274) );
  OAI211_X1 U16047 ( .C1(n14223), .C2(n14224), .A(n14222), .B(n14643), .ZN(
        n14228) );
  XNOR2_X1 U16048 ( .A(n14225), .B(n14224), .ZN(n14331) );
  NAND2_X1 U16049 ( .A1(n14331), .A2(n14723), .ZN(n14226) );
  NAND3_X1 U16050 ( .A1(n14228), .A2(n14227), .A3(n14226), .ZN(n14336) );
  AOI21_X1 U16051 ( .B1(n14229), .B2(n14645), .A(n14336), .ZN(n14237) );
  AOI21_X1 U16052 ( .B1(n14232), .B2(n14248), .A(n14683), .ZN(n14231) );
  NAND2_X1 U16053 ( .A1(n14231), .A2(n14230), .ZN(n14332) );
  AOI22_X1 U16054 ( .A1(n14232), .A2(n14647), .B1(n14646), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n14233) );
  OAI21_X1 U16055 ( .B1(n14332), .B2(n14234), .A(n14233), .ZN(n14235) );
  AOI21_X1 U16056 ( .B1(n14331), .B2(n14655), .A(n14235), .ZN(n14236) );
  OAI21_X1 U16057 ( .B1(n14237), .B2(n14646), .A(n14236), .ZN(P1_U3275) );
  XNOR2_X1 U16058 ( .A(n14238), .B(n14241), .ZN(n14342) );
  OAI211_X1 U16059 ( .C1(n14241), .C2(n14240), .A(n14239), .B(n14643), .ZN(
        n14244) );
  INV_X1 U16060 ( .A(n14242), .ZN(n14243) );
  NAND2_X1 U16061 ( .A1(n14244), .A2(n14243), .ZN(n14338) );
  OR2_X1 U16062 ( .A1(n14246), .A2(n14245), .ZN(n14247) );
  AND3_X1 U16063 ( .A1(n14248), .A2(n14651), .A3(n14247), .ZN(n14339) );
  NAND2_X1 U16064 ( .A1(n14339), .A2(n14654), .ZN(n14253) );
  OAI22_X1 U16065 ( .A1(n14671), .A2(n14250), .B1(n14249), .B2(n14662), .ZN(
        n14251) );
  AOI21_X1 U16066 ( .B1(n14340), .B2(n14647), .A(n14251), .ZN(n14252) );
  NAND2_X1 U16067 ( .A1(n14253), .A2(n14252), .ZN(n14254) );
  AOI21_X1 U16068 ( .B1(n14338), .B2(n14671), .A(n14254), .ZN(n14255) );
  OAI21_X1 U16069 ( .B1(n14342), .B2(n14256), .A(n14255), .ZN(P1_U3276) );
  OAI211_X1 U16070 ( .C1(n14258), .C2(n14698), .A(n14257), .B(n14259), .ZN(
        n14348) );
  MUX2_X1 U16071 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14348), .S(n14753), .Z(
        P1_U3559) );
  OAI211_X1 U16072 ( .C1(n14261), .C2(n14698), .A(n14260), .B(n14259), .ZN(
        n14349) );
  MUX2_X1 U16073 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14349), .S(n14753), .Z(
        P1_U3558) );
  NAND2_X1 U16074 ( .A1(n14263), .A2(n14262), .ZN(n14265) );
  OAI211_X1 U16075 ( .C1(n14269), .C2(n14677), .A(n14268), .B(n14267), .ZN(
        n14350) );
  MUX2_X1 U16076 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14350), .S(n14753), .Z(
        P1_U3557) );
  NAND2_X1 U16077 ( .A1(n14270), .A2(n14691), .ZN(n14271) );
  AND2_X1 U16078 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  MUX2_X1 U16079 ( .A(n14351), .B(P1_REG1_REG_28__SCAN_IN), .S(n14751), .Z(
        P1_U3556) );
  INV_X1 U16080 ( .A(n14708), .ZN(n14722) );
  NAND2_X1 U16081 ( .A1(n14276), .A2(n14722), .ZN(n14278) );
  MUX2_X1 U16082 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14352), .S(n14753), .Z(
        P1_U3555) );
  INV_X1 U16083 ( .A(n14280), .ZN(n14282) );
  AOI211_X1 U16084 ( .C1(n14691), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14284) );
  OAI211_X1 U16085 ( .C1(n14677), .C2(n14286), .A(n14285), .B(n14284), .ZN(
        n14353) );
  MUX2_X1 U16086 ( .A(n14353), .B(P1_REG1_REG_26__SCAN_IN), .S(n14751), .Z(
        P1_U3554) );
  NAND2_X1 U16087 ( .A1(n14287), .A2(n14643), .ZN(n14292) );
  AOI211_X1 U16088 ( .C1(n14691), .C2(n14290), .A(n14289), .B(n14288), .ZN(
        n14291) );
  OAI211_X1 U16089 ( .C1(n14677), .C2(n14293), .A(n14292), .B(n14291), .ZN(
        n14354) );
  MUX2_X1 U16090 ( .A(n14354), .B(P1_REG1_REG_25__SCAN_IN), .S(n14751), .Z(
        P1_U3553) );
  AOI21_X1 U16091 ( .B1(n14691), .B2(n14295), .A(n14294), .ZN(n14296) );
  OAI211_X1 U16092 ( .C1(n14677), .C2(n14298), .A(n14297), .B(n14296), .ZN(
        n14355) );
  MUX2_X1 U16093 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14355), .S(n14753), .Z(
        P1_U3552) );
  INV_X1 U16094 ( .A(n14677), .ZN(n14733) );
  OAI211_X1 U16095 ( .C1(n14301), .C2(n14698), .A(n14300), .B(n14299), .ZN(
        n14302) );
  AOI21_X1 U16096 ( .B1(n14303), .B2(n14733), .A(n14302), .ZN(n14304) );
  OAI21_X1 U16097 ( .B1(n14676), .B2(n14305), .A(n14304), .ZN(n14356) );
  MUX2_X1 U16098 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14356), .S(n14753), .Z(
        P1_U3551) );
  INV_X1 U16099 ( .A(n14306), .ZN(n14311) );
  AOI21_X1 U16100 ( .B1(n14691), .B2(n14308), .A(n14307), .ZN(n14309) );
  OAI211_X1 U16101 ( .C1(n14677), .C2(n14311), .A(n14310), .B(n14309), .ZN(
        n14357) );
  MUX2_X1 U16102 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14357), .S(n14753), .Z(
        P1_U3550) );
  AOI211_X1 U16103 ( .C1(n14691), .C2(n14314), .A(n14313), .B(n14312), .ZN(
        n14315) );
  OAI21_X1 U16104 ( .B1(n14677), .B2(n14316), .A(n14315), .ZN(n14358) );
  MUX2_X1 U16105 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14358), .S(n14753), .Z(
        P1_U3549) );
  INV_X1 U16106 ( .A(n14317), .ZN(n14318) );
  AOI21_X1 U16107 ( .B1(n14319), .B2(n14691), .A(n14318), .ZN(n14321) );
  OAI211_X1 U16108 ( .C1(n14322), .C2(n14677), .A(n14321), .B(n14320), .ZN(
        n14323) );
  INV_X1 U16109 ( .A(n14323), .ZN(n14324) );
  OAI21_X1 U16110 ( .B1(n14325), .B2(n14676), .A(n14324), .ZN(n14359) );
  MUX2_X1 U16111 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14359), .S(n14753), .Z(
        P1_U3548) );
  AOI21_X1 U16112 ( .B1(n14691), .B2(n14327), .A(n14326), .ZN(n14328) );
  OAI211_X1 U16113 ( .C1(n14677), .C2(n14330), .A(n14329), .B(n14328), .ZN(
        n14360) );
  MUX2_X1 U16114 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14360), .S(n14753), .Z(
        P1_U3547) );
  NAND2_X1 U16115 ( .A1(n14331), .A2(n14722), .ZN(n14333) );
  OAI211_X1 U16116 ( .C1(n14334), .C2(n14698), .A(n14333), .B(n14332), .ZN(
        n14335) );
  NOR2_X1 U16117 ( .A1(n14336), .A2(n14335), .ZN(n14361) );
  MUX2_X1 U16118 ( .A(n14615), .B(n14361), .S(n14753), .Z(n14337) );
  INV_X1 U16119 ( .A(n14337), .ZN(P1_U3546) );
  AOI211_X1 U16120 ( .C1(n14691), .C2(n14340), .A(n14339), .B(n14338), .ZN(
        n14341) );
  OAI21_X1 U16121 ( .B1(n14677), .B2(n14342), .A(n14341), .ZN(n14364) );
  MUX2_X1 U16122 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14364), .S(n14753), .Z(
        P1_U3545) );
  AOI211_X1 U16123 ( .C1(n14691), .C2(n14345), .A(n14344), .B(n14343), .ZN(
        n14346) );
  OAI21_X1 U16124 ( .B1(n14677), .B2(n14347), .A(n14346), .ZN(n14365) );
  MUX2_X1 U16125 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14365), .S(n14753), .Z(
        P1_U3543) );
  MUX2_X1 U16126 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14348), .S(n14742), .Z(
        P1_U3527) );
  MUX2_X1 U16127 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14349), .S(n14742), .Z(
        P1_U3526) );
  MUX2_X1 U16128 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14350), .S(n14742), .Z(
        P1_U3525) );
  MUX2_X1 U16129 ( .A(n14351), .B(P1_REG0_REG_28__SCAN_IN), .S(n14740), .Z(
        P1_U3524) );
  MUX2_X1 U16130 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14352), .S(n14742), .Z(
        P1_U3523) );
  MUX2_X1 U16131 ( .A(n14353), .B(P1_REG0_REG_26__SCAN_IN), .S(n14740), .Z(
        P1_U3522) );
  MUX2_X1 U16132 ( .A(n14354), .B(P1_REG0_REG_25__SCAN_IN), .S(n14740), .Z(
        P1_U3521) );
  MUX2_X1 U16133 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14355), .S(n14742), .Z(
        P1_U3520) );
  MUX2_X1 U16134 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14356), .S(n14742), .Z(
        P1_U3519) );
  MUX2_X1 U16135 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14357), .S(n14742), .Z(
        P1_U3518) );
  MUX2_X1 U16136 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14358), .S(n14742), .Z(
        P1_U3517) );
  MUX2_X1 U16137 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14359), .S(n14742), .Z(
        P1_U3516) );
  MUX2_X1 U16138 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14360), .S(n14742), .Z(
        P1_U3515) );
  INV_X1 U16139 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14362) );
  MUX2_X1 U16140 ( .A(n14362), .B(n14361), .S(n14742), .Z(n14363) );
  INV_X1 U16141 ( .A(n14363), .ZN(P1_U3513) );
  MUX2_X1 U16142 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14364), .S(n14742), .Z(
        P1_U3510) );
  MUX2_X1 U16143 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14365), .S(n14742), .Z(
        P1_U3504) );
  NOR4_X1 U16144 ( .A1(n14367), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n6493), .ZN(n14368) );
  AOI21_X1 U16145 ( .B1(n14369), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14368), 
        .ZN(n14370) );
  OAI21_X1 U16146 ( .B1(n14371), .B2(n14382), .A(n14370), .ZN(P1_U3324) );
  OAI222_X1 U16147 ( .A1(n14373), .A2(P1_U3086), .B1(n14382), .B2(n14372), 
        .C1(n14379), .C2(n11622), .ZN(P1_U3326) );
  OAI222_X1 U16148 ( .A1(P1_U3086), .A2(n14376), .B1(n14382), .B2(n14375), 
        .C1(n14374), .C2(n14379), .ZN(P1_U3327) );
  OAI222_X1 U16149 ( .A1(n14378), .A2(P1_U3086), .B1(n14382), .B2(n14377), 
        .C1(n7036), .C2(n14379), .ZN(P1_U3328) );
  OAI222_X1 U16150 ( .A1(n14383), .A2(P1_U3086), .B1(n14382), .B2(n14381), 
        .C1(n14380), .C2(n14379), .ZN(P1_U3329) );
  MUX2_X1 U16151 ( .A(n14385), .B(n14384), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16152 ( .A(n14386), .ZN(n14387) );
  MUX2_X1 U16153 ( .A(n14387), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16154 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14388), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16155 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14389) );
  OAI21_X1 U16156 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14389), 
        .ZN(U28) );
  AOI21_X1 U16157 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14390) );
  OAI21_X1 U16158 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14390), 
        .ZN(U29) );
  AOI21_X1 U16159 ( .B1(n14393), .B2(n14392), .A(n14391), .ZN(n14395) );
  XNOR2_X1 U16160 ( .A(n14395), .B(n14394), .ZN(SUB_1596_U61) );
  INV_X1 U16161 ( .A(n14396), .ZN(n14397) );
  AOI22_X1 U16162 ( .A1(n14397), .A2(n14413), .B1(SI_9_), .B2(n14412), .ZN(
        n14398) );
  OAI21_X1 U16163 ( .B1(P3_U3151), .B2(n14399), .A(n14398), .ZN(P3_U3286) );
  INV_X1 U16164 ( .A(n14400), .ZN(n14401) );
  AOI22_X1 U16165 ( .A1(n14401), .A2(n14413), .B1(SI_11_), .B2(n14412), .ZN(
        n14402) );
  OAI21_X1 U16166 ( .B1(P3_U3151), .B2(n14900), .A(n14402), .ZN(P3_U3284) );
  OAI22_X1 U16167 ( .A1(n14404), .A2(n13057), .B1(n14403), .B2(n13054), .ZN(
        n14405) );
  INV_X1 U16168 ( .A(n14405), .ZN(n14406) );
  OAI21_X1 U16169 ( .B1(P3_U3151), .B2(n14917), .A(n14406), .ZN(P3_U3282) );
  XOR2_X1 U16170 ( .A(n14408), .B(n14407), .Z(SUB_1596_U57) );
  AOI22_X1 U16171 ( .A1(n14409), .A2(n14413), .B1(SI_15_), .B2(n14412), .ZN(
        n14410) );
  OAI21_X1 U16172 ( .B1(P3_U3151), .B2(n14411), .A(n14410), .ZN(P3_U3280) );
  AOI22_X1 U16173 ( .A1(n14414), .A2(n14413), .B1(SI_16_), .B2(n14412), .ZN(
        n14415) );
  OAI21_X1 U16174 ( .B1(P3_U3151), .B2(n14416), .A(n14415), .ZN(P3_U3279) );
  XNOR2_X1 U16175 ( .A(n14417), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16176 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14418), .Z(SUB_1596_U54) );
  OAI21_X1 U16177 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14422) );
  XNOR2_X1 U16178 ( .A(n14422), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  AOI21_X1 U16179 ( .B1(n14691), .B2(n14424), .A(n14423), .ZN(n14425) );
  OAI21_X1 U16180 ( .B1(n14426), .B2(n14677), .A(n14425), .ZN(n14427) );
  NOR2_X1 U16181 ( .A1(n14428), .A2(n14427), .ZN(n14430) );
  INV_X1 U16182 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14429) );
  AOI22_X1 U16183 ( .A1(n14742), .A2(n14430), .B1(n14429), .B2(n14740), .ZN(
        P1_U3495) );
  AOI22_X1 U16184 ( .A1(n14753), .A2(n14430), .B1(n10545), .B2(n14751), .ZN(
        P1_U3540) );
  AOI21_X1 U16185 ( .B1(n14433), .B2(n14432), .A(n14431), .ZN(n14435) );
  XNOR2_X1 U16186 ( .A(n14435), .B(n14434), .ZN(SUB_1596_U63) );
  INV_X1 U16187 ( .A(n14436), .ZN(n14437) );
  AOI21_X1 U16188 ( .B1(n12488), .B2(n15001), .A(n14437), .ZN(n14453) );
  AOI22_X1 U16189 ( .A1(n15025), .A2(n14453), .B1(n12482), .B2(n15023), .ZN(
        P3_U3490) );
  AOI21_X1 U16190 ( .B1(n14438), .B2(n15001), .A(n14437), .ZN(n14455) );
  AOI22_X1 U16191 ( .A1(n15025), .A2(n14455), .B1(n14439), .B2(n15023), .ZN(
        P3_U3489) );
  OAI22_X1 U16192 ( .A1(n14441), .A2(n14449), .B1(n14440), .B2(n15004), .ZN(
        n14442) );
  NOR2_X1 U16193 ( .A1(n14443), .A2(n14442), .ZN(n14457) );
  AOI22_X1 U16194 ( .A1(n15025), .A2(n14457), .B1(n8731), .B2(n15023), .ZN(
        P3_U3472) );
  OAI22_X1 U16195 ( .A1(n14445), .A2(n14449), .B1(n14444), .B2(n15004), .ZN(
        n14446) );
  NOR2_X1 U16196 ( .A1(n14447), .A2(n14446), .ZN(n14459) );
  AOI22_X1 U16197 ( .A1(n15025), .A2(n14459), .B1(n11175), .B2(n15023), .ZN(
        P3_U3471) );
  OAI22_X1 U16198 ( .A1(n14450), .A2(n14449), .B1(n14448), .B2(n15004), .ZN(
        n14451) );
  NOR2_X1 U16199 ( .A1(n14452), .A2(n14451), .ZN(n14461) );
  AOI22_X1 U16200 ( .A1(n15025), .A2(n14461), .B1(n8693), .B2(n15023), .ZN(
        P3_U3470) );
  INV_X1 U16201 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U16202 ( .A1(n15012), .A2(n14454), .B1(n14453), .B2(n15010), .ZN(
        P3_U3458) );
  INV_X1 U16203 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U16204 ( .A1(n15012), .A2(n14456), .B1(n14455), .B2(n15010), .ZN(
        P3_U3457) );
  INV_X1 U16205 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U16206 ( .A1(n15012), .A2(n14458), .B1(n14457), .B2(n15010), .ZN(
        P3_U3429) );
  INV_X1 U16207 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U16208 ( .A1(n15012), .A2(n14460), .B1(n14459), .B2(n15010), .ZN(
        P3_U3426) );
  INV_X1 U16209 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U16210 ( .A1(n15012), .A2(n14462), .B1(n14461), .B2(n15010), .ZN(
        P3_U3423) );
  AND2_X1 U16211 ( .A1(n14488), .A2(n14463), .ZN(n14466) );
  OAI21_X1 U16212 ( .B1(n14466), .B2(n14465), .A(n14464), .ZN(n14467) );
  AOI222_X1 U16213 ( .A1(n14468), .A2(n14506), .B1(n14467), .B2(n14504), .C1(
        n14518), .C2(n14502), .ZN(n14469) );
  NAND2_X1 U16214 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14573)
         );
  OAI211_X1 U16215 ( .C1(n14511), .C2(n14470), .A(n14469), .B(n14573), .ZN(
        P1_U3215) );
  AND2_X1 U16216 ( .A1(n14471), .A2(n14691), .ZN(n14735) );
  INV_X1 U16217 ( .A(n14472), .ZN(n14479) );
  INV_X1 U16218 ( .A(n14498), .ZN(n14474) );
  AOI211_X1 U16219 ( .C1(n14477), .C2(n14476), .A(n14475), .B(n14474), .ZN(
        n14478) );
  AOI211_X1 U16220 ( .C1(n14480), .C2(n14735), .A(n14479), .B(n14478), .ZN(
        n14486) );
  AOI21_X1 U16221 ( .B1(n14483), .B2(n14482), .A(n14481), .ZN(n14484) );
  INV_X1 U16222 ( .A(n14484), .ZN(n14485) );
  OAI211_X1 U16223 ( .C1(n14511), .C2(n14487), .A(n14486), .B(n14485), .ZN(
        P1_U3217) );
  OAI211_X1 U16224 ( .C1(n14490), .C2(n14489), .A(n14488), .B(n14504), .ZN(
        n14494) );
  AOI22_X1 U16225 ( .A1(n14492), .A2(n14502), .B1(n14506), .B2(n14491), .ZN(
        n14493) );
  AND2_X1 U16226 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  NAND2_X1 U16227 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14558)
         );
  OAI211_X1 U16228 ( .C1(n14511), .C2(n14496), .A(n14495), .B(n14558), .ZN(
        P1_U3234) );
  AND2_X1 U16229 ( .A1(n14498), .A2(n14497), .ZN(n14501) );
  OAI21_X1 U16230 ( .B1(n14501), .B2(n14500), .A(n14499), .ZN(n14505) );
  AOI222_X1 U16231 ( .A1(n14507), .A2(n14506), .B1(n14505), .B2(n14504), .C1(
        n14503), .C2(n14502), .ZN(n14509) );
  OAI211_X1 U16232 ( .C1(n14511), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        P1_U3236) );
  OAI21_X1 U16233 ( .B1(n14513), .B2(n14698), .A(n14512), .ZN(n14515) );
  AOI211_X1 U16234 ( .C1(n14733), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        n14526) );
  INV_X1 U16235 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U16236 ( .A1(n14753), .A2(n14526), .B1(n14517), .B2(n14751), .ZN(
        P1_U3544) );
  AND2_X1 U16237 ( .A1(n14518), .A2(n14691), .ZN(n14519) );
  NOR2_X1 U16238 ( .A1(n14520), .A2(n14519), .ZN(n14523) );
  OR2_X1 U16239 ( .A1(n14521), .A2(n14677), .ZN(n14522) );
  AOI22_X1 U16240 ( .A1(n14753), .A2(n14527), .B1(n14023), .B2(n14751), .ZN(
        P1_U3542) );
  INV_X1 U16241 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U16242 ( .A1(n14742), .A2(n14526), .B1(n14525), .B2(n14740), .ZN(
        P1_U3507) );
  AOI22_X1 U16243 ( .A1(n14742), .A2(n14527), .B1(n11153), .B2(n14740), .ZN(
        P1_U3501) );
  AOI21_X1 U16244 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n14532) );
  XNOR2_X1 U16245 ( .A(n14532), .B(n14531), .ZN(SUB_1596_U69) );
  XNOR2_X1 U16246 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14533), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16247 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14537) );
  XNOR2_X1 U16248 ( .A(n14537), .B(n14775), .ZN(SUB_1596_U67) );
  AOI21_X1 U16249 ( .B1(n14540), .B2(n14539), .A(n14538), .ZN(n14541) );
  XNOR2_X1 U16250 ( .A(n14541), .B(n15193), .ZN(SUB_1596_U66) );
  NOR2_X1 U16251 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  XOR2_X1 U16252 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14544), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16253 ( .A1(n14546), .A2(n14545), .ZN(n14547) );
  XOR2_X1 U16254 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14547), .Z(SUB_1596_U64)
         );
  AOI211_X1 U16255 ( .C1(n14551), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        n14556) );
  AOI211_X1 U16256 ( .C1(n14554), .C2(n14553), .A(n14552), .B(n14566), .ZN(
        n14555) );
  AOI211_X1 U16257 ( .C1(n14625), .C2(n14557), .A(n14556), .B(n14555), .ZN(
        n14559) );
  OAI211_X1 U16258 ( .C1(n14560), .C2(n14633), .A(n14559), .B(n14558), .ZN(
        P1_U3256) );
  OAI21_X1 U16259 ( .B1(n14563), .B2(n14562), .A(n14561), .ZN(n14572) );
  INV_X1 U16260 ( .A(n14564), .ZN(n14565) );
  NOR2_X1 U16261 ( .A1(n14610), .A2(n14565), .ZN(n14571) );
  AOI211_X1 U16262 ( .C1(n14569), .C2(n14568), .A(n14567), .B(n14566), .ZN(
        n14570) );
  AOI211_X1 U16263 ( .C1(n14617), .C2(n14572), .A(n14571), .B(n14570), .ZN(
        n14574) );
  OAI211_X1 U16264 ( .C1(n14575), .C2(n14633), .A(n14574), .B(n14573), .ZN(
        P1_U3257) );
  OAI21_X1 U16265 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14584) );
  OAI21_X1 U16266 ( .B1(n14581), .B2(n14580), .A(n14579), .ZN(n14582) );
  AOI222_X1 U16267 ( .A1(n14584), .A2(n14620), .B1(n14583), .B2(n14625), .C1(
        n14582), .C2(n14617), .ZN(n14586) );
  OAI211_X1 U16268 ( .C1(n14587), .C2(n14633), .A(n14586), .B(n14585), .ZN(
        P1_U3258) );
  OAI211_X1 U16269 ( .C1(n14590), .C2(n14589), .A(n14588), .B(n14620), .ZN(
        n14595) );
  OAI211_X1 U16270 ( .C1(n14593), .C2(n14592), .A(n14591), .B(n14617), .ZN(
        n14594) );
  OAI211_X1 U16271 ( .C1(n14610), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        n14597) );
  INV_X1 U16272 ( .A(n14597), .ZN(n14599) );
  OAI211_X1 U16273 ( .C1(n14600), .C2(n14633), .A(n14599), .B(n14598), .ZN(
        P1_U3259) );
  INV_X1 U16274 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14614) );
  OAI211_X1 U16275 ( .C1(n14603), .C2(n14602), .A(n14601), .B(n14620), .ZN(
        n14608) );
  OAI211_X1 U16276 ( .C1(n14606), .C2(n14605), .A(n14604), .B(n14617), .ZN(
        n14607) );
  OAI211_X1 U16277 ( .C1(n14610), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        n14611) );
  INV_X1 U16278 ( .A(n14611), .ZN(n14613) );
  OAI211_X1 U16279 ( .C1(n14614), .C2(n14633), .A(n14613), .B(n14612), .ZN(
        P1_U3260) );
  NAND2_X1 U16280 ( .A1(n14616), .A2(n14615), .ZN(n14618) );
  NAND2_X1 U16281 ( .A1(n14618), .A2(n14617), .ZN(n14628) );
  NAND2_X1 U16282 ( .A1(n14619), .A2(n15192), .ZN(n14621) );
  NAND2_X1 U16283 ( .A1(n14621), .A2(n14620), .ZN(n14622) );
  OR2_X1 U16284 ( .A1(n14623), .A2(n14622), .ZN(n14627) );
  NAND2_X1 U16285 ( .A1(n14625), .A2(n14624), .ZN(n14626) );
  OAI211_X1 U16286 ( .C1(n14629), .C2(n14628), .A(n14627), .B(n14626), .ZN(
        n14630) );
  INV_X1 U16287 ( .A(n14630), .ZN(n14632) );
  OAI211_X1 U16288 ( .C1(n14634), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        P1_U3261) );
  OAI21_X1 U16289 ( .B1(n14636), .B2(n14638), .A(n14635), .ZN(n14642) );
  INV_X1 U16290 ( .A(n14637), .ZN(n14641) );
  XNOR2_X1 U16291 ( .A(n14639), .B(n14638), .ZN(n14649) );
  NOR2_X1 U16292 ( .A1(n14649), .A2(n14707), .ZN(n14640) );
  AOI211_X1 U16293 ( .C1(n14643), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        n14700) );
  AOI222_X1 U16294 ( .A1(n14648), .A2(n14647), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14646), .C1(n14645), .C2(n14644), .ZN(n14657) );
  INV_X1 U16295 ( .A(n14649), .ZN(n14703) );
  OAI211_X1 U16296 ( .C1(n14652), .C2(n14699), .A(n14651), .B(n14650), .ZN(
        n14697) );
  INV_X1 U16297 ( .A(n14697), .ZN(n14653) );
  AOI22_X1 U16298 ( .A1(n14703), .A2(n14655), .B1(n14654), .B2(n14653), .ZN(
        n14656) );
  OAI211_X1 U16299 ( .C1(n14646), .C2(n14700), .A(n14657), .B(n14656), .ZN(
        P1_U3287) );
  INV_X1 U16300 ( .A(n14658), .ZN(n14659) );
  NOR2_X1 U16301 ( .A1(n14660), .A2(n14659), .ZN(n14678) );
  INV_X1 U16302 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14661) );
  NOR2_X1 U16303 ( .A1(n14662), .A2(n14661), .ZN(n14664) );
  INV_X1 U16304 ( .A(n14663), .ZN(n14679) );
  AOI211_X1 U16305 ( .C1(n14678), .C2(n14665), .A(n14664), .B(n14679), .ZN(
        n14672) );
  OAI21_X1 U16306 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n14669) );
  OAI221_X1 U16307 ( .B1(n14646), .B2(n14672), .C1(n14671), .C2(n14670), .A(
        n14669), .ZN(P1_U3293) );
  AND2_X1 U16308 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14674), .ZN(P1_U3294) );
  AND2_X1 U16309 ( .A1(n14674), .A2(P1_D_REG_30__SCAN_IN), .ZN(P1_U3295) );
  AND2_X1 U16310 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14674), .ZN(P1_U3296) );
  AND2_X1 U16311 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14674), .ZN(P1_U3297) );
  AND2_X1 U16312 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14674), .ZN(P1_U3298) );
  AND2_X1 U16313 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14674), .ZN(P1_U3299) );
  AND2_X1 U16314 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14674), .ZN(P1_U3300) );
  INV_X1 U16315 ( .A(n14674), .ZN(n14673) );
  INV_X1 U16316 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15205) );
  NOR2_X1 U16317 ( .A1(n14673), .A2(n15205), .ZN(P1_U3301) );
  AND2_X1 U16318 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14674), .ZN(P1_U3302) );
  AND2_X1 U16319 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14674), .ZN(P1_U3303) );
  AND2_X1 U16320 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14674), .ZN(P1_U3304) );
  AND2_X1 U16321 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14674), .ZN(P1_U3305) );
  AND2_X1 U16322 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14674), .ZN(P1_U3306) );
  AND2_X1 U16323 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14674), .ZN(P1_U3307) );
  AND2_X1 U16324 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14674), .ZN(P1_U3308) );
  AND2_X1 U16325 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14674), .ZN(P1_U3309) );
  AND2_X1 U16326 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14674), .ZN(P1_U3310) );
  AND2_X1 U16327 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14674), .ZN(P1_U3311) );
  AND2_X1 U16328 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14674), .ZN(P1_U3312) );
  AND2_X1 U16329 ( .A1(n14674), .A2(P1_D_REG_12__SCAN_IN), .ZN(P1_U3313) );
  AND2_X1 U16330 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14674), .ZN(P1_U3314) );
  AND2_X1 U16331 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14674), .ZN(P1_U3315) );
  AND2_X1 U16332 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14674), .ZN(P1_U3316) );
  INV_X1 U16333 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15054) );
  NOR2_X1 U16334 ( .A1(n14673), .A2(n15054), .ZN(P1_U3317) );
  AND2_X1 U16335 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14674), .ZN(P1_U3318) );
  AND2_X1 U16336 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14674), .ZN(P1_U3319) );
  AND2_X1 U16337 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14674), .ZN(P1_U3320) );
  AND2_X1 U16338 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14674), .ZN(P1_U3321) );
  AND2_X1 U16339 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14674), .ZN(P1_U3322) );
  AND2_X1 U16340 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14674), .ZN(P1_U3323) );
  AOI21_X1 U16341 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14680) );
  NOR3_X1 U16342 ( .A1(n14680), .A2(n14679), .A3(n14678), .ZN(n14743) );
  INV_X1 U16343 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16344 ( .A1(n14742), .A2(n14743), .B1(n14681), .B2(n14740), .ZN(
        P1_U3459) );
  OAI21_X1 U16345 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n14686) );
  AOI211_X1 U16346 ( .C1(n14722), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14745) );
  INV_X1 U16347 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U16348 ( .A1(n14742), .A2(n14745), .B1(n14688), .B2(n14740), .ZN(
        P1_U3462) );
  AOI21_X1 U16349 ( .B1(n14691), .B2(n14690), .A(n14689), .ZN(n14692) );
  OAI211_X1 U16350 ( .C1(n14694), .C2(n14708), .A(n14693), .B(n14692), .ZN(
        n14695) );
  INV_X1 U16351 ( .A(n14695), .ZN(n14746) );
  INV_X1 U16352 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16353 ( .A1(n14742), .A2(n14746), .B1(n14696), .B2(n14740), .ZN(
        P1_U3474) );
  OAI21_X1 U16354 ( .B1(n14699), .B2(n14698), .A(n14697), .ZN(n14702) );
  INV_X1 U16355 ( .A(n14700), .ZN(n14701) );
  AOI211_X1 U16356 ( .C1(n14722), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14747) );
  INV_X1 U16357 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14704) );
  AOI22_X1 U16358 ( .A1(n14742), .A2(n14747), .B1(n14704), .B2(n14740), .ZN(
        P1_U3477) );
  INV_X1 U16359 ( .A(n14705), .ZN(n14713) );
  AOI21_X1 U16360 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14712) );
  INV_X1 U16361 ( .A(n14709), .ZN(n14711) );
  NOR4_X1 U16362 ( .A1(n14713), .A2(n14712), .A3(n14711), .A4(n14710), .ZN(
        n14748) );
  INV_X1 U16363 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14714) );
  AOI22_X1 U16364 ( .A1(n14742), .A2(n14748), .B1(n14714), .B2(n14740), .ZN(
        P1_U3480) );
  AND2_X1 U16365 ( .A1(n14715), .A2(n14733), .ZN(n14720) );
  INV_X1 U16366 ( .A(n14716), .ZN(n14718) );
  NOR4_X1 U16367 ( .A1(n14720), .A2(n14719), .A3(n14718), .A4(n14717), .ZN(
        n14749) );
  INV_X1 U16368 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14721) );
  AOI22_X1 U16369 ( .A1(n14742), .A2(n14749), .B1(n14721), .B2(n14740), .ZN(
        P1_U3483) );
  AND2_X1 U16370 ( .A1(n14724), .A2(n14722), .ZN(n14730) );
  AND2_X1 U16371 ( .A1(n14724), .A2(n14723), .ZN(n14729) );
  INV_X1 U16372 ( .A(n14725), .ZN(n14726) );
  NAND2_X1 U16373 ( .A1(n14727), .A2(n14726), .ZN(n14728) );
  NOR4_X1 U16374 ( .A1(n14731), .A2(n14730), .A3(n14729), .A4(n14728), .ZN(
        n14750) );
  INV_X1 U16375 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16376 ( .A1(n14742), .A2(n14750), .B1(n14732), .B2(n14740), .ZN(
        P1_U3486) );
  AND2_X1 U16377 ( .A1(n14734), .A2(n14733), .ZN(n14738) );
  OR2_X1 U16378 ( .A1(n14736), .A2(n14735), .ZN(n14737) );
  NOR3_X1 U16379 ( .A1(n14739), .A2(n14738), .A3(n14737), .ZN(n14752) );
  INV_X1 U16380 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14741) );
  AOI22_X1 U16381 ( .A1(n14742), .A2(n14752), .B1(n14741), .B2(n14740), .ZN(
        P1_U3489) );
  AOI22_X1 U16382 ( .A1(n14753), .A2(n14743), .B1(n9263), .B2(n14751), .ZN(
        P1_U3528) );
  AOI22_X1 U16383 ( .A1(n14753), .A2(n14745), .B1(n14744), .B2(n14751), .ZN(
        P1_U3529) );
  AOI22_X1 U16384 ( .A1(n14753), .A2(n14746), .B1(n9916), .B2(n14751), .ZN(
        P1_U3533) );
  AOI22_X1 U16385 ( .A1(n14753), .A2(n14747), .B1(n9229), .B2(n14751), .ZN(
        P1_U3534) );
  AOI22_X1 U16386 ( .A1(n14753), .A2(n14748), .B1(n9230), .B2(n14751), .ZN(
        P1_U3535) );
  AOI22_X1 U16387 ( .A1(n14753), .A2(n14749), .B1(n9319), .B2(n14751), .ZN(
        P1_U3536) );
  AOI22_X1 U16388 ( .A1(n14753), .A2(n14750), .B1(n9597), .B2(n14751), .ZN(
        P1_U3537) );
  AOI22_X1 U16389 ( .A1(n14753), .A2(n14752), .B1(n9932), .B2(n14751), .ZN(
        P1_U3538) );
  NOR2_X1 U16390 ( .A1(n15233), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI21_X1 U16391 ( .B1(n15223), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14754), .ZN(
        n14758) );
  AOI22_X1 U16392 ( .A1(n15233), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14757) );
  OAI22_X1 U16393 ( .A1(n15230), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14780), .ZN(n14755) );
  OAI21_X1 U16394 ( .B1(n15226), .B2(n14755), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14756) );
  OAI211_X1 U16395 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14758), .A(n14757), .B(
        n14756), .ZN(P2_U3214) );
  INV_X1 U16396 ( .A(n14759), .ZN(n14760) );
  OAI21_X1 U16397 ( .B1(n14824), .B2(n14761), .A(n14760), .ZN(n14762) );
  AOI21_X1 U16398 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15233), .A(n14762), .ZN(
        n14773) );
  AOI211_X1 U16399 ( .C1(n14765), .C2(n14764), .A(n14763), .B(n14780), .ZN(
        n14766) );
  INV_X1 U16400 ( .A(n14766), .ZN(n14772) );
  AOI211_X1 U16401 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n15230), .ZN(
        n14770) );
  INV_X1 U16402 ( .A(n14770), .ZN(n14771) );
  NAND3_X1 U16403 ( .A1(n14773), .A2(n14772), .A3(n14771), .ZN(P2_U3217) );
  NOR2_X1 U16404 ( .A1(n14775), .A2(n14774), .ZN(n14776) );
  AOI211_X1 U16405 ( .C1(n14778), .C2(n15226), .A(n14777), .B(n14776), .ZN(
        n14789) );
  AOI211_X1 U16406 ( .C1(n14782), .C2(n14781), .A(n14780), .B(n14779), .ZN(
        n14783) );
  INV_X1 U16407 ( .A(n14783), .ZN(n14788) );
  OAI211_X1 U16408 ( .C1(n14786), .C2(n14785), .A(n14784), .B(n14833), .ZN(
        n14787) );
  NAND3_X1 U16409 ( .A1(n14789), .A2(n14788), .A3(n14787), .ZN(P2_U3227) );
  AOI22_X1 U16410 ( .A1(n15233), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14799) );
  NAND2_X1 U16411 ( .A1(n15226), .A2(n14790), .ZN(n14798) );
  OAI211_X1 U16412 ( .C1(n14792), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14791), 
        .B(n14833), .ZN(n14797) );
  XOR2_X1 U16413 ( .A(n14794), .B(n14793), .Z(n14795) );
  NAND2_X1 U16414 ( .A1(n14795), .A2(n15223), .ZN(n14796) );
  NAND4_X1 U16415 ( .A1(n14799), .A2(n14798), .A3(n14797), .A4(n14796), .ZN(
        P2_U3228) );
  AOI22_X1 U16416 ( .A1(n15233), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14808) );
  NAND2_X1 U16417 ( .A1(n15226), .A2(n14800), .ZN(n14807) );
  OAI211_X1 U16418 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14802), .A(n14833), 
        .B(n14801), .ZN(n14806) );
  OAI211_X1 U16419 ( .C1(n14804), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15223), 
        .B(n14803), .ZN(n14805) );
  NAND4_X1 U16420 ( .A1(n14808), .A2(n14807), .A3(n14806), .A4(n14805), .ZN(
        P2_U3229) );
  INV_X1 U16421 ( .A(n14809), .ZN(n14811) );
  OAI21_X1 U16422 ( .B1(n14811), .B2(n14810), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14812) );
  OAI21_X1 U16423 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14812), .ZN(n14822) );
  XOR2_X1 U16424 ( .A(n14814), .B(n14813), .Z(n14815) );
  NAND2_X1 U16425 ( .A1(n14815), .A2(n14833), .ZN(n14821) );
  NAND2_X1 U16426 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n15233), .ZN(n14820) );
  XNOR2_X1 U16427 ( .A(n14817), .B(n14816), .ZN(n14818) );
  NAND2_X1 U16428 ( .A1(n14818), .A2(n15223), .ZN(n14819) );
  NAND4_X1 U16429 ( .A1(n14822), .A2(n14821), .A3(n14820), .A4(n14819), .ZN(
        P2_U3230) );
  NOR2_X1 U16430 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  AOI211_X1 U16431 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n15233), .A(n14826), 
        .B(n14825), .ZN(n14837) );
  OAI211_X1 U16432 ( .C1(n14829), .C2(n14828), .A(n14827), .B(n15223), .ZN(
        n14836) );
  NAND2_X1 U16433 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  NAND3_X1 U16434 ( .A1(n14834), .A2(n14833), .A3(n14832), .ZN(n14835) );
  NAND3_X1 U16435 ( .A1(n14837), .A2(n14836), .A3(n14835), .ZN(P2_U3231) );
  NOR2_X1 U16436 ( .A1(n14845), .A2(n14838), .ZN(n14839) );
  AND2_X1 U16437 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14840), .ZN(P2_U3266) );
  AND2_X1 U16438 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14840), .ZN(P2_U3267) );
  AND2_X1 U16439 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14840), .ZN(P2_U3268) );
  AND2_X1 U16440 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14840), .ZN(P2_U3269) );
  AND2_X1 U16441 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14840), .ZN(P2_U3270) );
  AND2_X1 U16442 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14840), .ZN(P2_U3271) );
  AND2_X1 U16443 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14840), .ZN(P2_U3272) );
  INV_X1 U16444 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15171) );
  NOR2_X1 U16445 ( .A1(n14839), .A2(n15171), .ZN(P2_U3273) );
  AND2_X1 U16446 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14840), .ZN(P2_U3274) );
  AND2_X1 U16447 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14840), .ZN(P2_U3275) );
  AND2_X1 U16448 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14840), .ZN(P2_U3276) );
  AND2_X1 U16449 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14840), .ZN(P2_U3277) );
  AND2_X1 U16450 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14840), .ZN(P2_U3278) );
  AND2_X1 U16451 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14840), .ZN(P2_U3279) );
  AND2_X1 U16452 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14840), .ZN(P2_U3280) );
  AND2_X1 U16453 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14840), .ZN(P2_U3281) );
  AND2_X1 U16454 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14840), .ZN(P2_U3282) );
  AND2_X1 U16455 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14840), .ZN(P2_U3283) );
  AND2_X1 U16456 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14840), .ZN(P2_U3284) );
  AND2_X1 U16457 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14840), .ZN(P2_U3285) );
  AND2_X1 U16458 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14840), .ZN(P2_U3286) );
  AND2_X1 U16459 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14840), .ZN(P2_U3287) );
  AND2_X1 U16460 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14840), .ZN(P2_U3288) );
  AND2_X1 U16461 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14840), .ZN(P2_U3289) );
  AND2_X1 U16462 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14840), .ZN(P2_U3290) );
  AND2_X1 U16463 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14840), .ZN(P2_U3291) );
  AND2_X1 U16464 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14840), .ZN(P2_U3292) );
  AND2_X1 U16465 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14840), .ZN(P2_U3293) );
  AND2_X1 U16466 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14840), .ZN(P2_U3294) );
  AND2_X1 U16467 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14840), .ZN(P2_U3295) );
  AOI22_X1 U16468 ( .A1(n14843), .A2(n14842), .B1(n14841), .B2(n14845), .ZN(
        P2_U3416) );
  AOI21_X1 U16469 ( .B1(n14846), .B2(n14845), .A(n14844), .ZN(P2_U3417) );
  OAI22_X1 U16470 ( .A1(n14850), .A2(n14849), .B1(n14848), .B2(n14847), .ZN(
        n14853) );
  INV_X1 U16471 ( .A(n14851), .ZN(n14852) );
  AOI211_X1 U16472 ( .C1(n14855), .C2(n14854), .A(n14853), .B(n14852), .ZN(
        n14888) );
  INV_X1 U16473 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U16474 ( .A1(n14886), .A2(n14888), .B1(n14856), .B2(n14884), .ZN(
        P2_U3430) );
  INV_X1 U16475 ( .A(n14857), .ZN(n14858) );
  OAI21_X1 U16476 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n14863) );
  INV_X1 U16477 ( .A(n14861), .ZN(n14862) );
  AOI211_X1 U16478 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14890) );
  INV_X1 U16479 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U16480 ( .A1(n14886), .A2(n14890), .B1(n14866), .B2(n14884), .ZN(
        P2_U3439) );
  AOI21_X1 U16481 ( .B1(n14877), .B2(n14868), .A(n14867), .ZN(n14869) );
  OAI211_X1 U16482 ( .C1(n14872), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        n14873) );
  INV_X1 U16483 ( .A(n14873), .ZN(n14892) );
  INV_X1 U16484 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U16485 ( .A1(n14886), .A2(n14892), .B1(n14874), .B2(n14884), .ZN(
        P2_U3445) );
  OR2_X1 U16486 ( .A1(n14876), .A2(n14875), .ZN(n14883) );
  AND2_X1 U16487 ( .A1(n14878), .A2(n14877), .ZN(n14879) );
  NOR2_X1 U16488 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  AND3_X1 U16489 ( .A1(n14883), .A2(n14882), .A3(n14881), .ZN(n14894) );
  INV_X1 U16490 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14885) );
  AOI22_X1 U16491 ( .A1(n14886), .A2(n14894), .B1(n14885), .B2(n14884), .ZN(
        P2_U3451) );
  AOI22_X1 U16492 ( .A1(n14895), .A2(n14888), .B1(n14887), .B2(n14893), .ZN(
        P2_U3499) );
  AOI22_X1 U16493 ( .A1(n14895), .A2(n14890), .B1(n14889), .B2(n14893), .ZN(
        P2_U3502) );
  AOI22_X1 U16494 ( .A1(n14895), .A2(n14892), .B1(n14891), .B2(n14893), .ZN(
        P2_U3504) );
  AOI22_X1 U16495 ( .A1(n14895), .A2(n14894), .B1(n9341), .B2(n14893), .ZN(
        P2_U3506) );
  NOR2_X1 U16496 ( .A1(P3_U3897), .A2(n14896), .ZN(P3_U3150) );
  AOI21_X1 U16497 ( .B1(n8692), .B2(n14898), .A(n14897), .ZN(n14912) );
  INV_X1 U16498 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14899) );
  OAI22_X1 U16499 ( .A1(n14918), .A2(n14900), .B1(n14916), .B2(n14899), .ZN(
        n14909) );
  AOI21_X1 U16500 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14907) );
  AOI21_X1 U16501 ( .B1(n8693), .B2(n14905), .A(n14904), .ZN(n14906) );
  OAI22_X1 U16502 ( .A1(n14907), .A2(n14928), .B1(n14906), .B2(n14926), .ZN(
        n14908) );
  NOR3_X1 U16503 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n14911) );
  OAI21_X1 U16504 ( .B1(n14912), .B2(n14934), .A(n14911), .ZN(P3_U3193) );
  AOI21_X1 U16505 ( .B1(n11383), .B2(n14914), .A(n14913), .ZN(n14935) );
  OAI22_X1 U16506 ( .A1(n14918), .A2(n14917), .B1(n14916), .B2(n14915), .ZN(
        n14931) );
  OR2_X1 U16507 ( .A1(n14920), .A2(n14919), .ZN(n14922) );
  AOI21_X1 U16508 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14929) );
  AOI21_X1 U16509 ( .B1(n8731), .B2(n14925), .A(n14924), .ZN(n14927) );
  OAI22_X1 U16510 ( .A1(n14929), .A2(n14928), .B1(n14927), .B2(n14926), .ZN(
        n14930) );
  NOR3_X1 U16511 ( .A1(n14932), .A2(n14931), .A3(n14930), .ZN(n14933) );
  OAI21_X1 U16512 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(P3_U3195) );
  XNOR2_X1 U16513 ( .A(n14936), .B(n14942), .ZN(n14950) );
  INV_X1 U16514 ( .A(n14950), .ZN(n14963) );
  NOR2_X1 U16515 ( .A1(n14937), .A2(n15004), .ZN(n14962) );
  NAND2_X1 U16516 ( .A1(n14962), .A2(n14938), .ZN(n14939) );
  OAI21_X1 U16517 ( .B1(n8563), .B2(n14940), .A(n14939), .ZN(n14951) );
  XNOR2_X1 U16518 ( .A(n14941), .B(n14942), .ZN(n14948) );
  OAI22_X1 U16519 ( .A1(n14945), .A2(n14944), .B1(n8559), .B2(n14943), .ZN(
        n14946) );
  AOI21_X1 U16520 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n14949) );
  OAI21_X1 U16521 ( .B1(n14997), .B2(n14950), .A(n14949), .ZN(n14961) );
  AOI211_X1 U16522 ( .C1(n14952), .C2(n14963), .A(n14951), .B(n14961), .ZN(
        n14954) );
  AOI22_X1 U16523 ( .A1(n14955), .A2(n9652), .B1(n14954), .B2(n14953), .ZN(
        P3_U3231) );
  INV_X1 U16524 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14960) );
  AOI211_X1 U16525 ( .C1(n14959), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n15013) );
  AOI22_X1 U16526 ( .A1(n15012), .A2(n14960), .B1(n15013), .B2(n15010), .ZN(
        P3_U3393) );
  INV_X1 U16527 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14964) );
  AOI211_X1 U16528 ( .C1(n14963), .C2(n15009), .A(n14962), .B(n14961), .ZN(
        n15014) );
  AOI22_X1 U16529 ( .A1(n15012), .A2(n14964), .B1(n15014), .B2(n15010), .ZN(
        P3_U3396) );
  INV_X1 U16530 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14969) );
  INV_X1 U16531 ( .A(n15009), .ZN(n14996) );
  OAI22_X1 U16532 ( .A1(n14966), .A2(n14996), .B1(n14965), .B2(n15004), .ZN(
        n14967) );
  NOR2_X1 U16533 ( .A1(n14968), .A2(n14967), .ZN(n15015) );
  AOI22_X1 U16534 ( .A1(n15012), .A2(n14969), .B1(n15015), .B2(n15010), .ZN(
        P3_U3399) );
  INV_X1 U16535 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14975) );
  INV_X1 U16536 ( .A(n14972), .ZN(n14974) );
  NAND2_X1 U16537 ( .A1(n6914), .A2(n15001), .ZN(n14970) );
  OAI211_X1 U16538 ( .C1(n14996), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        n14973) );
  AOI21_X1 U16539 ( .B1(n14974), .B2(n14993), .A(n14973), .ZN(n15017) );
  AOI22_X1 U16540 ( .A1(n15012), .A2(n14975), .B1(n15017), .B2(n15010), .ZN(
        P3_U3402) );
  INV_X1 U16541 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14982) );
  INV_X1 U16542 ( .A(n14979), .ZN(n14981) );
  NAND2_X1 U16543 ( .A1(n14976), .A2(n15001), .ZN(n14977) );
  OAI211_X1 U16544 ( .C1(n14996), .C2(n14979), .A(n14978), .B(n14977), .ZN(
        n14980) );
  AOI21_X1 U16545 ( .B1(n14981), .B2(n14993), .A(n14980), .ZN(n15018) );
  AOI22_X1 U16546 ( .A1(n15012), .A2(n14982), .B1(n15018), .B2(n15010), .ZN(
        P3_U3405) );
  INV_X1 U16547 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14987) );
  NOR2_X1 U16548 ( .A1(n14983), .A2(n15004), .ZN(n14985) );
  AOI211_X1 U16549 ( .C1(n15009), .C2(n14986), .A(n14985), .B(n14984), .ZN(
        n15020) );
  AOI22_X1 U16550 ( .A1(n15012), .A2(n14987), .B1(n15020), .B2(n15010), .ZN(
        P3_U3408) );
  INV_X1 U16551 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15201) );
  INV_X1 U16552 ( .A(n14991), .ZN(n14994) );
  NAND2_X1 U16553 ( .A1(n14988), .A2(n15001), .ZN(n14989) );
  OAI211_X1 U16554 ( .C1(n14996), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14992) );
  AOI21_X1 U16555 ( .B1(n14994), .B2(n14993), .A(n14992), .ZN(n15021) );
  AOI22_X1 U16556 ( .A1(n15012), .A2(n15201), .B1(n15021), .B2(n15010), .ZN(
        P3_U3411) );
  INV_X1 U16557 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15002) );
  AOI21_X1 U16558 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n14999) );
  AOI211_X1 U16559 ( .C1(n15001), .C2(n15000), .A(n14999), .B(n14998), .ZN(
        n15022) );
  AOI22_X1 U16560 ( .A1(n15012), .A2(n15002), .B1(n15022), .B2(n15010), .ZN(
        P3_U3414) );
  INV_X1 U16561 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15011) );
  INV_X1 U16562 ( .A(n15003), .ZN(n15008) );
  NOR2_X1 U16563 ( .A1(n15005), .A2(n15004), .ZN(n15007) );
  AOI211_X1 U16564 ( .C1(n15009), .C2(n15008), .A(n15007), .B(n15006), .ZN(
        n15024) );
  AOI22_X1 U16565 ( .A1(n15012), .A2(n15011), .B1(n15024), .B2(n15010), .ZN(
        P3_U3417) );
  AOI22_X1 U16566 ( .A1(n15025), .A2(n15013), .B1(n8542), .B2(n15023), .ZN(
        P3_U3460) );
  AOI22_X1 U16567 ( .A1(n15025), .A2(n15014), .B1(n9651), .B2(n15023), .ZN(
        P3_U3461) );
  AOI22_X1 U16568 ( .A1(n15025), .A2(n15015), .B1(n9703), .B2(n15023), .ZN(
        P3_U3462) );
  AOI22_X1 U16569 ( .A1(n15025), .A2(n15017), .B1(n15016), .B2(n15023), .ZN(
        P3_U3463) );
  AOI22_X1 U16570 ( .A1(n15025), .A2(n15018), .B1(n9712), .B2(n15023), .ZN(
        P3_U3464) );
  AOI22_X1 U16571 ( .A1(n15025), .A2(n15020), .B1(n15019), .B2(n15023), .ZN(
        P3_U3465) );
  AOI22_X1 U16572 ( .A1(n15025), .A2(n15021), .B1(n9779), .B2(n15023), .ZN(
        P3_U3466) );
  AOI22_X1 U16573 ( .A1(n15025), .A2(n15022), .B1(n9864), .B2(n15023), .ZN(
        P3_U3467) );
  AOI22_X1 U16574 ( .A1(n15025), .A2(n15024), .B1(n10308), .B2(n15023), .ZN(
        P3_U3468) );
  INV_X1 U16575 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15027) );
  AOI22_X1 U16576 ( .A1(n15157), .A2(keyinput98), .B1(keyinput125), .B2(n15027), .ZN(n15026) );
  OAI221_X1 U16577 ( .B1(n15157), .B2(keyinput98), .C1(n15027), .C2(
        keyinput125), .A(n15026), .ZN(n15038) );
  AOI22_X1 U16578 ( .A1(n15194), .A2(keyinput109), .B1(n15029), .B2(keyinput94), .ZN(n15028) );
  OAI221_X1 U16579 ( .B1(n15194), .B2(keyinput109), .C1(n15029), .C2(
        keyinput94), .A(n15028), .ZN(n15037) );
  AOI22_X1 U16580 ( .A1(n15032), .A2(keyinput86), .B1(keyinput79), .B2(n15031), 
        .ZN(n15030) );
  OAI221_X1 U16581 ( .B1(n15032), .B2(keyinput86), .C1(n15031), .C2(keyinput79), .A(n15030), .ZN(n15036) );
  XNOR2_X1 U16582 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput117), .ZN(n15034) );
  XNOR2_X1 U16583 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput91), .ZN(n15033) );
  NAND2_X1 U16584 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  NOR4_X1 U16585 ( .A1(n15038), .A2(n15037), .A3(n15036), .A4(n15035), .ZN(
        n15079) );
  AOI22_X1 U16586 ( .A1(n10478), .A2(keyinput118), .B1(keyinput89), .B2(n15159), .ZN(n15039) );
  OAI221_X1 U16587 ( .B1(n10478), .B2(keyinput118), .C1(n15159), .C2(
        keyinput89), .A(n15039), .ZN(n15051) );
  INV_X1 U16588 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U16589 ( .A1(n9172), .A2(keyinput66), .B1(keyinput70), .B2(n15041), 
        .ZN(n15040) );
  OAI221_X1 U16590 ( .B1(n9172), .B2(keyinput66), .C1(n15041), .C2(keyinput70), 
        .A(n15040), .ZN(n15050) );
  INV_X1 U16591 ( .A(SI_28_), .ZN(n15044) );
  AOI22_X1 U16592 ( .A1(n15044), .A2(keyinput100), .B1(n15043), .B2(keyinput97), .ZN(n15042) );
  OAI221_X1 U16593 ( .B1(n15044), .B2(keyinput100), .C1(n15043), .C2(
        keyinput97), .A(n15042), .ZN(n15049) );
  AOI22_X1 U16594 ( .A1(n15047), .A2(keyinput122), .B1(keyinput76), .B2(n15046), .ZN(n15045) );
  OAI221_X1 U16595 ( .B1(n15047), .B2(keyinput122), .C1(n15046), .C2(
        keyinput76), .A(n15045), .ZN(n15048) );
  NOR4_X1 U16596 ( .A1(n15051), .A2(n15050), .A3(n15049), .A4(n15048), .ZN(
        n15078) );
  AOI22_X1 U16597 ( .A1(n15054), .A2(keyinput65), .B1(n15053), .B2(keyinput73), 
        .ZN(n15052) );
  OAI221_X1 U16598 ( .B1(n15054), .B2(keyinput65), .C1(n15053), .C2(keyinput73), .A(n15052), .ZN(n15064) );
  AOI22_X1 U16599 ( .A1(n15056), .A2(keyinput96), .B1(n11432), .B2(keyinput127), .ZN(n15055) );
  OAI221_X1 U16600 ( .B1(n15056), .B2(keyinput96), .C1(n11432), .C2(
        keyinput127), .A(n15055), .ZN(n15063) );
  AOI22_X1 U16601 ( .A1(n15192), .A2(keyinput95), .B1(n15058), .B2(keyinput67), 
        .ZN(n15057) );
  OAI221_X1 U16602 ( .B1(n15192), .B2(keyinput95), .C1(n15058), .C2(keyinput67), .A(n15057), .ZN(n15062) );
  XOR2_X1 U16603 ( .A(n12737), .B(keyinput68), .Z(n15060) );
  XNOR2_X1 U16604 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput69), .ZN(n15059) );
  NAND2_X1 U16605 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  NOR4_X1 U16606 ( .A1(n15064), .A2(n15063), .A3(n15062), .A4(n15061), .ZN(
        n15077) );
  AOI22_X1 U16607 ( .A1(n15066), .A2(keyinput105), .B1(n15193), .B2(keyinput93), .ZN(n15065) );
  OAI221_X1 U16608 ( .B1(n15066), .B2(keyinput105), .C1(n15193), .C2(
        keyinput93), .A(n15065), .ZN(n15075) );
  INV_X1 U16609 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U16610 ( .A1(n15185), .A2(keyinput102), .B1(keyinput88), .B2(n15165), .ZN(n15067) );
  OAI221_X1 U16611 ( .B1(n15185), .B2(keyinput102), .C1(n15165), .C2(
        keyinput88), .A(n15067), .ZN(n15074) );
  AOI22_X1 U16612 ( .A1(n15069), .A2(keyinput71), .B1(n15201), .B2(keyinput81), 
        .ZN(n15068) );
  OAI221_X1 U16613 ( .B1(n15069), .B2(keyinput71), .C1(n15201), .C2(keyinput81), .A(n15068), .ZN(n15073) );
  INV_X1 U16614 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U16615 ( .A1(n15164), .A2(keyinput99), .B1(n15071), .B2(keyinput119), .ZN(n15070) );
  OAI221_X1 U16616 ( .B1(n15164), .B2(keyinput99), .C1(n15071), .C2(
        keyinput119), .A(n15070), .ZN(n15072) );
  NOR4_X1 U16617 ( .A1(n15075), .A2(n15074), .A3(n15073), .A4(n15072), .ZN(
        n15076) );
  AND4_X1 U16618 ( .A1(n15079), .A2(n15078), .A3(n15077), .A4(n15076), .ZN(
        n15219) );
  OAI22_X1 U16619 ( .A1(P1_D_REG_12__SCAN_IN), .A2(keyinput112), .B1(
        P2_REG0_REG_23__SCAN_IN), .B2(keyinput84), .ZN(n15080) );
  AOI221_X1 U16620 ( .B1(P1_D_REG_12__SCAN_IN), .B2(keyinput112), .C1(
        keyinput84), .C2(P2_REG0_REG_23__SCAN_IN), .A(n15080), .ZN(n15087) );
  OAI22_X1 U16621 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput110), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput115), .ZN(n15081) );
  AOI221_X1 U16622 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput110), .C1(
        keyinput115), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n15081), .ZN(n15086) );
  OAI22_X1 U16623 ( .A1(P3_REG2_REG_23__SCAN_IN), .A2(keyinput114), .B1(
        P1_REG2_REG_8__SCAN_IN), .B2(keyinput77), .ZN(n15082) );
  AOI221_X1 U16624 ( .B1(P3_REG2_REG_23__SCAN_IN), .B2(keyinput114), .C1(
        keyinput77), .C2(P1_REG2_REG_8__SCAN_IN), .A(n15082), .ZN(n15085) );
  OAI22_X1 U16625 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(keyinput78), .B1(
        keyinput124), .B2(P1_REG0_REG_14__SCAN_IN), .ZN(n15083) );
  AOI221_X1 U16626 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(keyinput78), .C1(
        P1_REG0_REG_14__SCAN_IN), .C2(keyinput124), .A(n15083), .ZN(n15084) );
  NAND4_X1 U16627 ( .A1(n15087), .A2(n15086), .A3(n15085), .A4(n15084), .ZN(
        n15119) );
  OAI22_X1 U16628 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput104), .B1(
        P1_REG0_REG_6__SCAN_IN), .B2(keyinput80), .ZN(n15088) );
  AOI221_X1 U16629 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput104), .C1(
        keyinput80), .C2(P1_REG0_REG_6__SCAN_IN), .A(n15088), .ZN(n15095) );
  OAI22_X1 U16630 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput116), .B1(
        P1_REG0_REG_4__SCAN_IN), .B2(keyinput103), .ZN(n15089) );
  AOI221_X1 U16631 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput116), .C1(
        keyinput103), .C2(P1_REG0_REG_4__SCAN_IN), .A(n15089), .ZN(n15094) );
  OAI22_X1 U16632 ( .A1(P1_D_REG_24__SCAN_IN), .A2(keyinput64), .B1(keyinput74), .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n15090) );
  AOI221_X1 U16633 ( .B1(P1_D_REG_24__SCAN_IN), .B2(keyinput64), .C1(
        P3_DATAO_REG_15__SCAN_IN), .C2(keyinput74), .A(n15090), .ZN(n15093) );
  OAI22_X1 U16634 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput82), .B1(
        P2_REG0_REG_31__SCAN_IN), .B2(keyinput90), .ZN(n15091) );
  AOI221_X1 U16635 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput82), .C1(
        keyinput90), .C2(P2_REG0_REG_31__SCAN_IN), .A(n15091), .ZN(n15092) );
  NAND4_X1 U16636 ( .A1(n15095), .A2(n15094), .A3(n15093), .A4(n15092), .ZN(
        n15118) );
  OAI22_X1 U16637 ( .A1(SI_14_), .A2(keyinput111), .B1(keyinput108), .B2(
        P1_REG3_REG_15__SCAN_IN), .ZN(n15096) );
  AOI221_X1 U16638 ( .B1(SI_14_), .B2(keyinput111), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput108), .A(n15096), .ZN(n15097) );
  INV_X1 U16639 ( .A(n15097), .ZN(n15104) );
  XNOR2_X1 U16640 ( .A(n15098), .B(keyinput72), .ZN(n15103) );
  XNOR2_X1 U16641 ( .A(n15186), .B(keyinput101), .ZN(n15100) );
  XNOR2_X1 U16642 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput92), .ZN(n15099) );
  NAND2_X1 U16643 ( .A1(n15100), .A2(n15099), .ZN(n15102) );
  XNOR2_X1 U16644 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(keyinput83), .ZN(n15101) );
  NOR4_X1 U16645 ( .A1(n15104), .A2(n15103), .A3(n15102), .A4(n15101), .ZN(
        n15107) );
  OAI22_X1 U16646 ( .A1(P3_REG2_REG_1__SCAN_IN), .A2(keyinput113), .B1(
        keyinput85), .B2(P1_REG1_REG_4__SCAN_IN), .ZN(n15105) );
  AOI221_X1 U16647 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(keyinput113), .C1(
        P1_REG1_REG_4__SCAN_IN), .C2(keyinput85), .A(n15105), .ZN(n15106) );
  NAND2_X1 U16648 ( .A1(n15107), .A2(n15106), .ZN(n15117) );
  OAI22_X1 U16649 ( .A1(P3_D_REG_5__SCAN_IN), .A2(keyinput121), .B1(keyinput87), .B2(P2_REG2_REG_10__SCAN_IN), .ZN(n15108) );
  AOI221_X1 U16650 ( .B1(P3_D_REG_5__SCAN_IN), .B2(keyinput121), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(keyinput87), .A(n15108), .ZN(n15115) );
  OAI22_X1 U16651 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput123), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput106), .ZN(n15109) );
  AOI221_X1 U16652 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput123), .C1(
        keyinput106), .C2(P3_REG3_REG_10__SCAN_IN), .A(n15109), .ZN(n15114) );
  OAI22_X1 U16653 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(keyinput126), .B1(
        keyinput75), .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n15110) );
  AOI221_X1 U16654 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput126), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput75), .A(n15110), .ZN(n15113) );
  OAI22_X1 U16655 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(keyinput120), .B1(
        keyinput107), .B2(P2_D_REG_24__SCAN_IN), .ZN(n15111) );
  AOI221_X1 U16656 ( .B1(P2_DATAO_REG_4__SCAN_IN), .B2(keyinput120), .C1(
        P2_D_REG_24__SCAN_IN), .C2(keyinput107), .A(n15111), .ZN(n15112) );
  NAND4_X1 U16657 ( .A1(n15115), .A2(n15114), .A3(n15113), .A4(n15112), .ZN(
        n15116) );
  NOR4_X1 U16658 ( .A1(n15119), .A2(n15118), .A3(n15117), .A4(n15116), .ZN(
        n15218) );
  AOI22_X1 U16659 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(keyinput41), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput51), .ZN(n15120) );
  OAI221_X1 U16660 ( .B1(P3_DATAO_REG_27__SCAN_IN), .B2(keyinput41), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput51), .A(n15120), .ZN(n15127) );
  AOI22_X1 U16661 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput60), .B1(
        P1_REG3_REG_16__SCAN_IN), .B2(keyinput63), .ZN(n15121) );
  OAI221_X1 U16662 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput60), .C1(
        P1_REG3_REG_16__SCAN_IN), .C2(keyinput63), .A(n15121), .ZN(n15126) );
  AOI22_X1 U16663 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput32), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(keyinput11), .ZN(n15122) );
  OAI221_X1 U16664 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput32), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput11), .A(n15122), .ZN(n15125) );
  AOI22_X1 U16665 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput13), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput42), .ZN(n15123) );
  OAI221_X1 U16666 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput13), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput42), .A(n15123), .ZN(n15124) );
  NOR4_X1 U16667 ( .A1(n15127), .A2(n15126), .A3(n15125), .A4(n15124), .ZN(
        n15155) );
  AOI22_X1 U16668 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(keyinput26), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(keyinput56), .ZN(n15128) );
  OAI221_X1 U16669 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(keyinput26), .C1(
        P2_DATAO_REG_4__SCAN_IN), .C2(keyinput56), .A(n15128), .ZN(n15135) );
  AOI22_X1 U16670 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(keyinput3), .B1(
        P3_D_REG_15__SCAN_IN), .B2(keyinput55), .ZN(n15129) );
  OAI221_X1 U16671 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(keyinput3), .C1(
        P3_D_REG_15__SCAN_IN), .C2(keyinput55), .A(n15129), .ZN(n15134) );
  AOI22_X1 U16672 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput19), .B1(
        P2_REG0_REG_14__SCAN_IN), .B2(keyinput6), .ZN(n15130) );
  OAI221_X1 U16673 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG0_REG_14__SCAN_IN), .C2(keyinput6), .A(n15130), .ZN(n15133) );
  AOI22_X1 U16674 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput23), .B1(
        P1_D_REG_30__SCAN_IN), .B2(keyinput40), .ZN(n15131) );
  OAI221_X1 U16675 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput23), .C1(
        P1_D_REG_30__SCAN_IN), .C2(keyinput40), .A(n15131), .ZN(n15132) );
  NOR4_X1 U16676 ( .A1(n15135), .A2(n15134), .A3(n15133), .A4(n15132), .ZN(
        n15154) );
  AOI22_X1 U16677 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(keyinput54), .B1(
        P3_IR_REG_14__SCAN_IN), .B2(keyinput5), .ZN(n15136) );
  OAI221_X1 U16678 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(keyinput54), .C1(
        P3_IR_REG_14__SCAN_IN), .C2(keyinput5), .A(n15136), .ZN(n15143) );
  AOI22_X1 U16679 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput28), .B1(
        P1_REG0_REG_6__SCAN_IN), .B2(keyinput16), .ZN(n15137) );
  OAI221_X1 U16680 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput28), .C1(
        P1_REG0_REG_6__SCAN_IN), .C2(keyinput16), .A(n15137), .ZN(n15142) );
  AOI22_X1 U16681 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput39), .B1(
        P3_D_REG_22__SCAN_IN), .B2(keyinput9), .ZN(n15138) );
  OAI221_X1 U16682 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput39), .C1(
        P3_D_REG_22__SCAN_IN), .C2(keyinput9), .A(n15138), .ZN(n15141) );
  AOI22_X1 U16683 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput12), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput48), .ZN(n15139) );
  OAI221_X1 U16684 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput12), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput48), .A(n15139), .ZN(n15140) );
  NOR4_X1 U16685 ( .A1(n15143), .A2(n15142), .A3(n15141), .A4(n15140), .ZN(
        n15153) );
  AOI22_X1 U16686 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput33), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput30), .ZN(n15144) );
  OAI221_X1 U16687 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput33), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput30), .A(n15144), .ZN(n15151) );
  AOI22_X1 U16688 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput61), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput46), .ZN(n15145) );
  OAI221_X1 U16689 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput61), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput46), .A(n15145), .ZN(n15150) );
  AOI22_X1 U16690 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(keyinput14), .B1(
        P1_D_REG_8__SCAN_IN), .B2(keyinput1), .ZN(n15146) );
  OAI221_X1 U16691 ( .B1(P1_REG2_REG_23__SCAN_IN), .B2(keyinput14), .C1(
        P1_D_REG_8__SCAN_IN), .C2(keyinput1), .A(n15146), .ZN(n15149) );
  AOI22_X1 U16692 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(keyinput58), .B1(SI_28_), 
        .B2(keyinput36), .ZN(n15147) );
  OAI221_X1 U16693 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(keyinput58), .C1(SI_28_), .C2(keyinput36), .A(n15147), .ZN(n15148) );
  NOR4_X1 U16694 ( .A1(n15151), .A2(n15150), .A3(n15149), .A4(n15148), .ZN(
        n15152) );
  NAND4_X1 U16695 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        n15217) );
  AOI22_X1 U16696 ( .A1(n15157), .A2(keyinput34), .B1(keyinput21), .B2(n9228), 
        .ZN(n15156) );
  OAI221_X1 U16697 ( .B1(n15157), .B2(keyinput34), .C1(n9228), .C2(keyinput21), 
        .A(n15156), .ZN(n15169) );
  AOI22_X1 U16698 ( .A1(n15160), .A2(keyinput20), .B1(keyinput25), .B2(n15159), 
        .ZN(n15158) );
  OAI221_X1 U16699 ( .B1(n15160), .B2(keyinput20), .C1(n15159), .C2(keyinput25), .A(n15158), .ZN(n15168) );
  AOI22_X1 U16700 ( .A1(n12737), .A2(keyinput4), .B1(n15162), .B2(keyinput57), 
        .ZN(n15161) );
  OAI221_X1 U16701 ( .B1(n12737), .B2(keyinput4), .C1(n15162), .C2(keyinput57), 
        .A(n15161), .ZN(n15167) );
  AOI22_X1 U16702 ( .A1(n15165), .A2(keyinput24), .B1(keyinput35), .B2(n15164), 
        .ZN(n15163) );
  OAI221_X1 U16703 ( .B1(n15165), .B2(keyinput24), .C1(n15164), .C2(keyinput35), .A(n15163), .ZN(n15166) );
  NOR4_X1 U16704 ( .A1(n15169), .A2(n15168), .A3(n15167), .A4(n15166), .ZN(
        n15215) );
  AOI22_X1 U16705 ( .A1(n15172), .A2(keyinput47), .B1(keyinput43), .B2(n15171), 
        .ZN(n15170) );
  OAI221_X1 U16706 ( .B1(n15172), .B2(keyinput47), .C1(n15171), .C2(keyinput43), .A(n15170), .ZN(n15180) );
  AOI22_X1 U16707 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput22), .B1(n9172), 
        .B2(keyinput2), .ZN(n15173) );
  OAI221_X1 U16708 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput22), .C1(n9172), 
        .C2(keyinput2), .A(n15173), .ZN(n15179) );
  AOI22_X1 U16709 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput7), .B1(SI_27_), 
        .B2(keyinput15), .ZN(n15174) );
  OAI221_X1 U16710 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput7), .C1(SI_27_), 
        .C2(keyinput15), .A(n15174), .ZN(n15178) );
  XOR2_X1 U16711 ( .A(n10834), .B(keyinput49), .Z(n15176) );
  XNOR2_X1 U16712 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput8), .ZN(n15175) );
  NAND2_X1 U16713 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  NOR4_X1 U16714 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15214) );
  AOI22_X1 U16715 ( .A1(n15183), .A2(keyinput10), .B1(n15182), .B2(keyinput59), 
        .ZN(n15181) );
  OAI221_X1 U16716 ( .B1(n15183), .B2(keyinput10), .C1(n15182), .C2(keyinput59), .A(n15181), .ZN(n15190) );
  AOI22_X1 U16717 ( .A1(n15186), .A2(keyinput37), .B1(keyinput38), .B2(n15185), 
        .ZN(n15184) );
  OAI221_X1 U16718 ( .B1(n15186), .B2(keyinput37), .C1(n15185), .C2(keyinput38), .A(n15184), .ZN(n15189) );
  XNOR2_X1 U16719 ( .A(n15187), .B(keyinput27), .ZN(n15188) );
  OR3_X1 U16720 ( .A1(n15190), .A2(n15189), .A3(n15188), .ZN(n15197) );
  AOI22_X1 U16721 ( .A1(n15193), .A2(keyinput29), .B1(n15192), .B2(keyinput31), 
        .ZN(n15191) );
  OAI221_X1 U16722 ( .B1(n15193), .B2(keyinput29), .C1(n15192), .C2(keyinput31), .A(n15191), .ZN(n15196) );
  XNOR2_X1 U16723 ( .A(n15194), .B(keyinput45), .ZN(n15195) );
  NOR3_X1 U16724 ( .A1(n15197), .A2(n15196), .A3(n15195), .ZN(n15213) );
  AOI22_X1 U16725 ( .A1(n15199), .A2(keyinput18), .B1(keyinput50), .B2(n12793), 
        .ZN(n15198) );
  OAI221_X1 U16726 ( .B1(n15199), .B2(keyinput18), .C1(n12793), .C2(keyinput50), .A(n15198), .ZN(n15211) );
  AOI22_X1 U16727 ( .A1(n15202), .A2(keyinput62), .B1(keyinput17), .B2(n15201), 
        .ZN(n15200) );
  OAI221_X1 U16728 ( .B1(n15202), .B2(keyinput62), .C1(n15201), .C2(keyinput17), .A(n15200), .ZN(n15210) );
  AOI22_X1 U16729 ( .A1(n15205), .A2(keyinput0), .B1(n15204), .B2(keyinput52), 
        .ZN(n15203) );
  OAI221_X1 U16730 ( .B1(n15205), .B2(keyinput0), .C1(n15204), .C2(keyinput52), 
        .A(n15203), .ZN(n15209) );
  XNOR2_X1 U16731 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput53), .ZN(n15207) );
  XNOR2_X1 U16732 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput44), .ZN(n15206)
         );
  NAND2_X1 U16733 ( .A1(n15207), .A2(n15206), .ZN(n15208) );
  NOR4_X1 U16734 ( .A1(n15211), .A2(n15210), .A3(n15209), .A4(n15208), .ZN(
        n15212) );
  NAND4_X1 U16735 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15216) );
  AOI211_X1 U16736 ( .C1(n15219), .C2(n15218), .A(n15217), .B(n15216), .ZN(
        n15235) );
  AND2_X1 U16737 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15232) );
  AOI21_X1 U16738 ( .B1(n15221), .B2(P2_REG2_REG_18__SCAN_IN), .A(n15220), 
        .ZN(n15229) );
  OAI211_X1 U16739 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n15224), .A(n15223), 
        .B(n15222), .ZN(n15228) );
  NAND2_X1 U16740 ( .A1(n15226), .A2(n15225), .ZN(n15227) );
  OAI211_X1 U16741 ( .C1(n15230), .C2(n15229), .A(n15228), .B(n15227), .ZN(
        n15231) );
  AOI211_X1 U16742 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15233), .A(n15232), 
        .B(n15231), .ZN(n15234) );
  XNOR2_X1 U16743 ( .A(n15235), .B(n15234), .ZN(P2_U3232) );
  XNOR2_X1 U16744 ( .A(n15237), .B(n15236), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16745 ( .A(n15238), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16746 ( .B1(n15240), .B2(n15239), .A(n15244), .ZN(SUB_1596_U53) );
  XOR2_X1 U16747 ( .A(n15241), .B(n15242), .Z(SUB_1596_U56) );
  XOR2_X1 U16748 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15243), .Z(SUB_1596_U60) );
  XOR2_X1 U16749 ( .A(n15245), .B(n15244), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7235 ( .A(n8928), .Z(n6484) );
  OR3_X1 U7306 ( .A1(n14085), .A2(n14100), .A3(n12087), .ZN(n12088) );
  NOR2_X1 U9332 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7425) );
  NOR2_X1 U9491 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9047) );
  AOI211_X1 U9585 ( .C1(n14691), .C2(n14266), .A(n14265), .B(n14264), .ZN(
        n14268) );
  AND4_X2 U11433 ( .A1(n9959), .A2(n9048), .A3(n9047), .A4(n9166), .ZN(n15253)
         );
endmodule

