

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9578, n9579, n9580, n9582, n9583, n9584, n9585, n9586, n9588, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9626, n9627, n9628, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915;

  OR2_X1 U11022 ( .A1(n15209), .A2(n10909), .ZN(n15210) );
  OR3_X1 U11023 ( .A1(n12362), .A2(n10402), .A3(n10953), .ZN(n14324) );
  NAND2_X1 U11024 ( .A1(n17588), .A2(n17912), .ZN(n17909) );
  AND2_X1 U11025 ( .A1(n10129), .A2(n10124), .ZN(n9653) );
  CLKBUF_X2 U11027 ( .A(n12174), .Z(n9633) );
  BUF_X1 U11028 ( .A(n10774), .Z(n10844) );
  NAND2_X1 U11029 ( .A1(n11170), .A2(n11169), .ZN(n13695) );
  BUF_X1 U11030 ( .A(n10027), .Z(n15676) );
  BUF_X1 U11031 ( .A(n11117), .Z(n14962) );
  CLKBUF_X2 U11032 ( .A(n9588), .Z(n9601) );
  INV_X1 U11033 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19716) );
  CLKBUF_X1 U11034 ( .A(n11114), .Z(n20078) );
  CLKBUF_X1 U11035 ( .A(n12507), .Z(n9594) );
  NOR2_X1 U11036 ( .A1(n13261), .A2(n14389), .ZN(n11083) );
  AND2_X2 U11038 ( .A1(n10145), .A2(n12491), .ZN(n10160) );
  AND2_X2 U11039 ( .A1(n12649), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10259) );
  CLKBUF_X2 U11040 ( .A(n12716), .Z(n17330) );
  CLKBUF_X1 U11041 ( .A(n12507), .Z(n9593) );
  CLKBUF_X2 U11042 ( .A(n12731), .Z(n17160) );
  INV_X1 U11043 ( .A(n15699), .ZN(n9965) );
  AND2_X2 U11044 ( .A1(n9930), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10300) );
  INV_X2 U11046 ( .A(n12760), .ZN(n17201) );
  NAND2_X2 U11047 ( .A1(n9781), .A2(n9780), .ZN(n19203) );
  INV_X1 U11048 ( .A(n11021), .ZN(n9590) );
  AOI22_X1 U11049 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n9971) );
  AND2_X4 U11050 ( .A1(n10494), .A2(n9897), .ZN(n9930) );
  INV_X2 U11052 ( .A(n9923), .ZN(n12632) );
  AND2_X2 U11053 ( .A1(n10143), .A2(n13794), .ZN(n12655) );
  INV_X1 U11054 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15659) );
  CLKBUF_X1 U11055 ( .A(n19178), .Z(n9578) );
  NOR2_X1 U11056 ( .A1(n13110), .A2(n19849), .ZN(n19178) );
  CLKBUF_X1 U11057 ( .A(n20033), .Z(n9579) );
  NOR2_X1 U11058 ( .A1(n20032), .A2(n20031), .ZN(n20033) );
  CLKBUF_X1 U11059 ( .A(n20083), .Z(n9580) );
  NOR2_X1 U11060 ( .A1(n20031), .A2(n20030), .ZN(n20083) );
  INV_X2 U11062 ( .A(n20913), .ZN(n9582) );
  INV_X1 U11066 ( .A(n12087), .ZN(n12035) );
  NAND2_X2 U11067 ( .A1(n10963), .A2(n13680), .ZN(n11021) );
  INV_X1 U11068 ( .A(n12096), .ZN(n11177) );
  INV_X1 U11069 ( .A(n9617), .ZN(n12060) );
  CLKBUF_X2 U11070 ( .A(n11126), .Z(n11860) );
  INV_X1 U11072 ( .A(n10477), .ZN(n10350) );
  OR2_X1 U11073 ( .A1(n15834), .A2(n16932), .ZN(n17188) );
  INV_X2 U11074 ( .A(n16052), .ZN(n14748) );
  XNOR2_X1 U11075 ( .A(n11395), .B(n20007), .ZN(n13609) );
  INV_X1 U11076 ( .A(n12882), .ZN(n17186) );
  NAND2_X1 U11077 ( .A1(n11738), .A2(n11737), .ZN(n14533) );
  AND2_X1 U11078 ( .A1(n10392), .A2(n10419), .ZN(n10418) );
  NAND2_X1 U11079 ( .A1(n10812), .A2(n10811), .ZN(n13985) );
  NOR2_X1 U11080 ( .A1(n15189), .A2(n15188), .ZN(n14328) );
  NAND2_X1 U11081 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16883) );
  CLKBUF_X3 U11082 ( .A(n12173), .Z(n20037) );
  NOR2_X1 U11084 ( .A1(n13614), .A2(n13615), .ZN(n15567) );
  INV_X1 U11085 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13794) );
  INV_X2 U11086 ( .A(n18274), .ZN(n17232) );
  INV_X1 U11087 ( .A(n15698), .ZN(n15696) );
  INV_X1 U11088 ( .A(n19902), .ZN(n19924) );
  INV_X1 U11090 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12933) );
  INV_X1 U11091 ( .A(n12083), .ZN(n11949) );
  MUX2_X1 U11092 ( .A(n14646), .B(n14645), .S(n16052), .Z(n14647) );
  OAI22_X1 U11093 ( .A1(n13370), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11392), 
        .B2(n11267), .ZN(n11192) );
  AND2_X1 U11095 ( .A1(n10143), .A2(n13794), .ZN(n9583) );
  AND2_X2 U11096 ( .A1(n10143), .A2(n13794), .ZN(n9584) );
  AND2_X2 U11097 ( .A1(n13694), .A2(n10964), .ZN(n11211) );
  OAI211_X2 U11098 ( .C1(n12994), .C2(n12993), .A(n12992), .B(n12991), .ZN(
        n17801) );
  AND2_X2 U11099 ( .A1(n11114), .A2(n9635), .ZN(n11526) );
  AND2_X2 U11100 ( .A1(n11108), .A2(n9835), .ZN(n13266) );
  AND2_X4 U11101 ( .A1(n10976), .A2(n10977), .ZN(n11108) );
  NAND2_X2 U11102 ( .A1(n9783), .A2(n9897), .ZN(n9923) );
  AND4_X2 U11103 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10976) );
  BUF_X4 U11106 ( .A(n10070), .Z(n10841) );
  NAND2_X1 U11107 ( .A1(n12189), .A2(n14380), .ZN(n13516) );
  XOR2_X2 U11108 ( .A(n12988), .B(n12987), .Z(n17831) );
  OR2_X2 U11109 ( .A1(n13383), .A2(n11139), .ZN(n13514) );
  XNOR2_X2 U11110 ( .A(n14647), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14790) );
  OAI21_X2 U11111 ( .B1(n14156), .B2(n11464), .A(n11463), .ZN(n11465) );
  INV_X1 U11112 ( .A(n10560), .ZN(n9585) );
  NAND2_X2 U11113 ( .A1(n9922), .A2(n9921), .ZN(n10017) );
  INV_X2 U11114 ( .A(n10017), .ZN(n10560) );
  INV_X1 U11115 ( .A(n12099), .ZN(n9586) );
  NAND2_X1 U11117 ( .A1(n10969), .A2(n13694), .ZN(n12057) );
  INV_X1 U11119 ( .A(n11775), .ZN(n9588) );
  INV_X2 U11120 ( .A(n14677), .ZN(n14666) );
  NAND2_X2 U11121 ( .A1(n11469), .A2(n14685), .ZN(n14677) );
  NAND2_X2 U11122 ( .A1(n13607), .A2(n11396), .ZN(n11401) );
  INV_X2 U11123 ( .A(n12083), .ZN(n9591) );
  INV_X1 U11124 ( .A(n9591), .ZN(n9592) );
  NAND2_X1 U11125 ( .A1(n10964), .A2(n10968), .ZN(n12083) );
  XOR2_X2 U11126 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12984), .Z(
        n17843) );
  NAND2_X2 U11127 ( .A1(n12983), .A2(n17854), .ZN(n12984) );
  AND2_X1 U11128 ( .A1(n9930), .A2(n9928), .ZN(n12507) );
  AND2_X4 U11129 ( .A1(n10963), .A2(n10964), .ZN(n11919) );
  NOR2_X4 U11130 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10964) );
  BUF_X2 U11132 ( .A(n12393), .Z(n9595) );
  XNOR2_X1 U11133 ( .A(n10086), .B(n10089), .ZN(n12393) );
  NAND2_X2 U11134 ( .A1(n9964), .A2(n9963), .ZN(n15699) );
  AND2_X4 U11135 ( .A1(n19849), .A2(n19240), .ZN(n10577) );
  INV_X1 U11136 ( .A(n17051), .ZN(n9596) );
  INV_X4 U11137 ( .A(n17051), .ZN(n17170) );
  AND2_X1 U11138 ( .A1(n12379), .A2(n13273), .ZN(n10125) );
  NAND2_X2 U11139 ( .A1(n13565), .A2(n11389), .ZN(n11395) );
  NAND2_X2 U11140 ( .A1(n10077), .A2(n10076), .ZN(n10749) );
  NAND2_X2 U11141 ( .A1(n11495), .A2(n20037), .ZN(n20744) );
  INV_X1 U11142 ( .A(n20054), .ZN(n11495) );
  AOI21_X1 U11143 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14667), .A(
        n14661), .ZN(n14662) );
  NAND2_X1 U11144 ( .A1(n9843), .A2(n9841), .ZN(n14156) );
  OAI21_X1 U11145 ( .B1(n14708), .B2(n9846), .A(n9844), .ZN(n14155) );
  NAND2_X1 U11146 ( .A1(n17570), .A2(n9807), .ZN(n12815) );
  AND2_X1 U11147 ( .A1(n15344), .A2(n16304), .ZN(n10892) );
  AOI21_X1 U11148 ( .B1(n9846), .B2(n9844), .A(n9842), .ZN(n9841) );
  NOR2_X2 U11149 ( .A1(n17718), .A2(n18058), .ZN(n18044) );
  NOR2_X1 U11150 ( .A1(n13586), .A2(n13592), .ZN(n13631) );
  OR2_X1 U11151 ( .A1(n13073), .A2(n13074), .ZN(n15023) );
  AND2_X1 U11152 ( .A1(n13571), .A2(n13572), .ZN(n13574) );
  NAND2_X1 U11153 ( .A1(n18143), .A2(n17811), .ZN(n17810) );
  NAND2_X1 U11155 ( .A1(n17817), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17816) );
  XNOR2_X1 U11156 ( .A(n12790), .B(n12789), .ZN(n17817) );
  NAND2_X1 U11157 ( .A1(n17832), .A2(n12787), .ZN(n12790) );
  NAND2_X1 U11158 ( .A1(n11171), .A2(n13695), .ZN(n13370) );
  NAND2_X1 U11159 ( .A1(n13462), .A2(n13227), .ZN(n20739) );
  INV_X4 U11160 ( .A(n16874), .ZN(n16903) );
  XNOR2_X1 U11161 ( .A(n10088), .B(n10087), .ZN(n10089) );
  NAND2_X2 U11162 ( .A1(n11523), .A2(n11524), .ZN(n13499) );
  OR2_X1 U11163 ( .A1(n10774), .A2(n13806), .ZN(n10084) );
  INV_X4 U11164 ( .A(n12329), .ZN(n12347) );
  NAND2_X1 U11165 ( .A1(n17872), .A2(n17871), .ZN(n17870) );
  XNOR2_X1 U11166 ( .A(n12776), .B(n12774), .ZN(n17872) );
  NAND2_X1 U11167 ( .A1(n10034), .A2(n13783), .ZN(n10855) );
  AND2_X1 U11168 ( .A1(n10272), .A2(n10273), .ZN(n10343) );
  AND2_X1 U11169 ( .A1(n9966), .A2(n10036), .ZN(n10927) );
  CLKBUF_X1 U11170 ( .A(n10745), .Z(n16341) );
  INV_X1 U11171 ( .A(n10705), .ZN(n9850) );
  NAND2_X1 U11172 ( .A1(n13512), .A2(n11362), .ZN(n11136) );
  NAND2_X1 U11173 ( .A1(n12156), .A2(n20054), .ZN(n13817) );
  AND3_X1 U11174 ( .A1(n15717), .A2(n15699), .A3(n9967), .ZN(n10019) );
  CLKBUF_X2 U11176 ( .A(n11107), .Z(n9634) );
  CLKBUF_X2 U11177 ( .A(n10584), .Z(n10725) );
  NAND4_X1 U11178 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(
        n11362) );
  AND2_X1 U11179 ( .A1(n9892), .A2(n9871), .ZN(n13506) );
  NAND2_X1 U11180 ( .A1(n9914), .A2(n9913), .ZN(n9922) );
  AND4_X1 U11181 ( .A1(n11013), .A2(n11012), .A3(n11011), .A4(n11010), .ZN(
        n11018) );
  CLKBUF_X2 U11182 ( .A(n11206), .Z(n12099) );
  AND4_X1 U11183 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10005) );
  AND3_X1 U11184 ( .A1(n9910), .A2(n9981), .A3(n9909), .ZN(n9914) );
  AND2_X1 U11185 ( .A1(n9982), .A2(n9981), .ZN(n9986) );
  AND2_X2 U11186 ( .A1(n12490), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10211) );
  INV_X1 U11187 ( .A(n12726), .ZN(n17022) );
  CLKBUF_X2 U11188 ( .A(n12904), .Z(n17155) );
  CLKBUF_X2 U11189 ( .A(n12716), .Z(n17094) );
  CLKBUF_X1 U11190 ( .A(n13681), .Z(n9617) );
  CLKBUF_X2 U11191 ( .A(n12731), .Z(n17331) );
  INV_X2 U11192 ( .A(n11021), .ZN(n12097) );
  OR2_X1 U11194 ( .A1(n18675), .A2(n12688), .ZN(n12848) );
  BUF_X2 U11195 ( .A(n9970), .Z(n12570) );
  NAND2_X1 U11196 ( .A1(n13682), .A2(n9759), .ZN(n13681) );
  AND2_X2 U11197 ( .A1(n10145), .A2(n13794), .ZN(n12658) );
  OR2_X1 U11198 ( .A1(n12689), .A2(n12688), .ZN(n17051) );
  INV_X4 U11199 ( .A(n17188), .ZN(n17341) );
  AND2_X2 U11200 ( .A1(n13682), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11126) );
  AND2_X2 U11201 ( .A1(n9623), .A2(n9981), .ZN(n10154) );
  NAND2_X1 U11202 ( .A1(n18849), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12689) );
  AND2_X1 U11204 ( .A1(n9894), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15662) );
  AND3_X2 U11205 ( .A1(n9782), .A2(n15659), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U11207 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12491) );
  AND2_X1 U11208 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10494) );
  AND2_X1 U11211 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13680) );
  OR2_X1 U11212 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16932) );
  AOI211_X1 U11213 ( .C1(n19198), .C2(n15528), .A(n15340), .B(n15339), .ZN(
        n15341) );
  AND3_X1 U11214 ( .A1(n10957), .A2(n10956), .A3(n10955), .ZN(n9882) );
  AOI21_X1 U11215 ( .B1(n14275), .B2(n16052), .A(n14274), .ZN(n14626) );
  NAND2_X1 U11216 ( .A1(n9709), .A2(n9708), .ZN(n15337) );
  AND2_X1 U11217 ( .A1(n12675), .A2(n12674), .ZN(n12676) );
  AOI211_X1 U11218 ( .C1(n15213), .C2(n19198), .A(n15212), .B(n15211), .ZN(
        n15214) );
  AOI211_X1 U11219 ( .C1(n15385), .C2(n15384), .A(n15383), .B(n15382), .ZN(
        n15386) );
  AOI211_X1 U11220 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15385), .A(
        n15370), .B(n15369), .ZN(n15373) );
  NOR2_X2 U11221 ( .A1(n15210), .A2(n15364), .ZN(n15194) );
  AND2_X1 U11222 ( .A1(n9610), .A2(n9883), .ZN(n14653) );
  AND2_X1 U11223 ( .A1(n14258), .A2(n10854), .ZN(n12673) );
  XNOR2_X1 U11224 ( .A(n14396), .B(n12162), .ZN(n14394) );
  NOR2_X1 U11225 ( .A1(n9734), .A2(n9673), .ZN(n15223) );
  NOR2_X2 U11226 ( .A1(n15064), .A2(n15065), .ZN(n15063) );
  AND2_X1 U11227 ( .A1(n15078), .A2(n15077), .ZN(n15080) );
  NOR2_X1 U11228 ( .A1(n15840), .A2(n16396), .ZN(n15890) );
  OR2_X1 U11229 ( .A1(n14155), .A2(n11466), .ZN(n14693) );
  NAND2_X1 U11230 ( .A1(n15249), .A2(n10464), .ZN(n15241) );
  OR2_X1 U11231 ( .A1(n14504), .A2(n14431), .ZN(n14498) );
  NAND2_X1 U11232 ( .A1(n14172), .A2(n14171), .ZN(n15263) );
  OR2_X1 U11233 ( .A1(n14506), .A2(n14507), .ZN(n14504) );
  NOR2_X1 U11234 ( .A1(n15083), .A2(n15082), .ZN(n15081) );
  OR2_X2 U11235 ( .A1(n15008), .A2(n15011), .ZN(n15009) );
  NAND2_X1 U11236 ( .A1(n14708), .A2(n9844), .ZN(n9843) );
  NOR2_X2 U11237 ( .A1(n16415), .A2(n12815), .ZN(n17563) );
  OAI21_X1 U11238 ( .B1(n9790), .B2(n9791), .A(n15072), .ZN(n15083) );
  XNOR2_X1 U11239 ( .A(n10469), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15225) );
  NAND2_X1 U11240 ( .A1(n9729), .A2(n9647), .ZN(n16218) );
  NAND2_X1 U11241 ( .A1(n9791), .A2(n9790), .ZN(n15072) );
  NOR2_X2 U11242 ( .A1(n15038), .A2(n13071), .ZN(n15020) );
  NAND2_X1 U11243 ( .A1(n17599), .A2(n17603), .ZN(n17598) );
  OR2_X1 U11244 ( .A1(n15274), .A2(n10436), .ZN(n15264) );
  AND2_X1 U11245 ( .A1(n15620), .A2(n15621), .ZN(n9778) );
  NAND2_X1 U11246 ( .A1(n11432), .A2(n11431), .ZN(n16065) );
  NOR2_X1 U11247 ( .A1(n17672), .A2(n13001), .ZN(n17604) );
  AND2_X1 U11248 ( .A1(n9847), .A2(n9845), .ZN(n9844) );
  INV_X1 U11249 ( .A(n13987), .ZN(n10812) );
  OR2_X1 U11250 ( .A1(n10738), .A2(n15136), .ZN(n16164) );
  CLKBUF_X1 U11251 ( .A(n10880), .Z(n10890) );
  NAND2_X1 U11252 ( .A1(n18044), .A2(n12997), .ZN(n17941) );
  OR2_X1 U11253 ( .A1(n10887), .A2(n10886), .ZN(n10901) );
  NAND2_X1 U11254 ( .A1(n13882), .A2(n13843), .ZN(n13987) );
  NAND2_X1 U11255 ( .A1(n10861), .A2(n15631), .ZN(n15620) );
  NAND2_X1 U11256 ( .A1(n11586), .A2(n11585), .ZN(n13968) );
  AND2_X1 U11257 ( .A1(n11461), .A2(n14712), .ZN(n14879) );
  AND2_X1 U11258 ( .A1(n14723), .A2(n11456), .ZN(n11461) );
  INV_X1 U11259 ( .A(n14154), .ZN(n9842) );
  NAND2_X1 U11260 ( .A1(n10316), .A2(n10315), .ZN(n10887) );
  OR2_X1 U11261 ( .A1(n14748), .A2(n16088), .ZN(n14723) );
  AND2_X1 U11262 ( .A1(n13087), .A2(n13837), .ZN(n13880) );
  NAND2_X1 U11263 ( .A1(n10432), .A2(n10467), .ZN(n10387) );
  NOR2_X2 U11264 ( .A1(n13599), .A2(n13088), .ZN(n13087) );
  NOR2_X1 U11265 ( .A1(n9825), .A2(n9824), .ZN(n14411) );
  XNOR2_X1 U11266 ( .A(n11435), .B(n11434), .ZN(n11584) );
  AND2_X1 U11267 ( .A1(n13574), .A2(n13405), .ZN(n13670) );
  NAND2_X1 U11268 ( .A1(n11361), .A2(n11360), .ZN(n11435) );
  AND2_X1 U11269 ( .A1(n10309), .A2(n10308), .ZN(n10315) );
  AND2_X1 U11270 ( .A1(n9755), .A2(n12347), .ZN(n14987) );
  OR2_X1 U11271 ( .A1(n10329), .A2(n10328), .ZN(n10341) );
  NOR2_X1 U11272 ( .A1(n19335), .A2(n19797), .ZN(n19326) );
  NAND2_X1 U11273 ( .A1(n9754), .A2(n9684), .ZN(n9755) );
  NAND2_X1 U11274 ( .A1(n9761), .A2(n11556), .ZN(n13587) );
  AND2_X1 U11275 ( .A1(n14508), .A2(n9826), .ZN(n14831) );
  NAND2_X1 U11276 ( .A1(n11342), .A2(n11341), .ZN(n11418) );
  AND2_X1 U11277 ( .A1(n13396), .A2(n12446), .ZN(n14049) );
  NOR2_X2 U11278 ( .A1(n14509), .A2(n14510), .ZN(n14508) );
  XNOR2_X1 U11279 ( .A(n11407), .B(n11403), .ZN(n11565) );
  AND2_X1 U11280 ( .A1(n15509), .A2(n15510), .ZN(n15512) );
  CLKBUF_X1 U11281 ( .A(n13704), .Z(n20034) );
  INV_X1 U11282 ( .A(n18096), .ZN(n16410) );
  INV_X1 U11283 ( .A(n10184), .ZN(n19593) );
  INV_X1 U11284 ( .A(n19632), .ZN(n19636) );
  NAND2_X1 U11285 ( .A1(n10760), .A2(n10759), .ZN(n13399) );
  CLKBUF_X1 U11286 ( .A(n14317), .Z(n14604) );
  AND2_X1 U11287 ( .A1(n15641), .A2(n19058), .ZN(n10130) );
  AND2_X1 U11288 ( .A1(n15665), .A2(n19058), .ZN(n10118) );
  INV_X2 U11289 ( .A(n15902), .ZN(n13739) );
  INV_X1 U11290 ( .A(n15665), .ZN(n15641) );
  NAND2_X1 U11291 ( .A1(n10099), .A2(n10091), .ZN(n15665) );
  NAND2_X1 U11292 ( .A1(n13334), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13333) );
  NOR2_X2 U11293 ( .A1(n19204), .A2(n19563), .ZN(n19205) );
  NOR2_X2 U11294 ( .A1(n19209), .A2(n19563), .ZN(n19210) );
  NAND2_X1 U11295 ( .A1(n12989), .A2(n17830), .ZN(n17824) );
  NOR2_X2 U11296 ( .A1(n19128), .A2(n19563), .ZN(n15716) );
  NOR2_X2 U11297 ( .A1(n19121), .A2(n19563), .ZN(n15706) );
  NOR2_X1 U11298 ( .A1(n14546), .A2(n14129), .ZN(n14528) );
  INV_X2 U11299 ( .A(n15123), .ZN(n13579) );
  OAI21_X1 U11300 ( .B1(n11536), .B2(n11409), .A(n11377), .ZN(n13334) );
  AOI221_X1 U11301 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16379), .C1(n19840), .C2(
        n16379), .A(n19634), .ZN(n19834) );
  AND2_X1 U11302 ( .A1(n11247), .A2(n11374), .ZN(n11278) );
  INV_X1 U11303 ( .A(n13400), .ZN(n10759) );
  OAI21_X1 U11304 ( .B1(n12329), .B2(n18936), .A(n18933), .ZN(n18917) );
  NAND2_X1 U11305 ( .A1(n12347), .A2(n12346), .ZN(n18933) );
  AND2_X2 U11306 ( .A1(n17457), .A2(n17490), .ZN(n17488) );
  NAND2_X1 U11307 ( .A1(n10095), .A2(n10094), .ZN(n10100) );
  AND2_X1 U11308 ( .A1(n11195), .A2(n11193), .ZN(n11271) );
  NOR2_X1 U11309 ( .A1(n10582), .A2(n9853), .ZN(n9856) );
  NAND2_X1 U11310 ( .A1(n10084), .A2(n10083), .ZN(n10751) );
  OR2_X1 U11311 ( .A1(n10369), .A2(n10477), .ZN(n10467) );
  INV_X2 U11312 ( .A(n20780), .ZN(n17258) );
  NAND2_X1 U11313 ( .A1(n10069), .A2(n10068), .ZN(n10087) );
  AOI21_X1 U11314 ( .B1(n10051), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10050), .ZN(n10058) );
  NAND2_X1 U11315 ( .A1(n9776), .A2(n10039), .ZN(n10042) );
  OR2_X1 U11316 ( .A1(n9834), .A2(n13869), .ZN(n9831) );
  NOR2_X2 U11317 ( .A1(n16578), .A2(n17584), .ZN(n17548) );
  NAND2_X1 U11318 ( .A1(n17881), .A2(n12773), .ZN(n12776) );
  NAND2_X1 U11319 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17583), .ZN(
        n16578) );
  OAI22_X1 U11320 ( .A1(n11504), .A2(n11503), .B1(n11513), .B2(n11505), .ZN(
        n9697) );
  NAND2_X1 U11321 ( .A1(n10561), .A2(n9849), .ZN(n13235) );
  NAND2_X1 U11322 ( .A1(n10743), .A2(n10925), .ZN(n13783) );
  AND2_X1 U11323 ( .A1(n12316), .A2(n12134), .ZN(n12314) );
  CLKBUF_X1 U11324 ( .A(n13243), .Z(n13815) );
  OR2_X1 U11325 ( .A1(n10070), .A2(n10052), .ZN(n10054) );
  NAND2_X1 U11327 ( .A1(n9732), .A2(n9730), .ZN(n10744) );
  NAND2_X1 U11328 ( .A1(n13244), .A2(n12174), .ZN(n12279) );
  AND2_X1 U11329 ( .A1(n11498), .A2(n13265), .ZN(n11512) );
  NAND2_X1 U11330 ( .A1(n12156), .A2(n11495), .ZN(n13353) );
  NOR2_X1 U11331 ( .A1(n17900), .A2(n17432), .ZN(n12976) );
  NOR2_X1 U11332 ( .A1(n17417), .A2(n12775), .ZN(n12778) );
  OR2_X1 U11333 ( .A1(n12176), .A2(n11136), .ZN(n13522) );
  INV_X2 U11334 ( .A(n11960), .ZN(n12161) );
  AND2_X1 U11335 ( .A1(n13817), .A2(n9760), .ZN(n11132) );
  NAND2_X2 U11336 ( .A1(n12175), .A2(n20037), .ZN(n12189) );
  AND2_X1 U11338 ( .A1(n9965), .A2(n15717), .ZN(n10925) );
  NAND2_X1 U11339 ( .A1(n10018), .A2(n10019), .ZN(n9732) );
  NAND2_X1 U11340 ( .A1(n11237), .A2(n11236), .ZN(n11375) );
  OR2_X1 U11341 ( .A1(n10204), .A2(n10203), .ZN(n10239) );
  INV_X1 U11342 ( .A(n13506), .ZN(n20059) );
  INV_X1 U11343 ( .A(n11108), .ZN(n11114) );
  INV_X4 U11344 ( .A(n10560), .ZN(n10477) );
  OR2_X1 U11345 ( .A1(n10166), .A2(n10165), .ZN(n10569) );
  BUF_X2 U11346 ( .A(n10559), .Z(n19849) );
  INV_X1 U11347 ( .A(n10559), .ZN(n10022) );
  NAND4_X1 U11348 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n12173) );
  NAND2_X2 U11349 ( .A1(n10008), .A2(n10007), .ZN(n15717) );
  NAND2_X2 U11350 ( .A1(n9937), .A2(n9936), .ZN(n19224) );
  INV_X1 U11351 ( .A(n10194), .ZN(n9628) );
  AND4_X1 U11352 ( .A1(n11009), .A2(n11008), .A3(n11007), .A4(n11006), .ZN(
        n11019) );
  AND4_X1 U11353 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(
        n10977) );
  AND4_X1 U11354 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10998) );
  AND4_X1 U11355 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11081) );
  NOR2_X1 U11356 ( .A1(n11094), .A2(n11093), .ZN(n11105) );
  AND4_X1 U11357 ( .A1(n11121), .A2(n11120), .A3(n11119), .A4(n11118), .ZN(
        n11131) );
  AND4_X1 U11358 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11057) );
  NAND2_X1 U11359 ( .A1(n10000), .A2(n9999), .ZN(n10008) );
  NAND3_X1 U11360 ( .A1(n9920), .A2(n9919), .A3(n9918), .ZN(n9921) );
  AND4_X1 U11361 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n11104) );
  INV_X2 U11362 ( .A(U214), .ZN(n16486) );
  AND4_X1 U11363 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11103) );
  AND4_X1 U11364 ( .A1(n11075), .A2(n11074), .A3(n11073), .A4(n11072), .ZN(
        n11080) );
  AND4_X1 U11365 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10997) );
  AND4_X1 U11366 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11056) );
  OR2_X1 U11367 ( .A1(n11775), .A2(n10978), .ZN(n10980) );
  INV_X2 U11368 ( .A(n20742), .ZN(n13766) );
  INV_X2 U11369 ( .A(n15808), .ZN(n17214) );
  AND4_X1 U11370 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  AND2_X1 U11371 ( .A1(n9912), .A2(n9911), .ZN(n9913) );
  AND4_X1 U11372 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10000)
         );
  NAND2_X2 U11373 ( .A1(n18822), .A2(n18756), .ZN(n18803) );
  INV_X2 U11374 ( .A(n16527), .ZN(U215) );
  NOR2_X1 U11375 ( .A1(n17845), .A2(n17844), .ZN(n17819) );
  NAND2_X1 U11376 ( .A1(n9616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10194) );
  NAND2_X2 U11377 ( .A1(n19867), .A2(n19742), .ZN(n19784) );
  AND2_X1 U11378 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n9806) );
  INV_X1 U11379 ( .A(n15808), .ZN(n9599) );
  INV_X1 U11380 ( .A(n11021), .ZN(n9624) );
  INV_X2 U11381 ( .A(n17457), .ZN(n9600) );
  OR2_X1 U11382 ( .A1(n11021), .A2(n11084), .ZN(n11085) );
  OR2_X1 U11384 ( .A1(n11979), .A2(n11122), .ZN(n11123) );
  INV_X2 U11385 ( .A(n16531), .ZN(n16533) );
  INV_X1 U11386 ( .A(n12677), .ZN(n18663) );
  OR2_X1 U11387 ( .A1(n12687), .A2(n12685), .ZN(n15797) );
  AND2_X2 U11388 ( .A1(n10970), .A2(n10969), .ZN(n9636) );
  NOR2_X1 U11389 ( .A1(n15834), .A2(n12689), .ZN(n12726) );
  AND2_X2 U11390 ( .A1(n13694), .A2(n13680), .ZN(n11172) );
  AND2_X1 U11391 ( .A1(n9896), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10145) );
  NAND2_X1 U11392 ( .A1(n9714), .A2(n18674), .ZN(n12688) );
  NAND2_X1 U11393 ( .A1(n18674), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12683) );
  NAND2_X1 U11394 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18675) );
  NAND2_X1 U11395 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15834) );
  INV_X1 U11396 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9714) );
  INV_X1 U11397 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18674) );
  NAND2_X1 U11398 ( .A1(n15622), .A2(n9778), .ZN(n15626) );
  NAND2_X1 U11399 ( .A1(n13941), .A2(n15630), .ZN(n15622) );
  NOR2_X1 U11400 ( .A1(n17909), .A2(n15892), .ZN(n9602) );
  NOR2_X1 U11401 ( .A1(n17909), .A2(n15892), .ZN(n16405) );
  AND2_X1 U11402 ( .A1(n11273), .A2(n11272), .ZN(n9603) );
  INV_X1 U11404 ( .A(n10028), .ZN(n13192) );
  AOI22_X1 U11405 ( .A1(n15676), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16369), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10025) );
  AND3_X1 U11406 ( .A1(n11108), .A2(n11486), .A3(n13512), .ZN(n13259) );
  AOI21_X1 U11407 ( .B1(n20078), .B2(n11486), .A(n14389), .ZN(n11151) );
  NAND2_X1 U11408 ( .A1(n15078), .A2(n9605), .ZN(n15064) );
  AND2_X1 U11409 ( .A1(n15077), .A2(n14973), .ZN(n9605) );
  NOR2_X2 U11411 ( .A1(n14398), .A2(n14399), .ZN(n14401) );
  INV_X1 U11412 ( .A(n9777), .ZN(n13238) );
  NAND2_X1 U11413 ( .A1(n13597), .A2(n13598), .ZN(n13599) );
  NOR2_X2 U11414 ( .A1(n14472), .A2(n14212), .ZN(n14211) );
  NAND2_X1 U11415 ( .A1(n15356), .A2(n15355), .ZN(n9607) );
  NAND2_X2 U11416 ( .A1(n10314), .A2(n10313), .ZN(n15356) );
  NAND4_X4 U11417 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11115) );
  INV_X1 U11418 ( .A(n9967), .ZN(n9608) );
  INV_X1 U11419 ( .A(n9967), .ZN(n10009) );
  OR2_X1 U11420 ( .A1(n19230), .A2(n9967), .ZN(n9948) );
  AND2_X1 U11421 ( .A1(n13574), .A2(n9609), .ZN(n13597) );
  AND2_X1 U11422 ( .A1(n13405), .A2(n10790), .ZN(n9609) );
  AND2_X1 U11423 ( .A1(n13880), .A2(n13879), .ZN(n13882) );
  NAND2_X1 U11424 ( .A1(n15020), .A2(n15019), .ZN(n15008) );
  NAND2_X1 U11425 ( .A1(n15063), .A2(n10851), .ZN(n14258) );
  NOR2_X2 U11426 ( .A1(n14439), .A2(n12299), .ZN(n15938) );
  NOR2_X2 U11427 ( .A1(n19940), .A2(n20661), .ZN(n19927) );
  NOR2_X2 U11428 ( .A1(n19917), .A2(n12159), .ZN(n19899) );
  NAND2_X1 U11429 ( .A1(n15575), .A2(n15493), .ZN(n14193) );
  AND2_X1 U11430 ( .A1(n15575), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15574) );
  AND2_X2 U11431 ( .A1(n15575), .A2(n9692), .ZN(n15226) );
  OR2_X2 U11432 ( .A1(n10208), .A2(n10209), .ZN(n10874) );
  INV_X1 U11433 ( .A(n14677), .ZN(n9610) );
  CLKBUF_X1 U11434 ( .A(n14118), .Z(n9611) );
  CLKBUF_X1 U11435 ( .A(n13998), .Z(n9612) );
  CLKBUF_X1 U11436 ( .A(n19977), .Z(n9613) );
  NAND2_X1 U11438 ( .A1(n19230), .A2(n19224), .ZN(n9777) );
  NOR2_X1 U11439 ( .A1(n9777), .A2(n10009), .ZN(n10011) );
  AND2_X1 U11440 ( .A1(n11115), .A2(n11107), .ZN(n9835) );
  NOR2_X1 U11441 ( .A1(n9626), .A2(n12007), .ZN(n11004) );
  NAND2_X2 U11442 ( .A1(n13511), .A2(n13514), .ZN(n11144) );
  NAND2_X1 U11443 ( .A1(n11273), .A2(n11272), .ZN(n20093) );
  NAND2_X1 U11444 ( .A1(n13251), .A2(n12157), .ZN(n11142) );
  INV_X1 U11445 ( .A(n11126), .ZN(n12064) );
  AND2_X1 U11446 ( .A1(n10927), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9615) );
  AND2_X1 U11447 ( .A1(n10145), .A2(n13794), .ZN(n9616) );
  INV_X2 U11448 ( .A(n9923), .ZN(n9618) );
  NAND2_X1 U11449 ( .A1(n9922), .A2(n9921), .ZN(n9619) );
  NAND4_X1 U11450 ( .A1(n9848), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n9759), .A4(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11775) );
  AND2_X1 U11451 ( .A1(n10969), .A2(n10968), .ZN(n9620) );
  AND2_X2 U11452 ( .A1(n10969), .A2(n10968), .ZN(n9621) );
  AND2_X2 U11453 ( .A1(n10969), .A2(n10968), .ZN(n12098) );
  AND2_X1 U11454 ( .A1(n10970), .A2(n10969), .ZN(n9622) );
  AND2_X1 U11455 ( .A1(n10970), .A2(n10969), .ZN(n11641) );
  AND3_X2 U11456 ( .A1(n9782), .A2(n15659), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9623) );
  INV_X1 U11457 ( .A(n11126), .ZN(n9626) );
  AND2_X4 U11458 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U11459 ( .A1(n20161), .A2(n11271), .ZN(n11274) );
  OR2_X1 U11460 ( .A1(n13333), .A2(n11379), .ZN(n11380) );
  OAI21_X2 U11461 ( .B1(n15263), .B2(n14173), .A(n15332), .ZN(n16201) );
  NOR2_X1 U11462 ( .A1(n12688), .A2(n16932), .ZN(n12684) );
  NOR2_X2 U11463 ( .A1(n15554), .A2(n15564), .ZN(n15335) );
  NAND2_X2 U11464 ( .A1(n13193), .A2(n9627), .ZN(n10511) );
  INV_X1 U11465 ( .A(n19203), .ZN(n9779) );
  INV_X1 U11467 ( .A(n10194), .ZN(n9630) );
  NOR2_X2 U11468 ( .A1(n16218), .A2(n16221), .ZN(n15557) );
  XNOR2_X1 U11469 ( .A(n11531), .B(n11277), .ZN(n13703) );
  NAND2_X1 U11470 ( .A1(n9837), .A2(n9836), .ZN(n11536) );
  NAND2_X1 U11471 ( .A1(n10101), .A2(n10100), .ZN(n19058) );
  AND2_X1 U11472 ( .A1(n20054), .A2(n12173), .ZN(n12174) );
  NAND2_X2 U11473 ( .A1(n13491), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13492) );
  XNOR2_X2 U11474 ( .A(n11378), .B(n13333), .ZN(n13491) );
  AOI211_X2 U11475 ( .C1(n15197), .C2(n15365), .A(n15198), .B(n10476), .ZN(
        n15189) );
  NOR2_X4 U11476 ( .A1(n15009), .A2(n14995), .ZN(n15078) );
  AOI21_X2 U11477 ( .B1(n15298), .B2(n14182), .A(n14181), .ZN(n14223) );
  OAI21_X2 U11478 ( .B1(n15305), .B2(n15306), .A(n14179), .ZN(n15298) );
  NAND4_X1 U11480 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11107) );
  OAI21_X1 U11481 ( .B1(n11165), .B2(n9848), .A(n11148), .ZN(n11195) );
  NOR2_X2 U11482 ( .A1(n13985), .A2(n10824), .ZN(n13058) );
  INV_X1 U11483 ( .A(n20914), .ZN(n9638) );
  NOR2_X2 U11484 ( .A1(n10033), .A2(n10032), .ZN(n10743) );
  NOR2_X4 U11485 ( .A1(n13968), .A2(n13969), .ZN(n13967) );
  NOR2_X1 U11486 ( .A1(n10559), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10563) );
  AND2_X1 U11487 ( .A1(n11404), .A2(n11403), .ZN(n11341) );
  NOR2_X1 U11488 ( .A1(n18239), .A2(n17232), .ZN(n12924) );
  OAI21_X1 U11489 ( .B1(n10239), .B2(n12350), .A(n10238), .ZN(n10498) );
  AND2_X1 U11490 ( .A1(n12444), .A2(n13847), .ZN(n13989) );
  NAND2_X1 U11491 ( .A1(n9738), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9737) );
  NOR2_X1 U11492 ( .A1(n15350), .A2(n9739), .ZN(n9738) );
  INV_X1 U11493 ( .A(n15541), .ZN(n9862) );
  AND3_X1 U11494 ( .A1(n10592), .A2(n10591), .A3(n10590), .ZN(n13423) );
  INV_X1 U11495 ( .A(n9648), .ZN(n9855) );
  OAI211_X1 U11496 ( .C1(n10014), .C2(n10013), .A(n10012), .B(n9627), .ZN(
        n10923) );
  NAND2_X1 U11497 ( .A1(n9949), .A2(n9948), .ZN(n10013) );
  NAND2_X1 U11498 ( .A1(n9703), .A2(n10018), .ZN(n12352) );
  AND2_X1 U11499 ( .A1(n10019), .A2(n19203), .ZN(n9703) );
  AND2_X1 U11500 ( .A1(n16345), .A2(n19849), .ZN(n13200) );
  NAND2_X1 U11501 ( .A1(n12927), .A2(n16537), .ZN(n16560) );
  NOR2_X1 U11502 ( .A1(n16412), .A2(n17732), .ZN(n12804) );
  OAI21_X1 U11503 ( .B1(n17723), .B2(n12795), .A(n12810), .ZN(n12807) );
  NOR2_X1 U11504 ( .A1(n12931), .A2(n17232), .ZN(n12950) );
  OR2_X1 U11505 ( .A1(n18665), .A2(n12966), .ZN(n12952) );
  NAND2_X1 U11506 ( .A1(n13499), .A2(n9702), .ZN(n13462) );
  AND2_X1 U11507 ( .A1(n12155), .A2(n13501), .ZN(n9702) );
  NAND2_X1 U11508 ( .A1(n14471), .A2(n14473), .ZN(n14472) );
  NAND2_X1 U11509 ( .A1(n13509), .A2(n13508), .ZN(n13524) );
  INV_X1 U11510 ( .A(n9632), .ZN(n20491) );
  NOR2_X1 U11511 ( .A1(n14066), .A2(n15112), .ZN(n15111) );
  AOI21_X1 U11512 ( .B1(n15665), .B2(n12394), .A(n12389), .ZN(n13247) );
  INV_X1 U11513 ( .A(n18264), .ZN(n17272) );
  INV_X1 U11514 ( .A(n18877), .ZN(n18248) );
  INV_X1 U11515 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11805) );
  INV_X1 U11516 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11894) );
  AND4_X1 U11517 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10227) );
  NAND2_X1 U11518 ( .A1(n11507), .A2(n9640), .ZN(n9696) );
  NAND2_X1 U11519 ( .A1(n10508), .A2(n9967), .ZN(n10518) );
  OR2_X1 U11520 ( .A1(n10265), .A2(n10264), .ZN(n10589) );
  INV_X1 U11521 ( .A(n15099), .ZN(n9795) );
  INV_X1 U11522 ( .A(n9732), .ZN(n9704) );
  AND2_X1 U11523 ( .A1(n9717), .A2(n9716), .ZN(n10192) );
  NAND2_X1 U11524 ( .A1(n19306), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n9716) );
  NAND2_X1 U11525 ( .A1(n10117), .A2(n10116), .ZN(n10123) );
  AND3_X1 U11526 ( .A1(n9917), .A2(n9916), .A3(n9956), .ZN(n9920) );
  OAI211_X1 U11528 ( .C1(n11546), .C2(n9763), .A(n9762), .B(n13587), .ZN(
        n13586) );
  OR2_X1 U11529 ( .A1(n11545), .A2(n9763), .ZN(n9762) );
  INV_X1 U11530 ( .A(n11547), .ZN(n9763) );
  AND2_X1 U11531 ( .A1(n11734), .A2(n11547), .ZN(n9766) );
  OR2_X1 U11532 ( .A1(n14748), .A2(n11460), .ZN(n14721) );
  INV_X1 U11533 ( .A(n13796), .ZN(n9834) );
  INV_X1 U11534 ( .A(n11417), .ZN(n11360) );
  INV_X1 U11535 ( .A(n11418), .ZN(n11361) );
  AND4_X1 U11536 ( .A1(n11235), .A2(n11234), .A3(n11233), .A4(n11232), .ZN(
        n11236) );
  INV_X1 U11537 ( .A(n11498), .ZN(n11519) );
  OR2_X1 U11538 ( .A1(n13374), .A2(n13500), .ZN(n13384) );
  OAI21_X1 U11539 ( .B1(n20745), .B2(n16147), .A(n15880), .ZN(n20036) );
  OR2_X1 U11540 ( .A1(n12329), .A2(n12322), .ZN(n9753) );
  NAND2_X1 U11541 ( .A1(n10404), .A2(n10382), .ZN(n10414) );
  AND2_X1 U11543 ( .A1(n10477), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U11544 ( .A1(n9792), .A2(n9664), .ZN(n9791) );
  NOR2_X1 U11545 ( .A1(n10566), .A2(n19716), .ZN(n12377) );
  AND2_X1 U11546 ( .A1(n12443), .A2(n13531), .ZN(n13847) );
  NAND2_X1 U11547 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U11548 ( .A1(n9881), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9747) );
  NAND2_X1 U11549 ( .A1(n10766), .A2(n10765), .ZN(n13480) );
  INV_X1 U11550 ( .A(n13481), .ZN(n10765) );
  INV_X1 U11551 ( .A(n13399), .ZN(n10766) );
  NAND2_X1 U11552 ( .A1(n15223), .A2(n15225), .ZN(n10472) );
  OR2_X1 U11553 ( .A1(n15546), .A2(n10445), .ZN(n14171) );
  INV_X1 U11554 ( .A(n14051), .ZN(n9865) );
  AND2_X1 U11555 ( .A1(n9644), .A2(n9860), .ZN(n9859) );
  INV_X1 U11556 ( .A(n13958), .ZN(n9860) );
  INV_X1 U11557 ( .A(n15540), .ZN(n9861) );
  INV_X1 U11558 ( .A(n13411), .ZN(n9868) );
  INV_X1 U11559 ( .A(n13451), .ZN(n9722) );
  AOI21_X1 U11560 ( .B1(n14320), .B2(n13451), .A(n13806), .ZN(n9728) );
  AND2_X1 U11561 ( .A1(n13801), .A2(n9725), .ZN(n9724) );
  NAND2_X1 U11562 ( .A1(n9726), .A2(n14320), .ZN(n9725) );
  OR2_X1 U11563 ( .A1(n10152), .A2(n10151), .ZN(n9851) );
  NAND2_X1 U11564 ( .A1(n16339), .A2(n9731), .ZN(n9730) );
  AND2_X1 U11565 ( .A1(n19849), .A2(n15717), .ZN(n9731) );
  AND2_X1 U11566 ( .A1(n12606), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12399) );
  AND2_X1 U11567 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n9951) );
  INV_X1 U11568 ( .A(n10539), .ZN(n10545) );
  NOR2_X1 U11569 ( .A1(n12685), .A2(n12688), .ZN(n12716) );
  NOR2_X1 U11570 ( .A1(n17409), .A2(n12780), .ZN(n12785) );
  NOR2_X1 U11571 ( .A1(n17689), .A2(n17631), .ZN(n17636) );
  XNOR2_X1 U11572 ( .A(n17432), .B(n17421), .ZN(n12772) );
  NAND2_X1 U11573 ( .A1(n12923), .A2(n12924), .ZN(n12932) );
  NAND3_X1 U11574 ( .A1(n17494), .A2(n16560), .A3(n12925), .ZN(n15825) );
  NOR2_X1 U11575 ( .A1(n12926), .A2(n18662), .ZN(n15741) );
  INV_X1 U11576 ( .A(n12950), .ZN(n12926) );
  NOR2_X1 U11577 ( .A1(n18665), .A2(n12930), .ZN(n15826) );
  NAND2_X1 U11578 ( .A1(n11287), .A2(n11286), .ZN(n20197) );
  INV_X1 U11579 ( .A(n14213), .ZN(n9824) );
  AND2_X1 U11580 ( .A1(n12224), .A2(n9874), .ZN(n14551) );
  OR2_X1 U11581 ( .A1(n13384), .A2(n13499), .ZN(n13728) );
  NAND2_X1 U11582 ( .A1(n13350), .A2(n13349), .ZN(n13359) );
  INV_X1 U11583 ( .A(n13772), .ZN(n13463) );
  AND2_X1 U11584 ( .A1(n20638), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12160) );
  NOR2_X2 U11585 ( .A1(n14395), .A2(n14397), .ZN(n14396) );
  AND2_X1 U11586 ( .A1(n11976), .A2(n14419), .ZN(n11977) );
  NOR2_X1 U11587 ( .A1(n11714), .A2(n14740), .ZN(n11719) );
  NOR2_X1 U11588 ( .A1(n11698), .A2(n9768), .ZN(n9767) );
  AND2_X1 U11589 ( .A1(n14136), .A2(n14554), .ZN(n9768) );
  INV_X1 U11590 ( .A(n11601), .ZN(n11605) );
  NAND2_X1 U11591 ( .A1(n11546), .A2(n11545), .ZN(n13558) );
  AND2_X1 U11592 ( .A1(n13499), .A2(n13501), .ZN(n13507) );
  AND2_X1 U11593 ( .A1(n20724), .A2(n20635), .ZN(n12119) );
  NAND2_X1 U11594 ( .A1(n13524), .A2(n13519), .ZN(n20018) );
  NAND2_X1 U11595 ( .A1(n12152), .A2(n12153), .ZN(n14311) );
  AND2_X1 U11596 ( .A1(n9631), .A2(n20491), .ZN(n20409) );
  INV_X1 U11598 ( .A(n10751), .ZN(n10085) );
  XNOR2_X1 U11599 ( .A(n12586), .B(n9889), .ZN(n15088) );
  OR2_X1 U11600 ( .A1(n15088), .A2(n15087), .ZN(n9792) );
  NOR2_X1 U11601 ( .A1(n15107), .A2(n15106), .ZN(n15105) );
  AND2_X1 U11602 ( .A1(n9798), .A2(n12477), .ZN(n9797) );
  AND3_X1 U11603 ( .A1(n10667), .A2(n10666), .A3(n10665), .ZN(n15541) );
  AND2_X1 U11604 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  XNOR2_X1 U11605 ( .A(n9743), .B(n9742), .ZN(n14372) );
  NAND2_X1 U11606 ( .A1(n12314), .A2(n9651), .ZN(n9743) );
  NOR2_X1 U11607 ( .A1(n9737), .A2(n16235), .ZN(n9736) );
  INV_X1 U11608 ( .A(n13988), .ZN(n10811) );
  NAND2_X1 U11609 ( .A1(n10347), .A2(n9641), .ZN(n9729) );
  NAND2_X1 U11610 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  INV_X1 U11611 ( .A(n13423), .ZN(n9854) );
  INV_X1 U11612 ( .A(n13810), .ZN(n10862) );
  AND2_X1 U11613 ( .A1(n10555), .A2(n19721), .ZN(n10936) );
  AOI21_X1 U11614 ( .B1(n13248), .B2(n13247), .A(n12392), .ZN(n13339) );
  NAND2_X1 U11615 ( .A1(n9789), .A2(n9787), .ZN(n13338) );
  NOR2_X1 U11616 ( .A1(n12399), .A2(n9788), .ZN(n9787) );
  INV_X1 U11617 ( .A(n12398), .ZN(n9788) );
  OR2_X1 U11618 ( .A1(n19810), .A2(n19820), .ZN(n19471) );
  NAND2_X1 U11619 ( .A1(n15692), .A2(n15691), .ZN(n15693) );
  NAND2_X1 U11620 ( .A1(n19810), .A2(n19817), .ZN(n19596) );
  NAND2_X1 U11621 ( .A1(n9979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9780) );
  NAND2_X1 U11622 ( .A1(n9980), .A2(n9999), .ZN(n9781) );
  NAND2_X1 U11623 ( .A1(n15727), .A2(n19827), .ZN(n19562) );
  NAND2_X1 U11624 ( .A1(n15727), .A2(n19063), .ZN(n19592) );
  INV_X1 U11625 ( .A(n19634), .ZN(n19563) );
  NOR2_X1 U11626 ( .A1(n18877), .A2(n18239), .ZN(n12927) );
  NAND2_X1 U11627 ( .A1(n17494), .A2(n12952), .ZN(n16537) );
  INV_X1 U11628 ( .A(n12791), .ZN(n12789) );
  NOR2_X1 U11629 ( .A1(n18877), .A2(n16544), .ZN(n13015) );
  NOR2_X1 U11630 ( .A1(n17605), .A2(n12808), .ZN(n17599) );
  NAND2_X1 U11631 ( .A1(n12807), .A2(n12806), .ZN(n17677) );
  NAND2_X1 U11632 ( .A1(n17810), .A2(n12798), .ZN(n17732) );
  XNOR2_X1 U11633 ( .A(n12782), .B(n12781), .ZN(n17848) );
  NAND2_X1 U11634 ( .A1(n12954), .A2(n18135), .ZN(n18684) );
  NOR2_X1 U11635 ( .A1(n14765), .A2(n19948), .ZN(n9698) );
  OR2_X1 U11636 ( .A1(n15913), .A2(n12304), .ZN(n14417) );
  NAND2_X1 U11637 ( .A1(n14876), .A2(n19936), .ZN(n9772) );
  AOI21_X1 U11638 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n12298), .A(n19905), 
        .ZN(n15957) );
  NAND2_X1 U11639 ( .A1(n15979), .A2(n9885), .ZN(n15975) );
  INV_X1 U11640 ( .A(n19953), .ZN(n19919) );
  AND2_X1 U11641 ( .A1(n14357), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19953) );
  XNOR2_X1 U11642 ( .A(n14504), .B(n14501), .ZN(n15955) );
  INV_X1 U11643 ( .A(n14741), .ZN(n19974) );
  AND2_X1 U11644 ( .A1(n15865), .A2(n13507), .ZN(n19981) );
  NAND2_X1 U11645 ( .A1(n9818), .A2(n9816), .ZN(n14300) );
  NAND2_X1 U11646 ( .A1(n14401), .A2(n9817), .ZN(n9816) );
  XNOR2_X1 U11647 ( .A(n12288), .B(n14381), .ZN(n9817) );
  OR2_X1 U11648 ( .A1(n14822), .A2(n14283), .ZN(n14798) );
  AND2_X1 U11649 ( .A1(n13524), .A2(n13515), .ZN(n20021) );
  AOI21_X1 U11650 ( .B1(n9838), .B2(n9840), .A(n9666), .ZN(n9836) );
  INV_X1 U11651 ( .A(n11374), .ZN(n9840) );
  CLKBUF_X1 U11652 ( .A(n13851), .Z(n20449) );
  CLKBUF_X1 U11653 ( .A(n13370), .Z(n20448) );
  NOR2_X1 U11654 ( .A1(n9748), .A2(n12329), .ZN(n13068) );
  INV_X1 U11655 ( .A(n19198), .ZN(n19185) );
  INV_X1 U11656 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19833) );
  INV_X1 U11657 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19824) );
  NAND2_X1 U11658 ( .A1(n19810), .A2(n19820), .ZN(n19794) );
  INV_X1 U11659 ( .A(n19526), .ZN(n19517) );
  NAND2_X1 U11660 ( .A1(n17276), .A2(n9682), .ZN(n9711) );
  NAND2_X1 U11661 ( .A1(n17277), .A2(n9582), .ZN(n17276) );
  NAND2_X1 U11662 ( .A1(n17282), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17277) );
  NOR2_X1 U11663 ( .A1(n17438), .A2(n17286), .ZN(n17282) );
  NOR2_X1 U11664 ( .A1(n17398), .A2(n17268), .ZN(n17269) );
  NOR2_X2 U11665 ( .A1(n17402), .A2(n17904), .ZN(n17812) );
  XNOR2_X1 U11666 ( .A(n17565), .B(n12810), .ZN(n17919) );
  OAI221_X2 U11667 ( .B1(n12967), .B2(n12966), .C1(n12967), .C2(n12965), .A(
        n18873), .ZN(n18182) );
  NAND2_X1 U11668 ( .A1(n18877), .A2(n18135), .ZN(n18201) );
  NOR2_X1 U11669 ( .A1(n11494), .A2(n11493), .ZN(n11504) );
  AOI211_X1 U11670 ( .C1(n13346), .C2(n20037), .A(n11507), .B(n11491), .ZN(
        n11494) );
  INV_X1 U11671 ( .A(n11172), .ZN(n12085) );
  AND4_X1 U11672 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11217) );
  NAND2_X1 U11673 ( .A1(n20037), .A2(n20059), .ZN(n9760) );
  INV_X1 U11674 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10958) );
  OR2_X1 U11675 ( .A1(n12940), .A2(n12941), .ZN(n12936) );
  NAND2_X1 U11676 ( .A1(n20037), .A2(n11115), .ZN(n11288) );
  OR2_X1 U11677 ( .A1(n13681), .A2(n10971), .ZN(n10972) );
  OR2_X1 U11678 ( .A1(n11115), .A2(n20635), .ZN(n11267) );
  NAND2_X1 U11679 ( .A1(n12152), .A2(n11113), .ZN(n13376) );
  INV_X1 U11680 ( .A(n13266), .ZN(n11109) );
  INV_X1 U11681 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11092) );
  OAI211_X1 U11682 ( .C1(n11177), .C2(n11805), .A(n11086), .B(n11085), .ZN(
        n11087) );
  NAND2_X1 U11683 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11086) );
  INV_X1 U11684 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12007) );
  NOR2_X1 U11685 ( .A1(n10984), .A2(n10983), .ZN(n10999) );
  NAND2_X1 U11686 ( .A1(n10009), .A2(n10556), .ZN(n10512) );
  CLKBUF_X1 U11687 ( .A(n9930), .Z(n12636) );
  INV_X1 U11688 ( .A(n19224), .ZN(n12376) );
  NAND2_X1 U11689 ( .A1(n10855), .A2(n9646), .ZN(n9776) );
  AND4_X1 U11690 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10225) );
  AOI22_X1 U11691 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19366), .B1(
        n10281), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10187) );
  NOR2_X1 U11692 ( .A1(n12350), .A2(n19716), .ZN(n10059) );
  NAND2_X1 U11693 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12933), .ZN(
        n12685) );
  AOI21_X1 U11694 ( .B1(n20892), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12934), .ZN(n12941) );
  AND2_X1 U11695 ( .A1(n12957), .A2(n12956), .ZN(n12934) );
  NAND2_X1 U11696 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12935), .ZN(
        n12687) );
  AND2_X1 U11697 ( .A1(n11288), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11502) );
  AND2_X1 U11698 ( .A1(n11484), .A2(n11483), .ZN(n12150) );
  OR2_X1 U11699 ( .A1(n11485), .A2(n11482), .ZN(n11484) );
  AOI21_X1 U11700 ( .B1(n9695), .B2(n11517), .A(n11516), .ZN(n11518) );
  AND2_X1 U11701 ( .A1(n11964), .A2(n14432), .ZN(n14420) );
  NAND2_X1 U11702 ( .A1(n13967), .A2(n9650), .ZN(n14137) );
  AND2_X1 U11703 ( .A1(n11621), .A2(n14034), .ZN(n9769) );
  INV_X1 U11704 ( .A(n14019), .ZN(n11621) );
  AND2_X1 U11705 ( .A1(n11190), .A2(n11189), .ZN(n11392) );
  NAND2_X1 U11706 ( .A1(n14833), .A2(n9820), .ZN(n9825) );
  NOR2_X1 U11707 ( .A1(n9821), .A2(n14474), .ZN(n9820) );
  INV_X1 U11708 ( .A(n9822), .ZN(n9821) );
  NOR2_X1 U11709 ( .A1(n14486), .A2(n9823), .ZN(n9822) );
  INV_X1 U11710 ( .A(n14423), .ZN(n9823) );
  OR2_X1 U11711 ( .A1(n11462), .A2(n14751), .ZN(n11463) );
  AND2_X1 U11712 ( .A1(n20054), .A2(n20073), .ZN(n13265) );
  NAND2_X1 U11713 ( .A1(n9633), .A2(n14380), .ZN(n12276) );
  AND2_X1 U11714 ( .A1(n20744), .A2(n13817), .ZN(n13255) );
  OR2_X1 U11715 ( .A1(n11266), .A2(n11265), .ZN(n11366) );
  NAND2_X1 U11716 ( .A1(n11274), .A2(n11164), .ZN(n11170) );
  OR2_X1 U11717 ( .A1(n12083), .A2(n11061), .ZN(n11062) );
  AND2_X1 U11718 ( .A1(n20634), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11525) );
  OR2_X1 U11719 ( .A1(n10178), .A2(n10177), .ZN(n10231) );
  INV_X1 U11720 ( .A(n10356), .ZN(n10353) );
  NOR2_X1 U11721 ( .A1(n10349), .A2(n10348), .ZN(n10359) );
  NAND2_X1 U11722 ( .A1(n10343), .A2(n10342), .ZN(n10349) );
  CLKBUF_X1 U11723 ( .A(n10343), .Z(n10310) );
  CLKBUF_X1 U11724 ( .A(n12649), .Z(n12659) );
  CLKBUF_X1 U11725 ( .A(n12490), .Z(n12654) );
  AOI21_X1 U11726 ( .B1(n12523), .B2(n9795), .A(n12547), .ZN(n9794) );
  AND2_X1 U11727 ( .A1(n14048), .A2(n15116), .ZN(n9798) );
  INV_X1 U11728 ( .A(n10231), .ZN(n10864) );
  AOI21_X1 U11729 ( .B1(n10807), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10071), .ZN(
        n10072) );
  NOR2_X1 U11730 ( .A1(n15202), .A2(n9673), .ZN(n9733) );
  NOR2_X1 U11731 ( .A1(n10907), .A2(n9785), .ZN(n9784) );
  OR2_X1 U11732 ( .A1(n15060), .A2(n10402), .ZN(n10447) );
  NAND2_X1 U11733 ( .A1(n15574), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15554) );
  OR2_X1 U11734 ( .A1(n13414), .A2(n10402), .ZN(n10363) );
  NAND2_X1 U11735 ( .A1(n10891), .A2(n10890), .ZN(n10895) );
  NAND2_X1 U11736 ( .A1(n10860), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15619) );
  NAND2_X1 U11737 ( .A1(n10874), .A2(n10875), .ZN(n9786) );
  NAND2_X1 U11738 ( .A1(n13811), .A2(n10873), .ZN(n10879) );
  NAND2_X1 U11739 ( .A1(n10245), .A2(n10251), .ZN(n10244) );
  NAND2_X1 U11740 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NAND2_X1 U11741 ( .A1(n10477), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10240) );
  AOI21_X1 U11742 ( .B1(n10807), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10056), .ZN(
        n10057) );
  NAND2_X1 U11743 ( .A1(n9851), .A2(n9850), .ZN(n9849) );
  OAI211_X1 U11744 ( .C1(n10566), .C2(n13790), .A(n10565), .B(n10564), .ZN(
        n13233) );
  NOR2_X1 U11745 ( .A1(n9884), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10564) );
  AND2_X1 U11746 ( .A1(n10509), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n9884) );
  INV_X1 U11747 ( .A(n16344), .ZN(n13183) );
  NAND2_X1 U11748 ( .A1(n10566), .A2(n10914), .ZN(n9705) );
  OR2_X1 U11749 ( .A1(n13397), .A2(n19213), .ZN(n12390) );
  NAND2_X1 U11751 ( .A1(n10022), .A2(n9779), .ZN(n10028) );
  NOR2_X1 U11752 ( .A1(n12379), .A2(n9595), .ZN(n10131) );
  AND2_X1 U11753 ( .A1(n10096), .A2(n10100), .ZN(n10124) );
  AND2_X1 U11754 ( .A1(n10105), .A2(n10104), .ZN(n10128) );
  AND2_X1 U11755 ( .A1(n12379), .A2(n9595), .ZN(n10119) );
  AOI22_X1 U11756 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n9933) );
  NAND3_X1 U11757 ( .A1(n19800), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19634), 
        .ZN(n15697) );
  INV_X1 U11758 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9782) );
  AND2_X1 U11759 ( .A1(n13108), .A2(n9706), .ZN(n10519) );
  INV_X1 U11760 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20867) );
  OR2_X1 U11761 ( .A1(n12687), .A2(n16932), .ZN(n12718) );
  INV_X1 U11762 ( .A(n12735), .ZN(n12882) );
  NOR2_X1 U11763 ( .A1(n12689), .A2(n12687), .ZN(n12871) );
  NAND2_X1 U11764 ( .A1(n17272), .A2(n12917), .ZN(n12922) );
  NAND2_X1 U11765 ( .A1(n12995), .A2(n17800), .ZN(n16411) );
  AND2_X1 U11766 ( .A1(n12929), .A2(n15909), .ZN(n12951) );
  INV_X1 U11767 ( .A(n12718), .ZN(n12905) );
  NAND2_X1 U11768 ( .A1(n20064), .A2(n20054), .ZN(n12176) );
  INV_X1 U11769 ( .A(n13353), .ZN(n13243) );
  NAND2_X1 U11770 ( .A1(n14128), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14446) );
  NAND2_X1 U11771 ( .A1(n19957), .A2(n12296), .ZN(n19940) );
  NAND2_X1 U11772 ( .A1(n12180), .A2(n12179), .ZN(n9815) );
  NOR2_X1 U11773 ( .A1(n13818), .A2(n12156), .ZN(n12293) );
  INV_X1 U11774 ( .A(n19957), .ZN(n14363) );
  OR3_X1 U11775 ( .A1(n20739), .A2(n19952), .A3(n12168), .ZN(n14357) );
  NOR2_X1 U11776 ( .A1(n14436), .A2(n9828), .ZN(n9826) );
  AND2_X1 U11777 ( .A1(n12216), .A2(n12215), .ZN(n13974) );
  OR3_X1 U11778 ( .A1(n13870), .A2(n9831), .A3(n9830), .ZN(n16106) );
  NAND2_X1 U11779 ( .A1(n13889), .A2(n9832), .ZN(n9830) );
  INV_X1 U11780 ( .A(n13974), .ZN(n9832) );
  OR3_X1 U11781 ( .A1(n13870), .A2(n9831), .A3(n9833), .ZN(n13975) );
  AND2_X1 U11782 ( .A1(n9814), .A2(n9815), .ZN(n13863) );
  NAND2_X1 U11783 ( .A1(n13517), .A2(n9633), .ZN(n9814) );
  INV_X1 U11784 ( .A(n20032), .ZN(n20030) );
  OR2_X1 U11785 ( .A1(n12051), .A2(n12050), .ZN(n12170) );
  AND2_X1 U11786 ( .A1(n11999), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12000) );
  AND2_X1 U11787 ( .A1(n11972), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U11788 ( .A1(n11839), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11998) );
  AND2_X1 U11789 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11838), .ZN(
        n11913) );
  INV_X1 U11790 ( .A(n11917), .ZN(n11838) );
  NAND2_X1 U11791 ( .A1(n11837), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11943) );
  AND2_X1 U11792 ( .A1(n11755), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11837) );
  NAND2_X1 U11793 ( .A1(n14515), .A2(n9775), .ZN(n9774) );
  INV_X1 U11794 ( .A(n14445), .ZN(n9775) );
  NOR2_X1 U11795 ( .A1(n11739), .A2(n15990), .ZN(n11755) );
  INV_X1 U11796 ( .A(n11694), .ZN(n11660) );
  AND2_X1 U11797 ( .A1(n11654), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11655) );
  NAND2_X1 U11798 ( .A1(n11655), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11694) );
  NOR2_X1 U11799 ( .A1(n11637), .A2(n14119), .ZN(n11654) );
  AND2_X1 U11800 ( .A1(n13967), .A2(n11621), .ZN(n14035) );
  NAND2_X1 U11801 ( .A1(n14751), .A2(n11447), .ZN(n13996) );
  AND3_X1 U11802 ( .A1(n11604), .A2(n11603), .A3(n11602), .ZN(n13969) );
  AOI21_X1 U11803 ( .B1(n11584), .B2(n11734), .A(n11583), .ZN(n13885) );
  INV_X1 U11804 ( .A(n13885), .ZN(n11585) );
  NOR2_X1 U11805 ( .A1(n11571), .A2(n19918), .ZN(n11580) );
  AOI21_X1 U11806 ( .B1(n11577), .B2(n11734), .A(n11576), .ZN(n13799) );
  INV_X1 U11807 ( .A(n11566), .ZN(n11567) );
  NAND2_X1 U11808 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11549) );
  NOR2_X1 U11809 ( .A1(n11549), .A2(n11548), .ZN(n11560) );
  INV_X1 U11810 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U11811 ( .A1(n11529), .A2(n11547), .ZN(n9764) );
  XNOR2_X1 U11812 ( .A(n12288), .B(n14380), .ZN(n9819) );
  NAND2_X1 U11813 ( .A1(n14833), .A2(n9822), .ZN(n14483) );
  AND2_X1 U11814 ( .A1(n14831), .A2(n14830), .ZN(n14833) );
  NAND2_X1 U11815 ( .A1(n14833), .A2(n14423), .ZN(n14485) );
  NAND2_X1 U11816 ( .A1(n14508), .A2(n9827), .ZN(n14495) );
  NAND2_X1 U11817 ( .A1(n9813), .A2(n9812), .ZN(n14509) );
  INV_X1 U11818 ( .A(n14158), .ZN(n9812) );
  INV_X1 U11819 ( .A(n14522), .ZN(n9813) );
  NAND2_X1 U11820 ( .A1(n16052), .A2(n9694), .ZN(n9845) );
  INV_X1 U11821 ( .A(n14710), .ZN(n9847) );
  OR2_X1 U11822 ( .A1(n14520), .A2(n14519), .ZN(n14522) );
  NAND2_X1 U11823 ( .A1(n14530), .A2(n14449), .ZN(n14520) );
  AND2_X1 U11824 ( .A1(n14528), .A2(n14527), .ZN(n14530) );
  OR2_X1 U11825 ( .A1(n14140), .A2(n12234), .ZN(n14546) );
  OR2_X1 U11826 ( .A1(n16106), .A2(n16105), .ZN(n16108) );
  NOR2_X1 U11827 ( .A1(n16108), .A2(n14042), .ZN(n14552) );
  OR2_X1 U11828 ( .A1(n11444), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16062) );
  AND2_X1 U11829 ( .A1(n12195), .A2(n12194), .ZN(n13733) );
  NAND2_X1 U11830 ( .A1(n12197), .A2(n12196), .ZN(n13870) );
  INV_X1 U11831 ( .A(n13733), .ZN(n12196) );
  INV_X1 U11832 ( .A(n13736), .ZN(n12197) );
  NAND2_X1 U11833 ( .A1(n19977), .A2(n19976), .ZN(n19975) );
  AND2_X1 U11834 ( .A1(n13862), .A2(n13863), .ZN(n13865) );
  NAND2_X1 U11835 ( .A1(n13865), .A2(n9654), .ZN(n13736) );
  OR2_X1 U11836 ( .A1(n11519), .A2(n11803), .ZN(n11246) );
  AOI21_X1 U11837 ( .B1(n11374), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9839), 
        .ZN(n9838) );
  XNOR2_X1 U11838 ( .A(n11278), .B(n11279), .ZN(n11530) );
  INV_X1 U11839 ( .A(n9631), .ZN(n20318) );
  OAI211_X1 U11840 ( .C1(n13369), .C2(n13368), .A(n13367), .B(n13366), .ZN(
        n15854) );
  CLKBUF_X1 U11841 ( .A(n11362), .Z(n20073) );
  AND3_X1 U11842 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20635), .A3(n20036), 
        .ZN(n20084) );
  INV_X1 U11843 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20572) );
  NOR2_X1 U11844 ( .A1(n20525), .A2(n9631), .ZN(n20492) );
  OR2_X1 U11845 ( .A1(n20034), .A2(n13709), .ZN(n20525) );
  AOI21_X1 U11846 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20493), .A(n20095), 
        .ZN(n20580) );
  NAND2_X1 U11847 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13499), .ZN(n15880) );
  MUX2_X1 U11848 ( .A(n10231), .B(n10524), .S(n12350), .Z(n10503) );
  OR2_X1 U11849 ( .A1(n19837), .A2(n10910), .ZN(n10506) );
  NAND2_X1 U11850 ( .A1(n12314), .A2(n9649), .ZN(n12312) );
  NAND2_X1 U11851 ( .A1(n15016), .A2(n12347), .ZN(n9754) );
  INV_X1 U11852 ( .A(n15235), .ZN(n9752) );
  AND2_X1 U11853 ( .A1(n10466), .A2(n10385), .ZN(n13069) );
  OR2_X1 U11854 ( .A1(n10428), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U11855 ( .A1(n10387), .A2(n10430), .ZN(n10434) );
  NAND2_X1 U11856 ( .A1(n10418), .A2(n15122), .ZN(n10428) );
  NOR2_X1 U11857 ( .A1(n12343), .A2(n15307), .ZN(n12344) );
  INV_X1 U11858 ( .A(n15072), .ZN(n12624) );
  XNOR2_X1 U11859 ( .A(n9796), .B(n12567), .ZN(n15094) );
  AND2_X1 U11860 ( .A1(n12445), .A2(n13989), .ZN(n12446) );
  AND2_X1 U11861 ( .A1(n13204), .A2(n13203), .ZN(n19139) );
  INV_X1 U11862 ( .A(n13050), .ZN(n15698) );
  OR2_X1 U11863 ( .A1(n9741), .A2(n15290), .ZN(n9740) );
  NOR2_X1 U11864 ( .A1(n12332), .A2(n9747), .ZN(n12342) );
  NOR2_X1 U11865 ( .A1(n9747), .A2(n9745), .ZN(n9744) );
  AND2_X1 U11866 ( .A1(n10798), .A2(n10797), .ZN(n13088) );
  NAND2_X1 U11867 ( .A1(n9746), .A2(n9881), .ZN(n12340) );
  INV_X1 U11868 ( .A(n9737), .ZN(n9735) );
  AND2_X1 U11869 ( .A1(n10770), .A2(n10769), .ZN(n13577) );
  OR2_X1 U11870 ( .A1(n10844), .A2(n15357), .ZN(n10770) );
  AND2_X1 U11871 ( .A1(n10764), .A2(n10763), .ZN(n13481) );
  OR2_X1 U11872 ( .A1(n10844), .A2(n15631), .ZN(n10764) );
  INV_X1 U11873 ( .A(n12338), .ZN(n12131) );
  INV_X1 U11874 ( .A(n13401), .ZN(n10760) );
  INV_X1 U11875 ( .A(n10074), .ZN(n10088) );
  INV_X1 U11876 ( .A(n16322), .ZN(n14342) );
  INV_X1 U11877 ( .A(n10841), .ZN(n14252) );
  INV_X1 U11878 ( .A(n15135), .ZN(n9866) );
  AND2_X1 U11879 ( .A1(n15458), .A2(n10932), .ZN(n15405) );
  INV_X1 U11880 ( .A(n15241), .ZN(n9734) );
  XNOR2_X1 U11881 ( .A(n10386), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15268) );
  NAND2_X1 U11882 ( .A1(n13069), .A2(n14320), .ZN(n10386) );
  AND2_X1 U11883 ( .A1(n14200), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15458) );
  NAND2_X1 U11884 ( .A1(n13058), .A2(n13059), .ZN(n15036) );
  NAND2_X1 U11885 ( .A1(n9864), .A2(n13061), .ZN(n9863) );
  INV_X1 U11886 ( .A(n14238), .ZN(n9864) );
  NOR3_X1 U11887 ( .A1(n14027), .A2(n9678), .A3(n14238), .ZN(n14239) );
  OR2_X1 U11888 ( .A1(n16268), .A2(n10943), .ZN(n15480) );
  OR3_X1 U11889 ( .A1(n18930), .A2(n10402), .A3(n10930), .ZN(n15296) );
  NAND2_X1 U11890 ( .A1(n9859), .A2(n16267), .ZN(n9858) );
  OR2_X1 U11891 ( .A1(n18966), .A2(n10453), .ZN(n15321) );
  AND3_X1 U11892 ( .A1(n10692), .A2(n10691), .A3(n10690), .ZN(n13958) );
  INV_X1 U11893 ( .A(n15337), .ZN(n15529) );
  INV_X1 U11894 ( .A(n15335), .ZN(n15555) );
  AND2_X1 U11895 ( .A1(n13534), .A2(n13535), .ZN(n10790) );
  AND2_X1 U11896 ( .A1(n9645), .A2(n15581), .ZN(n9867) );
  AND2_X1 U11897 ( .A1(n15589), .A2(n9645), .ZN(n15582) );
  NAND2_X1 U11898 ( .A1(n15358), .A2(n10888), .ZN(n15345) );
  NAND2_X1 U11899 ( .A1(n9667), .A2(n9857), .ZN(n15627) );
  NAND2_X1 U11900 ( .A1(n9857), .A2(n9683), .ZN(n13424) );
  INV_X1 U11901 ( .A(n10582), .ZN(n9852) );
  NOR2_X1 U11902 ( .A1(n14342), .A2(n13805), .ZN(n15602) );
  AOI21_X1 U11903 ( .B1(n9724), .B2(n9727), .A(n9721), .ZN(n9720) );
  NOR2_X1 U11904 ( .A1(n9724), .A2(n9728), .ZN(n9723) );
  AND2_X1 U11905 ( .A1(n9728), .A2(n9722), .ZN(n9721) );
  INV_X1 U11906 ( .A(n9851), .ZN(n13306) );
  NAND2_X1 U11907 ( .A1(n10092), .A2(n10093), .ZN(n10101) );
  XNOR2_X1 U11908 ( .A(n9658), .B(n10573), .ZN(n13543) );
  INV_X1 U11909 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9896) );
  CLKBUF_X1 U11910 ( .A(n10494), .Z(n15669) );
  NAND2_X1 U11911 ( .A1(n12402), .A2(n12401), .ZN(n13443) );
  NAND2_X1 U11912 ( .A1(n13338), .A2(n13339), .ZN(n12402) );
  AND2_X1 U11913 ( .A1(n12406), .A2(n12385), .ZN(n13444) );
  INV_X1 U11914 ( .A(n19274), .ZN(n19270) );
  NAND2_X1 U11915 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19634), .ZN(n19220) );
  NOR2_X2 U11916 ( .A1(n15696), .A2(n15697), .ZN(n19234) );
  NOR2_X2 U11917 ( .A1(n15698), .A2(n15697), .ZN(n19233) );
  INV_X1 U11918 ( .A(n19220), .ZN(n19229) );
  NAND2_X1 U11919 ( .A1(n10547), .A2(n10546), .ZN(n16345) );
  AOI21_X1 U11920 ( .B1(n12959), .B2(n12962), .A(n12958), .ZN(n18682) );
  OAI22_X1 U11921 ( .A1(n13013), .A2(n18684), .B1(n18688), .B2(n18201), .ZN(
        n18690) );
  NAND2_X1 U11922 ( .A1(n18890), .A2(n18239), .ZN(n16567) );
  CLKBUF_X1 U11923 ( .A(n12726), .Z(n17217) );
  NOR2_X1 U11924 ( .A1(n15834), .A2(n18675), .ZN(n12677) );
  NOR2_X1 U11925 ( .A1(n12723), .A2(n9806), .ZN(n9805) );
  NAND2_X1 U11926 ( .A1(n15742), .A2(n15828), .ZN(n15906) );
  AND2_X1 U11927 ( .A1(n16564), .A2(n13098), .ZN(n15831) );
  NAND2_X1 U11928 ( .A1(n12950), .A2(n9715), .ZN(n17494) );
  INV_X1 U11929 ( .A(n12922), .ZN(n9715) );
  OAI21_X1 U11930 ( .B1(n17894), .B2(n17678), .A(n18278), .ZN(n17694) );
  NOR2_X1 U11931 ( .A1(n17720), .A2(n17695), .ZN(n17691) );
  NOR2_X1 U11932 ( .A1(n18086), .A2(n18098), .ZN(n17746) );
  INV_X1 U11933 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17844) );
  NOR2_X1 U11934 ( .A1(n15892), .A2(n17908), .ZN(n16394) );
  NAND2_X1 U11935 ( .A1(n17563), .A2(n12816), .ZN(n15840) );
  AND2_X1 U11936 ( .A1(n17589), .A2(n9681), .ZN(n9807) );
  NAND2_X1 U11937 ( .A1(n12785), .A2(n12969), .ZN(n12788) );
  AOI21_X1 U11938 ( .B1(n17598), .B2(n12810), .A(n12809), .ZN(n12813) );
  NOR2_X1 U11939 ( .A1(n12810), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12809) );
  NOR2_X1 U11940 ( .A1(n12799), .A2(n12804), .ZN(n17689) );
  NOR2_X1 U11941 ( .A1(n18096), .A2(n16412), .ZN(n18045) );
  NAND2_X1 U11942 ( .A1(n12794), .A2(n12793), .ZN(n17723) );
  NAND2_X1 U11943 ( .A1(n17719), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17718) );
  NOR2_X1 U11944 ( .A1(n17772), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17762) );
  NAND2_X1 U11945 ( .A1(n17792), .A2(n18122), .ZN(n17772) );
  NAND2_X1 U11946 ( .A1(n18100), .A2(n18670), .ZN(n18073) );
  NOR2_X1 U11947 ( .A1(n18684), .A2(n16419), .ZN(n18097) );
  INV_X1 U11948 ( .A(n16411), .ZN(n18098) );
  OAI21_X1 U11949 ( .B1(n18661), .B2(n15825), .A(n18660), .ZN(n18668) );
  AND2_X1 U11950 ( .A1(n9809), .A2(n17816), .ZN(n17792) );
  NOR2_X1 U11951 ( .A1(n9810), .A2(n17811), .ZN(n9809) );
  INV_X1 U11952 ( .A(n9810), .ZN(n9808) );
  NOR2_X1 U11953 ( .A1(n17825), .A2(n17824), .ZN(n17823) );
  INV_X1 U11954 ( .A(n18251), .ZN(n12966) );
  XNOR2_X1 U11955 ( .A(n12772), .B(n12759), .ZN(n17883) );
  XNOR2_X1 U11956 ( .A(n17432), .B(n18836), .ZN(n17891) );
  NOR2_X1 U11957 ( .A1(n15826), .A2(n15825), .ZN(n18100) );
  NAND2_X1 U11958 ( .A1(n12915), .A2(n12918), .ZN(n18665) );
  NAND2_X1 U11959 ( .A1(n15741), .A2(n18888), .ZN(n18670) );
  INV_X1 U11960 ( .A(n17433), .ZN(n18239) );
  NOR2_X1 U11961 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18238), .ZN(n18579) );
  NAND3_X1 U11962 ( .A1(n12902), .A2(n12901), .A3(n12900), .ZN(n18264) );
  AOI211_X1 U11963 ( .C1(n17334), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n12899), .B(n12898), .ZN(n12900) );
  NOR2_X2 U11964 ( .A1(n12837), .A2(n12836), .ZN(n18877) );
  INV_X1 U11965 ( .A(n18725), .ZN(n18873) );
  INV_X1 U11966 ( .A(n17494), .ZN(n18718) );
  NOR2_X1 U11967 ( .A1(n15997), .A2(n20675), .ZN(n14128) );
  NAND2_X1 U11968 ( .A1(n16007), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15997) );
  NOR2_X1 U11969 ( .A1(n16020), .A2(n20669), .ZN(n16007) );
  INV_X1 U11970 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19918) );
  INV_X1 U11971 ( .A(n19909), .ZN(n19965) );
  XNOR2_X1 U11972 ( .A(n9815), .B(n13517), .ZN(n13852) );
  INV_X1 U11973 ( .A(n14300), .ZN(n14466) );
  CLKBUF_X1 U11974 ( .A(n14550), .Z(n19968) );
  INV_X1 U11975 ( .A(n19967), .ZN(n16021) );
  OR2_X1 U11976 ( .A1(n13726), .A2(n13729), .ZN(n13727) );
  INV_X1 U11977 ( .A(n14577), .ZN(n14603) );
  INV_X1 U11978 ( .A(n14614), .ZN(n14618) );
  OR2_X1 U11979 ( .A1(n14618), .A2(n13356), .ZN(n14617) );
  NOR2_X1 U11980 ( .A1(n13463), .A2(n20742), .ZN(n15902) );
  OR2_X1 U11981 ( .A1(n13462), .A2(n13461), .ZN(n13772) );
  INV_X1 U11982 ( .A(n14071), .ZN(n14116) );
  AOI21_X1 U11983 ( .B1(n14435), .B2(n14498), .A(n14576), .ZN(n14691) );
  NAND2_X1 U11984 ( .A1(n13558), .A2(n11547), .ZN(n13588) );
  INV_X1 U11985 ( .A(n19985), .ZN(n16048) );
  OR2_X1 U11986 ( .A1(n19981), .A2(n12116), .ZN(n14741) );
  OR2_X1 U11987 ( .A1(n16145), .A2(n20574), .ZN(n20031) );
  AND2_X1 U11988 ( .A1(n14818), .A2(n14294), .ZN(n14809) );
  AOI21_X1 U11989 ( .B1(n14936), .B2(n20018), .A(n20015), .ZN(n20003) );
  AND2_X1 U11990 ( .A1(n20011), .A2(n14955), .ZN(n20009) );
  INV_X1 U11991 ( .A(n16120), .ZN(n20013) );
  INV_X1 U11992 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20493) );
  INV_X1 U11993 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20320) );
  NAND2_X1 U11994 ( .A1(n11407), .A2(n11391), .ZN(n20035) );
  INV_X1 U11995 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20029) );
  NAND2_X1 U11996 ( .A1(n13702), .A2(n20095), .ZN(n20028) );
  INV_X1 U11997 ( .A(n20120), .ZN(n20111) );
  OAI21_X1 U11998 ( .B1(n9875), .B2(n20203), .A(n20530), .ZN(n20221) );
  INV_X1 U11999 ( .A(n20218), .ZN(n20220) );
  OAI211_X1 U12000 ( .C1(n9879), .C2(n20451), .A(n20377), .B(n20325), .ZN(
        n20342) );
  INV_X1 U12001 ( .A(n20408), .ZN(n20367) );
  INV_X1 U12002 ( .A(n20442), .ZN(n20576) );
  INV_X1 U12003 ( .A(n20463), .ZN(n20593) );
  INV_X1 U12004 ( .A(n20467), .ZN(n20599) );
  INV_X1 U12005 ( .A(n20475), .ZN(n20611) );
  INV_X1 U12006 ( .A(n20479), .ZN(n20617) );
  INV_X1 U12007 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20893) );
  NOR2_X1 U12008 ( .A1(n14974), .A2(n12329), .ZN(n16155) );
  OAI21_X1 U12009 ( .B1(n16167), .B2(n9757), .A(n9756), .ZN(n14974) );
  NAND2_X1 U12010 ( .A1(n15208), .A2(n9758), .ZN(n9757) );
  NAND2_X1 U12011 ( .A1(n12329), .A2(n15208), .ZN(n9756) );
  INV_X1 U12012 ( .A(n16166), .ZN(n9758) );
  NOR2_X1 U12013 ( .A1(n16167), .A2(n16166), .ZN(n16165) );
  INV_X1 U12014 ( .A(n9755), .ZN(n15002) );
  NOR2_X1 U12015 ( .A1(n15017), .A2(n12329), .ZN(n15003) );
  NOR2_X1 U12016 ( .A1(n15016), .A2(n15256), .ZN(n15017) );
  NAND2_X1 U12017 ( .A1(n9750), .A2(n15282), .ZN(n9749) );
  OR2_X1 U12018 ( .A1(n12329), .A2(n9751), .ZN(n9750) );
  INV_X1 U12019 ( .A(n14192), .ZN(n9751) );
  NOR2_X1 U12020 ( .A1(n13054), .A2(n12329), .ZN(n15032) );
  NOR2_X1 U12021 ( .A1(n13055), .A2(n14192), .ZN(n13054) );
  AND2_X1 U12022 ( .A1(n10406), .A2(n10413), .ZN(n13954) );
  NAND2_X1 U12023 ( .A1(n12366), .A2(n12354), .ZN(n19030) );
  AND2_X1 U12024 ( .A1(n19030), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19036) );
  AND2_X1 U12025 ( .A1(n19858), .A2(n12351), .ZN(n19041) );
  INV_X1 U12026 ( .A(n19724), .ZN(n19042) );
  INV_X1 U12027 ( .A(n15063), .ZN(n10853) );
  INV_X1 U12028 ( .A(n19801), .ZN(n15727) );
  INV_X1 U12029 ( .A(n15130), .ZN(n15118) );
  AND2_X1 U12030 ( .A1(n12672), .A2(n19721), .ZN(n15123) );
  OR2_X1 U12031 ( .A1(n13579), .A2(n10509), .ZN(n15130) );
  INV_X1 U12032 ( .A(n9792), .ZN(n15086) );
  NOR2_X1 U12033 ( .A1(n15100), .A2(n15099), .ZN(n15098) );
  NOR2_X1 U12034 ( .A1(n15105), .A2(n12523), .ZN(n15100) );
  NOR2_X1 U12035 ( .A1(n14027), .A2(n14026), .ZN(n14050) );
  AND2_X1 U12036 ( .A1(n14006), .A2(n15696), .ZN(n19072) );
  AND2_X1 U12037 ( .A1(n14006), .A2(n15698), .ZN(n19073) );
  NOR2_X1 U12038 ( .A1(n15540), .A2(n15541), .ZN(n13090) );
  NOR2_X1 U12039 ( .A1(n19108), .A2(n19130), .ZN(n19114) );
  INV_X1 U12040 ( .A(n16191), .ZN(n19130) );
  INV_X1 U12041 ( .A(n19134), .ZN(n19108) );
  NOR2_X1 U12042 ( .A1(n13219), .A2(n13223), .ZN(n19063) );
  INV_X1 U12043 ( .A(n19103), .ZN(n19129) );
  CLKBUF_X1 U12044 ( .A(n19172), .Z(n19162) );
  NOR2_X1 U12046 ( .A1(n19139), .A2(n19860), .ZN(n19172) );
  INV_X1 U12048 ( .A(n16258), .ZN(n19191) );
  AND2_X1 U12049 ( .A1(n19202), .A2(n19816), .ZN(n19198) );
  AND2_X1 U12050 ( .A1(n19202), .A2(n13310), .ZN(n16258) );
  OR2_X1 U12051 ( .A1(n15127), .A2(n15126), .ZN(n18919) );
  INV_X1 U12052 ( .A(n15327), .ZN(n18972) );
  NAND2_X1 U12053 ( .A1(n9729), .A2(n10364), .ZN(n15577) );
  OAI21_X1 U12054 ( .B1(n10862), .B2(n14320), .A(n13451), .ZN(n13803) );
  INV_X1 U12055 ( .A(n16326), .ZN(n16299) );
  INV_X1 U12056 ( .A(n16318), .ZN(n16307) );
  INV_X1 U12057 ( .A(n16330), .ZN(n16295) );
  NAND2_X1 U12058 ( .A1(n10936), .A2(n10747), .ZN(n16318) );
  NAND2_X1 U12059 ( .A1(n15490), .A2(n15495), .ZN(n16322) );
  INV_X1 U12060 ( .A(n19063), .ZN(n19827) );
  INV_X1 U12061 ( .A(n19817), .ZN(n19820) );
  XNOR2_X1 U12062 ( .A(n13341), .B(n13340), .ZN(n19810) );
  INV_X1 U12063 ( .A(n16371), .ZN(n15692) );
  OAI21_X1 U12064 ( .B1(n19339), .B2(n19355), .A(n19338), .ZN(n19357) );
  NOR2_X1 U12065 ( .A1(n19335), .A2(n19596), .ZN(n19386) );
  NOR2_X1 U12066 ( .A1(n19361), .A2(n19794), .ZN(n19462) );
  OAI21_X1 U12067 ( .B1(n19465), .B2(n19445), .A(n19634), .ZN(n19467) );
  INV_X1 U12068 ( .A(n19498), .ZN(n19491) );
  OAI21_X1 U12069 ( .B1(n19504), .B2(n19521), .A(n19634), .ZN(n19523) );
  INV_X1 U12070 ( .A(n19683), .ZN(n19643) );
  INV_X1 U12071 ( .A(n19611), .ZN(n19653) );
  INV_X1 U12072 ( .A(n19255), .ZN(n19652) );
  INV_X1 U12073 ( .A(n19672), .ZN(n19657) );
  INV_X1 U12074 ( .A(n19689), .ZN(n19658) );
  OAI21_X1 U12075 ( .B1(n19639), .B2(n19638), .A(n19637), .ZN(n19668) );
  INV_X1 U12076 ( .A(n19617), .ZN(n19692) );
  INV_X1 U12077 ( .A(n19714), .ZN(n19700) );
  INV_X1 U12078 ( .A(n19620), .ZN(n19698) );
  INV_X1 U12079 ( .A(n19666), .ZN(n19699) );
  INV_X1 U12080 ( .A(n19627), .ZN(n19709) );
  AND2_X1 U12081 ( .A1(n16345), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16371) );
  CLKBUF_X1 U12082 ( .A(n19781), .Z(n19778) );
  INV_X1 U12083 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18741) );
  INV_X1 U12084 ( .A(n16897), .ZN(n16934) );
  NOR2_X2 U12085 ( .A1(n16567), .A2(n18720), .ZN(n16926) );
  INV_X1 U12086 ( .A(n16926), .ZN(n16937) );
  INV_X1 U12087 ( .A(n16933), .ZN(n16946) );
  NAND3_X1 U12088 ( .A1(n12880), .A2(n12879), .A3(n12878), .ZN(n18274) );
  NAND4_X1 U12089 ( .A1(n18873), .A2(n18248), .A3(n18239), .A4(n15906), .ZN(
        n17263) );
  NAND2_X1 U12090 ( .A1(n17287), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17286) );
  NOR3_X1 U12091 ( .A1(n17302), .A2(n17442), .A3(n9713), .ZN(n17287) );
  NOR2_X1 U12092 ( .A1(n17302), .A2(n17442), .ZN(n17296) );
  NOR2_X1 U12093 ( .A1(n18274), .A2(n17306), .ZN(n17303) );
  NOR3_X1 U12094 ( .A1(n17366), .A2(n17313), .A3(n17448), .ZN(n17307) );
  NAND2_X1 U12095 ( .A1(n17307), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17306) );
  NAND2_X1 U12096 ( .A1(n17370), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17366) );
  INV_X1 U12097 ( .A(n17318), .ZN(n17365) );
  NOR2_X1 U12098 ( .A1(n17375), .A2(n17544), .ZN(n17370) );
  NAND2_X1 U12099 ( .A1(n17426), .A2(n9712), .ZN(n17398) );
  AND2_X1 U12100 ( .A1(n17267), .A2(n9693), .ZN(n9712) );
  NOR2_X1 U12101 ( .A1(n12705), .A2(n12704), .ZN(n17409) );
  NAND2_X1 U12102 ( .A1(n17266), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17427) );
  NOR2_X1 U12103 ( .A1(n17427), .A2(n17516), .ZN(n17426) );
  NAND2_X1 U12104 ( .A1(n15909), .A2(n17266), .ZN(n17431) );
  INV_X1 U12105 ( .A(n17431), .ZN(n17397) );
  NOR3_X1 U12106 ( .A1(n18248), .A2(n17494), .A3(n17493), .ZN(n17503) );
  CLKBUF_X1 U12107 ( .A(n17540), .Z(n17533) );
  INV_X1 U12108 ( .A(n17503), .ZN(n17543) );
  NOR2_X1 U12109 ( .A1(n17533), .A2(n18877), .ZN(n17541) );
  NAND2_X1 U12110 ( .A1(n18013), .A2(n17795), .ZN(n17704) );
  INV_X1 U12111 ( .A(n17754), .ZN(n17741) );
  INV_X1 U12112 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17806) );
  INV_X1 U12113 ( .A(n17895), .ZN(n17885) );
  NAND2_X1 U12114 ( .A1(n17858), .A2(n17901), .ZN(n17896) );
  NAND2_X1 U12115 ( .A1(n17741), .A2(n17678), .ZN(n17895) );
  INV_X1 U12116 ( .A(n17893), .ZN(n17905) );
  NAND2_X1 U12117 ( .A1(n12815), .A2(n16415), .ZN(n16426) );
  NOR2_X1 U12118 ( .A1(n18182), .A2(n17983), .ZN(n18036) );
  NOR2_X1 U12119 ( .A1(n18073), .A2(n18668), .ZN(n18135) );
  NAND2_X1 U12120 ( .A1(n17870), .A2(n12777), .ZN(n17861) );
  INV_X1 U12121 ( .A(n18670), .ZN(n18689) );
  INV_X1 U12122 ( .A(n18182), .ZN(n18218) );
  INV_X1 U12123 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18240) );
  CLKBUF_X1 U12124 ( .A(n18816), .Z(n18810) );
  INV_X1 U12126 ( .A(U212), .ZN(n16489) );
  AOI211_X1 U12127 ( .C1(n9699), .C2(n9659), .A(n14387), .B(n9698), .ZN(n14388) );
  OAI21_X1 U12128 ( .B1(n14408), .B2(n20702), .A(n14383), .ZN(n9699) );
  AOI211_X1 U12129 ( .C1(P1_REIP_REG_28__SCAN_IN), .C2(n14417), .A(n14416), 
        .B(n14415), .ZN(n14418) );
  OAI21_X1 U12130 ( .B1(n15955), .B2(n19924), .A(n9770), .ZN(P1_U2820) );
  AOI21_X1 U12131 ( .B1(n9773), .B2(n15957), .A(n9771), .ZN(n9770) );
  OR2_X1 U12132 ( .A1(n15956), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n9773) );
  AOI21_X1 U12133 ( .B1(n14300), .B2(n20021), .A(n14299), .ZN(n14301) );
  OAI21_X1 U12134 ( .B1(n15061), .B2(n19185), .A(n14374), .ZN(n14375) );
  AOI21_X1 U12135 ( .B1(n9711), .B2(P3_EAX_REG_31__SCAN_IN), .A(n9710), .ZN(
        n17270) );
  AND2_X1 U12136 ( .A1(n17364), .A2(BUF2_REG_31__SCAN_IN), .ZN(n9710) );
  AOI21_X1 U12137 ( .B1(n13026), .B2(n17893), .A(n13025), .ZN(n13027) );
  OAI21_X1 U12138 ( .B1(n13024), .B2(n17745), .A(n13023), .ZN(n13025) );
  OAI21_X1 U12139 ( .B1(n17919), .B2(n17778), .A(n9802), .ZN(P3_U2803) );
  AOI21_X1 U12140 ( .B1(n9804), .B2(n17568), .A(n9803), .ZN(n9802) );
  OR2_X1 U12141 ( .A1(n17567), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9804) );
  AOI21_X1 U12142 ( .B1(n13026), .B2(n18225), .A(n13010), .ZN(n13011) );
  OAI21_X1 U12143 ( .B1(n13024), .B2(n18139), .A(n13009), .ZN(n13010) );
  CLKBUF_X3 U12144 ( .A(n12904), .Z(n17329) );
  INV_X1 U12145 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10266) );
  INV_X2 U12146 ( .A(n13081), .ZN(n12329) );
  INV_X1 U12147 ( .A(n12684), .ZN(n15808) );
  NAND2_X1 U12148 ( .A1(n12337), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12335) );
  OR2_X1 U12149 ( .A1(n14027), .A2(n9678), .ZN(n9639) );
  INV_X2 U12150 ( .A(n12057), .ZN(n11206) );
  NOR3_X1 U12151 ( .A1(n14027), .A2(n9678), .A3(n9863), .ZN(n13060) );
  NOR2_X1 U12152 ( .A1(n14988), .A2(n9691), .ZN(n10738) );
  AND2_X1 U12153 ( .A1(n11502), .A2(n11511), .ZN(n9640) );
  AND2_X1 U12154 ( .A1(n10346), .A2(n9675), .ZN(n9641) );
  INV_X1 U12155 ( .A(n11183), .ZN(n12089) );
  NOR3_X1 U12156 ( .A1(n14988), .A2(n15149), .A3(n14978), .ZN(n14977) );
  OR2_X1 U12157 ( .A1(n17566), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9642) );
  NOR2_X1 U12158 ( .A1(n12343), .A2(n9740), .ZN(n12324) );
  NAND3_X1 U12159 ( .A1(n12131), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U12160 ( .A1(n9746), .A2(n9744), .ZN(n12330) );
  NAND2_X1 U12161 ( .A1(n12337), .A2(n9735), .ZN(n12333) );
  AND2_X1 U12162 ( .A1(n9861), .A2(n9859), .ZN(n9643) );
  AND2_X1 U12163 ( .A1(n9862), .A2(n13091), .ZN(n9644) );
  AND2_X1 U12164 ( .A1(n9868), .A2(n15588), .ZN(n9645) );
  NAND2_X1 U12165 ( .A1(n11579), .A2(n11578), .ZN(n13798) );
  AND2_X1 U12166 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n9646) );
  AND2_X1 U12167 ( .A1(n10364), .A2(n9685), .ZN(n9647) );
  NOR2_X1 U12168 ( .A1(n12323), .A2(n15262), .ZN(n12316) );
  AND4_X1 U12169 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n10585), .ZN(
        n9648) );
  AND2_X1 U12170 ( .A1(n12135), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9649) );
  INV_X1 U12171 ( .A(n13276), .ZN(n9857) );
  AND2_X1 U12172 ( .A1(n9769), .A2(n11659), .ZN(n9650) );
  AND2_X1 U12173 ( .A1(n9649), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9651) );
  AND2_X2 U12174 ( .A1(n9584), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10153) );
  AND2_X2 U12175 ( .A1(n10143), .A2(n12491), .ZN(n10159) );
  AND2_X1 U12176 ( .A1(n11130), .A2(n9891), .ZN(n9652) );
  INV_X1 U12177 ( .A(n9930), .ZN(n12653) );
  AND2_X1 U12178 ( .A1(n12188), .A2(n12187), .ZN(n9654) );
  NAND2_X1 U12179 ( .A1(n9607), .A2(n10346), .ZN(n15348) );
  NOR2_X1 U12180 ( .A1(n14533), .A2(n14445), .ZN(n14444) );
  NAND2_X1 U12181 ( .A1(n15575), .A2(n9784), .ZN(n9655) );
  AND2_X1 U12182 ( .A1(n13967), .A2(n9769), .ZN(n9656) );
  INV_X1 U12183 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9928) );
  INV_X1 U12184 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9956) );
  INV_X1 U12185 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9999) );
  OR4_X1 U12186 ( .A1(n14408), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14383), .A4(
        n20702), .ZN(n9657) );
  AND2_X2 U12187 ( .A1(n10129), .A2(n10130), .ZN(n10290) );
  AND2_X1 U12188 ( .A1(n17816), .A2(n9808), .ZN(n12797) );
  AND2_X1 U12189 ( .A1(n13233), .A2(n13235), .ZN(n9658) );
  OR2_X1 U12190 ( .A1(n14417), .A2(n12306), .ZN(n9659) );
  AND4_X1 U12191 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n9660) );
  AND2_X1 U12192 ( .A1(n14880), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9661) );
  OR2_X1 U12193 ( .A1(n14394), .A2(n20031), .ZN(n9662) );
  OR2_X1 U12194 ( .A1(n10919), .A2(n10023), .ZN(n9663) );
  NAND2_X1 U12195 ( .A1(n12586), .A2(n9889), .ZN(n9664) );
  INV_X1 U12196 ( .A(n11373), .ZN(n9839) );
  AND4_X1 U12197 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n9665) );
  AND2_X1 U12198 ( .A1(n9839), .A2(n11374), .ZN(n9666) );
  NAND2_X1 U12199 ( .A1(n9793), .A2(n9794), .ZN(n9796) );
  AND2_X1 U12200 ( .A1(n9856), .A2(n15628), .ZN(n9667) );
  AND2_X1 U12201 ( .A1(n14516), .A2(n11977), .ZN(n14471) );
  NAND2_X1 U12202 ( .A1(n13353), .A2(n9700), .ZN(n11507) );
  INV_X1 U12203 ( .A(n13889), .ZN(n9833) );
  AND2_X1 U12204 ( .A1(n12210), .A2(n12209), .ZN(n13889) );
  NAND2_X1 U12205 ( .A1(n14411), .A2(n14410), .ZN(n14398) );
  AND2_X1 U12206 ( .A1(n15268), .A2(n10437), .ZN(n9668) );
  AND2_X1 U12207 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12779), .ZN(
        n9669) );
  NOR2_X1 U12208 ( .A1(n13920), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11425) );
  AND2_X1 U12209 ( .A1(n12812), .A2(n12813), .ZN(n9670) );
  INV_X1 U12210 ( .A(n11362), .ZN(n11486) );
  AND2_X1 U12211 ( .A1(n10341), .A2(n10340), .ZN(n10885) );
  INV_X1 U12212 ( .A(n10885), .ZN(n10886) );
  NAND2_X1 U12213 ( .A1(n13442), .A2(n12407), .ZN(n13396) );
  NAND2_X1 U12214 ( .A1(n10563), .A2(n10560), .ZN(n10705) );
  INV_X1 U12215 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12935) );
  OR2_X1 U12216 ( .A1(n12343), .A2(n9741), .ZN(n9671) );
  NAND2_X1 U12217 ( .A1(n13810), .A2(n13809), .ZN(n13811) );
  NOR2_X1 U12218 ( .A1(n12336), .A2(n16256), .ZN(n12337) );
  NOR2_X1 U12219 ( .A1(n12330), .A2(n10801), .ZN(n12331) );
  NAND2_X1 U12220 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  AND2_X1 U12221 ( .A1(n12337), .A2(n9736), .ZN(n12334) );
  AND2_X1 U12222 ( .A1(n14508), .A2(n14502), .ZN(n9672) );
  NAND2_X1 U12223 ( .A1(n10465), .A2(n15240), .ZN(n9673) );
  OAI21_X1 U12224 ( .B1(n19058), .B2(n12387), .A(n12386), .ZN(n13219) );
  OAI21_X1 U12225 ( .B1(n10862), .B2(n9723), .A(n9720), .ZN(n13942) );
  INV_X1 U12226 ( .A(n12332), .ZN(n9746) );
  XNOR2_X1 U12227 ( .A(n14266), .B(n14265), .ZN(n19066) );
  INV_X1 U12228 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20635) );
  OR2_X1 U12229 ( .A1(n14988), .A2(n15149), .ZN(n9674) );
  AND2_X1 U12230 ( .A1(n10362), .A2(n10361), .ZN(n9675) );
  INV_X1 U12231 ( .A(n9727), .ZN(n9726) );
  NAND2_X1 U12232 ( .A1(n13451), .A2(n13806), .ZN(n9727) );
  INV_X1 U12233 ( .A(n13798), .ZN(n11586) );
  AND2_X1 U12234 ( .A1(n10397), .A2(n10930), .ZN(n15295) );
  NAND2_X1 U12235 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12338) );
  OR2_X1 U12236 ( .A1(n20078), .A2(n20638), .ZN(n11717) );
  NOR2_X1 U12237 ( .A1(n16165), .A2(n12329), .ZN(n9676) );
  AND2_X1 U12238 ( .A1(n12337), .A2(n9738), .ZN(n9677) );
  INV_X1 U12239 ( .A(n11184), .ZN(n12087) );
  AND2_X2 U12240 ( .A1(n10970), .A2(n13680), .ZN(n11184) );
  INV_X1 U12241 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12395) );
  INV_X1 U12242 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9739) );
  OR2_X1 U12243 ( .A1(n9865), .A2(n14026), .ZN(n9678) );
  NAND2_X1 U12244 ( .A1(n10601), .A2(n10600), .ZN(n15589) );
  NOR2_X1 U12245 ( .A1(n13870), .A2(n13869), .ZN(n9679) );
  NAND2_X1 U12246 ( .A1(n12324), .A2(n9887), .ZN(n12323) );
  NAND2_X1 U12247 ( .A1(n14049), .A2(n9797), .ZN(n14066) );
  NAND2_X1 U12248 ( .A1(n9861), .A2(n9644), .ZN(n13089) );
  NAND2_X1 U12249 ( .A1(n15589), .A2(n15588), .ZN(n13410) );
  NOR2_X1 U12250 ( .A1(n15540), .A2(n9858), .ZN(n15509) );
  NAND2_X1 U12251 ( .A1(n15589), .A2(n9867), .ZN(n13614) );
  INV_X1 U12252 ( .A(n19936), .ZN(n19948) );
  AND2_X1 U12253 ( .A1(n12293), .A2(n12290), .ZN(n19936) );
  NAND2_X1 U12254 ( .A1(n14049), .A2(n9798), .ZN(n14065) );
  NOR2_X1 U12255 ( .A1(n13870), .A2(n9831), .ZN(n9680) );
  NAND2_X1 U12256 ( .A1(n10511), .A2(n12352), .ZN(n10745) );
  INV_X1 U12257 ( .A(n12608), .ZN(n9790) );
  NOR2_X1 U12258 ( .A1(n13276), .A2(n10582), .ZN(n13449) );
  NAND2_X1 U12259 ( .A1(n15627), .A2(n10597), .ZN(n15605) );
  OR2_X1 U12260 ( .A1(n12810), .A2(n17912), .ZN(n9681) );
  NOR2_X2 U12261 ( .A1(n13480), .A2(n13577), .ZN(n13571) );
  AND2_X1 U12262 ( .A1(n9765), .A2(n9764), .ZN(n13557) );
  OR2_X1 U12263 ( .A1(n17401), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9682) );
  AND2_X1 U12264 ( .A1(n9852), .A2(n9855), .ZN(n9683) );
  INV_X1 U12265 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15350) );
  AND2_X1 U12266 ( .A1(n9753), .A2(n9752), .ZN(n9684) );
  NAND2_X1 U12267 ( .A1(n10441), .A2(n15563), .ZN(n9685) );
  INV_X1 U12268 ( .A(n9828), .ZN(n9827) );
  OR2_X1 U12269 ( .A1(n14494), .A2(n9829), .ZN(n9828) );
  AND2_X1 U12270 ( .A1(n14049), .A2(n14048), .ZN(n9686) );
  AOI21_X1 U12271 ( .B1(n13055), .B2(n12347), .A(n9749), .ZN(n9748) );
  AND2_X1 U12272 ( .A1(n9857), .A2(n9856), .ZN(n9687) );
  AND2_X1 U12273 ( .A1(n9769), .A2(n9767), .ZN(n9688) );
  OR2_X1 U12274 ( .A1(n15959), .A2(n19919), .ZN(n9689) );
  OAI22_X1 U12275 ( .A1(n19716), .A2(n14341), .B1(n14372), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U12276 ( .A1(n12314), .A2(n12135), .ZN(n12311) );
  INV_X1 U12277 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9811) );
  OR2_X1 U12278 ( .A1(n18175), .A2(n18806), .ZN(n9690) );
  INV_X1 U12279 ( .A(n16340), .ZN(n9707) );
  INV_X1 U12280 ( .A(n14502), .ZN(n9829) );
  OR3_X1 U12281 ( .A1(n15149), .A2(n14978), .A3(n9866), .ZN(n9691) );
  INV_X1 U12282 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9745) );
  AND2_X1 U12283 ( .A1(n9784), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9692) );
  AND2_X1 U12284 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .ZN(n9693) );
  INV_X1 U12285 ( .A(n15493), .ZN(n9785) );
  OR3_X1 U12286 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n9694) );
  INV_X1 U12287 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9742) );
  INV_X1 U12288 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n9713) );
  INV_X1 U12289 ( .A(n12165), .ZN(n12079) );
  AND2_X1 U12290 ( .A1(n15693), .A2(n19716), .ZN(n19634) );
  AOI22_X2 U12291 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9580), .B1(DATAI_30_), 
        .B2(n9579), .ZN(n20559) );
  AOI22_X2 U12292 ( .A1(DATAI_17_), .A2(n9579), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9580), .ZN(n20592) );
  AOI22_X2 U12293 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9580), .B1(DATAI_23_), 
        .B2(n9579), .ZN(n20633) );
  AOI22_X2 U12294 ( .A1(DATAI_18_), .A2(n9579), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n9580), .ZN(n20598) );
  AOI22_X2 U12295 ( .A1(DATAI_19_), .A2(n9579), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9580), .ZN(n20604) );
  AOI22_X2 U12296 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9580), .B1(DATAI_29_), 
        .B2(n9579), .ZN(n20555) );
  AOI22_X2 U12297 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9580), .B1(DATAI_28_), 
        .B2(n9579), .ZN(n20551) );
  NOR3_X2 U12298 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20493), .A3(
        n20571), .ZN(n20514) );
  AOI22_X2 U12299 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9580), .B1(DATAI_16_), 
        .B2(n9579), .ZN(n20586) );
  NOR3_X4 U12300 ( .A1(n18416), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18477) );
  NOR2_X2 U12301 ( .A1(n14428), .A2(n20694), .ZN(n15925) );
  NAND2_X1 U12302 ( .A1(n15938), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U12303 ( .A1(n15956), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14439) );
  NAND3_X1 U12304 ( .A1(n9697), .A2(n11506), .A3(n9696), .ZN(n9695) );
  NOR2_X2 U12305 ( .A1(n14446), .A2(n20678), .ZN(n15979) );
  NAND2_X1 U12306 ( .A1(n20073), .A2(n11495), .ZN(n9700) );
  NAND2_X4 U12307 ( .A1(n9652), .A2(n11131), .ZN(n20054) );
  AND2_X2 U12308 ( .A1(n9701), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10963) );
  INV_X2 U12309 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9701) );
  AND2_X2 U12310 ( .A1(n12293), .A2(n12158), .ZN(n19957) );
  AND3_X1 U12311 ( .A1(n10512), .A2(n19230), .A3(n10518), .ZN(n10916) );
  XNOR2_X1 U12312 ( .A(n19224), .B(n10017), .ZN(n10508) );
  OR2_X2 U12313 ( .A1(n19224), .A2(n9619), .ZN(n10556) );
  AND2_X2 U12314 ( .A1(n10874), .A2(n10210), .ZN(n13810) );
  NAND2_X1 U12315 ( .A1(n10059), .A2(n9704), .ZN(n10070) );
  OAI21_X1 U12316 ( .B1(n10566), .B2(n9732), .A(n9705), .ZN(n10520) );
  NOR2_X1 U12317 ( .A1(n9707), .A2(n9732), .ZN(n9706) );
  NAND2_X1 U12318 ( .A1(n15335), .A2(n16282), .ZN(n9709) );
  NAND2_X1 U12319 ( .A1(n15536), .A2(n10411), .ZN(n9708) );
  OR2_X2 U12320 ( .A1(n10895), .A2(n10896), .ZN(n15344) );
  NAND2_X2 U12321 ( .A1(n15626), .A2(n15619), .ZN(n10891) );
  NAND2_X2 U12322 ( .A1(n10904), .A2(n10903), .ZN(n15575) );
  INV_X1 U12323 ( .A(n17287), .ZN(n17292) );
  INV_X2 U12324 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18849) );
  NAND2_X1 U12325 ( .A1(n9653), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10127) );
  NAND2_X1 U12326 ( .A1(n9653), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n9717) );
  NAND3_X2 U12327 ( .A1(n9719), .A2(n9718), .A3(n10589), .ZN(n10876) );
  INV_X1 U12328 ( .A(n10208), .ZN(n9718) );
  INV_X1 U12329 ( .A(n10209), .ZN(n9719) );
  NAND2_X1 U12330 ( .A1(n13942), .A2(n13943), .ZN(n10280) );
  XNOR2_X2 U12331 ( .A(n10749), .B(n10748), .ZN(n12379) );
  NAND3_X1 U12332 ( .A1(n10019), .A2(n13238), .A3(n10560), .ZN(n16339) );
  NAND3_X1 U12333 ( .A1(n15241), .A2(n15225), .A3(n9733), .ZN(n9890) );
  AND2_X2 U12334 ( .A1(n9759), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11022) );
  INV_X2 U12335 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9759) );
  NAND3_X1 U12336 ( .A1(n13264), .A2(n13263), .A3(n9760), .ZN(n13374) );
  AOI21_X1 U12337 ( .B1(n11565), .B2(n11734), .A(n11564), .ZN(n13592) );
  NAND3_X1 U12338 ( .A1(n11407), .A2(n11391), .A3(n11734), .ZN(n9761) );
  NAND3_X1 U12339 ( .A1(n11390), .A2(n11383), .A3(n9766), .ZN(n9765) );
  NAND2_X1 U12340 ( .A1(n11390), .A2(n11383), .ZN(n13704) );
  OR2_X2 U12341 ( .A1(n11382), .A2(n11381), .ZN(n11390) );
  AND2_X2 U12342 ( .A1(n13967), .A2(n9688), .ZN(n14540) );
  NAND3_X1 U12343 ( .A1(n15958), .A2(n9689), .A3(n9772), .ZN(n9771) );
  NOR2_X4 U12344 ( .A1(n14533), .A2(n9774), .ZN(n14516) );
  NAND2_X1 U12345 ( .A1(n14516), .A2(n14432), .ZN(n14506) );
  AND2_X2 U12346 ( .A1(n10855), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10051) );
  INV_X1 U12347 ( .A(n10051), .ZN(n10774) );
  NOR2_X2 U12348 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U12349 ( .A1(n15669), .A2(n9783), .ZN(n13785) );
  NAND2_X1 U12350 ( .A1(n9786), .A2(n10876), .ZN(n10878) );
  AND2_X2 U12351 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10143) );
  NAND3_X1 U12352 ( .A1(n9949), .A2(n9948), .A3(n10509), .ZN(n10035) );
  NAND2_X1 U12353 ( .A1(n9595), .A2(n12394), .ZN(n9789) );
  NAND2_X1 U12354 ( .A1(n9789), .A2(n12398), .ZN(n12400) );
  NAND2_X1 U12355 ( .A1(n15105), .A2(n9795), .ZN(n9793) );
  OAI21_X2 U12356 ( .B1(n17870), .B2(n9801), .A(n9799), .ZN(n12782) );
  AOI21_X1 U12357 ( .B1(n9800), .B2(n17862), .A(n9669), .ZN(n9799) );
  INV_X1 U12358 ( .A(n12777), .ZN(n9800) );
  INV_X1 U12359 ( .A(n17862), .ZN(n9801) );
  NAND2_X1 U12360 ( .A1(n17861), .A2(n17862), .ZN(n17860) );
  NAND3_X1 U12361 ( .A1(n9642), .A2(n17569), .A3(n9690), .ZN(n9803) );
  NAND4_X1 U12362 ( .A1(n9665), .A2(n12724), .A3(n12725), .A4(n9805), .ZN(
        n17421) );
  NAND3_X1 U12363 ( .A1(n12812), .A2(n12813), .A3(n20800), .ZN(n17570) );
  NOR2_X2 U12364 ( .A1(n17676), .A2(n17811), .ZN(n17605) );
  NOR2_X2 U12365 ( .A1(n17677), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17676) );
  NAND2_X1 U12366 ( .A1(n17816), .A2(n12792), .ZN(n12796) );
  NAND2_X1 U12367 ( .A1(n12792), .A2(n9811), .ZN(n9810) );
  NOR2_X4 U12368 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13694) );
  OR2_X1 U12369 ( .A1(n14401), .A2(n9819), .ZN(n9818) );
  INV_X1 U12370 ( .A(n9825), .ZN(n14475) );
  NAND3_X1 U12371 ( .A1(n11108), .A2(n9835), .A3(n11362), .ZN(n11117) );
  NAND2_X1 U12372 ( .A1(n11117), .A2(n20064), .ZN(n11111) );
  NAND2_X1 U12373 ( .A1(n11537), .A2(n9838), .ZN(n9837) );
  NAND2_X1 U12374 ( .A1(n11537), .A2(n20635), .ZN(n11372) );
  NOR2_X2 U12375 ( .A1(n9661), .A2(n16052), .ZN(n9846) );
  OAI21_X2 U12376 ( .B1(n13998), .B2(n11449), .A(n11448), .ZN(n14118) );
  OAI21_X2 U12377 ( .B1(n16065), .B2(n16061), .A(n16062), .ZN(n13998) );
  INV_X2 U12378 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9848) );
  NOR2_X2 U12379 ( .A1(n9701), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U12380 ( .A1(n10291), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10116) );
  AND2_X2 U12381 ( .A1(n10125), .A2(n10124), .ZN(n19527) );
  INV_X1 U12382 ( .A(n11390), .ZN(n11305) );
  NAND2_X1 U12383 ( .A1(n10289), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10117) );
  AND2_X1 U12384 ( .A1(n14533), .A2(n14532), .ZN(n16042) );
  XNOR2_X2 U12385 ( .A(n10312), .B(n15631), .ZN(n15618) );
  NAND2_X2 U12386 ( .A1(n10311), .A2(n19033), .ZN(n10312) );
  XNOR2_X1 U12387 ( .A(n10879), .B(n10878), .ZN(n13941) );
  NAND2_X1 U12388 ( .A1(n14552), .A2(n14551), .ZN(n14140) );
  NAND2_X1 U12389 ( .A1(n10035), .A2(n9994), .ZN(n10045) );
  INV_X1 U12390 ( .A(n10859), .ZN(n10957) );
  NAND2_X2 U12391 ( .A1(n13564), .A2(n13563), .ZN(n13565) );
  INV_X1 U12392 ( .A(n13629), .ZN(n11579) );
  INV_X1 U12393 ( .A(n15626), .ZN(n10882) );
  NAND2_X1 U12394 ( .A1(n15512), .A2(n14004), .ZN(n14027) );
  AOI22_X1 U12395 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n9958) );
  AOI22_X1 U12396 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n9942) );
  AND2_X1 U12397 ( .A1(n15111), .A2(n12543), .ZN(n12523) );
  OAI21_X2 U12398 ( .B1(n16201), .B2(n14174), .A(n16200), .ZN(n15323) );
  INV_X1 U12399 ( .A(n14124), .ZN(n11738) );
  INV_X1 U12400 ( .A(n12295), .ZN(n12308) );
  OR2_X1 U12401 ( .A1(n11144), .A2(n11143), .ZN(n11145) );
  NAND2_X1 U12402 ( .A1(n10131), .A2(n10130), .ZN(n10322) );
  NAND2_X1 U12403 ( .A1(n10131), .A2(n10128), .ZN(n10183) );
  NAND2_X1 U12404 ( .A1(n10131), .A2(n10118), .ZN(n19274) );
  AND2_X2 U12405 ( .A1(n10131), .A2(n10124), .ZN(n19306) );
  OAI211_X1 U12406 ( .C1(n16319), .C2(n15061), .A(n14345), .B(n14344), .ZN(
        n14346) );
  NAND2_X1 U12407 ( .A1(n14540), .A2(n14125), .ZN(n14124) );
  CLKBUF_X1 U12408 ( .A(n11537), .Z(n20160) );
  XNOR2_X1 U12409 ( .A(n11195), .B(n11194), .ZN(n11537) );
  INV_X1 U12410 ( .A(n15955), .ZN(n14706) );
  OAI21_X2 U12411 ( .B1(n15314), .B2(n15313), .A(n14177), .ZN(n15305) );
  AND2_X1 U12412 ( .A1(n12128), .A2(n9578), .ZN(n9869) );
  OR2_X1 U12413 ( .A1(n14751), .A2(n16115), .ZN(n9870) );
  INV_X1 U12414 ( .A(n14535), .ZN(n14548) );
  INV_X1 U12415 ( .A(n20739), .ZN(n13818) );
  INV_X1 U12416 ( .A(n20095), .ZN(n20202) );
  AND2_X1 U12417 ( .A1(n11304), .A2(n11303), .ZN(n13709) );
  INV_X1 U12419 ( .A(n12686), .ZN(n12870) );
  INV_X1 U12420 ( .A(n13967), .ZN(n14020) );
  AND4_X1 U12421 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n9871) );
  NAND2_X1 U12422 ( .A1(n10477), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n9872) );
  INV_X1 U12423 ( .A(n17811), .ZN(n12810) );
  INV_X1 U12424 ( .A(n17755), .ZN(n17731) );
  AND4_X1 U12425 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n9873) );
  OR2_X1 U12426 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9874) );
  NOR2_X1 U12427 ( .A1(n20441), .A2(n20251), .ZN(n9875) );
  AND3_X1 U12428 ( .A1(n12734), .A2(n12733), .A3(n12732), .ZN(n9876) );
  AND4_X1 U12429 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n9877) );
  AND2_X1 U12430 ( .A1(n10881), .A2(n10886), .ZN(n9878) );
  NOR2_X1 U12431 ( .A1(n20441), .A2(n20410), .ZN(n9879) );
  NOR2_X1 U12432 ( .A1(n20448), .A2(n20197), .ZN(n9880) );
  NOR2_X1 U12433 ( .A1(n10791), .A2(n10778), .ZN(n9881) );
  INV_X1 U12434 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14279) );
  AND3_X1 U12435 ( .A1(n11468), .A2(n11467), .A3(n20806), .ZN(n9883) );
  NOR2_X1 U12436 ( .A1(n12689), .A2(n12683), .ZN(n12731) );
  INV_X1 U12437 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12009) );
  INV_X1 U12438 ( .A(n15619), .ZN(n10881) );
  INV_X1 U12439 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11468) );
  INV_X1 U12440 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20805) );
  AND2_X1 U12441 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n9885) );
  INV_X1 U12442 ( .A(n12393), .ZN(n13273) );
  AND2_X1 U12443 ( .A1(n14327), .A2(n14324), .ZN(n9886) );
  INV_X1 U12444 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12774) );
  AND2_X1 U12445 ( .A1(n12132), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9887) );
  OR2_X1 U12446 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9888) );
  INV_X1 U12447 ( .A(n14633), .ZN(n11471) );
  AND2_X1 U12448 ( .A1(n12585), .A2(n12606), .ZN(n9889) );
  INV_X1 U12449 ( .A(n12678), .ZN(n12893) );
  INV_X1 U12450 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11166) );
  AND2_X2 U12451 ( .A1(n10119), .A2(n10130), .ZN(n10291) );
  AND3_X1 U12452 ( .A1(n11129), .A2(n11128), .A3(n11127), .ZN(n9891) );
  INV_X1 U12453 ( .A(n12176), .ZN(n13244) );
  AND4_X1 U12454 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n9892) );
  NAND2_X1 U12455 ( .A1(n13444), .A2(n13443), .ZN(n13442) );
  OR2_X1 U12456 ( .A1(n9658), .A2(n10573), .ZN(n9893) );
  INV_X1 U12457 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19240) );
  NOR3_X1 U12458 ( .A1(n11502), .A2(n11495), .A3(n11501), .ZN(n11513) );
  NAND2_X1 U12459 ( .A1(n19527), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10126) );
  NAND2_X1 U12460 ( .A1(n11513), .A2(n12146), .ZN(n11514) );
  NAND2_X1 U12461 ( .A1(n10127), .A2(n10126), .ZN(n10134) );
  NAND2_X1 U12462 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  AOI22_X1 U12463 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10290), .B1(
        n10291), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10190) );
  AND2_X1 U12464 ( .A1(n12649), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9950) );
  AND2_X1 U12465 ( .A1(n20493), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11496) );
  INV_X1 U12466 ( .A(n12098), .ZN(n12008) );
  INV_X1 U12467 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11667) );
  AND4_X1 U12468 ( .A1(n11215), .A2(n11214), .A3(n11213), .A4(n11212), .ZN(
        n11216) );
  AND4_X1 U12469 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n11189) );
  OR2_X1 U12470 ( .A1(n11321), .A2(n11320), .ZN(n11420) );
  AND4_X1 U12471 ( .A1(n11224), .A2(n11223), .A3(n11222), .A4(n11221), .ZN(
        n11228) );
  AND2_X1 U12472 ( .A1(n11270), .A2(n11269), .ZN(n11279) );
  INV_X1 U12473 ( .A(n15264), .ZN(n10437) );
  NAND2_X1 U12474 ( .A1(n10029), .A2(n9965), .ZN(n10031) );
  AOI21_X1 U12475 ( .B1(n11519), .B2(n12146), .A(n11518), .ZN(n11520) );
  INV_X1 U12476 ( .A(n11259), .ZN(n12092) );
  INV_X1 U12477 ( .A(n13799), .ZN(n11578) );
  NAND2_X1 U12478 ( .A1(n11340), .A2(n11339), .ZN(n11403) );
  INV_X1 U12479 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U12480 ( .A1(n13506), .A2(n20064), .ZN(n13261) );
  AND4_X1 U12481 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n11237) );
  NAND2_X1 U12482 ( .A1(n12350), .A2(n10534), .ZN(n10238) );
  NAND2_X1 U12483 ( .A1(n10079), .A2(n10078), .ZN(n10750) );
  INV_X1 U12484 ( .A(n12567), .ZN(n12568) );
  INV_X1 U12485 ( .A(n10266), .ZN(n9981) );
  INV_X1 U12486 ( .A(n16236), .ZN(n10361) );
  INV_X1 U12487 ( .A(n16240), .ZN(n10362) );
  INV_X1 U12488 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9894) );
  INV_X1 U12489 ( .A(n10045), .ZN(n10046) );
  CLKBUF_X1 U12490 ( .A(n12658), .Z(n10146) );
  OAI21_X1 U12491 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n9714), .A(
        n12936), .ZN(n12937) );
  NOR2_X1 U12492 ( .A1(n11067), .A2(n11066), .ZN(n11082) );
  NOR2_X1 U12493 ( .A1(n13681), .A2(n11092), .ZN(n11093) );
  OR2_X1 U12494 ( .A1(n12049), .A2(n14637), .ZN(n12051) );
  NOR2_X1 U12495 ( .A1(n11912), .A2(n11871), .ZN(n11851) );
  AND2_X1 U12496 ( .A1(n11359), .A2(n11358), .ZN(n11417) );
  OR2_X1 U12497 ( .A1(n14316), .A2(n20638), .ZN(n11554) );
  OR2_X1 U12498 ( .A1(n11242), .A2(n20635), .ZN(n11363) );
  NAND2_X1 U12499 ( .A1(n11246), .A2(n11245), .ZN(n11374) );
  NAND2_X1 U12500 ( .A1(n20319), .A2(n20635), .ZN(n11304) );
  INV_X1 U12501 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10367) );
  AND2_X1 U12502 ( .A1(n12606), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12380) );
  NAND2_X1 U12503 ( .A1(n9796), .A2(n12568), .ZN(n12569) );
  INV_X1 U12504 ( .A(n14068), .ZN(n12477) );
  NAND2_X1 U12505 ( .A1(n12673), .A2(n16294), .ZN(n10858) );
  OR2_X1 U12507 ( .A1(n15480), .A2(n10930), .ZN(n14242) );
  AND2_X1 U12508 ( .A1(n13621), .A2(n13669), .ZN(n13535) );
  INV_X1 U12509 ( .A(n15620), .ZN(n15624) );
  INV_X1 U12510 ( .A(n12379), .ZN(n13450) );
  INV_X1 U12511 ( .A(n10183), .ZN(n10281) );
  NAND2_X1 U12512 ( .A1(n10119), .A2(n10128), .ZN(n10184) );
  NAND2_X1 U12513 ( .A1(n9962), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9963) );
  NOR2_X1 U12514 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12933), .ZN(
        n12956) );
  INV_X1 U12515 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12793) );
  INV_X1 U12516 ( .A(n12783), .ZN(n12781) );
  INV_X1 U12517 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20851) );
  OAI211_X1 U12518 ( .C1(n9614), .C2(n11166), .A(n11168), .B(n11167), .ZN(
        n11169) );
  AND2_X1 U12519 ( .A1(n12238), .A2(n12237), .ZN(n14129) );
  INV_X1 U12520 ( .A(n14136), .ZN(n11659) );
  AND2_X1 U12521 ( .A1(n11851), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U12522 ( .A1(n11913), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11912) );
  INV_X1 U12523 ( .A(n11717), .ZN(n11734) );
  OR2_X1 U12524 ( .A1(n11425), .A2(n11430), .ZN(n11431) );
  XNOR2_X1 U12525 ( .A(n11401), .B(n19999), .ZN(n19977) );
  AND3_X1 U12526 ( .A1(n13373), .A2(n13258), .A3(n11475), .ZN(n13363) );
  OR2_X1 U12527 ( .A1(n10823), .A2(n14230), .ZN(n10824) );
  AND2_X1 U12528 ( .A1(n10758), .A2(n10757), .ZN(n13400) );
  AND2_X1 U12529 ( .A1(n12377), .A2(n12376), .ZN(n12606) );
  OR2_X1 U12530 ( .A1(n10306), .A2(n10305), .ZN(n10593) );
  AND2_X1 U12531 ( .A1(n10539), .A2(n10491), .ZN(n16340) );
  OR2_X1 U12532 ( .A1(n10844), .A2(n10411), .ZN(n10798) );
  OAI211_X1 U12533 ( .C1(n14352), .C2(n16318), .A(n10858), .B(n12137), .ZN(
        n10859) );
  INV_X1 U12534 ( .A(n15295), .ZN(n14180) );
  AOI21_X1 U12535 ( .B1(n10882), .B2(n10884), .A(n9878), .ZN(n10883) );
  INV_X1 U12536 ( .A(n10189), .ZN(n15725) );
  INV_X1 U12537 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20794) );
  AOI21_X1 U12538 ( .B1(n17402), .B2(n12788), .A(n17811), .ZN(n12791) );
  AND2_X1 U12539 ( .A1(n17811), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12816) );
  NOR2_X1 U12540 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17637), .ZN(
        n17627) );
  OAI22_X1 U12541 ( .A1(n12804), .A2(n17703), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n12810), .ZN(n12805) );
  NOR2_X1 U12542 ( .A1(n17823), .A2(n18130), .ZN(n12990) );
  INV_X1 U12543 ( .A(n12882), .ZN(n17340) );
  AND2_X1 U12544 ( .A1(n12223), .A2(n12222), .ZN(n14042) );
  AND2_X1 U12545 ( .A1(n14420), .A2(n11975), .ZN(n14419) );
  OR2_X1 U12546 ( .A1(n9635), .A2(n20638), .ZN(n11960) );
  NAND2_X1 U12547 ( .A1(n12000), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12049) );
  NOR2_X1 U12548 ( .A1(n11943), .A2(n15968), .ZN(n11916) );
  INV_X1 U12549 ( .A(n12079), .ZN(n12112) );
  NAND2_X1 U12550 ( .A1(n11660), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U12551 ( .A1(n11605), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11637) );
  INV_X2 U12552 ( .A(n16052), .ZN(n14751) );
  NAND2_X1 U12553 ( .A1(n14935), .A2(n20003), .ZN(n16123) );
  NAND2_X1 U12554 ( .A1(n19987), .A2(n20009), .ZN(n14936) );
  NAND2_X1 U12555 ( .A1(n13524), .A2(n13685), .ZN(n14914) );
  NAND2_X1 U12556 ( .A1(n20093), .A2(n11274), .ZN(n13851) );
  OR2_X1 U12557 ( .A1(n20034), .A2(n13710), .ZN(n20290) );
  AND2_X1 U12558 ( .A1(n20521), .A2(n20202), .ZN(n20377) );
  AND2_X1 U12559 ( .A1(n20379), .A2(n20202), .ZN(n20530) );
  NAND2_X1 U12560 ( .A1(n20635), .A2(n20036), .ZN(n20095) );
  OR2_X1 U12561 ( .A1(n13693), .A2(n13692), .ZN(n15864) );
  OR2_X1 U12562 ( .A1(n10912), .A2(n10911), .ZN(n16344) );
  INV_X1 U12563 ( .A(n19052), .ZN(n12367) );
  INV_X1 U12564 ( .A(n12350), .ZN(n12364) );
  INV_X1 U12565 ( .A(n12606), .ZN(n13397) );
  AND2_X1 U12566 ( .A1(n16340), .A2(n19721), .ZN(n13099) );
  INV_X1 U12567 ( .A(n10954), .ZN(n10955) );
  NAND2_X1 U12568 ( .A1(n15287), .A2(n14180), .ZN(n14181) );
  NOR2_X1 U12569 ( .A1(n16302), .A2(n16301), .ZN(n15579) );
  AND3_X1 U12570 ( .A1(n10617), .A2(n10616), .A3(n10615), .ZN(n13411) );
  AND2_X1 U12571 ( .A1(n12401), .A2(n13338), .ZN(n13341) );
  NAND2_X1 U12572 ( .A1(n19801), .A2(n19827), .ZN(n19335) );
  NAND2_X1 U12573 ( .A1(n19801), .A2(n19063), .ZN(n19361) );
  OR3_X1 U12574 ( .A1(n19593), .A2(n19630), .A3(n19852), .ZN(n19598) );
  INV_X1 U12575 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19852) );
  NAND2_X1 U12576 ( .A1(n16573), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16572) );
  NOR2_X1 U12577 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16792), .ZN(n16772) );
  NOR2_X1 U12578 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16843), .ZN(n16821) );
  NOR2_X1 U12579 ( .A1(n16574), .A2(n17546), .ZN(n16573) );
  NOR2_X1 U12580 ( .A1(n17750), .A2(n17742), .ZN(n17736) );
  NOR2_X1 U12581 ( .A1(n17820), .A2(n17806), .ZN(n17802) );
  NAND2_X1 U12582 ( .A1(n13097), .A2(n17901), .ZN(n17678) );
  OAI21_X1 U12583 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18872), .A(n16544), 
        .ZN(n17901) );
  INV_X1 U12584 ( .A(n17746), .ZN(n18078) );
  INV_X1 U12585 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12759) );
  INV_X1 U12586 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20892) );
  NOR2_X1 U12587 ( .A1(n12868), .A2(n12867), .ZN(n17433) );
  AOI211_X1 U12588 ( .C1(n17334), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n12877), .B(n12876), .ZN(n12878) );
  AND2_X1 U12589 ( .A1(n14357), .A2(n12172), .ZN(n19902) );
  NAND2_X1 U12590 ( .A1(n13359), .A2(n13501), .ZN(n13355) );
  AND2_X1 U12591 ( .A1(n14434), .A2(n14433), .ZN(n14576) );
  NAND2_X1 U12592 ( .A1(n11916), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U12593 ( .A1(n11567), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11571) );
  INV_X1 U12594 ( .A(n20499), .ZN(n20574) );
  OR3_X1 U12595 ( .A1(n20010), .A2(n14288), .A3(n14287), .ZN(n16073) );
  NOR2_X1 U12596 ( .A1(n16123), .A2(n14157), .ZN(n14927) );
  AND2_X1 U12597 ( .A1(n12119), .A2(n20638), .ZN(n19973) );
  OR2_X1 U12598 ( .A1(n13934), .A2(n14920), .ZN(n20010) );
  OR2_X1 U12599 ( .A1(n14291), .A2(n14848), .ZN(n16118) );
  NOR2_X1 U12600 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20724) );
  OAI211_X1 U12601 ( .C1(n20047), .C2(n20451), .A(n20377), .B(n20046), .ZN(
        n20089) );
  AND2_X1 U12602 ( .A1(n20156), .A2(n20318), .ZN(n20092) );
  AND2_X1 U12603 ( .A1(n20035), .A2(n20034), .ZN(n20156) );
  INV_X1 U12604 ( .A(n20244), .ZN(n20247) );
  NOR2_X1 U12605 ( .A1(n20290), .A2(n9631), .ZN(n20228) );
  NOR2_X1 U12606 ( .A1(n20290), .A2(n20318), .ZN(n20287) );
  INV_X1 U12607 ( .A(n20307), .ZN(n20341) );
  AND2_X1 U12608 ( .A1(n9631), .A2(n9632), .ZN(n20523) );
  NOR2_X1 U12609 ( .A1(n20035), .A2(n13708), .ZN(n20413) );
  AND2_X1 U12610 ( .A1(n20492), .A2(n9632), .ZN(n20516) );
  OAI211_X1 U12611 ( .C1(n20560), .C2(n20531), .A(n20530), .B(n20529), .ZN(
        n20563) );
  INV_X1 U12612 ( .A(n20459), .ZN(n20587) );
  INV_X1 U12613 ( .A(n20471), .ZN(n20605) );
  INV_X1 U12614 ( .A(n20484), .ZN(n20624) );
  AND2_X1 U12615 ( .A1(n10372), .A2(n10374), .ZN(n13626) );
  OR2_X1 U12616 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  OR2_X1 U12617 ( .A1(n13776), .A2(n13532), .ZN(n13833) );
  AND2_X1 U12618 ( .A1(n19103), .A2(n13237), .ZN(n19071) );
  OR2_X1 U12619 ( .A1(n19071), .A2(n14006), .ZN(n19105) );
  INV_X1 U12620 ( .A(n13141), .ZN(n13196) );
  INV_X1 U12621 ( .A(n19202), .ZN(n19177) );
  AOI21_X1 U12622 ( .B1(n14223), .B2(n14221), .A(n14183), .ZN(n14188) );
  OR2_X1 U12623 ( .A1(n15562), .A2(n10946), .ZN(n15479) );
  INV_X1 U12624 ( .A(n14176), .ZN(n15313) );
  INV_X1 U12625 ( .A(n10856), .ZN(n19176) );
  INV_X1 U12626 ( .A(n15263), .ZN(n15334) );
  AND2_X1 U12627 ( .A1(n10936), .A2(n19839), .ZN(n16326) );
  OAI21_X1 U12628 ( .B1(n15705), .B2(n15704), .A(n15703), .ZN(n19235) );
  NOR2_X2 U12629 ( .A1(n19471), .A2(n19335), .ZN(n19266) );
  NOR2_X1 U12630 ( .A1(n19471), .A2(n19361), .ZN(n19287) );
  NOR2_X1 U12631 ( .A1(n19361), .A2(n19797), .ZN(n19348) );
  NOR2_X1 U12632 ( .A1(n19361), .A2(n19596), .ZN(n19393) );
  NOR2_X2 U12633 ( .A1(n19794), .A2(n19335), .ZN(n19437) );
  OAI21_X1 U12634 ( .B1(n19449), .B2(n19448), .A(n19447), .ZN(n19466) );
  NOR2_X2 U12635 ( .A1(n19562), .A2(n19797), .ZN(n19554) );
  OR2_X1 U12636 ( .A1(n19810), .A2(n19817), .ZN(n19797) );
  NOR2_X2 U12637 ( .A1(n19562), .A2(n19596), .ZN(n19623) );
  INV_X1 U12638 ( .A(n19577), .ZN(n19648) );
  INV_X1 U12639 ( .A(n19642), .ZN(n19675) );
  NOR2_X2 U12640 ( .A1(n19592), .A2(n19794), .ZN(n19710) );
  AND2_X1 U12641 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10554), .ZN(n19721) );
  AND3_X1 U12642 ( .A1(n17494), .A2(n16560), .A3(n16559), .ZN(n18683) );
  NAND2_X1 U12643 ( .A1(n12948), .A2(n12947), .ZN(n18688) );
  NOR2_X1 U12644 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16696), .ZN(n16682) );
  NOR2_X1 U12645 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16721), .ZN(n16704) );
  NOR2_X1 U12646 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16746), .ZN(n16726) );
  NOR2_X1 U12647 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16764), .ZN(n16753) );
  NOR2_X1 U12648 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16813), .ZN(n16795) );
  NOR2_X1 U12649 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16862), .ZN(n16847) );
  AOI211_X2 U12650 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(n18722), .A(n18890), 
        .B(n16563), .ZN(n16933) );
  NOR2_X1 U12651 ( .A1(n20777), .A2(n20776), .ZN(n20775) );
  OR2_X1 U12652 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16931) );
  NAND2_X1 U12653 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17303), .ZN(n17302) );
  INV_X1 U12654 ( .A(n17349), .ZN(n17364) );
  INV_X1 U12656 ( .A(n17543), .ZN(n17534) );
  NAND2_X1 U12657 ( .A1(n17912), .A2(n17580), .ZN(n17908) );
  NOR2_X1 U12658 ( .A1(n18853), .A2(n17896), .ZN(n17754) );
  OAI22_X1 U12659 ( .A1(n18098), .A2(n17905), .B1(n17745), .B2(n18096), .ZN(
        n17795) );
  INV_X1 U12660 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17820) );
  INV_X1 U12661 ( .A(n18278), .ZN(n18607) );
  INV_X1 U12662 ( .A(n17901), .ZN(n17888) );
  NOR2_X1 U12663 ( .A1(n12770), .A2(n12769), .ZN(n17900) );
  NOR2_X1 U12664 ( .A1(n17603), .A2(n17940), .ZN(n17580) );
  NOR2_X1 U12665 ( .A1(n18078), .A2(n17734), .ZN(n17719) );
  NOR2_X1 U12666 ( .A1(n18085), .A2(n18182), .ZN(n18123) );
  NAND2_X1 U12667 ( .A1(n17831), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17830) );
  INV_X1 U12668 ( .A(n18221), .ZN(n18204) );
  INV_X1 U12669 ( .A(n18579), .ZN(n18285) );
  NAND2_X1 U12670 ( .A1(n9659), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U12671 ( .A1(n14315), .A2(n19902), .ZN(n12309) );
  NAND2_X1 U12672 ( .A1(n14535), .A2(n9634), .ZN(n14550) );
  INV_X1 U12673 ( .A(n16042), .ZN(n14612) );
  NAND2_X1 U12674 ( .A1(n13355), .A2(n13354), .ZN(n14614) );
  NAND2_X1 U12675 ( .A1(n13463), .A2(n20037), .ZN(n13769) );
  INV_X1 U12676 ( .A(n13894), .ZN(n14114) );
  INV_X1 U12677 ( .A(n19981), .ZN(n19877) );
  NAND2_X1 U12678 ( .A1(n14741), .A2(n12118), .ZN(n19985) );
  INV_X1 U12679 ( .A(n20021), .ZN(n19993) );
  NAND2_X1 U12680 ( .A1(n13524), .A2(n13513), .ZN(n16120) );
  NAND2_X1 U12681 ( .A1(n20092), .A2(n9632), .ZN(n20120) );
  NAND2_X1 U12682 ( .A1(n20092), .A2(n20491), .ZN(n20150) );
  NAND2_X1 U12683 ( .A1(n20156), .A2(n20523), .ZN(n20191) );
  NAND2_X1 U12684 ( .A1(n20156), .A2(n20409), .ZN(n20218) );
  NAND2_X1 U12685 ( .A1(n20228), .A2(n9632), .ZN(n20244) );
  NAND2_X1 U12686 ( .A1(n20228), .A2(n20491), .ZN(n20286) );
  NAND2_X1 U12687 ( .A1(n20287), .A2(n9632), .ZN(n20317) );
  OR2_X1 U12688 ( .A1(n20350), .A2(n20491), .ZN(n20371) );
  OR2_X1 U12689 ( .A1(n20350), .A2(n9632), .ZN(n20408) );
  NAND2_X1 U12690 ( .A1(n20413), .A2(n20523), .ZN(n20432) );
  NAND2_X1 U12691 ( .A1(n20413), .A2(n20409), .ZN(n20490) );
  NAND2_X1 U12692 ( .A1(n20492), .A2(n20491), .ZN(n20566) );
  NAND2_X1 U12693 ( .A1(n20578), .A2(n20409), .ZN(n20632) );
  INV_X1 U12694 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20634) );
  INV_X1 U12695 ( .A(n20721), .ZN(n20717) );
  OR2_X1 U12696 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19868), .ZN(n20737) );
  AND2_X1 U12697 ( .A1(n12370), .A2(n12369), .ZN(n12371) );
  OR2_X1 U12698 ( .A1(n12366), .A2(n12365), .ZN(n19052) );
  INV_X1 U12699 ( .A(n19041), .ZN(n19057) );
  NAND2_X1 U12700 ( .A1(n13442), .A2(n13445), .ZN(n19801) );
  XNOR2_X1 U12701 ( .A(n13249), .B(n13248), .ZN(n19817) );
  AND2_X1 U12702 ( .A1(n13231), .A2(n19721), .ZN(n19103) );
  INV_X1 U12703 ( .A(n19105), .ZN(n19138) );
  INV_X1 U12704 ( .A(n19139), .ZN(n19174) );
  INV_X1 U12705 ( .A(n13161), .ZN(n13201) );
  INV_X1 U12706 ( .A(n9578), .ZN(n19192) );
  INV_X1 U12707 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16256) );
  NAND2_X1 U12708 ( .A1(n13110), .A2(n12129), .ZN(n19202) );
  AND2_X1 U12709 ( .A1(n13945), .A2(n10941), .ZN(n16316) );
  INV_X1 U12710 ( .A(n16294), .ZN(n16319) );
  INV_X1 U12711 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16358) );
  AOI211_X2 U12712 ( .C1(n15695), .C2(n15704), .A(n15694), .B(n19563), .ZN(
        n19239) );
  INV_X1 U12713 ( .A(n19287), .ZN(n19299) );
  INV_X1 U12714 ( .A(n19326), .ZN(n19318) );
  INV_X1 U12715 ( .A(n19348), .ZN(n19360) );
  INV_X1 U12716 ( .A(n19386), .ZN(n19384) );
  INV_X1 U12717 ( .A(n19393), .ZN(n19420) );
  INV_X1 U12718 ( .A(n19438), .ZN(n19435) );
  INV_X1 U12719 ( .A(n19462), .ZN(n19470) );
  OR2_X1 U12720 ( .A1(n19562), .A2(n19471), .ZN(n19498) );
  OR2_X1 U12721 ( .A1(n19592), .A2(n19471), .ZN(n19526) );
  OR2_X1 U12722 ( .A1(n19592), .A2(n19797), .ZN(n19591) );
  OR2_X1 U12723 ( .A1(n19592), .A2(n19596), .ZN(n19672) );
  INV_X1 U12724 ( .A(n19711), .ZN(n19704) );
  OR2_X1 U12725 ( .A1(n19562), .A2(n19794), .ZN(n19714) );
  NOR2_X1 U12726 ( .A1(n18683), .A2(n17493), .ZN(n18890) );
  NAND2_X1 U12727 ( .A1(n18873), .A2(n18690), .ZN(n16544) );
  INV_X1 U12728 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17742) );
  INV_X1 U12729 ( .A(n16921), .ZN(n16943) );
  INV_X1 U12730 ( .A(n16890), .ZN(n16944) );
  AND2_X1 U12731 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17236), .ZN(n17231) );
  NOR2_X2 U12732 ( .A1(n12695), .A2(n12694), .ZN(n17402) );
  NOR2_X1 U12733 ( .A1(n12715), .A2(n12714), .ZN(n17417) );
  AOI21_X1 U12734 ( .B1(n15908), .B2(n15907), .A(n18725), .ZN(n17266) );
  INV_X1 U12735 ( .A(n17453), .ZN(n17460) );
  NAND2_X1 U12736 ( .A1(n17492), .A2(n15831), .ZN(n17490) );
  INV_X1 U12737 ( .A(n17541), .ZN(n17536) );
  NAND2_X1 U12738 ( .A1(n17402), .A2(n13015), .ZN(n17745) );
  NOR2_X1 U12739 ( .A1(n17715), .A2(n17714), .ZN(n17702) );
  INV_X1 U12740 ( .A(n17812), .ZN(n17778) );
  INV_X1 U12741 ( .A(n13015), .ZN(n17904) );
  INV_X1 U12742 ( .A(n18141), .ZN(n18127) );
  INV_X1 U12743 ( .A(n18225), .ZN(n18187) );
  NAND2_X1 U12744 ( .A1(n18175), .A2(n18182), .ZN(n18221) );
  INV_X1 U12745 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18830) );
  INV_X1 U12746 ( .A(n16484), .ZN(n16491) );
  OAI211_X1 U12747 ( .C1(n14768), .C2(n19877), .A(n9662), .B(n12124), .ZN(
        P1_U2969) );
  AND2_X4 U12748 ( .A1(n15662), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12490) );
  INV_X2 U12749 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9897) );
  AND3_X4 U12750 ( .A1(n15659), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n9897), .ZN(n12649) );
  AOI22_X1 U12751 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n9895) );
  AND2_X1 U12752 ( .A1(n9895), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9901) );
  AOI22_X1 U12753 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n9900) );
  AOI22_X1 U12754 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U12755 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n9898) );
  NAND4_X1 U12756 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(n9908)
         );
  AOI22_X1 U12757 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n9902) );
  AND2_X1 U12758 ( .A1(n9902), .A2(n10266), .ZN(n9906) );
  AOI22_X1 U12759 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U12760 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U12761 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9623), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9903) );
  NAND4_X1 U12762 ( .A1(n9906), .A2(n9905), .A3(n9904), .A4(n9903), .ZN(n9907)
         );
  NAND2_X2 U12763 ( .A1(n9908), .A2(n9907), .ZN(n9967) );
  AOI22_X1 U12764 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U12765 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U12766 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U12767 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U12768 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U12769 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U12770 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9583), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U12771 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U12772 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U12773 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n9926) );
  INV_X2 U12774 ( .A(n9923), .ZN(n10001) );
  AOI22_X1 U12775 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U12776 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n9924) );
  NAND4_X1 U12777 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9929)
         );
  NAND2_X1 U12778 ( .A1(n9929), .A2(n9928), .ZN(n9937) );
  AOI22_X1 U12779 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U12780 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U12781 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n9931) );
  NAND4_X1 U12782 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9935)
         );
  NAND2_X1 U12783 ( .A1(n9935), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9936) );
  MUX2_X1 U12784 ( .A(n9608), .B(n10017), .S(n19224), .Z(n9949) );
  AOI22_X1 U12785 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U12786 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9970), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U12787 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U12788 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n9938) );
  NAND4_X1 U12789 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9947)
         );
  AOI22_X1 U12790 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n9945) );
  AOI22_X1 U12791 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U12792 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n9943) );
  NAND4_X1 U12793 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9946)
         );
  MUX2_X2 U12794 ( .A(n9947), .B(n9946), .S(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19230) );
  INV_X1 U12795 ( .A(n19230), .ZN(n10509) );
  INV_X1 U12796 ( .A(n10035), .ZN(n9966) );
  AOI22_X1 U12797 ( .A1(n9970), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9584), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U12798 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U12799 ( .A1(n9951), .A2(n9950), .ZN(n9953) );
  AOI22_X1 U12800 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n9952) );
  NAND4_X1 U12801 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9957)
         );
  NAND2_X1 U12802 ( .A1(n9957), .A2(n9956), .ZN(n9964) );
  AOI22_X1 U12803 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n9961) );
  AOI22_X1 U12804 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U12805 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n9959) );
  NAND4_X1 U12806 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9962)
         );
  NAND2_X1 U12807 ( .A1(n9966), .A2(n9965), .ZN(n9969) );
  NAND2_X1 U12808 ( .A1(n10916), .A2(n15699), .ZN(n9968) );
  NAND2_X1 U12809 ( .A1(n9969), .A2(n9968), .ZN(n10047) );
  AOI22_X1 U12810 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U12811 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U12812 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9972) );
  NAND4_X1 U12813 ( .A1(n9971), .A2(n9973), .A3(n9972), .A4(n9974), .ZN(n9980)
         );
  AOI22_X1 U12814 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9970), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U12815 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U12816 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U12817 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n9975) );
  NAND4_X1 U12818 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n9979)
         );
  AOI22_X1 U12819 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U12820 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U12821 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U12822 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n9983) );
  NAND4_X1 U12823 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9993)
         );
  AOI22_X1 U12824 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U12825 ( .A1(n9584), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9989) );
  AOI22_X1 U12826 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9970), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U12827 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U12828 ( .A1(n9991), .A2(n10266), .ZN(n9992) );
  AND2_X2 U12829 ( .A1(n9993), .A2(n9992), .ZN(n10559) );
  NOR2_X1 U12830 ( .A1(n10047), .A2(n12350), .ZN(n10016) );
  AND2_X1 U12831 ( .A1(n10022), .A2(n10556), .ZN(n9994) );
  NAND2_X1 U12832 ( .A1(n10045), .A2(n9627), .ZN(n10015) );
  NAND2_X1 U12833 ( .A1(n10556), .A2(n15699), .ZN(n10030) );
  AOI22_X1 U12834 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U12835 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U12836 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U12837 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U12838 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U12839 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12649), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10004) );
  AOI22_X1 U12840 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U12841 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9583), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12842 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  NAND2_X1 U12843 ( .A1(n10030), .A2(n15717), .ZN(n10014) );
  NOR2_X1 U12844 ( .A1(n10017), .A2(n15699), .ZN(n10010) );
  AND3_X2 U12845 ( .A1(n10011), .A2(n10010), .A3(n10914), .ZN(n13193) );
  INV_X1 U12846 ( .A(n13193), .ZN(n10012) );
  NAND2_X1 U12847 ( .A1(n10015), .A2(n10923), .ZN(n10048) );
  OAI21_X1 U12848 ( .B1(n10016), .B2(n10048), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10021) );
  NAND2_X1 U12849 ( .A1(n10017), .A2(n19230), .ZN(n10562) );
  NOR2_X1 U12850 ( .A1(n10562), .A2(n19224), .ZN(n10018) );
  NAND2_X1 U12851 ( .A1(n19203), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U12853 ( .A1(n10021), .A2(n20915), .ZN(n10066) );
  NAND2_X1 U12854 ( .A1(n10066), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10026) );
  INV_X1 U12855 ( .A(n10745), .ZN(n10024) );
  NAND2_X1 U12856 ( .A1(n13192), .A2(n10925), .ZN(n10919) );
  NAND2_X1 U12857 ( .A1(n13238), .A2(n9585), .ZN(n10023) );
  NAND2_X1 U12858 ( .A1(n10024), .A2(n9663), .ZN(n10027) );
  NOR2_X1 U12859 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16369) );
  NAND2_X1 U12860 ( .A1(n10026), .A2(n10025), .ZN(n10043) );
  INV_X1 U12861 ( .A(n10043), .ZN(n10041) );
  INV_X2 U12862 ( .A(n19849), .ZN(n10566) );
  NAND2_X1 U12863 ( .A1(n10027), .A2(n10566), .ZN(n10034) );
  NAND3_X1 U12864 ( .A1(n13107), .A2(n10009), .A3(n19230), .ZN(n10033) );
  NAND3_X1 U12865 ( .A1(n10022), .A2(n10017), .A3(n12376), .ZN(n10029) );
  NAND2_X1 U12866 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  INV_X1 U12867 ( .A(n10925), .ZN(n10913) );
  NOR2_X1 U12868 ( .A1(n10913), .A2(n12350), .ZN(n10036) );
  AND2_X4 U12869 ( .A1(n10927), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10807) );
  INV_X1 U12870 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10037) );
  INV_X2 U12871 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13789) );
  OAI22_X1 U12872 ( .A1(n10070), .A2(n10037), .B1(n13789), .B2(n13547), .ZN(
        n10038) );
  AOI21_X1 U12873 ( .B1(n9615), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10038), .ZN(
        n10039) );
  INV_X1 U12874 ( .A(n10042), .ZN(n10040) );
  NAND2_X1 U12875 ( .A1(n10041), .A2(n10040), .ZN(n10065) );
  NAND2_X1 U12876 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  AND2_X2 U12877 ( .A1(n10065), .A2(n10044), .ZN(n10097) );
  NOR2_X1 U12878 ( .A1(n10047), .A2(n10046), .ZN(n10926) );
  OAI21_X1 U12879 ( .B1(n10926), .B2(n10048), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10049) );
  INV_X1 U12880 ( .A(n10049), .ZN(n10050) );
  INV_X1 U12881 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U12882 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10053) );
  INV_X1 U12883 ( .A(n16369), .ZN(n10061) );
  NAND4_X1 U12884 ( .A1(n20915), .A2(n10054), .A3(n10053), .A4(n10061), .ZN(
        n10056) );
  NAND2_X1 U12885 ( .A1(n10058), .A2(n10057), .ZN(n10092) );
  AND2_X1 U12886 ( .A1(n10059), .A2(n10925), .ZN(n10060) );
  OAI22_X1 U12887 ( .A1(n10066), .A2(n10060), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10807), .ZN(n10064) );
  OAI22_X1 U12888 ( .A1(n13783), .A2(n19716), .B1(n10061), .B2(n19833), .ZN(
        n10062) );
  INV_X1 U12889 ( .A(n10062), .ZN(n10063) );
  NAND2_X1 U12890 ( .A1(n10064), .A2(n10063), .ZN(n10093) );
  NAND2_X1 U12891 ( .A1(n10097), .A2(n10101), .ZN(n10090) );
  NAND2_X1 U12892 ( .A1(n10090), .A2(n10065), .ZN(n10086) );
  NAND2_X1 U12894 ( .A1(n10067), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10069) );
  AOI21_X1 U12895 ( .B1(n19716), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10068) );
  INV_X1 U12896 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10934) );
  INV_X1 U12897 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n13281) );
  INV_X1 U12898 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19201) );
  OAI22_X1 U12899 ( .A1(n10841), .A2(n13281), .B1(n13789), .B2(n19201), .ZN(
        n10071) );
  OAI21_X2 U12900 ( .B1(n10774), .B2(n10934), .A(n10072), .ZN(n10074) );
  NAND2_X1 U12901 ( .A1(n10087), .A2(n10074), .ZN(n10073) );
  NAND2_X1 U12902 ( .A1(n10086), .A2(n10073), .ZN(n10077) );
  INV_X1 U12903 ( .A(n10087), .ZN(n10075) );
  NAND2_X1 U12904 ( .A1(n10075), .A2(n10088), .ZN(n10076) );
  NAND2_X1 U12905 ( .A1(n10067), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10079) );
  NAND2_X1 U12906 ( .A1(n16369), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10078) );
  INV_X1 U12907 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13806) );
  INV_X1 U12908 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10081) );
  INV_X1 U12909 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10080) );
  OAI22_X1 U12910 ( .A1(n10841), .A2(n10081), .B1(n13789), .B2(n10080), .ZN(
        n10082) );
  AOI21_X1 U12911 ( .B1(n10807), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10082), .ZN(
        n10083) );
  XNOR2_X2 U12912 ( .A(n10750), .B(n10085), .ZN(n10748) );
  INV_X1 U12914 ( .A(n10091), .ZN(n10096) );
  INV_X1 U12915 ( .A(n10092), .ZN(n10095) );
  INV_X1 U12916 ( .A(n10093), .ZN(n10094) );
  INV_X1 U12917 ( .A(n19306), .ZN(n19303) );
  INV_X1 U12918 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10103) );
  INV_X1 U12919 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10102) );
  INV_X1 U12920 ( .A(n10101), .ZN(n10098) );
  INV_X1 U12921 ( .A(n9606), .ZN(n10104) );
  NAND2_X1 U12922 ( .A1(n10098), .A2(n10104), .ZN(n10099) );
  OAI22_X1 U12923 ( .A1(n19303), .A2(n10103), .B1(n10102), .B2(n19274), .ZN(
        n10109) );
  INV_X1 U12924 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10107) );
  INV_X1 U12925 ( .A(n19058), .ZN(n10105) );
  INV_X1 U12926 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10106) );
  OAI22_X1 U12927 ( .A1(n10107), .A2(n10183), .B1(n10184), .B2(n10106), .ZN(
        n10108) );
  NOR2_X1 U12928 ( .A1(n10109), .A2(n10108), .ZN(n10138) );
  INV_X1 U12929 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10111) );
  AND2_X2 U12930 ( .A1(n13450), .A2(n9595), .ZN(n10129) );
  AND2_X2 U12931 ( .A1(n10129), .A2(n10118), .ZN(n10283) );
  INV_X1 U12932 ( .A(n10283), .ZN(n19398) );
  AND2_X2 U12933 ( .A1(n10125), .A2(n10130), .ZN(n10181) );
  NAND2_X1 U12934 ( .A1(n10181), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10110) );
  OAI211_X1 U12935 ( .C1(n10111), .C2(n19398), .A(n10110), .B(n19849), .ZN(
        n10115) );
  INV_X1 U12936 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10113) );
  INV_X1 U12937 ( .A(n10290), .ZN(n19334) );
  NAND2_X1 U12938 ( .A1(n10125), .A2(n10118), .ZN(n19503) );
  INV_X1 U12939 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10112) );
  OAI22_X1 U12940 ( .A1(n10113), .A2(n19334), .B1(n19503), .B2(n10112), .ZN(
        n10114) );
  NOR2_X1 U12941 ( .A1(n10115), .A2(n10114), .ZN(n10137) );
  AND2_X2 U12942 ( .A1(n10125), .A2(n10128), .ZN(n10289) );
  INV_X1 U12943 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12944 ( .A1(n10119), .A2(n10118), .ZN(n19632) );
  NAND2_X1 U12945 ( .A1(n10119), .A2(n10124), .ZN(n10189) );
  INV_X1 U12946 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10120) );
  OAI22_X1 U12947 ( .A1(n10121), .A2(n19632), .B1(n10189), .B2(n10120), .ZN(
        n10122) );
  NOR2_X1 U12948 ( .A1(n10123), .A2(n10122), .ZN(n10136) );
  INV_X1 U12949 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12950 ( .A1(n10129), .A2(n10128), .ZN(n10182) );
  INV_X1 U12951 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19213) );
  OAI22_X1 U12952 ( .A1(n10132), .A2(n10182), .B1(n10322), .B2(n19213), .ZN(
        n10133) );
  NOR2_X1 U12953 ( .A1(n10134), .A2(n10133), .ZN(n10135) );
  NAND4_X1 U12954 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10180) );
  AND2_X2 U12955 ( .A1(n12649), .A2(n9956), .ZN(n12512) );
  AOI22_X1 U12956 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n9593), .B1(
        n12512), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10142) );
  AND2_X2 U12957 ( .A1(n20914), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10604) );
  AOI22_X1 U12958 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10604), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10141) );
  AND2_X2 U12959 ( .A1(n12490), .A2(n10266), .ZN(n12478) );
  AOI22_X1 U12960 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U12961 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10139) );
  NAND4_X1 U12962 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10152) );
  NOR2_X1 U12963 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10144) );
  AND2_X2 U12964 ( .A1(n12491), .A2(n10144), .ZN(n12513) );
  AOI22_X1 U12965 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10159), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10150) );
  AND2_X2 U12966 ( .A1(n15662), .A2(n12491), .ZN(n12514) );
  AOI22_X1 U12967 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U12968 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n10259), .ZN(n10148) );
  AND2_X2 U12969 ( .A1(n10001), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10168) );
  AND2_X2 U12970 ( .A1(n20914), .A2(n10266), .ZN(n15682) );
  AOI22_X1 U12971 ( .A1(n10168), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10147) );
  NAND4_X1 U12972 ( .A1(n10150), .A2(n10149), .A3(n10148), .A4(n10147), .ZN(
        n10151) );
  AOI22_X1 U12973 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12478), .B1(
        n10211), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U12974 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U12975 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10168), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U12976 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10604), .B1(
        n9593), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U12977 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10166) );
  AOI22_X1 U12978 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n15682), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U12979 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U12980 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12514), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U12981 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10160), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10161) );
  NAND4_X1 U12982 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10165) );
  NAND2_X1 U12983 ( .A1(n10566), .A2(n10569), .ZN(n10167) );
  OR2_X1 U12984 ( .A1(n13306), .A2(n10167), .ZN(n10863) );
  AOI22_X1 U12985 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10211), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U12986 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U12987 ( .A1(n10168), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U12988 ( .A1(n12507), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10169) );
  NAND4_X1 U12989 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10178) );
  AOI22_X1 U12990 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U12991 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U12992 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U12993 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U12994 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NAND2_X1 U12995 ( .A1(n10863), .A2(n10864), .ZN(n10179) );
  NAND2_X1 U12996 ( .A1(n10180), .A2(n10179), .ZN(n10208) );
  INV_X1 U12997 ( .A(n10322), .ZN(n10282) );
  AOI22_X1 U12998 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10181), .B1(
        n10282), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10188) );
  INV_X1 U12999 ( .A(n10182), .ZN(n19366) );
  AOI22_X1 U13000 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19593), .B1(
        n10289), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10186) );
  INV_X1 U13001 ( .A(n19503), .ZN(n10288) );
  AOI22_X1 U13002 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19270), .B1(
        n10288), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10185) );
  NAND4_X1 U13003 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10207) );
  AOI22_X1 U13004 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n15725), .B1(
        n10283), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U13005 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19636), .B1(
        n19527), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10191) );
  NAND4_X1 U13006 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10206) );
  AOI22_X1 U13007 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13008 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13009 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13010 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n9593), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10195) );
  NAND4_X1 U13011 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10204) );
  AOI22_X1 U13012 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10300), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13013 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13014 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10159), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13015 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10199) );
  NAND4_X1 U13016 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  INV_X1 U13017 ( .A(n10239), .ZN(n10583) );
  NAND2_X1 U13018 ( .A1(n10583), .A2(n10566), .ZN(n10205) );
  OAI21_X2 U13019 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(n10209) );
  NAND2_X1 U13020 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NAND2_X1 U13021 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10215) );
  NAND2_X1 U13022 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10214) );
  NAND2_X1 U13023 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10213) );
  NAND2_X1 U13024 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10212) );
  AOI22_X1 U13025 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U13026 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U13027 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U13028 ( .A1(n10259), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10216) );
  AND4_X1 U13029 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10226) );
  NAND2_X1 U13030 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10223) );
  NAND2_X1 U13031 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13032 ( .A1(n10168), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U13033 ( .A1(n10153), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10220) );
  AOI22_X1 U13034 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U13035 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10351) );
  INV_X1 U13036 ( .A(n10351), .ZN(n10402) );
  INV_X2 U13037 ( .A(n10402), .ZN(n14320) );
  XNOR2_X1 U13038 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10501) );
  NAND2_X1 U13039 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19833), .ZN(
        n10489) );
  INV_X1 U13040 ( .A(n10489), .ZN(n10228) );
  NAND2_X1 U13041 ( .A1(n10501), .A2(n10228), .ZN(n10230) );
  NAND2_X1 U13042 ( .A1(n19824), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U13043 ( .A1(n10230), .A2(n10229), .ZN(n10235) );
  MUX2_X1 U13044 ( .A(n12395), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10234) );
  XNOR2_X1 U13045 ( .A(n10235), .B(n10234), .ZN(n10484) );
  INV_X1 U13046 ( .A(n10484), .ZN(n10524) );
  INV_X1 U13047 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13434) );
  MUX2_X1 U13048 ( .A(n10503), .B(n13434), .S(n10477), .Z(n10245) );
  NOR2_X1 U13049 ( .A1(n10560), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10247) );
  INV_X1 U13050 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13548) );
  NAND2_X1 U13051 ( .A1(n10247), .A2(n13548), .ZN(n10233) );
  NAND2_X1 U13052 ( .A1(n10569), .A2(n10560), .ZN(n10232) );
  NAND2_X1 U13053 ( .A1(n10233), .A2(n10232), .ZN(n10251) );
  NAND2_X1 U13054 ( .A1(n10235), .A2(n10234), .ZN(n10237) );
  NAND2_X1 U13055 ( .A1(n12395), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10236) );
  NAND2_X1 U13056 ( .A1(n10237), .A2(n10236), .ZN(n10269) );
  XNOR2_X1 U13057 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10268) );
  XNOR2_X1 U13058 ( .A(n10269), .B(n10268), .ZN(n10534) );
  NAND2_X1 U13059 ( .A1(n10498), .A2(n10350), .ZN(n10241) );
  NOR2_X2 U13060 ( .A1(n10244), .A2(n10242), .ZN(n10272) );
  INV_X1 U13061 ( .A(n10272), .ZN(n10275) );
  NAND2_X1 U13062 ( .A1(n10244), .A2(n10242), .ZN(n10243) );
  NAND2_X1 U13063 ( .A1(n10275), .A2(n10243), .ZN(n13451) );
  OAI21_X1 U13064 ( .B1(n10245), .B2(n10251), .A(n10244), .ZN(n13438) );
  OAI21_X1 U13065 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19833), .A(
        n10489), .ZN(n10526) );
  MUX2_X1 U13066 ( .A(n13306), .B(n10526), .S(n12350), .Z(n10246) );
  NAND2_X1 U13067 ( .A1(n10246), .A2(n10350), .ZN(n10249) );
  INV_X1 U13068 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U13069 ( .A1(n10249), .A2(n10248), .ZN(n19051) );
  INV_X1 U13070 ( .A(n19051), .ZN(n10250) );
  NAND2_X1 U13071 ( .A1(n10250), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13305) );
  INV_X1 U13072 ( .A(n10251), .ZN(n10253) );
  NAND3_X1 U13073 ( .A1(n10477), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U13074 ( .A1(n10253), .A2(n10252), .ZN(n13544) );
  NOR2_X1 U13075 ( .A1(n13305), .A2(n13544), .ZN(n10254) );
  NAND2_X1 U13076 ( .A1(n13305), .A2(n13544), .ZN(n13296) );
  OAI21_X1 U13077 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10254), .A(
        n13296), .ZN(n13285) );
  XNOR2_X1 U13078 ( .A(n13438), .B(n10934), .ZN(n13284) );
  OR2_X1 U13079 ( .A1(n13285), .A2(n13284), .ZN(n13287) );
  OAI21_X1 U13080 ( .B1(n13438), .B2(n10934), .A(n13287), .ZN(n13801) );
  AOI22_X1 U13081 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13082 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13083 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13084 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U13085 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10265) );
  AOI22_X1 U13086 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13087 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13088 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13089 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10260) );
  NAND4_X1 U13090 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n10264) );
  NOR2_X1 U13091 ( .A1(n10266), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10267) );
  AOI21_X1 U13092 ( .B1(n10269), .B2(n10268), .A(n10267), .ZN(n10486) );
  NOR2_X1 U13093 ( .A1(n16358), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10270) );
  AND2_X1 U13094 ( .A1(n10486), .A2(n10270), .ZN(n10540) );
  INV_X1 U13095 ( .A(n10540), .ZN(n10271) );
  MUX2_X1 U13096 ( .A(n10589), .B(n10271), .S(n12350), .Z(n10499) );
  INV_X1 U13097 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13403) );
  MUX2_X1 U13098 ( .A(n10499), .B(n13403), .S(n10477), .Z(n10273) );
  INV_X1 U13099 ( .A(n10310), .ZN(n10277) );
  INV_X1 U13100 ( .A(n10273), .ZN(n10274) );
  NAND2_X1 U13101 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NAND2_X1 U13102 ( .A1(n10277), .A2(n10276), .ZN(n13428) );
  XNOR2_X1 U13103 ( .A(n13428), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13943) );
  INV_X1 U13104 ( .A(n13428), .ZN(n10278) );
  NAND2_X1 U13105 ( .A1(n10278), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10279) );
  NAND2_X1 U13106 ( .A1(n10280), .A2(n10279), .ZN(n15617) );
  AOI22_X1 U13107 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19366), .B1(
        n10281), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13108 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19270), .B1(
        n19593), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U13109 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10282), .B1(
        n10181), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13110 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10283), .B1(
        n15725), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13111 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19306), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13112 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19527), .B1(
        n19636), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13113 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n10288), .B1(
        n10289), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13114 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10290), .B1(
        n10291), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U13115 ( .A1(n9877), .A2(n9660), .ZN(n10309) );
  AOI22_X1 U13116 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13117 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13118 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13119 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10296) );
  NAND4_X1 U13120 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10306) );
  AOI22_X1 U13121 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13122 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13123 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13124 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10301) );
  NAND4_X1 U13125 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  INV_X1 U13126 ( .A(n10593), .ZN(n10307) );
  NAND2_X1 U13127 ( .A1(n10307), .A2(n10566), .ZN(n10308) );
  XNOR2_X2 U13128 ( .A(n10876), .B(n10315), .ZN(n10860) );
  NAND2_X1 U13129 ( .A1(n10860), .A2(n10402), .ZN(n10311) );
  INV_X1 U13130 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19031) );
  MUX2_X1 U13131 ( .A(n19031), .B(n10593), .S(n10350), .Z(n10342) );
  XNOR2_X1 U13132 ( .A(n10310), .B(n10342), .ZN(n19033) );
  INV_X1 U13133 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U13134 ( .A1(n15617), .A2(n15618), .ZN(n10314) );
  NAND2_X1 U13135 ( .A1(n10312), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10313) );
  INV_X1 U13136 ( .A(n10876), .ZN(n10316) );
  AOI22_X1 U13137 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19527), .B1(
        n19636), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13138 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19306), .B1(
        n9653), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13139 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10290), .B1(
        n10291), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13140 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10283), .B1(
        n15725), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10317) );
  NAND4_X1 U13141 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10329) );
  AOI22_X1 U13142 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19593), .B1(
        n10289), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13143 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19270), .B1(
        n10288), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13144 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19366), .B1(
        n10281), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10325) );
  INV_X1 U13145 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19228) );
  INV_X1 U13146 ( .A(n10181), .ZN(n19444) );
  INV_X1 U13147 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10321) );
  OAI22_X1 U13148 ( .A1(n19228), .A2(n10322), .B1(n19444), .B2(n10321), .ZN(
        n10323) );
  INV_X1 U13149 ( .A(n10323), .ZN(n10324) );
  NAND4_X1 U13150 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10328) );
  AOI22_X1 U13151 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13152 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13153 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13154 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10330) );
  NAND4_X1 U13155 ( .A1(n10333), .A2(n10332), .A3(n10331), .A4(n10330), .ZN(
        n10339) );
  AOI22_X1 U13156 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13157 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13158 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13159 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10334) );
  NAND4_X1 U13160 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  NOR2_X1 U13161 ( .A1(n10339), .A2(n10338), .ZN(n10596) );
  NAND2_X1 U13162 ( .A1(n10596), .A2(n10566), .ZN(n10340) );
  XNOR2_X1 U13163 ( .A(n10887), .B(n10885), .ZN(n10880) );
  NAND2_X1 U13164 ( .A1(n10880), .A2(n10402), .ZN(n10344) );
  MUX2_X1 U13165 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n10596), .S(n10350), .Z(
        n10348) );
  XNOR2_X1 U13166 ( .A(n10349), .B(n10348), .ZN(n19018) );
  NAND2_X1 U13167 ( .A1(n10344), .A2(n19018), .ZN(n10345) );
  INV_X1 U13168 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15357) );
  XNOR2_X1 U13169 ( .A(n10345), .B(n15357), .ZN(n15355) );
  NAND2_X1 U13170 ( .A1(n15356), .A2(n15355), .ZN(n10347) );
  NAND2_X1 U13171 ( .A1(n10345), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10346) );
  INV_X1 U13172 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10352) );
  MUX2_X1 U13173 ( .A(n10352), .B(n10351), .S(n10350), .Z(n10358) );
  NAND2_X1 U13174 ( .A1(n10359), .A2(n10358), .ZN(n10355) );
  INV_X1 U13175 ( .A(n10355), .ZN(n10354) );
  NAND2_X1 U13176 ( .A1(n10354), .A2(n10353), .ZN(n10366) );
  NAND2_X1 U13177 ( .A1(n10369), .A2(n10356), .ZN(n10357) );
  NAND2_X1 U13178 ( .A1(n10366), .A2(n10357), .ZN(n13414) );
  INV_X1 U13179 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16315) );
  NOR2_X1 U13180 ( .A1(n10363), .A2(n16315), .ZN(n16240) );
  OR2_X1 U13181 ( .A1(n10359), .A2(n10358), .ZN(n10360) );
  NAND2_X1 U13182 ( .A1(n10369), .A2(n10360), .ZN(n19010) );
  INV_X1 U13183 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16304) );
  NOR2_X1 U13184 ( .A1(n19010), .A2(n16304), .ZN(n16236) );
  NAND2_X1 U13185 ( .A1(n10363), .A2(n16315), .ZN(n16238) );
  NAND2_X1 U13186 ( .A1(n19010), .A2(n16304), .ZN(n16237) );
  AND2_X1 U13187 ( .A1(n16238), .A2(n16237), .ZN(n10364) );
  NAND2_X1 U13188 ( .A1(n10477), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10365) );
  XNOR2_X1 U13189 ( .A(n10366), .B(n10365), .ZN(n19000) );
  NAND2_X1 U13190 ( .A1(n19000), .A2(n14320), .ZN(n10441) );
  INV_X1 U13191 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15563) );
  AND2_X1 U13192 ( .A1(n10477), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10370) );
  INV_X1 U13193 ( .A(n10366), .ZN(n10368) );
  NAND2_X1 U13194 ( .A1(n10368), .A2(n10367), .ZN(n10371) );
  INV_X1 U13195 ( .A(n10467), .ZN(n10424) );
  AOI21_X1 U13196 ( .B1(n10370), .B2(n10371), .A(n10424), .ZN(n10372) );
  NOR2_X2 U13197 ( .A1(n10371), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10373) );
  INV_X1 U13198 ( .A(n10373), .ZN(n10374) );
  AOI21_X1 U13199 ( .B1(n13626), .B2(n14320), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16221) );
  INV_X1 U13200 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U13201 ( .A1(n13541), .A2(n10373), .ZN(n10377) );
  NAND2_X1 U13202 ( .A1(n10377), .A2(n10467), .ZN(n10376) );
  AND3_X1 U13203 ( .A1(n10477), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10374), .ZN(
        n10375) );
  OR2_X1 U13204 ( .A1(n10376), .A2(n10375), .ZN(n10442) );
  INV_X1 U13205 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15564) );
  OAI21_X1 U13206 ( .B1(n10442), .B2(n10402), .A(n15564), .ZN(n15559) );
  NAND2_X1 U13207 ( .A1(n10477), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10379) );
  AND2_X2 U13208 ( .A1(n10376), .A2(n10379), .ZN(n10408) );
  INV_X1 U13209 ( .A(n10377), .ZN(n10378) );
  NOR2_X1 U13210 ( .A1(n10379), .A2(n10378), .ZN(n10380) );
  OR2_X1 U13211 ( .A1(n10408), .A2(n10380), .ZN(n18977) );
  NOR2_X1 U13212 ( .A1(n18977), .A2(n10402), .ZN(n10444) );
  INV_X1 U13213 ( .A(n10444), .ZN(n10381) );
  NAND2_X1 U13214 ( .A1(n10381), .A2(n15539), .ZN(n10439) );
  AND2_X1 U13215 ( .A1(n15559), .A2(n10439), .ZN(n14170) );
  NAND2_X1 U13216 ( .A1(n10477), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10407) );
  OAI21_X1 U13217 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n10477), .ZN(n10382) );
  INV_X1 U13218 ( .A(n10414), .ZN(n10383) );
  NAND2_X1 U13219 ( .A1(n10383), .A2(n9872), .ZN(n10399) );
  AND2_X1 U13220 ( .A1(n10477), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10398) );
  NOR2_X2 U13221 ( .A1(n10399), .A2(n10398), .ZN(n10393) );
  NAND2_X1 U13222 ( .A1(n10477), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10394) );
  AND2_X2 U13223 ( .A1(n10393), .A2(n10394), .ZN(n10392) );
  NAND2_X1 U13224 ( .A1(n10477), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10419) );
  INV_X1 U13225 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U13226 ( .A1(n10477), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10430) );
  AND2_X1 U13227 ( .A1(n10477), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10384) );
  OR2_X2 U13228 ( .A1(n10434), .A2(n10384), .ZN(n10466) );
  NAND2_X1 U13229 ( .A1(n10434), .A2(n10384), .ZN(n10385) );
  INV_X1 U13230 ( .A(n10387), .ZN(n10389) );
  NAND3_X1 U13231 ( .A1(n10428), .A2(n10477), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n10388) );
  NAND2_X1 U13232 ( .A1(n10389), .A2(n10388), .ZN(n13057) );
  INV_X1 U13233 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14199) );
  OAI21_X1 U13234 ( .B1(n13057), .B2(n10402), .A(n14199), .ZN(n14185) );
  NAND3_X1 U13235 ( .A1(n10414), .A2(n10477), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n10390) );
  OAI211_X1 U13236 ( .C1(n10414), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10467), .B(
        n10390), .ZN(n18958) );
  OR2_X1 U13237 ( .A1(n18958), .A2(n10402), .ZN(n10391) );
  XNOR2_X1 U13238 ( .A(n10391), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14176) );
  INV_X1 U13239 ( .A(n10392), .ZN(n10421) );
  INV_X1 U13240 ( .A(n10393), .ZN(n10401) );
  INV_X1 U13241 ( .A(n10394), .ZN(n10395) );
  NAND2_X1 U13242 ( .A1(n10401), .A2(n10395), .ZN(n10396) );
  NAND2_X1 U13243 ( .A1(n10421), .A2(n10396), .ZN(n18930) );
  OR2_X1 U13244 ( .A1(n18930), .A2(n10402), .ZN(n10397) );
  INV_X1 U13245 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U13246 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  NAND2_X1 U13247 ( .A1(n10401), .A2(n10400), .ZN(n18947) );
  OR2_X1 U13248 ( .A1(n18947), .A2(n10402), .ZN(n10403) );
  INV_X1 U13249 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U13250 ( .A1(n10403), .A2(n15507), .ZN(n14179) );
  NAND2_X1 U13251 ( .A1(n10477), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10405) );
  MUX2_X1 U13252 ( .A(n10405), .B(n10477), .S(n10410), .Z(n10406) );
  INV_X1 U13253 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13842) );
  NAND2_X1 U13254 ( .A1(n10410), .A2(n13842), .ZN(n10413) );
  NAND2_X1 U13255 ( .A1(n13954), .A2(n14320), .ZN(n10456) );
  INV_X1 U13256 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16198) );
  NAND2_X1 U13257 ( .A1(n10456), .A2(n16198), .ZN(n16199) );
  NOR2_X1 U13258 ( .A1(n10408), .A2(n10407), .ZN(n10409) );
  OR2_X1 U13259 ( .A1(n10410), .A2(n10409), .ZN(n13086) );
  INV_X1 U13260 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10411) );
  OAI21_X1 U13261 ( .B1(n13086), .B2(n10402), .A(n10411), .ZN(n15332) );
  AND2_X1 U13262 ( .A1(n10477), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U13263 ( .A1(n10413), .A2(n10412), .ZN(n10415) );
  NAND2_X1 U13264 ( .A1(n10415), .A2(n10414), .ZN(n18966) );
  OR2_X1 U13265 ( .A1(n18966), .A2(n10402), .ZN(n10416) );
  INV_X1 U13266 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U13267 ( .A1(n10416), .A2(n14226), .ZN(n15322) );
  NAND4_X1 U13268 ( .A1(n14179), .A2(n16199), .A3(n15332), .A4(n15322), .ZN(
        n10417) );
  NOR2_X1 U13269 ( .A1(n15295), .A2(n10417), .ZN(n10423) );
  INV_X1 U13270 ( .A(n10418), .ZN(n10426) );
  INV_X1 U13271 ( .A(n10419), .ZN(n10420) );
  NAND2_X1 U13272 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  NAND2_X1 U13273 ( .A1(n10426), .A2(n10422), .ZN(n18918) );
  INV_X1 U13274 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15471) );
  OAI21_X1 U13275 ( .B1(n18918), .B2(n10402), .A(n15471), .ZN(n15287) );
  AND2_X1 U13276 ( .A1(n10423), .A2(n15287), .ZN(n10429) );
  AND2_X1 U13277 ( .A1(n10477), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10425) );
  AOI21_X1 U13278 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n10427) );
  NAND2_X1 U13279 ( .A1(n10428), .A2(n10427), .ZN(n15060) );
  INV_X1 U13280 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13281 ( .A1(n10447), .A2(n10816), .ZN(n14221) );
  NAND4_X1 U13282 ( .A1(n14185), .A2(n14176), .A3(n10429), .A4(n14221), .ZN(
        n15274) );
  INV_X1 U13283 ( .A(n10430), .ZN(n10431) );
  NAND2_X1 U13284 ( .A1(n10432), .A2(n10431), .ZN(n10433) );
  NAND2_X1 U13285 ( .A1(n10434), .A2(n10433), .ZN(n15048) );
  OR2_X1 U13286 ( .A1(n15048), .A2(n10402), .ZN(n10435) );
  INV_X1 U13287 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15461) );
  NAND2_X1 U13288 ( .A1(n10435), .A2(n15461), .ZN(n15273) );
  INV_X1 U13289 ( .A(n15273), .ZN(n10436) );
  AND2_X1 U13290 ( .A1(n14170), .A2(n9668), .ZN(n10438) );
  NAND2_X1 U13291 ( .A1(n15557), .A2(n10438), .ZN(n15249) );
  NAND2_X1 U13292 ( .A1(n10467), .A2(n14320), .ZN(n15250) );
  INV_X1 U13293 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15402) );
  NOR2_X1 U13294 ( .A1(n15250), .A2(n15402), .ZN(n10463) );
  INV_X1 U13295 ( .A(n10439), .ZN(n15546) );
  AND2_X1 U13296 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U13297 ( .A1(n13626), .A2(n10440), .ZN(n16219) );
  OR2_X1 U13298 ( .A1(n10441), .A2(n15563), .ZN(n16217) );
  INV_X1 U13299 ( .A(n10442), .ZN(n18989) );
  AND2_X1 U13300 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13301 ( .A1(n18989), .A2(n10443), .ZN(n15558) );
  NAND3_X1 U13302 ( .A1(n16219), .A2(n16217), .A3(n15558), .ZN(n15543) );
  AND2_X1 U13303 ( .A1(n10444), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15547) );
  NOR2_X1 U13304 ( .A1(n15543), .A2(n15547), .ZN(n10445) );
  NAND2_X1 U13305 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10446) );
  NOR2_X1 U13306 ( .A1(n13057), .A2(n10446), .ZN(n14184) );
  INV_X1 U13307 ( .A(n10447), .ZN(n10448) );
  NAND2_X1 U13308 ( .A1(n10448), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14222) );
  INV_X1 U13309 ( .A(n18918), .ZN(n10450) );
  AND2_X1 U13310 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10449) );
  NAND2_X1 U13311 ( .A1(n10450), .A2(n10449), .ZN(n15286) );
  AND2_X1 U13312 ( .A1(n15286), .A2(n15296), .ZN(n14182) );
  NAND2_X1 U13313 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10451) );
  OR2_X1 U13314 ( .A1(n18947), .A2(n10451), .ZN(n14178) );
  NAND2_X1 U13315 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10452) );
  OR2_X1 U13316 ( .A1(n18958), .A2(n10452), .ZN(n14177) );
  NAND2_X1 U13317 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10453) );
  INV_X1 U13318 ( .A(n13086), .ZN(n10455) );
  AND2_X1 U13319 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13320 ( .A1(n10455), .A2(n10454), .ZN(n15331) );
  AND4_X1 U13321 ( .A1(n14178), .A2(n14177), .A3(n15321), .A4(n15331), .ZN(
        n10458) );
  INV_X1 U13322 ( .A(n10456), .ZN(n10457) );
  NAND2_X1 U13323 ( .A1(n10457), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16200) );
  NAND4_X1 U13324 ( .A1(n14222), .A2(n14182), .A3(n10458), .A4(n16200), .ZN(
        n10459) );
  NOR2_X1 U13325 ( .A1(n14184), .A2(n10459), .ZN(n15275) );
  NAND2_X1 U13326 ( .A1(n14320), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10460) );
  OR2_X1 U13327 ( .A1(n15048), .A2(n10460), .ZN(n15272) );
  AND2_X1 U13328 ( .A1(n15275), .A2(n15272), .ZN(n15265) );
  AND2_X1 U13329 ( .A1(n14171), .A2(n15265), .ZN(n10462) );
  NAND3_X1 U13330 ( .A1(n13069), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14320), .ZN(n10461) );
  NAND2_X1 U13331 ( .A1(n10462), .A2(n10461), .ZN(n15247) );
  NOR2_X1 U13332 ( .A1(n10463), .A2(n15247), .ZN(n10464) );
  INV_X1 U13333 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15426) );
  AND2_X1 U13334 ( .A1(n15250), .A2(n15426), .ZN(n15238) );
  INV_X1 U13335 ( .A(n15238), .ZN(n10465) );
  NAND2_X1 U13336 ( .A1(n15250), .A2(n15402), .ZN(n15240) );
  NOR2_X2 U13337 ( .A1(n10466), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15018) );
  INV_X1 U13338 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U13339 ( .A1(n15018), .A2(n15005), .ZN(n15004) );
  OR2_X2 U13340 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n15004), .ZN(n16172) );
  NAND2_X2 U13341 ( .A1(n10467), .A2(n16172), .ZN(n14261) );
  AND3_X1 U13342 ( .A1(n10477), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n15004), .ZN(
        n10468) );
  NOR2_X1 U13343 ( .A1(n14261), .A2(n10468), .ZN(n14992) );
  NAND2_X1 U13344 ( .A1(n14992), .A2(n14320), .ZN(n10469) );
  INV_X1 U13345 ( .A(n10472), .ZN(n15197) );
  AND2_X1 U13346 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15365) );
  INV_X1 U13347 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15413) );
  OR2_X1 U13348 ( .A1(n10469), .A2(n15413), .ZN(n10471) );
  INV_X1 U13349 ( .A(n15250), .ZN(n10470) );
  NAND2_X1 U13350 ( .A1(n10470), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15222) );
  NAND2_X1 U13351 ( .A1(n10471), .A2(n15222), .ZN(n15198) );
  NAND2_X1 U13352 ( .A1(n9585), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16169) );
  NAND2_X2 U13353 ( .A1(n14261), .A2(n16169), .ZN(n16170) );
  NAND2_X1 U13354 ( .A1(n16170), .A2(n14320), .ZN(n15202) );
  NOR2_X1 U13355 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10475) );
  INV_X1 U13356 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14981) );
  NOR2_X1 U13357 ( .A1(n10350), .A2(n14981), .ZN(n10473) );
  NOR2_X2 U13358 ( .A1(n16170), .A2(n10473), .ZN(n10481) );
  AND2_X1 U13359 ( .A1(n16170), .A2(n10473), .ZN(n10474) );
  NOR2_X1 U13360 ( .A1(n10481), .A2(n10474), .ZN(n14983) );
  NAND2_X1 U13361 ( .A1(n14983), .A2(n14320), .ZN(n15204) );
  AOI21_X1 U13362 ( .B1(n9890), .B2(n10475), .A(n15204), .ZN(n10476) );
  NAND2_X1 U13363 ( .A1(n10477), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10480) );
  INV_X1 U13364 ( .A(n10480), .ZN(n10478) );
  XNOR2_X1 U13365 ( .A(n10481), .B(n10478), .ZN(n10479) );
  AOI21_X1 U13366 ( .B1(n10479), .B2(n14320), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15188) );
  INV_X1 U13367 ( .A(n14328), .ZN(n14332) );
  INV_X1 U13368 ( .A(n10479), .ZN(n16160) );
  INV_X1 U13369 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15364) );
  OR3_X2 U13370 ( .A1(n16160), .A2(n10402), .A3(n15364), .ZN(n15186) );
  NAND2_X1 U13371 ( .A1(n14332), .A2(n15186), .ZN(n10483) );
  NAND2_X1 U13372 ( .A1(n10481), .A2(n10480), .ZN(n14262) );
  INV_X1 U13373 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10849) );
  NOR2_X1 U13374 ( .A1(n10350), .A2(n10849), .ZN(n10482) );
  XNOR2_X1 U13375 ( .A(n14262), .B(n10482), .ZN(n12362) );
  INV_X1 U13376 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10953) );
  OAI21_X1 U13377 ( .B1(n12362), .B2(n10402), .A(n10953), .ZN(n14327) );
  XNOR2_X1 U13378 ( .A(n10483), .B(n9886), .ZN(n12142) );
  OR3_X1 U13379 ( .A1(n10540), .A2(n10534), .A3(n10484), .ZN(n10492) );
  NAND2_X1 U13380 ( .A1(n16358), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10485) );
  NAND2_X1 U13381 ( .A1(n10486), .A2(n10485), .ZN(n10488) );
  INV_X1 U13382 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13195) );
  NAND2_X1 U13383 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13195), .ZN(
        n10487) );
  NAND2_X1 U13384 ( .A1(n10488), .A2(n10487), .ZN(n10539) );
  XNOR2_X1 U13385 ( .A(n10501), .B(n10489), .ZN(n10527) );
  INV_X1 U13386 ( .A(n10492), .ZN(n10490) );
  NAND2_X1 U13387 ( .A1(n10527), .A2(n10490), .ZN(n10491) );
  OAI21_X1 U13388 ( .B1(n10526), .B2(n10492), .A(n16340), .ZN(n10493) );
  INV_X1 U13389 ( .A(n10493), .ZN(n10496) );
  NAND2_X1 U13390 ( .A1(n15669), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13391 ( .A1(n10495), .A2(n13195), .ZN(n13191) );
  INV_X1 U13392 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13111) );
  OAI21_X1 U13393 ( .B1(n10211), .B2(n13191), .A(n13111), .ZN(n19829) );
  MUX2_X1 U13394 ( .A(n10496), .B(n19829), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15905) );
  NOR2_X1 U13395 ( .A1(n16339), .A2(n10566), .ZN(n10497) );
  NAND2_X1 U13396 ( .A1(n15905), .A2(n10497), .ZN(n10507) );
  INV_X1 U13397 ( .A(n10498), .ZN(n10500) );
  NAND2_X1 U13398 ( .A1(n10500), .A2(n10499), .ZN(n10522) );
  INV_X1 U13399 ( .A(n10501), .ZN(n10525) );
  NOR2_X1 U13400 ( .A1(n10525), .A2(n10526), .ZN(n10502) );
  NOR2_X1 U13401 ( .A1(n10503), .A2(n10502), .ZN(n10504) );
  OAI21_X1 U13402 ( .B1(n10522), .B2(n10504), .A(n10539), .ZN(n19837) );
  INV_X1 U13403 ( .A(n16339), .ZN(n10505) );
  AND2_X1 U13404 ( .A1(n10566), .A2(n19203), .ZN(n10510) );
  NAND2_X1 U13405 ( .A1(n10505), .A2(n10510), .ZN(n10910) );
  NAND2_X1 U13406 ( .A1(n10507), .A2(n10506), .ZN(n12126) );
  INV_X1 U13407 ( .A(n12126), .ZN(n10553) );
  OAI21_X1 U13408 ( .B1(n10508), .B2(n10509), .A(n10510), .ZN(n10917) );
  NAND2_X1 U13409 ( .A1(n10512), .A2(n15717), .ZN(n10513) );
  NAND2_X1 U13410 ( .A1(n10511), .A2(n10513), .ZN(n10517) );
  NAND2_X1 U13411 ( .A1(n10009), .A2(n10566), .ZN(n10911) );
  NAND2_X1 U13412 ( .A1(n10911), .A2(n9627), .ZN(n10514) );
  NAND3_X1 U13413 ( .A1(n10514), .A2(n15699), .A3(n19230), .ZN(n10515) );
  NAND2_X1 U13414 ( .A1(n10515), .A2(n15717), .ZN(n10516) );
  NAND4_X1 U13415 ( .A1(n10518), .A2(n10917), .A3(n10517), .A4(n10516), .ZN(
        n10912) );
  NAND2_X1 U13416 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19861) );
  INV_X1 U13417 ( .A(n19861), .ZN(n19853) );
  NAND2_X1 U13418 ( .A1(n20893), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19864) );
  INV_X2 U13419 ( .A(n19864), .ZN(n19867) );
  NAND2_X1 U13420 ( .A1(n19867), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19781) );
  NOR2_X1 U13421 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19727) );
  INV_X1 U13422 ( .A(n19727), .ZN(n19736) );
  NAND3_X1 U13423 ( .A1(n20893), .A2(n19778), .A3(n19736), .ZN(n19848) );
  NOR2_X1 U13424 ( .A1(n19853), .A2(n19848), .ZN(n13108) );
  OR2_X1 U13425 ( .A1(n10912), .A2(n10519), .ZN(n13184) );
  AND3_X1 U13426 ( .A1(n10520), .A2(n16340), .A3(n19861), .ZN(n10521) );
  NOR2_X1 U13427 ( .A1(n13184), .A2(n10521), .ZN(n10552) );
  NAND2_X1 U13428 ( .A1(n10522), .A2(n12350), .ZN(n10538) );
  NAND2_X1 U13429 ( .A1(n19849), .A2(n10544), .ZN(n10523) );
  MUX2_X1 U13430 ( .A(n10523), .B(n12350), .S(n10524), .Z(n10533) );
  NAND2_X1 U13431 ( .A1(n13192), .A2(n10524), .ZN(n10531) );
  OAI21_X1 U13432 ( .B1(n10525), .B2(n10526), .A(n12364), .ZN(n10530) );
  NAND2_X1 U13433 ( .A1(n10566), .A2(n10526), .ZN(n10528) );
  NAND3_X1 U13434 ( .A1(n10528), .A2(n9627), .A3(n10527), .ZN(n10529) );
  NAND3_X1 U13435 ( .A1(n10531), .A2(n10530), .A3(n10529), .ZN(n10532) );
  NAND2_X1 U13436 ( .A1(n10533), .A2(n10532), .ZN(n10536) );
  INV_X1 U13437 ( .A(n10534), .ZN(n10535) );
  NAND2_X1 U13438 ( .A1(n10536), .A2(n10535), .ZN(n10537) );
  NAND2_X1 U13439 ( .A1(n10538), .A2(n10537), .ZN(n10542) );
  AOI21_X1 U13440 ( .B1(n12364), .B2(n10540), .A(n10545), .ZN(n10541) );
  NAND2_X1 U13441 ( .A1(n10542), .A2(n10541), .ZN(n10543) );
  MUX2_X1 U13442 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10543), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10547) );
  INV_X1 U13443 ( .A(n10544), .ZN(n19846) );
  NAND2_X1 U13444 ( .A1(n19846), .A2(n10545), .ZN(n10546) );
  NAND3_X1 U13445 ( .A1(n13200), .A2(n10914), .A3(n13108), .ZN(n10551) );
  INV_X1 U13446 ( .A(n10547), .ZN(n10549) );
  INV_X1 U13447 ( .A(n13200), .ZN(n10548) );
  OAI211_X1 U13448 ( .C1(n10549), .C2(n19203), .A(n10548), .B(n10009), .ZN(
        n10550) );
  NAND4_X1 U13449 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10555) );
  NAND2_X1 U13450 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13789), .ZN(n13103) );
  INV_X1 U13451 ( .A(n13103), .ZN(n10554) );
  NOR2_X1 U13452 ( .A1(n16339), .A2(n12350), .ZN(n19839) );
  INV_X1 U13453 ( .A(n10556), .ZN(n13232) );
  NAND2_X1 U13454 ( .A1(n13232), .A2(n10577), .ZN(n10575) );
  OAI22_X1 U13455 ( .A1(n19230), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19833), 
        .B2(n19240), .ZN(n10557) );
  INV_X1 U13456 ( .A(n10557), .ZN(n10558) );
  AND2_X1 U13457 ( .A1(n10575), .A2(n10558), .ZN(n10561) );
  INV_X1 U13458 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13790) );
  INV_X1 U13459 ( .A(n10562), .ZN(n13237) );
  AND2_X2 U13460 ( .A1(n13237), .A2(n10563), .ZN(n10712) );
  NAND2_X1 U13461 ( .A1(n10712), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U13462 ( .A1(n10712), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10568) );
  NOR2_X1 U13463 ( .A1(n19230), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13464 ( .A1(n10584), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13465 ( .A1(n10568), .A2(n10567), .ZN(n10573) );
  INV_X1 U13466 ( .A(n10569), .ZN(n10866) );
  OR2_X1 U13467 ( .A1(n10705), .A2(n10866), .ZN(n10572) );
  AND2_X1 U13468 ( .A1(n19230), .A2(n19240), .ZN(n10570) );
  AOI22_X1 U13469 ( .A1(n10556), .A2(n10570), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U13470 ( .A1(n10572), .A2(n10571), .ZN(n13542) );
  OAI21_X1 U13471 ( .B1(n13543), .B2(n13542), .A(n9893), .ZN(n10574) );
  INV_X1 U13472 ( .A(n10574), .ZN(n10581) );
  NAND2_X1 U13473 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10576) );
  OAI211_X1 U13474 ( .C1(n10705), .C2(n10864), .A(n10576), .B(n10575), .ZN(
        n10580) );
  XNOR2_X1 U13475 ( .A(n10581), .B(n10580), .ZN(n13275) );
  NAND2_X1 U13476 ( .A1(n10712), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13477 ( .A1(n10725), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10578) );
  NAND2_X1 U13478 ( .A1(n10579), .A2(n10578), .ZN(n13274) );
  NOR2_X1 U13479 ( .A1(n13275), .A2(n13274), .ZN(n13276) );
  NOR2_X1 U13480 ( .A1(n10581), .A2(n10580), .ZN(n10582) );
  NAND2_X1 U13481 ( .A1(n10712), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10588) );
  OR2_X1 U13482 ( .A1(n10705), .A2(n10583), .ZN(n10587) );
  AOI22_X1 U13483 ( .A1(n10577), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10586) );
  NAND2_X1 U13484 ( .A1(n10725), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13485 ( .A1(n10712), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13486 ( .A1(n10725), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10591) );
  INV_X1 U13487 ( .A(n10589), .ZN(n10875) );
  OR2_X1 U13488 ( .A1(n10705), .A2(n10875), .ZN(n10590) );
  AOI22_X1 U13489 ( .A1(n10712), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n10577), .ZN(n10595) );
  AOI22_X1 U13490 ( .A1(n9850), .A2(n10593), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n10725), .ZN(n10594) );
  NAND2_X1 U13491 ( .A1(n10595), .A2(n10594), .ZN(n15628) );
  OR2_X1 U13492 ( .A1(n10705), .A2(n10596), .ZN(n10597) );
  NAND2_X1 U13493 ( .A1(n10712), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13494 ( .A1(n10725), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10598) );
  NAND2_X1 U13495 ( .A1(n10599), .A2(n10598), .ZN(n15606) );
  NAND2_X1 U13496 ( .A1(n15605), .A2(n15606), .ZN(n10601) );
  OR2_X1 U13497 ( .A1(n10705), .A2(n10402), .ZN(n10600) );
  NAND2_X1 U13498 ( .A1(n10712), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13499 ( .A1(n10725), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13500 ( .A1(n10603), .A2(n10602), .ZN(n15588) );
  NAND2_X1 U13501 ( .A1(n10712), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13502 ( .A1(n10725), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13503 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n9628), .B1(
        n10211), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13504 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12478), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13505 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13506 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10604), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10605) );
  NAND4_X1 U13507 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .ZN(
        n10614) );
  AOI22_X1 U13508 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10300), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13509 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13510 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10159), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13511 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13512 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10613) );
  OR2_X1 U13513 ( .A1(n10614), .A2(n10613), .ZN(n13722) );
  INV_X1 U13514 ( .A(n13722), .ZN(n13668) );
  OR2_X1 U13515 ( .A1(n10705), .A2(n13668), .ZN(n10615) );
  AOI22_X1 U13516 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13517 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13518 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10604), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13520 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10627) );
  AOI22_X1 U13521 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10300), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12513), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10622) );
  NAND4_X1 U13525 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10626) );
  OR2_X1 U13526 ( .A1(n10627), .A2(n10626), .ZN(n13774) );
  AOI22_X1 U13527 ( .A1(n9850), .A2(n13774), .B1(n10712), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13528 ( .A1(n10725), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10577), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13529 ( .A1(n10629), .A2(n10628), .ZN(n15581) );
  AOI22_X1 U13530 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10211), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13531 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13532 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13533 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10630) );
  NAND4_X1 U13534 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10639) );
  AOI22_X1 U13535 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13536 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13537 ( .A1(n12514), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13538 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10634) );
  NAND4_X1 U13539 ( .A1(n10637), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n10638) );
  OR2_X1 U13540 ( .A1(n10639), .A2(n10638), .ZN(n13777) );
  INV_X1 U13541 ( .A(n13777), .ZN(n10641) );
  AOI22_X1 U13542 ( .A1(n10725), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10640) );
  OAI21_X1 U13543 ( .B1(n10641), .B2(n10705), .A(n10640), .ZN(n10642) );
  AOI21_X1 U13544 ( .B1(n10712), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10642), 
        .ZN(n13615) );
  AOI22_X1 U13545 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13546 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13547 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n9593), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13549 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10652) );
  AOI22_X1 U13550 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13551 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13552 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10159), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13554 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10651) );
  NOR2_X1 U13555 ( .A1(n10652), .A2(n10651), .ZN(n13532) );
  NAND2_X1 U13556 ( .A1(n10712), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13557 ( .A1(n10725), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10653) );
  OAI211_X1 U13558 ( .C1(n10705), .C2(n13532), .A(n10654), .B(n10653), .ZN(
        n15568) );
  NAND2_X1 U13559 ( .A1(n15567), .A2(n15568), .ZN(n15540) );
  NAND2_X1 U13560 ( .A1(n10712), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13561 ( .A1(n10725), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13562 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13563 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13564 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13565 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9593), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13566 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10664) );
  AOI22_X1 U13567 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13568 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13569 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13570 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10659) );
  NAND4_X1 U13571 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10663) );
  NOR2_X1 U13572 ( .A1(n10664), .A2(n10663), .ZN(n13601) );
  OR2_X1 U13573 ( .A1(n10705), .A2(n13601), .ZN(n10665) );
  AOI22_X1 U13574 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13575 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13576 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13577 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10668) );
  NAND4_X1 U13578 ( .A1(n10671), .A2(n10670), .A3(n10669), .A4(n10668), .ZN(
        n10677) );
  AOI22_X1 U13579 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13580 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13581 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13582 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13583 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10676) );
  NOR2_X1 U13584 ( .A1(n10677), .A2(n10676), .ZN(n13663) );
  NAND2_X1 U13585 ( .A1(n10712), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13586 ( .A1(n10725), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10678) );
  OAI211_X1 U13587 ( .C1(n10705), .C2(n13663), .A(n10679), .B(n10678), .ZN(
        n13091) );
  NAND2_X1 U13588 ( .A1(n10712), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13589 ( .A1(n10725), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13590 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10211), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13591 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13592 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13593 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9593), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13594 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10689) );
  AOI22_X1 U13595 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13596 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13597 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13598 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U13599 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  OR2_X1 U13600 ( .A1(n10689), .A2(n10688), .ZN(n13835) );
  INV_X1 U13601 ( .A(n13835), .ZN(n12438) );
  OR2_X1 U13602 ( .A1(n10705), .A2(n12438), .ZN(n10690) );
  AOI22_X1 U13603 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13604 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13605 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13606 ( .A1(n9593), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13607 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10702) );
  AOI22_X1 U13608 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13609 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13610 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13611 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U13612 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  OR2_X1 U13613 ( .A1(n10702), .A2(n10701), .ZN(n13877) );
  INV_X1 U13614 ( .A(n13877), .ZN(n12439) );
  NAND2_X1 U13615 ( .A1(n10712), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13616 ( .A1(n10725), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10703) );
  OAI211_X1 U13617 ( .C1(n10705), .C2(n12439), .A(n10704), .B(n10703), .ZN(
        n16267) );
  NAND2_X1 U13618 ( .A1(n10712), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13619 ( .A1(n10725), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U13620 ( .A1(n10707), .A2(n10706), .ZN(n15510) );
  NAND2_X1 U13621 ( .A1(n10712), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13622 ( .A1(n10725), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U13623 ( .A1(n10709), .A2(n10708), .ZN(n14004) );
  NAND2_X1 U13624 ( .A1(n10712), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13625 ( .A1(n10725), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10710) );
  AND2_X1 U13626 ( .A1(n10711), .A2(n10710), .ZN(n14026) );
  NAND2_X1 U13627 ( .A1(n10712), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13628 ( .A1(n10725), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U13629 ( .A1(n10714), .A2(n10713), .ZN(n14051) );
  NAND2_X1 U13630 ( .A1(n10712), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13631 ( .A1(n10725), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10715) );
  AND2_X1 U13632 ( .A1(n10716), .A2(n10715), .ZN(n14238) );
  NAND2_X1 U13633 ( .A1(n10712), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13634 ( .A1(n10725), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13635 ( .A1(n10718), .A2(n10717), .ZN(n13061) );
  NAND2_X1 U13636 ( .A1(n10712), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13637 ( .A1(n10725), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U13638 ( .A1(n10720), .A2(n10719), .ZN(n15039) );
  NAND2_X1 U13639 ( .A1(n13060), .A2(n15039), .ZN(n13073) );
  NAND2_X1 U13640 ( .A1(n10712), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13641 ( .A1(n10725), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10721) );
  AND2_X1 U13642 ( .A1(n10722), .A2(n10721), .ZN(n13074) );
  NAND2_X1 U13643 ( .A1(n10712), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13644 ( .A1(n10725), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10723) );
  AND2_X1 U13645 ( .A1(n10724), .A2(n10723), .ZN(n15022) );
  OR2_X2 U13646 ( .A1(n15023), .A2(n15022), .ZN(n15025) );
  NAND2_X1 U13647 ( .A1(n10712), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13648 ( .A1(n10725), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10726) );
  AND2_X1 U13649 ( .A1(n10727), .A2(n10726), .ZN(n15012) );
  NAND2_X1 U13651 ( .A1(n10712), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13652 ( .A1(n10725), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U13653 ( .A1(n10729), .A2(n10728), .ZN(n14989) );
  NAND2_X1 U13654 ( .A1(n10712), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13655 ( .A1(n10725), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10730) );
  AND2_X1 U13656 ( .A1(n10731), .A2(n10730), .ZN(n15149) );
  NAND2_X1 U13657 ( .A1(n10712), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13658 ( .A1(n10725), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10732) );
  AND2_X1 U13659 ( .A1(n10733), .A2(n10732), .ZN(n14978) );
  NAND2_X1 U13660 ( .A1(n10712), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13661 ( .A1(n10725), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13662 ( .A1(n10735), .A2(n10734), .ZN(n15135) );
  NAND2_X1 U13663 ( .A1(n10712), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13664 ( .A1(n10725), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10577), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13665 ( .A1(n10737), .A2(n10736), .ZN(n10739) );
  NAND2_X1 U13666 ( .A1(n10738), .A2(n10739), .ZN(n14266) );
  INV_X1 U13667 ( .A(n10738), .ZN(n10741) );
  INV_X1 U13668 ( .A(n10739), .ZN(n10740) );
  NAND2_X1 U13669 ( .A1(n10741), .A2(n10740), .ZN(n10742) );
  NAND2_X1 U13670 ( .A1(n14266), .A2(n10742), .ZN(n14352) );
  NAND2_X1 U13671 ( .A1(n10744), .A2(n10743), .ZN(n13782) );
  NAND2_X1 U13672 ( .A1(n16341), .A2(n19849), .ZN(n10746) );
  NAND2_X1 U13673 ( .A1(n13782), .A2(n10746), .ZN(n10747) );
  NAND2_X1 U13674 ( .A1(n10749), .A2(n10748), .ZN(n10753) );
  OR2_X1 U13675 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  NAND2_X1 U13676 ( .A1(n10753), .A2(n10752), .ZN(n13401) );
  INV_X1 U13677 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15630) );
  OR2_X1 U13678 ( .A1(n10844), .A2(n15630), .ZN(n10758) );
  INV_X1 U13679 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10755) );
  INV_X1 U13680 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10754) );
  OAI22_X1 U13681 ( .A1(n10841), .A2(n10755), .B1(n13789), .B2(n10754), .ZN(
        n10756) );
  AOI21_X1 U13682 ( .B1(n10807), .B2(P2_EBX_REG_4__SCAN_IN), .A(n10756), .ZN(
        n10757) );
  INV_X1 U13683 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10761) );
  OAI22_X1 U13684 ( .A1(n10841), .A2(n10761), .B1(n13789), .B2(n16256), .ZN(
        n10762) );
  AOI21_X1 U13685 ( .B1(n10807), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10762), .ZN(
        n10763) );
  INV_X1 U13686 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10767) );
  OAI22_X1 U13687 ( .A1(n10841), .A2(n10767), .B1(n13789), .B2(n9739), .ZN(
        n10768) );
  AOI21_X1 U13688 ( .B1(n10807), .B2(P2_EBX_REG_6__SCAN_IN), .A(n10768), .ZN(
        n10769) );
  INV_X1 U13689 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10771) );
  OAI22_X1 U13690 ( .A1(n10841), .A2(n10771), .B1(n13789), .B2(n15350), .ZN(
        n10772) );
  AOI21_X1 U13691 ( .B1(n10807), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10772), .ZN(
        n10773) );
  OAI21_X1 U13692 ( .B1(n10774), .B2(n16304), .A(n10773), .ZN(n13572) );
  INV_X1 U13693 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13413) );
  INV_X1 U13694 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10775) );
  OAI22_X1 U13695 ( .A1(n10841), .A2(n13413), .B1(n13789), .B2(n10775), .ZN(
        n10776) );
  AOI21_X1 U13696 ( .B1(n10807), .B2(P2_EBX_REG_8__SCAN_IN), .A(n10776), .ZN(
        n10777) );
  OAI21_X1 U13697 ( .B1(n10844), .B2(n16315), .A(n10777), .ZN(n13405) );
  OR2_X1 U13698 ( .A1(n10844), .A2(n15564), .ZN(n10782) );
  INV_X1 U13699 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10779) );
  INV_X1 U13700 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10778) );
  OAI22_X1 U13701 ( .A1(n10841), .A2(n10779), .B1(n13789), .B2(n10778), .ZN(
        n10780) );
  AOI21_X1 U13702 ( .B1(n10807), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10780), .ZN(
        n10781) );
  NAND2_X1 U13703 ( .A1(n10782), .A2(n10781), .ZN(n13534) );
  INV_X1 U13704 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16289) );
  OR2_X1 U13705 ( .A1(n10844), .A2(n16289), .ZN(n10786) );
  INV_X1 U13706 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13620) );
  INV_X1 U13707 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10783) );
  OAI22_X1 U13708 ( .A1(n10841), .A2(n13620), .B1(n13789), .B2(n10783), .ZN(
        n10784) );
  AOI21_X1 U13709 ( .B1(n10807), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10784), .ZN(
        n10785) );
  NAND2_X1 U13710 ( .A1(n10786), .A2(n10785), .ZN(n13621) );
  INV_X1 U13711 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10787) );
  OAI22_X1 U13712 ( .A1(n10841), .A2(n10787), .B1(n13789), .B2(n16235), .ZN(
        n10788) );
  AOI21_X1 U13713 ( .B1(n10807), .B2(P2_EBX_REG_9__SCAN_IN), .A(n10788), .ZN(
        n10789) );
  OAI21_X1 U13714 ( .B1(n10844), .B2(n15563), .A(n10789), .ZN(n13669) );
  INV_X1 U13715 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10792) );
  INV_X1 U13716 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10791) );
  OAI22_X1 U13717 ( .A1(n10841), .A2(n10792), .B1(n13789), .B2(n10791), .ZN(
        n10793) );
  AOI21_X1 U13718 ( .B1(n10807), .B2(P2_EBX_REG_12__SCAN_IN), .A(n10793), .ZN(
        n10794) );
  OAI21_X1 U13719 ( .B1(n10844), .B2(n15539), .A(n10794), .ZN(n13598) );
  INV_X1 U13720 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15336) );
  INV_X1 U13721 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10795) );
  OAI22_X1 U13722 ( .A1(n10841), .A2(n15336), .B1(n13789), .B2(n10795), .ZN(
        n10796) );
  AOI21_X1 U13723 ( .B1(n10807), .B2(P2_EBX_REG_13__SCAN_IN), .A(n10796), .ZN(
        n10797) );
  INV_X1 U13724 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13960) );
  OAI22_X1 U13725 ( .A1(n10841), .A2(n13960), .B1(n13789), .B2(n9745), .ZN(
        n10799) );
  AOI21_X1 U13726 ( .B1(n10807), .B2(P2_EBX_REG_14__SCAN_IN), .A(n10799), .ZN(
        n10800) );
  OAI21_X1 U13727 ( .B1(n10844), .B2(n16198), .A(n10800), .ZN(n13837) );
  INV_X1 U13728 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15326) );
  INV_X1 U13729 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10801) );
  OAI22_X1 U13730 ( .A1(n10841), .A2(n15326), .B1(n13789), .B2(n10801), .ZN(
        n10802) );
  AOI21_X1 U13731 ( .B1(n10807), .B2(P2_EBX_REG_15__SCAN_IN), .A(n10802), .ZN(
        n10803) );
  OAI21_X1 U13732 ( .B1(n10844), .B2(n14226), .A(n10803), .ZN(n13879) );
  INV_X1 U13733 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15502) );
  INV_X1 U13734 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15513) );
  INV_X1 U13735 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10804) );
  OAI22_X1 U13736 ( .A1(n10841), .A2(n15513), .B1(n13789), .B2(n10804), .ZN(
        n10805) );
  AOI21_X1 U13737 ( .B1(n10807), .B2(P2_EBX_REG_16__SCAN_IN), .A(n10805), .ZN(
        n10806) );
  OAI21_X1 U13738 ( .B1(n10844), .B2(n15502), .A(n10806), .ZN(n13843) );
  INV_X1 U13739 ( .A(n10844), .ZN(n14256) );
  INV_X1 U13740 ( .A(n10807), .ZN(n14254) );
  INV_X1 U13741 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13742 ( .A1(n14252), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10808) );
  OAI21_X1 U13743 ( .B1(n14254), .B2(n10809), .A(n10808), .ZN(n10810) );
  AOI21_X1 U13744 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10810), .ZN(n13988) );
  INV_X1 U13745 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19763) );
  INV_X1 U13746 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10813) );
  OAI22_X1 U13747 ( .A1(n10841), .A2(n19763), .B1(n13789), .B2(n10813), .ZN(
        n10814) );
  AOI21_X1 U13748 ( .B1(n10807), .B2(P2_EBX_REG_20__SCAN_IN), .A(n10814), .ZN(
        n10815) );
  OAI21_X1 U13749 ( .B1(n10844), .B2(n10816), .A(n10815), .ZN(n14231) );
  INV_X1 U13750 ( .A(n14231), .ZN(n10823) );
  INV_X1 U13751 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13752 ( .A1(n14252), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10817) );
  OAI21_X1 U13753 ( .B1(n14254), .B2(n10818), .A(n10817), .ZN(n10819) );
  AOI21_X1 U13754 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10819), .ZN(n15124) );
  INV_X1 U13755 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13756 ( .A1(n14252), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10820) );
  OAI21_X1 U13757 ( .B1(n14254), .B2(n10821), .A(n10820), .ZN(n10822) );
  AOI21_X1 U13758 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10822), .ZN(n14013) );
  OR2_X1 U13759 ( .A1(n15124), .A2(n14013), .ZN(n14230) );
  INV_X1 U13760 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19765) );
  INV_X1 U13761 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14189) );
  OAI22_X1 U13762 ( .A1(n10841), .A2(n19765), .B1(n13789), .B2(n14189), .ZN(
        n10825) );
  AOI21_X1 U13763 ( .B1(n10807), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10825), .ZN(
        n10826) );
  OAI21_X1 U13764 ( .B1(n10844), .B2(n14199), .A(n10826), .ZN(n13059) );
  INV_X1 U13765 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U13766 ( .A1(n14252), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10827) );
  OAI21_X1 U13767 ( .B1(n14254), .B2(n15115), .A(n10827), .ZN(n10828) );
  AOI21_X1 U13768 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10828), .ZN(n15035) );
  OR2_X2 U13769 ( .A1(n15036), .A2(n15035), .ZN(n15038) );
  INV_X1 U13770 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13771 ( .A1(n14252), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10829) );
  OAI21_X1 U13772 ( .B1(n14254), .B2(n10830), .A(n10829), .ZN(n10831) );
  AOI21_X1 U13773 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10831), .ZN(n13071) );
  INV_X1 U13774 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15253) );
  INV_X1 U13775 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15254) );
  OAI22_X1 U13776 ( .A1(n10841), .A2(n15253), .B1(n13789), .B2(n15254), .ZN(
        n10832) );
  AOI21_X1 U13777 ( .B1(n10807), .B2(P2_EBX_REG_24__SCAN_IN), .A(n10832), .ZN(
        n10833) );
  OAI21_X1 U13778 ( .B1(n10844), .B2(n15402), .A(n10833), .ZN(n15019) );
  AOI22_X1 U13779 ( .A1(n14252), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10834) );
  OAI21_X1 U13780 ( .B1(n14254), .B2(n15005), .A(n10834), .ZN(n10835) );
  AOI21_X1 U13781 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10835), .ZN(n15011) );
  INV_X1 U13782 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15091) );
  AOI22_X1 U13783 ( .A1(n14252), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10836) );
  OAI21_X1 U13784 ( .B1(n14254), .B2(n15091), .A(n10836), .ZN(n10837) );
  AOI21_X1 U13785 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10837), .ZN(n14995) );
  INV_X1 U13786 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15391) );
  INV_X1 U13787 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19775) );
  INV_X1 U13788 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15216) );
  OAI22_X1 U13789 ( .A1(n10841), .A2(n19775), .B1(n13789), .B2(n15216), .ZN(
        n10838) );
  AOI21_X1 U13790 ( .B1(n10807), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10838), .ZN(
        n10839) );
  OAI21_X1 U13791 ( .B1(n10844), .B2(n15391), .A(n10839), .ZN(n15077) );
  INV_X1 U13792 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15375) );
  INV_X1 U13793 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19776) );
  INV_X1 U13794 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10840) );
  OAI22_X1 U13795 ( .A1(n10841), .A2(n19776), .B1(n13789), .B2(n10840), .ZN(
        n10842) );
  AOI21_X1 U13796 ( .B1(n10807), .B2(P2_EBX_REG_28__SCAN_IN), .A(n10842), .ZN(
        n10843) );
  OAI21_X1 U13797 ( .B1(n10844), .B2(n15375), .A(n10843), .ZN(n14973) );
  INV_X1 U13798 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13799 ( .A1(n14252), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10845) );
  OAI21_X1 U13800 ( .B1(n14254), .B2(n10846), .A(n10845), .ZN(n10847) );
  AOI21_X1 U13801 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10847), .ZN(n15065) );
  AOI22_X1 U13802 ( .A1(n14252), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10848) );
  OAI21_X1 U13803 ( .B1(n14254), .B2(n10849), .A(n10848), .ZN(n10850) );
  AOI21_X1 U13804 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10850), .ZN(n10852) );
  INV_X1 U13805 ( .A(n10852), .ZN(n10851) );
  NAND2_X1 U13806 ( .A1(n10853), .A2(n10852), .ZN(n10854) );
  AND2_X1 U13807 ( .A1(n10855), .A2(n10936), .ZN(n16294) );
  NOR2_X1 U13808 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19799) );
  NAND2_X1 U13809 ( .A1(n19799), .A2(n19852), .ZN(n13101) );
  OR2_X1 U13810 ( .A1(n13101), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10856) );
  INV_X1 U13811 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n10857) );
  OR2_X1 U13812 ( .A1(n10856), .A2(n10857), .ZN(n12137) );
  INV_X1 U13813 ( .A(n10860), .ZN(n10861) );
  XOR2_X1 U13814 ( .A(n10864), .B(n10863), .Z(n13289) );
  OR2_X1 U13815 ( .A1(n13306), .A2(n19849), .ZN(n10865) );
  NAND2_X1 U13816 ( .A1(n10865), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13308) );
  XNOR2_X1 U13817 ( .A(n13306), .B(n10866), .ZN(n10867) );
  NOR2_X1 U13818 ( .A1(n13308), .A2(n10867), .ZN(n10868) );
  INV_X1 U13819 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15642) );
  XNOR2_X1 U13820 ( .A(n13308), .B(n10867), .ZN(n13299) );
  NOR2_X1 U13821 ( .A1(n15642), .A2(n13299), .ZN(n13298) );
  NOR2_X1 U13822 ( .A1(n10868), .A2(n13298), .ZN(n10869) );
  XNOR2_X1 U13823 ( .A(n10934), .B(n10869), .ZN(n13288) );
  NOR2_X1 U13824 ( .A1(n13289), .A2(n13288), .ZN(n10871) );
  NOR2_X1 U13825 ( .A1(n10869), .A2(n10934), .ZN(n10870) );
  OR2_X1 U13826 ( .A1(n10871), .A2(n10870), .ZN(n10872) );
  XNOR2_X1 U13827 ( .A(n10872), .B(n13806), .ZN(n13809) );
  NAND2_X1 U13828 ( .A1(n10872), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10873) );
  INV_X1 U13829 ( .A(n10879), .ZN(n10877) );
  NAND2_X1 U13830 ( .A1(n10877), .A2(n10878), .ZN(n15621) );
  INV_X1 U13831 ( .A(n10890), .ZN(n10884) );
  OAI21_X2 U13832 ( .B1(n10891), .B2(n10884), .A(n10883), .ZN(n15358) );
  XNOR2_X1 U13833 ( .A(n10901), .B(n14320), .ZN(n10889) );
  AND2_X1 U13834 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10889), .ZN(
        n10888) );
  INV_X1 U13835 ( .A(n10889), .ZN(n10896) );
  NAND2_X1 U13836 ( .A1(n15345), .A2(n10892), .ZN(n16244) );
  NOR2_X1 U13837 ( .A1(n10901), .A2(n10402), .ZN(n10893) );
  XNOR2_X1 U13838 ( .A(n10893), .B(n16315), .ZN(n16246) );
  AND2_X1 U13839 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16246), .ZN(
        n10894) );
  NAND2_X1 U13840 ( .A1(n15358), .A2(n10894), .ZN(n10899) );
  INV_X1 U13841 ( .A(n16246), .ZN(n10897) );
  AND2_X2 U13842 ( .A1(n10896), .A2(n10895), .ZN(n15342) );
  OR2_X2 U13843 ( .A1(n10897), .A2(n15342), .ZN(n10898) );
  NAND2_X1 U13844 ( .A1(n10899), .A2(n10898), .ZN(n10900) );
  NAND2_X1 U13845 ( .A1(n16244), .A2(n10900), .ZN(n10904) );
  INV_X1 U13846 ( .A(n10901), .ZN(n10902) );
  NAND3_X1 U13847 ( .A1(n10902), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n14320), .ZN(n10903) );
  INV_X1 U13848 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15539) );
  NOR2_X1 U13849 ( .A1(n15539), .A2(n10411), .ZN(n16282) );
  NAND2_X1 U13850 ( .A1(n16282), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16280) );
  AND3_X1 U13851 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15522) );
  INV_X1 U13852 ( .A(n15522), .ZN(n15524) );
  NOR2_X1 U13853 ( .A1(n16280), .A2(n15524), .ZN(n15493) );
  AND2_X1 U13854 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10931) );
  AND2_X1 U13855 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14227) );
  NAND2_X1 U13856 ( .A1(n10931), .A2(n14227), .ZN(n10905) );
  OR2_X1 U13857 ( .A1(n10905), .A2(n15502), .ZN(n10906) );
  OR2_X1 U13858 ( .A1(n10906), .A2(n14226), .ZN(n14195) );
  OR2_X1 U13859 ( .A1(n14199), .A2(n14195), .ZN(n14194) );
  NAND2_X1 U13860 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15444) );
  OR2_X1 U13861 ( .A1(n14194), .A2(n15444), .ZN(n10907) );
  AND2_X1 U13862 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U13863 ( .A1(n15226), .A2(n10908), .ZN(n15209) );
  INV_X1 U13864 ( .A(n15365), .ZN(n10909) );
  XNOR2_X1 U13865 ( .A(n15194), .B(n10953), .ZN(n12128) );
  INV_X1 U13866 ( .A(n10910), .ZN(n19838) );
  NAND2_X1 U13867 ( .A1(n10936), .A2(n19838), .ZN(n16330) );
  NAND2_X1 U13868 ( .A1(n12128), .A2(n16295), .ZN(n10956) );
  NAND2_X1 U13869 ( .A1(n10936), .A2(n13183), .ZN(n15490) );
  NAND2_X1 U13870 ( .A1(n10913), .A2(n9967), .ZN(n10915) );
  INV_X1 U13871 ( .A(n13107), .ZN(n13104) );
  AOI22_X1 U13872 ( .A1(n10915), .A2(n13104), .B1(n19203), .B2(n10914), .ZN(
        n10922) );
  OR2_X1 U13873 ( .A1(n10916), .A2(n10566), .ZN(n15653) );
  NAND2_X1 U13874 ( .A1(n15653), .A2(n10917), .ZN(n10918) );
  NAND2_X1 U13875 ( .A1(n10918), .A2(n15699), .ZN(n10921) );
  INV_X1 U13876 ( .A(n10919), .ZN(n10920) );
  NAND2_X1 U13877 ( .A1(n9966), .A2(n10920), .ZN(n13229) );
  NAND4_X1 U13878 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n13229), .ZN(
        n10924) );
  AOI21_X1 U13879 ( .B1(n10926), .B2(n10925), .A(n10924), .ZN(n15651) );
  INV_X1 U13880 ( .A(n10927), .ZN(n13784) );
  NAND2_X1 U13881 ( .A1(n15651), .A2(n13784), .ZN(n10928) );
  NAND2_X1 U13882 ( .A1(n10936), .A2(n10928), .ZN(n15495) );
  NOR2_X1 U13883 ( .A1(n13790), .A2(n15642), .ZN(n13293) );
  INV_X1 U13884 ( .A(n15490), .ZN(n10929) );
  INV_X1 U13885 ( .A(n13293), .ZN(n15647) );
  NOR2_X1 U13886 ( .A1(n10934), .A2(n15647), .ZN(n13280) );
  OAI22_X1 U13887 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13293), .B1(
        n10929), .B2(n13280), .ZN(n13805) );
  NAND3_X1 U13888 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15603) );
  NOR2_X1 U13889 ( .A1(n15357), .A2(n15603), .ZN(n10939) );
  NAND2_X1 U13890 ( .A1(n15602), .A2(n10939), .ZN(n16302) );
  NAND2_X1 U13891 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16301) );
  NAND2_X1 U13892 ( .A1(n15493), .A2(n15579), .ZN(n16268) );
  NAND3_X1 U13893 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10943) );
  INV_X1 U13894 ( .A(n10931), .ZN(n14243) );
  NOR2_X1 U13895 ( .A1(n14242), .A2(n14243), .ZN(n14200) );
  INV_X1 U13896 ( .A(n15444), .ZN(n10932) );
  NAND2_X1 U13897 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15406) );
  NOR2_X1 U13898 ( .A1(n15402), .A2(n15406), .ZN(n10933) );
  NAND2_X1 U13899 ( .A1(n15405), .A2(n10933), .ZN(n15376) );
  NAND2_X1 U13900 ( .A1(n15365), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10951) );
  NOR2_X1 U13901 ( .A1(n15376), .A2(n10951), .ZN(n14337) );
  INV_X1 U13902 ( .A(n14337), .ZN(n10952) );
  INV_X1 U13903 ( .A(n10933), .ZN(n10950) );
  INV_X1 U13904 ( .A(n15495), .ZN(n10935) );
  NAND2_X1 U13905 ( .A1(n10935), .A2(n10934), .ZN(n13279) );
  OR3_X1 U13906 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13293), .A3(
        n15490), .ZN(n13282) );
  NAND2_X1 U13907 ( .A1(n13279), .A2(n13282), .ZN(n10938) );
  INV_X1 U13908 ( .A(n10936), .ZN(n10937) );
  INV_X1 U13909 ( .A(n19176), .ZN(n18941) );
  NAND2_X1 U13910 ( .A1(n10937), .A2(n18941), .ZN(n16320) );
  OAI21_X1 U13911 ( .B1(n15495), .B2(n13293), .A(n16320), .ZN(n13278) );
  NOR2_X1 U13912 ( .A1(n10938), .A2(n13278), .ZN(n13945) );
  INV_X1 U13913 ( .A(n10939), .ZN(n10940) );
  NAND2_X1 U13914 ( .A1(n16322), .A2(n10940), .ZN(n10941) );
  NAND2_X1 U13915 ( .A1(n16322), .A2(n16301), .ZN(n10942) );
  NAND2_X1 U13916 ( .A1(n16316), .A2(n10942), .ZN(n15562) );
  INV_X1 U13917 ( .A(n10943), .ZN(n10944) );
  NAND3_X1 U13918 ( .A1(n15493), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n10944), .ZN(n10945) );
  AND2_X1 U13919 ( .A1(n16322), .A2(n10945), .ZN(n10946) );
  AND2_X1 U13920 ( .A1(n16322), .A2(n14243), .ZN(n10947) );
  OR2_X1 U13921 ( .A1(n15479), .A2(n10947), .ZN(n14206) );
  AND2_X1 U13922 ( .A1(n16322), .A2(n14199), .ZN(n10948) );
  NOR2_X1 U13923 ( .A1(n14206), .A2(n10948), .ZN(n15462) );
  NAND2_X1 U13924 ( .A1(n16322), .A2(n15444), .ZN(n10949) );
  NAND2_X1 U13925 ( .A1(n15462), .A2(n10949), .ZN(n15440) );
  AOI21_X1 U13926 ( .B1(n10950), .B2(n16322), .A(n15440), .ZN(n15363) );
  INV_X1 U13927 ( .A(n15363), .ZN(n15397) );
  AOI211_X1 U13928 ( .C1(n16322), .C2(n10951), .A(n10953), .B(n15397), .ZN(
        n14340) );
  AOI21_X1 U13929 ( .B1(n10953), .B2(n10952), .A(n14340), .ZN(n10954) );
  OAI21_X1 U13930 ( .B1(n12142), .B2(n16299), .A(n9882), .ZN(P2_U3016) );
  AOI22_X1 U13931 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11919), .B1(
        n11641), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10962) );
  AND2_X2 U13932 ( .A1(n10963), .A2(n11022), .ZN(n11183) );
  AOI22_X1 U13933 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9588), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10961) );
  AND2_X4 U13934 ( .A1(n11022), .A2(n13694), .ZN(n12096) );
  AOI22_X1 U13935 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13936 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10959) );
  AND2_X2 U13937 ( .A1(n10968), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13682) );
  INV_X1 U13938 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11699) );
  AND2_X2 U13939 ( .A1(n10969), .A2(n10963), .ZN(n11332) );
  NAND2_X1 U13940 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U13941 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10965) );
  OAI211_X1 U13942 ( .C1(n12064), .C2(n11699), .A(n10966), .B(n10965), .ZN(
        n10967) );
  INV_X1 U13943 ( .A(n10967), .ZN(n10975) );
  AOI22_X1 U13944 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n9621), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10974) );
  AND2_X2 U13945 ( .A1(n10970), .A2(n10964), .ZN(n11173) );
  AOI22_X1 U13946 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11173), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10973) );
  INV_X1 U13947 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U13948 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10982) );
  NAND2_X1 U13949 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10981) );
  INV_X1 U13950 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13951 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10979) );
  NAND4_X1 U13952 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10984) );
  NOR2_X1 U13953 ( .A1(n13681), .A2(n11894), .ZN(n10983) );
  NAND2_X1 U13954 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U13955 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10987) );
  NAND2_X1 U13956 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10986) );
  NAND2_X1 U13957 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U13958 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U13959 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10991) );
  NAND2_X1 U13960 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U13961 ( .A1(n9591), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U13963 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10994) );
  NAND2_X1 U13964 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10993) );
  OAI211_X1 U13965 ( .C1(n12064), .C2(n11667), .A(n10994), .B(n10993), .ZN(
        n10995) );
  INV_X1 U13966 ( .A(n10995), .ZN(n10996) );
  NAND2_X1 U13967 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11003) );
  NAND2_X1 U13968 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U13969 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11001) );
  NAND2_X1 U13970 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11000) );
  NAND4_X1 U13971 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11005) );
  NOR2_X2 U13972 ( .A1(n11005), .A2(n11004), .ZN(n11020) );
  NAND2_X1 U13973 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U13974 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11008) );
  NAND2_X1 U13975 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U13976 ( .A1(n9588), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11006) );
  NAND2_X1 U13977 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U13978 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U13979 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U13980 ( .A1(n9591), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U13981 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U13982 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11014) );
  OAI211_X1 U13983 ( .C1(n13681), .C2(n12009), .A(n11015), .B(n11014), .ZN(
        n11016) );
  INV_X1 U13984 ( .A(n11016), .ZN(n11017) );
  INV_X2 U13985 ( .A(n11115), .ZN(n13512) );
  AOI22_X1 U13986 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9588), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11029) );
  INV_X1 U13987 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11024) );
  NAND2_X2 U13988 ( .A1(n11022), .A2(n13694), .ZN(n11979) );
  INV_X1 U13989 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11023) );
  OAI22_X1 U13990 ( .A1(n11021), .A2(n11024), .B1(n11979), .B2(n11023), .ZN(
        n11025) );
  INV_X1 U13991 ( .A(n11025), .ZN(n11028) );
  AOI22_X1 U13992 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13993 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11026) );
  INV_X1 U13994 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U13995 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U13996 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11030) );
  OAI211_X1 U13997 ( .C1(n13681), .C2(n11032), .A(n11031), .B(n11030), .ZN(
        n11033) );
  INV_X1 U13998 ( .A(n11033), .ZN(n11037) );
  AOI22_X1 U13999 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11173), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14000 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U14001 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14002 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U14003 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14004 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U14005 ( .A1(n9591), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11038) );
  NAND4_X1 U14006 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11038), .ZN(
        n11043) );
  INV_X1 U14007 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11928) );
  NOR2_X1 U14008 ( .A1(n13681), .A2(n11928), .ZN(n11042) );
  NOR2_X1 U14009 ( .A1(n11043), .A2(n11042), .ZN(n11059) );
  INV_X1 U14010 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11046) );
  NAND2_X1 U14011 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14012 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11044) );
  OAI211_X1 U14013 ( .C1(n11979), .C2(n11046), .A(n11045), .B(n11044), .ZN(
        n11047) );
  INV_X1 U14014 ( .A(n11047), .ZN(n11058) );
  NAND2_X1 U14015 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11051) );
  NAND2_X1 U14016 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14017 ( .A1(n9588), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11049) );
  NAND2_X1 U14018 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U14019 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11055) );
  NAND2_X1 U14020 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U14021 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11053) );
  NAND2_X1 U14022 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11052) );
  NAND4_X2 U14023 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n20064) );
  NAND2_X1 U14024 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11065) );
  NAND2_X1 U14025 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14026 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11063) );
  INV_X1 U14027 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11061) );
  NAND4_X1 U14028 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11067) );
  INV_X1 U14029 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11720) );
  NOR2_X1 U14030 ( .A1(n9626), .A2(n11720), .ZN(n11066) );
  NAND2_X1 U14031 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14032 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U14033 ( .A1(n9588), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11069) );
  NAND2_X1 U14034 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14035 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U14036 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U14037 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14038 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11072) );
  INV_X1 U14039 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U14040 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14041 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11076) );
  OAI211_X1 U14042 ( .C1(n13681), .C2(n12082), .A(n11077), .B(n11076), .ZN(
        n11078) );
  INV_X1 U14043 ( .A(n11078), .ZN(n11079) );
  NAND2_X1 U14044 ( .A1(n13259), .A2(n11083), .ZN(n13343) );
  INV_X1 U14045 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11084) );
  INV_X1 U14046 ( .A(n11087), .ZN(n11106) );
  NAND2_X1 U14047 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11091) );
  NAND2_X1 U14048 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11090) );
  NAND2_X1 U14049 ( .A1(n11172), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14050 ( .A1(n9591), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11088) );
  NAND4_X1 U14051 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n11094) );
  NAND2_X1 U14052 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U14053 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14054 ( .A1(n9588), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14055 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14056 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U14057 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U14058 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11100) );
  NAND2_X1 U14059 ( .A1(n11211), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11099) );
  OR2_X2 U14060 ( .A1(n13343), .A2(n12156), .ZN(n12154) );
  INV_X2 U14061 ( .A(n12154), .ZN(n13251) );
  INV_X1 U14062 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19868) );
  XNOR2_X1 U14063 ( .A(n19868), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12157) );
  NAND2_X1 U14064 ( .A1(n13506), .A2(n11362), .ZN(n11368) );
  NAND2_X1 U14065 ( .A1(n11526), .A2(n11368), .ZN(n11110) );
  NAND2_X1 U14066 ( .A1(n11110), .A2(n11109), .ZN(n11112) );
  AND2_X2 U14067 ( .A1(n11112), .A2(n11111), .ZN(n12152) );
  NAND2_X1 U14068 ( .A1(n11136), .A2(n20059), .ZN(n11113) );
  NAND2_X1 U14069 ( .A1(n13376), .A2(n12156), .ZN(n11135) );
  INV_X2 U14070 ( .A(n9634), .ZN(n14389) );
  NAND2_X1 U14071 ( .A1(n11108), .A2(n11362), .ZN(n13360) );
  OR2_X1 U14072 ( .A1(n13360), .A2(n11115), .ZN(n11116) );
  NAND2_X1 U14073 ( .A1(n13373), .A2(n13512), .ZN(n11149) );
  NAND2_X1 U14074 ( .A1(n11149), .A2(n14962), .ZN(n11134) );
  AOI22_X1 U14075 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14076 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9588), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14077 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14078 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11211), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11118) );
  INV_X1 U14079 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14080 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11124) );
  INV_X1 U14081 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11122) );
  OAI211_X1 U14082 ( .C1(n13681), .C2(n11760), .A(n11124), .B(n11123), .ZN(
        n11125) );
  INV_X1 U14083 ( .A(n11125), .ZN(n11130) );
  AOI22_X1 U14084 ( .A1(n11173), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11172), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14085 ( .A1(n11206), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U14086 ( .A1(n11126), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11127) );
  OAI211_X1 U14087 ( .C1(n20744), .C2(n13512), .A(n11132), .B(n13522), .ZN(
        n11154) );
  NOR2_X2 U14088 ( .A1(n20064), .A2(n20059), .ZN(n13371) );
  NOR2_X1 U14089 ( .A1(n11154), .A2(n13371), .ZN(n11133) );
  NAND4_X1 U14090 ( .A1(n11142), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(
        n11140) );
  NOR2_X1 U14091 ( .A1(n11136), .A2(n20037), .ZN(n11137) );
  NAND2_X2 U14092 ( .A1(n12152), .A2(n11137), .ZN(n12143) );
  NAND2_X1 U14093 ( .A1(n12143), .A2(n12154), .ZN(n11138) );
  NAND2_X1 U14094 ( .A1(n11138), .A2(n13255), .ZN(n13511) );
  NAND2_X1 U14095 ( .A1(n13243), .A2(n13371), .ZN(n13383) );
  NAND2_X1 U14096 ( .A1(n11526), .A2(n11486), .ZN(n11139) );
  OAI21_X2 U14097 ( .B1(n11140), .B2(n11144), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11165) );
  NAND2_X1 U14098 ( .A1(n20572), .A2(n20493), .ZN(n20441) );
  NAND2_X1 U14099 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20568) );
  NAND2_X1 U14100 ( .A1(n20441), .A2(n20568), .ZN(n20375) );
  INV_X1 U14101 ( .A(n20375), .ZN(n20126) );
  INV_X1 U14102 ( .A(n11525), .ZN(n15874) );
  AND2_X1 U14103 ( .A1(n15874), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11160) );
  AOI21_X1 U14104 ( .B1(n20126), .B2(n12119), .A(n11160), .ZN(n11141) );
  OAI21_X2 U14105 ( .B1(n11165), .B2(n9701), .A(n11141), .ZN(n11146) );
  INV_X1 U14106 ( .A(n11142), .ZN(n11143) );
  NAND2_X2 U14107 ( .A1(n11145), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11159) );
  XNOR2_X2 U14108 ( .A(n11146), .B(n11159), .ZN(n20161) );
  INV_X1 U14109 ( .A(n12119), .ZN(n11147) );
  MUX2_X1 U14110 ( .A(n11525), .B(n11147), .S(n20493), .Z(n11148) );
  INV_X1 U14111 ( .A(n11149), .ZN(n11158) );
  NAND2_X1 U14112 ( .A1(n14962), .A2(n20054), .ZN(n11157) );
  NAND3_X1 U14113 ( .A1(n13353), .A2(n13360), .A3(n20064), .ZN(n11150) );
  NAND2_X1 U14114 ( .A1(n13376), .A2(n11150), .ZN(n11156) );
  OR2_X1 U14115 ( .A1(n11151), .A2(n20744), .ZN(n11152) );
  NAND2_X1 U14116 ( .A1(n13371), .A2(n11108), .ZN(n13520) );
  NAND4_X1 U14117 ( .A1(n11152), .A2(n13520), .A3(n20724), .A4(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11153) );
  NOR2_X1 U14118 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  OAI211_X1 U14119 ( .C1(n11158), .C2(n11157), .A(n11156), .B(n11155), .ZN(
        n11193) );
  INV_X1 U14120 ( .A(n11159), .ZN(n11163) );
  INV_X1 U14121 ( .A(n11160), .ZN(n11161) );
  NAND2_X1 U14122 ( .A1(n11161), .A2(n9701), .ZN(n11162) );
  NAND2_X1 U14123 ( .A1(n11163), .A2(n11162), .ZN(n11164) );
  XNOR2_X1 U14124 ( .A(n20568), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20049) );
  NAND2_X1 U14125 ( .A1(n12119), .A2(n20049), .ZN(n11168) );
  NAND2_X1 U14126 ( .A1(n15874), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11167) );
  INV_X2 U14128 ( .A(n12085), .ZN(n12029) );
  AOI22_X1 U14129 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11176) );
  INV_X1 U14130 ( .A(n11173), .ZN(n11260) );
  AOI22_X1 U14131 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U14132 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11174) );
  NAND3_X1 U14133 ( .A1(n11176), .A2(n11175), .A3(n11174), .ZN(n11182) );
  INV_X1 U14134 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U14135 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U14136 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11178) );
  OAI211_X1 U14137 ( .C1(n11180), .C2(n11177), .A(n11179), .B(n11178), .ZN(
        n11181) );
  NOR2_X1 U14138 ( .A1(n11182), .A2(n11181), .ZN(n11190) );
  INV_X2 U14139 ( .A(n12089), .ZN(n12065) );
  AOI22_X1 U14140 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14141 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14142 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11186) );
  INV_X1 U14143 ( .A(n11211), .ZN(n11259) );
  AOI22_X1 U14144 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11185) );
  INV_X1 U14145 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20854) );
  NAND2_X1 U14146 ( .A1(n12156), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11248) );
  OAI22_X1 U14147 ( .A1(n11519), .A2(n20854), .B1(n11392), .B2(n11248), .ZN(
        n11191) );
  XNOR2_X1 U14148 ( .A(n11192), .B(n11191), .ZN(n11382) );
  INV_X1 U14149 ( .A(n11193), .ZN(n11194) );
  NAND2_X1 U14150 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U14151 ( .A(n11260), .ZN(n11220) );
  NAND2_X1 U14152 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U14153 ( .A1(n12029), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11197) );
  NAND2_X1 U14154 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11196) );
  NAND4_X1 U14155 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11202) );
  INV_X1 U14156 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11200) );
  NOR2_X1 U14157 ( .A1(n9617), .A2(n11200), .ZN(n11201) );
  NOR2_X1 U14158 ( .A1(n11202), .A2(n11201), .ZN(n11219) );
  INV_X1 U14159 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U14160 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14161 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11203) );
  OAI211_X1 U14162 ( .C1(n11790), .C2(n11979), .A(n11204), .B(n11203), .ZN(
        n11205) );
  INV_X1 U14163 ( .A(n11205), .ZN(n11218) );
  NAND2_X1 U14164 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14165 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U14166 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11208) );
  NAND2_X1 U14167 ( .A1(n12035), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14168 ( .A1(n9622), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11215) );
  NAND2_X1 U14169 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11214) );
  NAND2_X1 U14170 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11213) );
  NAND2_X1 U14171 ( .A1(n12036), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11212) );
  NAND4_X1 U14172 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11439) );
  NAND2_X1 U14173 ( .A1(n13512), .A2(n11439), .ZN(n11242) );
  INV_X1 U14174 ( .A(n11439), .ZN(n11445) );
  NAND2_X1 U14175 ( .A1(n11445), .A2(n13512), .ZN(n11238) );
  NAND2_X1 U14176 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14177 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11223) );
  NAND2_X1 U14178 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14179 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11221) );
  AOI22_X1 U14180 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U14181 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U14182 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11225) );
  INV_X1 U14183 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11230) );
  INV_X1 U14184 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11229) );
  OAI22_X1 U14185 ( .A1(n12028), .A2(n11230), .B1(n11177), .B2(n11229), .ZN(
        n11231) );
  INV_X1 U14186 ( .A(n11231), .ZN(n11235) );
  AOI22_X1 U14187 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14188 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14189 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11232) );
  MUX2_X1 U14190 ( .A(n11242), .B(n11238), .S(n11375), .Z(n11239) );
  INV_X1 U14191 ( .A(n11239), .ZN(n11240) );
  NAND2_X1 U14192 ( .A1(n11240), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11373) );
  AND2_X1 U14193 ( .A1(n11373), .A2(n11363), .ZN(n11241) );
  NAND2_X1 U14194 ( .A1(n11372), .A2(n11241), .ZN(n11247) );
  INV_X1 U14195 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11803) );
  INV_X1 U14196 ( .A(n11375), .ZN(n11243) );
  OAI211_X1 U14197 ( .C1(n11243), .C2(n20037), .A(n11242), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11244) );
  INV_X1 U14198 ( .A(n11244), .ZN(n11245) );
  INV_X1 U14199 ( .A(n11248), .ZN(n11268) );
  INV_X1 U14200 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14201 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11250) );
  NAND2_X1 U14202 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11249) );
  OAI211_X1 U14203 ( .C1(n9617), .C2(n11824), .A(n11250), .B(n11249), .ZN(
        n11251) );
  INV_X1 U14204 ( .A(n11251), .ZN(n11255) );
  AOI22_X1 U14205 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14206 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U14207 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11252) );
  NAND4_X1 U14208 ( .A1(n11255), .A2(n11254), .A3(n11253), .A4(n11252), .ZN(
        n11266) );
  INV_X1 U14209 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11257) );
  INV_X1 U14210 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11256) );
  OAI22_X1 U14211 ( .A1(n12028), .A2(n11257), .B1(n11979), .B2(n11256), .ZN(
        n11258) );
  INV_X1 U14212 ( .A(n11258), .ZN(n11264) );
  AOI22_X1 U14213 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11263) );
  INV_X1 U14214 ( .A(n11259), .ZN(n12036) );
  AOI22_X1 U14215 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11262) );
  INV_X1 U14216 ( .A(n11260), .ZN(n11789) );
  AOI22_X1 U14217 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11261) );
  NAND4_X1 U14218 ( .A1(n11264), .A2(n11263), .A3(n11262), .A4(n11261), .ZN(
        n11265) );
  INV_X1 U14219 ( .A(n11267), .ZN(n11275) );
  AOI22_X1 U14220 ( .A1(n11268), .A2(n11366), .B1(n11275), .B2(n11445), .ZN(
        n11270) );
  NAND2_X1 U14221 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11269) );
  INV_X1 U14222 ( .A(n20161), .ZN(n11273) );
  INV_X1 U14223 ( .A(n11271), .ZN(n11272) );
  NAND2_X1 U14224 ( .A1(n11275), .A2(n11366), .ZN(n11276) );
  OAI21_X2 U14225 ( .B1(n13851), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11276), 
        .ZN(n11277) );
  INV_X1 U14226 ( .A(n11277), .ZN(n11365) );
  NAND2_X1 U14227 ( .A1(n11530), .A2(n11365), .ZN(n11282) );
  INV_X1 U14228 ( .A(n11278), .ZN(n11280) );
  NAND2_X1 U14229 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  NAND2_X1 U14230 ( .A1(n11282), .A2(n11281), .ZN(n11381) );
  INV_X1 U14231 ( .A(n9614), .ZN(n11283) );
  NAND2_X1 U14232 ( .A1(n11283), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11287) );
  INV_X1 U14233 ( .A(n20568), .ZN(n20157) );
  INV_X1 U14234 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20125) );
  NAND2_X1 U14235 ( .A1(n20125), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20251) );
  INV_X1 U14236 ( .A(n20251), .ZN(n11284) );
  NAND2_X1 U14237 ( .A1(n20157), .A2(n11284), .ZN(n20288) );
  OAI21_X1 U14238 ( .B1(n20568), .B2(n20320), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U14239 ( .A1(n20288), .A2(n11285), .ZN(n20321) );
  AOI22_X1 U14240 ( .A1(n20321), .A2(n12119), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15874), .ZN(n11286) );
  XNOR2_X2 U14241 ( .A(n13695), .B(n20197), .ZN(n20319) );
  AOI22_X1 U14242 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14243 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14244 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14245 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11289) );
  AND4_X1 U14246 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11302) );
  INV_X1 U14247 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U14248 ( .A1(n9621), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14249 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11293) );
  OAI211_X1 U14250 ( .C1(n9617), .C2(n11978), .A(n11294), .B(n11293), .ZN(
        n11295) );
  INV_X1 U14251 ( .A(n11295), .ZN(n11301) );
  INV_X1 U14252 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U14253 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14254 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11296) );
  OAI211_X1 U14255 ( .C1(n11298), .C2(n11177), .A(n11297), .B(n11296), .ZN(
        n11299) );
  INV_X1 U14256 ( .A(n11299), .ZN(n11300) );
  NAND3_X1 U14257 ( .A1(n11302), .A2(n11301), .A3(n11300), .ZN(n11411) );
  AOI22_X1 U14258 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11502), .B2(n11411), .ZN(n11303) );
  NAND2_X2 U14259 ( .A1(n11305), .A2(n13710), .ZN(n11407) );
  INV_X1 U14260 ( .A(n11407), .ZN(n11342) );
  NAND2_X1 U14261 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11323) );
  INV_X1 U14262 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14263 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U14264 ( .A1(n12092), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11306) );
  OAI211_X1 U14265 ( .C1(n9617), .C2(n12026), .A(n11307), .B(n11306), .ZN(
        n11308) );
  INV_X1 U14266 ( .A(n11308), .ZN(n11312) );
  AOI22_X1 U14267 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14268 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14269 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11309) );
  NAND4_X1 U14270 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n11321) );
  AOI22_X1 U14271 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11319) );
  INV_X1 U14272 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11314) );
  INV_X1 U14273 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11313) );
  OAI22_X1 U14274 ( .A1(n12028), .A2(n11314), .B1(n11177), .B2(n11313), .ZN(
        n11315) );
  INV_X1 U14275 ( .A(n11315), .ZN(n11318) );
  AOI22_X1 U14276 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14277 ( .A1(n9620), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11316) );
  NAND4_X1 U14278 ( .A1(n11319), .A2(n11318), .A3(n11317), .A4(n11316), .ZN(
        n11320) );
  NAND2_X1 U14279 ( .A1(n11502), .A2(n11420), .ZN(n11322) );
  NAND2_X1 U14280 ( .A1(n11323), .A2(n11322), .ZN(n11404) );
  INV_X1 U14281 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12006) );
  OR2_X1 U14282 ( .A1(n11519), .A2(n12006), .ZN(n11340) );
  AOI22_X1 U14283 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14284 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14285 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11324) );
  NAND3_X1 U14286 ( .A1(n11326), .A2(n11325), .A3(n11324), .ZN(n11331) );
  INV_X1 U14287 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14288 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14289 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11327) );
  OAI211_X1 U14290 ( .C1(n11329), .C2(n11979), .A(n11328), .B(n11327), .ZN(
        n11330) );
  NOR2_X1 U14291 ( .A1(n11331), .A2(n11330), .ZN(n11338) );
  AOI22_X1 U14292 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14293 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14294 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14295 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11333) );
  AND4_X1 U14296 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11337) );
  NAND2_X1 U14297 ( .A1(n11338), .A2(n11337), .ZN(n11410) );
  NAND2_X1 U14298 ( .A1(n11502), .A2(n11410), .ZN(n11339) );
  NAND2_X1 U14299 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11359) );
  AOI22_X1 U14300 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14301 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11344) );
  NAND2_X1 U14302 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11343) );
  NAND3_X1 U14303 ( .A1(n11345), .A2(n11344), .A3(n11343), .ZN(n11351) );
  INV_X1 U14304 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14305 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11348) );
  INV_X1 U14306 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11346) );
  OR2_X1 U14307 ( .A1(n12028), .A2(n11346), .ZN(n11347) );
  OAI211_X1 U14308 ( .C1(n11177), .C2(n11349), .A(n11348), .B(n11347), .ZN(
        n11350) );
  NOR2_X1 U14309 ( .A1(n11351), .A2(n11350), .ZN(n11357) );
  AOI22_X1 U14310 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14311 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14312 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14313 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11352) );
  AND4_X1 U14314 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11356) );
  NAND2_X1 U14315 ( .A1(n11357), .A2(n11356), .ZN(n11437) );
  NAND2_X1 U14316 ( .A1(n11502), .A2(n11437), .ZN(n11358) );
  INV_X1 U14317 ( .A(n13265), .ZN(n11409) );
  NOR2_X1 U14318 ( .A1(n11409), .A2(n11363), .ZN(n11364) );
  AND2_X4 U14319 ( .A1(n11435), .A2(n11364), .ZN(n16052) );
  INV_X1 U14320 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14760) );
  NAND2_X1 U14321 ( .A1(n16052), .A2(n14760), .ZN(n14625) );
  NAND2_X1 U14322 ( .A1(n11365), .A2(n20054), .ZN(n11371) );
  INV_X1 U14323 ( .A(n20744), .ZN(n11440) );
  NAND2_X1 U14324 ( .A1(n11375), .A2(n11366), .ZN(n11393) );
  OAI21_X1 U14325 ( .B1(n11366), .B2(n11375), .A(n11393), .ZN(n11367) );
  INV_X1 U14326 ( .A(n11367), .ZN(n11369) );
  AOI21_X1 U14327 ( .B1(n11440), .B2(n11369), .A(n11368), .ZN(n11370) );
  NAND2_X1 U14328 ( .A1(n11371), .A2(n11370), .ZN(n11378) );
  NAND2_X1 U14329 ( .A1(n12156), .A2(n20064), .ZN(n11384) );
  OAI21_X1 U14330 ( .B1(n20744), .B2(n11375), .A(n11384), .ZN(n11376) );
  INV_X1 U14331 ( .A(n11376), .ZN(n11377) );
  INV_X1 U14332 ( .A(n11378), .ZN(n11379) );
  NAND2_X2 U14333 ( .A1(n13492), .A2(n11380), .ZN(n11388) );
  INV_X1 U14334 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20026) );
  XNOR2_X2 U14335 ( .A(n11388), .B(n20026), .ZN(n13564) );
  NAND2_X1 U14336 ( .A1(n11382), .A2(n11381), .ZN(n11383) );
  XNOR2_X1 U14337 ( .A(n11393), .B(n11392), .ZN(n11386) );
  INV_X1 U14338 ( .A(n11384), .ZN(n11385) );
  AOI21_X1 U14339 ( .B1(n11386), .B2(n11440), .A(n11385), .ZN(n11387) );
  OAI21_X2 U14340 ( .B1(n13704), .B2(n11409), .A(n11387), .ZN(n13563) );
  NAND2_X1 U14341 ( .A1(n11388), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11389) );
  INV_X1 U14342 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20007) );
  NAND2_X1 U14343 ( .A1(n11390), .A2(n13709), .ZN(n11391) );
  NAND2_X1 U14344 ( .A1(n11393), .A2(n11392), .ZN(n11413) );
  XNOR2_X1 U14345 ( .A(n11413), .B(n11411), .ZN(n11394) );
  OAI22_X1 U14346 ( .A1(n20035), .A2(n11409), .B1(n20744), .B2(n11394), .ZN(
        n13608) );
  NAND2_X1 U14347 ( .A1(n13609), .A2(n13608), .ZN(n13607) );
  NAND2_X1 U14348 ( .A1(n11395), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11396) );
  INV_X1 U14349 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19999) );
  NAND2_X1 U14350 ( .A1(n11565), .A2(n13265), .ZN(n11400) );
  NAND2_X1 U14351 ( .A1(n11413), .A2(n11411), .ZN(n11397) );
  XNOR2_X1 U14352 ( .A(n11397), .B(n11410), .ZN(n11398) );
  NAND2_X1 U14353 ( .A1(n11398), .A2(n11440), .ZN(n11399) );
  NAND2_X1 U14354 ( .A1(n11400), .A2(n11399), .ZN(n19976) );
  NAND2_X1 U14355 ( .A1(n11401), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11402) );
  NAND2_X1 U14356 ( .A1(n19975), .A2(n11402), .ZN(n13918) );
  INV_X1 U14357 ( .A(n11403), .ZN(n11406) );
  INV_X1 U14358 ( .A(n11404), .ZN(n11405) );
  OAI21_X1 U14359 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n11408) );
  NAND2_X1 U14360 ( .A1(n11418), .A2(n11408), .ZN(n11570) );
  OR2_X1 U14361 ( .A1(n11570), .A2(n11409), .ZN(n11416) );
  AND2_X1 U14362 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  NAND2_X1 U14363 ( .A1(n11413), .A2(n11412), .ZN(n11419) );
  XNOR2_X1 U14364 ( .A(n11419), .B(n11420), .ZN(n11414) );
  NAND2_X1 U14365 ( .A1(n11414), .A2(n11440), .ZN(n11415) );
  NAND2_X1 U14366 ( .A1(n11416), .A2(n11415), .ZN(n11428) );
  INV_X1 U14367 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16138) );
  XNOR2_X1 U14368 ( .A(n11428), .B(n16138), .ZN(n16069) );
  NAND2_X1 U14369 ( .A1(n11418), .A2(n11417), .ZN(n11577) );
  NAND3_X1 U14370 ( .A1(n11435), .A2(n11577), .A3(n13265), .ZN(n11424) );
  INV_X1 U14371 ( .A(n11419), .ZN(n11421) );
  NAND2_X1 U14372 ( .A1(n11421), .A2(n11420), .ZN(n11436) );
  XNOR2_X1 U14373 ( .A(n11436), .B(n11437), .ZN(n11422) );
  NAND2_X1 U14374 ( .A1(n11422), .A2(n11440), .ZN(n11423) );
  NAND2_X1 U14375 ( .A1(n11424), .A2(n11423), .ZN(n13920) );
  INV_X1 U14376 ( .A(n11425), .ZN(n11427) );
  AND2_X1 U14377 ( .A1(n16069), .A2(n11427), .ZN(n11426) );
  NAND2_X1 U14378 ( .A1(n13918), .A2(n11426), .ZN(n11432) );
  NAND2_X1 U14379 ( .A1(n11428), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13919) );
  NAND2_X1 U14380 ( .A1(n13920), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11429) );
  AND2_X1 U14381 ( .A1(n13919), .A2(n11429), .ZN(n11430) );
  INV_X1 U14382 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U14383 ( .A1(n11502), .A2(n11439), .ZN(n11433) );
  OAI21_X1 U14384 ( .B1(n11519), .B2(n12084), .A(n11433), .ZN(n11434) );
  NAND2_X1 U14385 ( .A1(n11584), .A2(n13265), .ZN(n11443) );
  INV_X1 U14386 ( .A(n11436), .ZN(n11438) );
  NAND2_X1 U14387 ( .A1(n11438), .A2(n11437), .ZN(n11446) );
  XNOR2_X1 U14388 ( .A(n11446), .B(n11439), .ZN(n11441) );
  NAND2_X1 U14389 ( .A1(n11441), .A2(n11440), .ZN(n11442) );
  NAND2_X1 U14390 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  AND2_X1 U14391 ( .A1(n11444), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16061) );
  OR3_X1 U14392 ( .A1(n11446), .A2(n11445), .A3(n20744), .ZN(n11447) );
  NOR2_X1 U14393 ( .A1(n13996), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U14394 ( .A1(n13996), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11448) );
  INV_X1 U14395 ( .A(n14118), .ZN(n11450) );
  INV_X1 U14396 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16115) );
  NAND2_X1 U14397 ( .A1(n11450), .A2(n9870), .ZN(n14746) );
  NAND2_X1 U14398 ( .A1(n14748), .A2(n16115), .ZN(n11451) );
  NAND2_X2 U14399 ( .A1(n14746), .A2(n11451), .ZN(n14708) );
  INV_X1 U14400 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16088) );
  NAND2_X1 U14401 ( .A1(n14748), .A2(n16088), .ZN(n11452) );
  NAND2_X1 U14402 ( .A1(n14723), .A2(n11452), .ZN(n14739) );
  INV_X1 U14403 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11459) );
  AND2_X1 U14404 ( .A1(n14748), .A2(n11459), .ZN(n14737) );
  NOR2_X1 U14405 ( .A1(n14739), .A2(n14737), .ZN(n14722) );
  NAND2_X1 U14406 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14407 ( .A1(n14748), .A2(n11453), .ZN(n14735) );
  INV_X1 U14408 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U14409 ( .A1(n14748), .A2(n14926), .ZN(n11454) );
  AND2_X1 U14410 ( .A1(n14735), .A2(n11454), .ZN(n11455) );
  NAND2_X1 U14411 ( .A1(n14722), .A2(n11455), .ZN(n14709) );
  OR2_X1 U14412 ( .A1(n14748), .A2(n14926), .ZN(n11456) );
  INV_X1 U14413 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11457) );
  OR2_X1 U14414 ( .A1(n14748), .A2(n11457), .ZN(n14712) );
  XNOR2_X1 U14415 ( .A(n14751), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14715) );
  NAND2_X1 U14416 ( .A1(n14748), .A2(n11457), .ZN(n14713) );
  NAND2_X1 U14417 ( .A1(n14715), .A2(n14713), .ZN(n11458) );
  AOI21_X1 U14418 ( .B1(n14709), .B2(n14879), .A(n11458), .ZN(n14880) );
  INV_X1 U14419 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14747) );
  INV_X1 U14420 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14733) );
  AND3_X1 U14421 ( .A1(n11459), .A2(n14747), .A3(n14733), .ZN(n11460) );
  NAND2_X1 U14422 ( .A1(n11461), .A2(n14721), .ZN(n14710) );
  XNOR2_X1 U14423 ( .A(n14751), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14154) );
  NAND2_X1 U14424 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14850) );
  NAND2_X1 U14425 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14856) );
  NOR2_X1 U14426 ( .A1(n14850), .A2(n14856), .ZN(n14817) );
  INV_X1 U14427 ( .A(n14817), .ZN(n11464) );
  INV_X1 U14428 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11462) );
  INV_X1 U14429 ( .A(n11465), .ZN(n11469) );
  INV_X1 U14430 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14700) );
  INV_X1 U14431 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14699) );
  INV_X1 U14432 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14868) );
  NAND3_X1 U14433 ( .A1(n14700), .A2(n14699), .A3(n14868), .ZN(n11466) );
  OAI21_X2 U14434 ( .B1(n14693), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16052), .ZN(n14685) );
  NAND2_X1 U14435 ( .A1(n11469), .A2(n14751), .ZN(n14659) );
  NAND2_X1 U14436 ( .A1(n14659), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11470) );
  NOR2_X1 U14437 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14781) );
  NAND3_X1 U14438 ( .A1(n14653), .A2(n9604), .A3(n14781), .ZN(n14275) );
  INV_X1 U14439 ( .A(n11470), .ZN(n11472) );
  AND2_X1 U14440 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U14441 ( .A1(n14801), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14633) );
  NAND2_X1 U14442 ( .A1(n11472), .A2(n11471), .ZN(n14646) );
  NAND2_X1 U14443 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14780) );
  NOR2_X2 U14444 ( .A1(n14646), .A2(n14780), .ZN(n14274) );
  NAND2_X1 U14445 ( .A1(n14748), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14624) );
  INV_X1 U14446 ( .A(n14624), .ZN(n11473) );
  NAND2_X1 U14447 ( .A1(n14274), .A2(n11473), .ZN(n14276) );
  OAI21_X1 U14448 ( .B1(n14625), .B2(n14275), .A(n14276), .ZN(n11474) );
  XNOR2_X1 U14449 ( .A(n11474), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14768) );
  INV_X1 U14450 ( .A(n13261), .ZN(n13258) );
  NAND2_X1 U14451 ( .A1(n14962), .A2(n12156), .ZN(n11475) );
  INV_X1 U14452 ( .A(n11136), .ZN(n13346) );
  AND2_X1 U14453 ( .A1(n13363), .A2(n13346), .ZN(n15865) );
  XNOR2_X1 U14454 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14455 ( .A1(n11496), .A2(n11497), .ZN(n11477) );
  NAND2_X1 U14456 ( .A1(n20572), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11476) );
  NAND2_X1 U14457 ( .A1(n11477), .A2(n11476), .ZN(n11488) );
  XNOR2_X1 U14458 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U14459 ( .A1(n11488), .A2(n11487), .ZN(n11479) );
  NAND2_X1 U14460 ( .A1(n20320), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11478) );
  NAND2_X1 U14461 ( .A1(n11479), .A2(n11478), .ZN(n11509) );
  MUX2_X1 U14462 ( .A(n20125), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11508) );
  NAND2_X1 U14463 ( .A1(n11509), .A2(n11508), .ZN(n11481) );
  NAND2_X1 U14464 ( .A1(n20125), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14465 ( .A1(n11481), .A2(n11480), .ZN(n11485) );
  INV_X1 U14466 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16141) );
  NOR2_X1 U14467 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16141), .ZN(
        n11482) );
  OR2_X1 U14468 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20029), .ZN(
        n11483) );
  NAND2_X1 U14469 ( .A1(n11512), .A2(n12150), .ZN(n11524) );
  NAND2_X1 U14470 ( .A1(n12150), .A2(n11502), .ZN(n11522) );
  NOR3_X1 U14471 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20029), .A3(
        n11485), .ZN(n12146) );
  XNOR2_X1 U14472 ( .A(n11488), .B(n11487), .ZN(n12145) );
  INV_X1 U14473 ( .A(n12145), .ZN(n11511) );
  INV_X1 U14474 ( .A(n11496), .ZN(n11490) );
  NAND2_X1 U14475 ( .A1(n9848), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11489) );
  NAND2_X1 U14476 ( .A1(n11490), .A2(n11489), .ZN(n11491) );
  INV_X1 U14477 ( .A(n11491), .ZN(n11492) );
  AOI21_X1 U14478 ( .B1(n11502), .B2(n11492), .A(n11512), .ZN(n11493) );
  INV_X1 U14479 ( .A(n11502), .ZN(n11500) );
  XNOR2_X1 U14480 ( .A(n11497), .B(n11496), .ZN(n12148) );
  NOR2_X1 U14481 ( .A1(n20635), .A2(n20073), .ZN(n11501) );
  AOI21_X1 U14482 ( .B1(n12148), .B2(n11498), .A(n11501), .ZN(n11499) );
  OAI21_X1 U14483 ( .B1(n11495), .B2(n11500), .A(n11499), .ZN(n11503) );
  NAND2_X1 U14484 ( .A1(n11504), .A2(n11503), .ZN(n11506) );
  INV_X1 U14485 ( .A(n12148), .ZN(n11505) );
  NOR2_X1 U14486 ( .A1(n9640), .A2(n11507), .ZN(n11510) );
  XNOR2_X1 U14487 ( .A(n11509), .B(n11508), .ZN(n12144) );
  OAI22_X1 U14488 ( .A1(n11511), .A2(n11519), .B1(n11510), .B2(n12144), .ZN(
        n11517) );
  NAND2_X1 U14489 ( .A1(n11512), .A2(n12144), .ZN(n11515) );
  AOI21_X1 U14490 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20635), .A(
        n11520), .ZN(n11521) );
  NAND2_X1 U14491 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  AND2_X1 U14492 ( .A1(n11525), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13501) );
  INV_X2 U14493 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20638) );
  INV_X1 U14494 ( .A(n11526), .ZN(n14316) );
  NOR2_X1 U14495 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12165) );
  XNOR2_X1 U14496 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14361) );
  AOI21_X1 U14497 ( .B1(n12112), .B2(n14361), .A(n12160), .ZN(n11528) );
  NAND2_X1 U14498 ( .A1(n12161), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11527) );
  OAI211_X1 U14499 ( .C1(n11554), .C2(n11166), .A(n11528), .B(n11527), .ZN(
        n11529) );
  NAND2_X1 U14500 ( .A1(n12160), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11547) );
  INV_X1 U14501 ( .A(n13557), .ZN(n11546) );
  INV_X1 U14502 ( .A(n11530), .ZN(n11531) );
  NAND2_X1 U14503 ( .A1(n13703), .A2(n11734), .ZN(n11535) );
  INV_X1 U14504 ( .A(n11554), .ZN(n11557) );
  INV_X1 U14505 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11532) );
  INV_X1 U14506 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13853) );
  OAI22_X1 U14507 ( .A1(n11960), .A2(n11532), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13853), .ZN(n11533) );
  AOI21_X1 U14508 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11557), .A(
        n11533), .ZN(n11534) );
  NAND2_X1 U14509 ( .A1(n11535), .A2(n11534), .ZN(n13489) );
  AOI21_X1 U14510 ( .B1(n9632), .B2(n11108), .A(n20638), .ZN(n13331) );
  NAND2_X1 U14511 ( .A1(n20160), .A2(n11734), .ZN(n11542) );
  NAND2_X1 U14512 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20638), .ZN(
        n11539) );
  NAND2_X1 U14513 ( .A1(n12161), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11538) );
  OAI211_X1 U14514 ( .C1(n11554), .C2(n9848), .A(n11539), .B(n11538), .ZN(
        n11540) );
  INV_X1 U14515 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U14516 ( .A1(n11542), .A2(n11541), .ZN(n13330) );
  NAND2_X1 U14517 ( .A1(n13331), .A2(n13330), .ZN(n13329) );
  INV_X1 U14518 ( .A(n13330), .ZN(n11543) );
  NAND2_X1 U14519 ( .A1(n11543), .A2(n12112), .ZN(n11544) );
  NAND2_X1 U14520 ( .A1(n13329), .A2(n11544), .ZN(n13488) );
  NAND2_X1 U14521 ( .A1(n13489), .A2(n13488), .ZN(n13560) );
  INV_X1 U14522 ( .A(n13560), .ZN(n11545) );
  INV_X1 U14523 ( .A(n11549), .ZN(n11551) );
  INV_X1 U14524 ( .A(n11560), .ZN(n11550) );
  OAI21_X1 U14525 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11551), .A(
        n11550), .ZN(n13821) );
  AOI22_X1 U14526 ( .A1(n12112), .A2(n13821), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14527 ( .A1(n12161), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14528 ( .C1(n11554), .C2(n9759), .A(n11553), .B(n11552), .ZN(
        n11555) );
  INV_X1 U14529 ( .A(n11555), .ZN(n11556) );
  NAND2_X1 U14530 ( .A1(n11557), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11563) );
  INV_X1 U14531 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11558) );
  AOI21_X1 U14532 ( .B1(n11558), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11559) );
  AOI21_X1 U14533 ( .B1(n12161), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11559), .ZN(
        n11562) );
  NAND2_X1 U14534 ( .A1(n11560), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11566) );
  OAI21_X1 U14535 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11560), .A(
        n11566), .ZN(n19984) );
  NOR2_X1 U14536 ( .A1(n19984), .A2(n12079), .ZN(n11561) );
  AOI21_X1 U14537 ( .B1(n11563), .B2(n11562), .A(n11561), .ZN(n11564) );
  OAI21_X1 U14538 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11567), .A(
        n11571), .ZN(n19947) );
  AOI22_X1 U14539 ( .A1(n12112), .A2(n19947), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14540 ( .A1(n12161), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11568) );
  OAI211_X1 U14541 ( .C1(n11570), .C2(n11717), .A(n11569), .B(n11568), .ZN(
        n13630) );
  NAND2_X1 U14542 ( .A1(n13631), .A2(n13630), .ZN(n13629) );
  INV_X1 U14543 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11575) );
  INV_X1 U14544 ( .A(n11571), .ZN(n11573) );
  INV_X1 U14545 ( .A(n11580), .ZN(n11572) );
  OAI21_X1 U14546 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11573), .A(
        n11572), .ZN(n19923) );
  AOI22_X1 U14547 ( .A1(n12112), .A2(n19923), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11574) );
  OAI21_X1 U14548 ( .B1(n11960), .B2(n11575), .A(n11574), .ZN(n11576) );
  INV_X1 U14549 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14550 ( .A1(n11580), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11601) );
  OAI21_X1 U14551 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11580), .A(
        n11601), .ZN(n19907) );
  AOI22_X1 U14552 ( .A1(n12165), .A2(n19907), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11581) );
  OAI21_X1 U14553 ( .B1(n11960), .B2(n11582), .A(n11581), .ZN(n11583) );
  NAND2_X1 U14554 ( .A1(n12161), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14555 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11592) );
  INV_X1 U14556 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11587) );
  INV_X1 U14557 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11804) );
  OAI22_X1 U14558 ( .A1(n12028), .A2(n11587), .B1(n11979), .B2(n11804), .ZN(
        n11588) );
  INV_X1 U14559 ( .A(n11588), .ZN(n11591) );
  AOI22_X1 U14560 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14561 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11589) );
  AND4_X1 U14562 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11599) );
  AOI22_X1 U14563 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14564 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14565 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U14566 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11593) );
  AND3_X1 U14567 ( .A1(n11595), .A2(n11594), .A3(n11593), .ZN(n11597) );
  NAND2_X1 U14568 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11596) );
  NAND4_X1 U14569 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11600) );
  NAND2_X1 U14570 ( .A1(n11734), .A2(n11600), .ZN(n11603) );
  XNOR2_X1 U14571 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11605), .ZN(
        n14000) );
  AOI22_X1 U14572 ( .A1(n12165), .A2(n14000), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11602) );
  XNOR2_X1 U14573 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11637), .ZN(
        n14121) );
  INV_X1 U14574 ( .A(n14121), .ZN(n19893) );
  INV_X1 U14575 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U14576 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14577 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14578 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14579 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11606) );
  AND4_X1 U14580 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11616) );
  AOI22_X1 U14581 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14582 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11611) );
  NAND2_X1 U14583 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11610) );
  AND3_X1 U14584 ( .A1(n11612), .A2(n11611), .A3(n11610), .ZN(n11615) );
  AOI22_X1 U14585 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11614) );
  NAND2_X1 U14586 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11613) );
  NAND4_X1 U14587 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11617) );
  NAND2_X1 U14588 ( .A1(n11734), .A2(n11617), .ZN(n11619) );
  NAND2_X1 U14589 ( .A1(n12160), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11618) );
  OAI211_X1 U14590 ( .C1(n14024), .C2(n11960), .A(n11619), .B(n11618), .ZN(
        n11620) );
  AOI21_X1 U14591 ( .B1(n19893), .B2(n12165), .A(n11620), .ZN(n14019) );
  INV_X1 U14592 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U14593 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U14594 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11622) );
  OAI211_X1 U14595 ( .C1(n9617), .C2(n11776), .A(n11623), .B(n11622), .ZN(
        n11624) );
  INV_X1 U14596 ( .A(n11624), .ZN(n11628) );
  AOI22_X1 U14597 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14598 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11626) );
  NAND2_X1 U14599 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11625) );
  NAND4_X1 U14600 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11636) );
  INV_X1 U14601 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11773) );
  INV_X1 U14602 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11629) );
  OAI22_X1 U14603 ( .A1(n12028), .A2(n11773), .B1(n11177), .B2(n11629), .ZN(
        n11630) );
  INV_X1 U14604 ( .A(n11630), .ZN(n11634) );
  AOI22_X1 U14605 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14606 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14607 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11631) );
  NAND4_X1 U14608 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11631), .ZN(
        n11635) );
  NOR2_X1 U14609 ( .A1(n11636), .A2(n11635), .ZN(n11640) );
  XNOR2_X1 U14610 ( .A(n11654), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14755) );
  NAND2_X1 U14611 ( .A1(n14755), .A2(n12165), .ZN(n11639) );
  AOI22_X1 U14612 ( .A1(n12161), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12160), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11638) );
  OAI211_X1 U14613 ( .C1(n11640), .C2(n11717), .A(n11639), .B(n11638), .ZN(
        n14034) );
  AOI22_X1 U14614 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14615 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14616 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14617 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11642) );
  AND4_X1 U14618 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11652) );
  AOI22_X1 U14619 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14620 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14621 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14622 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11646) );
  AND3_X1 U14623 ( .A1(n11648), .A2(n11647), .A3(n11646), .ZN(n11650) );
  NAND2_X1 U14624 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11649) );
  NAND4_X1 U14625 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11653) );
  NAND2_X1 U14626 ( .A1(n11734), .A2(n11653), .ZN(n14554) );
  INV_X1 U14627 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11657) );
  INV_X1 U14628 ( .A(n12160), .ZN(n11675) );
  OAI21_X1 U14629 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11655), .A(
        n11694), .ZN(n16060) );
  NAND2_X1 U14630 ( .A1(n16060), .A2(n12165), .ZN(n11656) );
  OAI21_X1 U14631 ( .B1(n11657), .B2(n11675), .A(n11656), .ZN(n11658) );
  AOI21_X1 U14632 ( .B1(n12161), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11658), .ZN(
        n14136) );
  XNOR2_X1 U14633 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11714), .ZN(
        n16001) );
  AOI22_X1 U14634 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14635 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11661) );
  AND2_X1 U14636 ( .A1(n11662), .A2(n11661), .ZN(n11666) );
  AOI22_X1 U14637 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14638 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14639 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11663) );
  NAND4_X1 U14640 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11674) );
  AOI22_X1 U14641 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11672) );
  OAI22_X1 U14642 ( .A1(n12028), .A2(n11667), .B1(n11979), .B2(n10978), .ZN(
        n11668) );
  INV_X1 U14643 ( .A(n11668), .ZN(n11671) );
  AOI22_X1 U14644 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14645 ( .A1(n12035), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14646 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  NOR2_X1 U14647 ( .A1(n11674), .A2(n11673), .ZN(n11676) );
  INV_X1 U14648 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14740) );
  OAI22_X1 U14649 ( .A1(n11717), .A2(n11676), .B1(n11675), .B2(n14740), .ZN(
        n11678) );
  INV_X1 U14650 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14615) );
  NOR2_X1 U14651 ( .A1(n11960), .A2(n14615), .ZN(n11677) );
  NOR2_X1 U14652 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  OAI21_X1 U14653 ( .B1(n16001), .B2(n12079), .A(n11679), .ZN(n14539) );
  INV_X1 U14654 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U14655 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11685) );
  INV_X1 U14656 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11680) );
  OAI22_X1 U14657 ( .A1(n12028), .A2(n12007), .B1(n11177), .B2(n11680), .ZN(
        n11681) );
  INV_X1 U14658 ( .A(n11681), .ZN(n11684) );
  AOI22_X1 U14659 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14660 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11682) );
  AND4_X1 U14661 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11692) );
  AOI22_X1 U14662 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14663 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14664 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11687) );
  NAND2_X1 U14665 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11686) );
  AND3_X1 U14666 ( .A1(n11688), .A2(n11687), .A3(n11686), .ZN(n11690) );
  NAND2_X1 U14667 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11689) );
  NAND4_X1 U14668 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11693) );
  NAND2_X1 U14669 ( .A1(n11734), .A2(n11693), .ZN(n11697) );
  XNOR2_X1 U14670 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11694), .ZN(
        n16047) );
  INV_X1 U14671 ( .A(n16047), .ZN(n11695) );
  AOI22_X1 U14672 ( .A1(n12160), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12112), .B2(n11695), .ZN(n11696) );
  OAI211_X1 U14673 ( .C1(n14147), .C2(n11960), .A(n11697), .B(n11696), .ZN(
        n14138) );
  NAND2_X1 U14674 ( .A1(n14539), .A2(n14138), .ZN(n11698) );
  INV_X1 U14675 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11702) );
  OR2_X1 U14676 ( .A1(n12028), .A2(n11699), .ZN(n11701) );
  NAND2_X1 U14677 ( .A1(n12100), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11700) );
  OAI211_X1 U14678 ( .C1(n9617), .C2(n11702), .A(n11701), .B(n11700), .ZN(
        n11703) );
  INV_X1 U14679 ( .A(n11703), .ZN(n11707) );
  AOI22_X1 U14680 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11789), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14681 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11705) );
  NAND2_X1 U14682 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11704) );
  NAND4_X1 U14683 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11713) );
  AOI22_X1 U14684 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12096), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14685 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14686 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14687 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14688 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  NOR2_X1 U14689 ( .A1(n11713), .A2(n11712), .ZN(n11718) );
  XNOR2_X1 U14690 ( .A(n11719), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14727) );
  NAND2_X1 U14691 ( .A1(n14727), .A2(n12112), .ZN(n11716) );
  AOI22_X1 U14692 ( .A1(n12161), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12160), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11715) );
  OAI211_X1 U14693 ( .C1(n11718), .C2(n11717), .A(n11716), .B(n11715), .ZN(
        n14125) );
  NAND2_X1 U14694 ( .A1(n11719), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11739) );
  XNOR2_X1 U14695 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11739), .ZN(
        n16041) );
  AOI22_X1 U14696 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11725) );
  INV_X1 U14697 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11788) );
  OAI22_X1 U14698 ( .A1(n12028), .A2(n11720), .B1(n11979), .B2(n11788), .ZN(
        n11721) );
  INV_X1 U14699 ( .A(n11721), .ZN(n11724) );
  AOI22_X1 U14700 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14701 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11722) );
  AND4_X1 U14702 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11732) );
  AOI22_X1 U14703 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14704 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14705 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U14706 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11726) );
  AND3_X1 U14707 ( .A1(n11728), .A2(n11727), .A3(n11726), .ZN(n11730) );
  NAND2_X1 U14708 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11729) );
  NAND4_X1 U14709 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11733) );
  AOI22_X1 U14710 ( .A1(n11734), .A2(n11733), .B1(n12160), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11736) );
  NAND2_X1 U14711 ( .A1(n12161), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11735) );
  OAI211_X1 U14712 ( .C1(n16041), .C2(n12079), .A(n11736), .B(n11735), .ZN(
        n11737) );
  INV_X1 U14713 ( .A(n11737), .ZN(n14531) );
  INV_X1 U14714 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15990) );
  XNOR2_X1 U14715 ( .A(n11755), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14717) );
  NOR2_X1 U14716 ( .A1(n14962), .A2(n20635), .ZN(n12109) );
  AOI22_X1 U14717 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14718 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14719 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14720 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11740) );
  AND4_X1 U14721 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11750) );
  AOI22_X1 U14722 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14723 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14724 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11745) );
  NAND2_X1 U14725 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11744) );
  AND3_X1 U14726 ( .A1(n11746), .A2(n11745), .A3(n11744), .ZN(n11748) );
  NAND2_X1 U14727 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11747) );
  NAND4_X1 U14728 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  NAND2_X1 U14729 ( .A1(n12109), .A2(n11751), .ZN(n11753) );
  AOI22_X1 U14730 ( .A1(n12161), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20638), .ZN(n11752) );
  AOI21_X1 U14731 ( .B1(n11753), .B2(n11752), .A(n12112), .ZN(n11754) );
  AOI21_X1 U14732 ( .B1(n14717), .B2(n12112), .A(n11754), .ZN(n14445) );
  XOR2_X1 U14733 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11837), .Z(
        n16036) );
  AOI22_X1 U14734 ( .A1(n12161), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12160), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14735 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14736 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14737 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14738 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14739 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11769) );
  AND2_X1 U14740 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11763) );
  INV_X1 U14741 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11761) );
  OAI22_X1 U14742 ( .A1(n12028), .A2(n11761), .B1(n11979), .B2(n11760), .ZN(
        n11762) );
  NOR2_X1 U14743 ( .A1(n11763), .A2(n11762), .ZN(n11767) );
  AOI22_X1 U14744 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14745 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U14746 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11764) );
  NAND4_X1 U14747 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(
        n11768) );
  OAI21_X1 U14748 ( .B1(n11769), .B2(n11768), .A(n12109), .ZN(n11770) );
  OAI211_X1 U14749 ( .C1(n16036), .C2(n12079), .A(n11771), .B(n11770), .ZN(
        n14515) );
  INV_X1 U14750 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11781) );
  INV_X1 U14751 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11772) );
  OAI22_X1 U14752 ( .A1(n12008), .A2(n11773), .B1(n12087), .B2(n11772), .ZN(
        n11778) );
  INV_X1 U14753 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11774) );
  OAI22_X1 U14754 ( .A1(n12089), .A2(n11776), .B1(n11775), .B2(n11774), .ZN(
        n11777) );
  AOI211_X1 U14755 ( .C1(n12060), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11778), .B(n11777), .ZN(n11780) );
  AOI22_X1 U14756 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11779) );
  OAI211_X1 U14757 ( .C1(n12064), .C2(n11781), .A(n11780), .B(n11779), .ZN(
        n11787) );
  AOI22_X1 U14758 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14759 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14760 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14761 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11782) );
  NAND4_X1 U14762 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n11786) );
  NOR2_X1 U14763 ( .A1(n11787), .A2(n11786), .ZN(n11993) );
  INV_X1 U14764 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11796) );
  INV_X1 U14765 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U14766 ( .A1(n9586), .A2(n12095), .B1(n9592), .B2(n11788), .ZN(
        n11793) );
  INV_X1 U14767 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11791) );
  OAI22_X1 U14768 ( .A1(n12008), .A2(n11791), .B1(n11260), .B2(n11790), .ZN(
        n11792) );
  AOI211_X1 U14769 ( .C1(n11860), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11793), .B(n11792), .ZN(n11795) );
  AOI22_X1 U14770 ( .A1(n12035), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11794) );
  OAI211_X1 U14771 ( .C1(n9617), .C2(n11796), .A(n11795), .B(n11794), .ZN(
        n11802) );
  AOI22_X1 U14772 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14773 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14774 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14775 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11797) );
  NAND4_X1 U14776 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11801) );
  NOR2_X1 U14777 ( .A1(n11802), .A2(n11801), .ZN(n11845) );
  INV_X1 U14778 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11811) );
  OAI22_X1 U14779 ( .A1(n11260), .A2(n11804), .B1(n12085), .B2(n11803), .ZN(
        n11808) );
  INV_X1 U14780 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11806) );
  OAI22_X1 U14781 ( .A1(n12087), .A2(n11806), .B1(n11259), .B2(n11805), .ZN(
        n11807) );
  AOI211_X1 U14782 ( .C1(n11860), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11808), .B(n11807), .ZN(n11810) );
  AOI22_X1 U14783 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11809) );
  OAI211_X1 U14784 ( .C1(n9617), .C2(n11811), .A(n11810), .B(n11809), .ZN(
        n11817) );
  AOI22_X1 U14785 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14786 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14787 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14788 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U14789 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11816) );
  NOR2_X1 U14790 ( .A1(n11817), .A2(n11816), .ZN(n11846) );
  NOR2_X1 U14791 ( .A1(n11845), .A2(n11846), .ZN(n11966) );
  AOI22_X1 U14792 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14793 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U14794 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11818) );
  NAND3_X1 U14795 ( .A1(n11820), .A2(n11819), .A3(n11818), .ZN(n11826) );
  NAND2_X1 U14796 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11823) );
  INV_X1 U14797 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11821) );
  OR2_X1 U14798 ( .A1(n12028), .A2(n11821), .ZN(n11822) );
  OAI211_X1 U14799 ( .C1(n11824), .C2(n11177), .A(n11823), .B(n11822), .ZN(
        n11825) );
  NOR2_X1 U14800 ( .A1(n11826), .A2(n11825), .ZN(n11832) );
  AOI22_X1 U14801 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14802 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14803 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14804 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11827) );
  AND4_X1 U14805 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11831) );
  NAND2_X1 U14806 ( .A1(n11832), .A2(n11831), .ZN(n11965) );
  NAND2_X1 U14807 ( .A1(n11966), .A2(n11965), .ZN(n11992) );
  XNOR2_X1 U14808 ( .A(n11993), .B(n11992), .ZN(n11836) );
  INV_X1 U14809 ( .A(n12109), .ZN(n12076) );
  NAND2_X1 U14810 ( .A1(n20638), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11833) );
  NAND2_X1 U14811 ( .A1(n12079), .A2(n11833), .ZN(n11834) );
  AOI21_X1 U14812 ( .B1(n12161), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11834), .ZN(
        n11835) );
  OAI21_X1 U14813 ( .B1(n11836), .B2(n12076), .A(n11835), .ZN(n11844) );
  INV_X1 U14814 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15968) );
  INV_X1 U14815 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11871) );
  INV_X1 U14816 ( .A(n11839), .ZN(n11841) );
  INV_X1 U14817 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14818 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  NAND2_X1 U14819 ( .A1(n11998), .A2(n11842), .ZN(n15922) );
  OR2_X1 U14820 ( .A1(n15922), .A2(n12079), .ZN(n11843) );
  NAND2_X1 U14821 ( .A1(n11844), .A2(n11843), .ZN(n14480) );
  INV_X1 U14822 ( .A(n14480), .ZN(n11976) );
  XNOR2_X1 U14823 ( .A(n11846), .B(n11845), .ZN(n11850) );
  NAND2_X1 U14824 ( .A1(n20638), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11847) );
  NAND2_X1 U14825 ( .A1(n12079), .A2(n11847), .ZN(n11848) );
  AOI21_X1 U14826 ( .B1(n12161), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11848), .ZN(
        n11849) );
  OAI21_X1 U14827 ( .B1(n12076), .B2(n11850), .A(n11849), .ZN(n11855) );
  NOR2_X1 U14828 ( .A1(n11851), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11852) );
  OR2_X1 U14829 ( .A1(n11972), .A2(n11852), .ZN(n15932) );
  INV_X1 U14830 ( .A(n15932), .ZN(n11853) );
  NAND2_X1 U14831 ( .A1(n11853), .A2(n12112), .ZN(n11854) );
  AND2_X1 U14832 ( .A1(n11855), .A2(n11854), .ZN(n14575) );
  INV_X1 U14833 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11858) );
  OR2_X1 U14834 ( .A1(n11979), .A2(n10971), .ZN(n11857) );
  NAND2_X1 U14835 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11856) );
  OAI211_X1 U14836 ( .C1(n9617), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n11859) );
  INV_X1 U14837 ( .A(n11859), .ZN(n11864) );
  AOI22_X1 U14838 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12098), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14839 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11789), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11862) );
  NAND2_X1 U14840 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11861) );
  NAND4_X1 U14841 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11870) );
  AOI22_X1 U14842 ( .A1(n12097), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11919), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14843 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14844 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14845 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U14846 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11869) );
  NOR2_X1 U14847 ( .A1(n11870), .A2(n11869), .ZN(n11874) );
  AOI21_X1 U14848 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n11871), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11872) );
  AOI21_X1 U14849 ( .B1(n12161), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11872), .ZN(
        n11873) );
  OAI21_X1 U14850 ( .B1(n12076), .B2(n11874), .A(n11873), .ZN(n11876) );
  XNOR2_X1 U14851 ( .A(n11912), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14687) );
  NAND2_X1 U14852 ( .A1(n14687), .A2(n12165), .ZN(n11875) );
  NAND2_X1 U14853 ( .A1(n11876), .A2(n11875), .ZN(n14435) );
  AOI22_X1 U14854 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11944), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14855 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14856 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14857 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11877) );
  AND4_X1 U14858 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11887) );
  AOI22_X1 U14859 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14860 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14861 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11882) );
  NAND2_X1 U14862 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11881) );
  AND3_X1 U14863 ( .A1(n11883), .A2(n11882), .A3(n11881), .ZN(n11885) );
  NAND2_X1 U14864 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11884) );
  NAND4_X1 U14865 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n11888) );
  NAND2_X1 U14866 ( .A1(n12109), .A2(n11888), .ZN(n11891) );
  INV_X1 U14867 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15959) );
  OAI21_X1 U14868 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15959), .A(n12079), 
        .ZN(n11889) );
  AOI21_X1 U14869 ( .B1(n12161), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11889), .ZN(
        n11890) );
  NAND2_X1 U14870 ( .A1(n11891), .A2(n11890), .ZN(n11893) );
  XNOR2_X1 U14871 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11917), .ZN(
        n15953) );
  NAND2_X1 U14872 ( .A1(n12112), .A2(n15953), .ZN(n11892) );
  NAND2_X1 U14873 ( .A1(n11893), .A2(n11892), .ZN(n14501) );
  AND2_X1 U14874 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11897) );
  INV_X1 U14875 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11895) );
  OAI22_X1 U14876 ( .A1(n12028), .A2(n11895), .B1(n11979), .B2(n11894), .ZN(
        n11896) );
  NOR2_X1 U14877 ( .A1(n11897), .A2(n11896), .ZN(n11901) );
  AOI22_X1 U14878 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14879 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U14880 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11898) );
  NAND4_X1 U14881 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11907) );
  AOI22_X1 U14882 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14883 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14884 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14885 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U14886 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11906) );
  NOR2_X1 U14887 ( .A1(n11907), .A2(n11906), .ZN(n11911) );
  NAND2_X1 U14888 ( .A1(n20638), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U14889 ( .A1(n12079), .A2(n11908), .ZN(n11909) );
  AOI21_X1 U14890 ( .B1(n12161), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11909), .ZN(
        n11910) );
  OAI21_X1 U14891 ( .B1(n12076), .B2(n11911), .A(n11910), .ZN(n11915) );
  OAI21_X1 U14892 ( .B1(n11913), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11912), .ZN(n15942) );
  OR2_X1 U14893 ( .A1(n15942), .A2(n12079), .ZN(n11914) );
  NAND2_X1 U14894 ( .A1(n11915), .A2(n11914), .ZN(n14497) );
  OR2_X1 U14895 ( .A1(n14501), .A2(n14497), .ZN(n14431) );
  OR2_X1 U14896 ( .A1(n14435), .A2(n14431), .ZN(n11942) );
  OR2_X1 U14897 ( .A1(n11916), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U14898 ( .A1(n11918), .A2(n11917), .ZN(n16035) );
  INV_X1 U14899 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11922) );
  NAND2_X1 U14900 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U14901 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11920) );
  OAI211_X1 U14902 ( .C1(n9617), .C2(n11922), .A(n11921), .B(n11920), .ZN(
        n11923) );
  INV_X1 U14903 ( .A(n11923), .ZN(n11927) );
  AOI22_X1 U14904 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14905 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U14906 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11924) );
  NAND4_X1 U14907 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11936) );
  INV_X1 U14908 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11929) );
  OAI22_X1 U14909 ( .A1(n12028), .A2(n11929), .B1(n11177), .B2(n11928), .ZN(
        n11930) );
  INV_X1 U14910 ( .A(n11930), .ZN(n11934) );
  AOI22_X1 U14911 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11789), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14912 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14913 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U14914 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  NOR2_X1 U14915 ( .A1(n11936), .A2(n11935), .ZN(n11940) );
  NAND2_X1 U14916 ( .A1(n20638), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U14917 ( .A1(n12079), .A2(n11937), .ZN(n11938) );
  AOI21_X1 U14918 ( .B1(n12161), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11938), .ZN(
        n11939) );
  OAI21_X1 U14919 ( .B1(n12076), .B2(n11940), .A(n11939), .ZN(n11941) );
  OAI21_X1 U14920 ( .B1(n16035), .B2(n12079), .A(n11941), .ZN(n14507) );
  NOR2_X1 U14921 ( .A1(n11942), .A2(n14507), .ZN(n14433) );
  AND2_X1 U14922 ( .A1(n14575), .A2(n14433), .ZN(n11964) );
  XNOR2_X1 U14923 ( .A(n11943), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15973) );
  AOI22_X1 U14924 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14925 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14926 ( .A1(n9601), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U14927 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11945) );
  AND4_X1 U14928 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11956) );
  AOI22_X1 U14929 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U14930 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14931 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U14932 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11950) );
  AND3_X1 U14933 ( .A1(n11952), .A2(n11951), .A3(n11950), .ZN(n11954) );
  NAND2_X1 U14934 ( .A1(n12060), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11953) );
  NAND4_X1 U14935 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(
        n11962) );
  INV_X1 U14936 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n11959) );
  AOI21_X1 U14937 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15968), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11957) );
  INV_X1 U14938 ( .A(n11957), .ZN(n11958) );
  OAI21_X1 U14939 ( .B1(n11960), .B2(n11959), .A(n11958), .ZN(n11961) );
  AOI21_X1 U14940 ( .B1(n12109), .B2(n11962), .A(n11961), .ZN(n11963) );
  AOI21_X1 U14941 ( .B1(n15973), .B2(n12112), .A(n11963), .ZN(n14432) );
  XNOR2_X1 U14942 ( .A(n11966), .B(n11965), .ZN(n11970) );
  NAND2_X1 U14943 ( .A1(n20638), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U14944 ( .A1(n12079), .A2(n11967), .ZN(n11968) );
  AOI21_X1 U14945 ( .B1(n12161), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11968), .ZN(
        n11969) );
  OAI21_X1 U14946 ( .B1(n11970), .B2(n12076), .A(n11969), .ZN(n11974) );
  INV_X1 U14947 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11971) );
  XNOR2_X1 U14948 ( .A(n11972), .B(n11971), .ZN(n14670) );
  NAND2_X1 U14949 ( .A1(n14670), .A2(n12112), .ZN(n11973) );
  NAND2_X1 U14950 ( .A1(n11974), .A2(n11973), .ZN(n14421) );
  INV_X1 U14951 ( .A(n14421), .ZN(n11975) );
  INV_X1 U14952 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11980) );
  OAI22_X1 U14953 ( .A1(n12028), .A2(n11980), .B1(n11979), .B2(n11978), .ZN(
        n11985) );
  INV_X1 U14954 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U14955 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U14956 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11981) );
  OAI211_X1 U14957 ( .C1(n9617), .C2(n11983), .A(n11982), .B(n11981), .ZN(
        n11984) );
  AOI211_X1 U14958 ( .C1(n11860), .C2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11985), .B(n11984), .ZN(n11991) );
  AOI22_X1 U14959 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U14960 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U14961 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U14962 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11986) );
  AND4_X1 U14963 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11990) );
  NAND2_X1 U14964 ( .A1(n11991), .A2(n11990), .ZN(n12004) );
  NOR2_X1 U14965 ( .A1(n11993), .A2(n11992), .ZN(n12005) );
  XOR2_X1 U14966 ( .A(n12004), .B(n12005), .Z(n11994) );
  NAND2_X1 U14967 ( .A1(n11994), .A2(n12109), .ZN(n11997) );
  INV_X1 U14968 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14655) );
  NOR2_X1 U14969 ( .A1(n14655), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11995) );
  AOI211_X1 U14970 ( .C1(n12161), .C2(P1_EAX_REG_26__SCAN_IN), .A(n12112), .B(
        n11995), .ZN(n11996) );
  XNOR2_X1 U14971 ( .A(n11998), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15912) );
  AOI22_X1 U14972 ( .A1(n11997), .A2(n11996), .B1(n12112), .B2(n15912), .ZN(
        n14473) );
  INV_X1 U14973 ( .A(n11998), .ZN(n11999) );
  INV_X1 U14974 ( .A(n12000), .ZN(n12002) );
  INV_X1 U14975 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U14976 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  NAND2_X1 U14977 ( .A1(n12049), .A2(n12003), .ZN(n14643) );
  NAND2_X1 U14978 ( .A1(n12005), .A2(n12004), .ZN(n12043) );
  INV_X1 U14979 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12015) );
  OAI22_X1 U14980 ( .A1(n12008), .A2(n12007), .B1(n12085), .B2(n12006), .ZN(
        n12012) );
  INV_X1 U14981 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12010) );
  OAI22_X1 U14982 ( .A1(n12087), .A2(n12010), .B1(n9592), .B2(n12009), .ZN(
        n12011) );
  AOI211_X1 U14983 ( .C1(n12060), .C2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n12012), .B(n12011), .ZN(n12014) );
  AOI22_X1 U14984 ( .A1(n9590), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12013) );
  OAI211_X1 U14985 ( .C1(n12064), .C2(n12015), .A(n12014), .B(n12013), .ZN(
        n12021) );
  AOI22_X1 U14986 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U14987 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U14988 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U14989 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U14990 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  NOR2_X1 U14991 ( .A1(n12021), .A2(n12020), .ZN(n12044) );
  XNOR2_X1 U14992 ( .A(n12043), .B(n12044), .ZN(n12024) );
  AOI21_X1 U14993 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20638), .A(
        n12165), .ZN(n12023) );
  NAND2_X1 U14994 ( .A1(n12161), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12022) );
  OAI211_X1 U14995 ( .C1(n12024), .C2(n12076), .A(n12023), .B(n12022), .ZN(
        n12025) );
  OAI21_X1 U14996 ( .B1(n12079), .B2(n14643), .A(n12025), .ZN(n14212) );
  INV_X1 U14997 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12027) );
  OAI22_X1 U14998 ( .A1(n12028), .A2(n12027), .B1(n11177), .B2(n12026), .ZN(
        n12034) );
  INV_X1 U14999 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15000 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12029), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15001 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12030) );
  OAI211_X1 U15002 ( .C1(n9617), .C2(n12032), .A(n12031), .B(n12030), .ZN(
        n12033) );
  AOI211_X1 U15003 ( .C1(n11860), .C2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12034), .B(n12033), .ZN(n12042) );
  AOI22_X1 U15004 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15005 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15006 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12035), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15007 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12036), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12037) );
  AND4_X1 U15008 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12041) );
  NAND2_X1 U15009 ( .A1(n12042), .A2(n12041), .ZN(n12072) );
  NOR2_X1 U15010 ( .A1(n12044), .A2(n12043), .ZN(n12073) );
  XOR2_X1 U15011 ( .A(n12072), .B(n12073), .Z(n12045) );
  NAND2_X1 U15012 ( .A1(n12045), .A2(n12109), .ZN(n12048) );
  INV_X1 U15013 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14637) );
  NOR2_X1 U15014 ( .A1(n14637), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12046) );
  AOI211_X1 U15015 ( .C1(n12161), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12165), .B(
        n12046), .ZN(n12047) );
  XNOR2_X1 U15016 ( .A(n12049), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14641) );
  AOI22_X1 U15017 ( .A1(n12048), .A2(n12047), .B1(n12112), .B2(n14641), .ZN(
        n14409) );
  NAND2_X1 U15018 ( .A1(n14211), .A2(n14409), .ZN(n14395) );
  INV_X1 U15019 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U15020 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  NAND2_X1 U15021 ( .A1(n12170), .A2(n12052), .ZN(n14629) );
  INV_X1 U15022 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12063) );
  INV_X1 U15023 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12054) );
  INV_X1 U15024 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12053) );
  OAI22_X1 U15025 ( .A1(n12054), .A2(n11260), .B1(n12085), .B2(n12053), .ZN(
        n12059) );
  INV_X1 U15026 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12056) );
  INV_X1 U15027 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12055) );
  OAI22_X1 U15028 ( .A1(n9586), .A2(n12056), .B1(n12087), .B2(n12055), .ZN(
        n12058) );
  AOI211_X1 U15029 ( .C1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .C2(n12060), .A(
        n12059), .B(n12058), .ZN(n12062) );
  AOI22_X1 U15030 ( .A1(n12096), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12061) );
  OAI211_X1 U15031 ( .C1(n9626), .C2(n12063), .A(n12062), .B(n12061), .ZN(
        n12071) );
  AOI22_X1 U15032 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9636), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15033 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15034 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12065), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15035 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9591), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U15036 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12070) );
  NOR2_X1 U15037 ( .A1(n12071), .A2(n12070), .ZN(n12081) );
  NAND2_X1 U15038 ( .A1(n12073), .A2(n12072), .ZN(n12080) );
  XNOR2_X1 U15039 ( .A(n12081), .B(n12080), .ZN(n12077) );
  AOI21_X1 U15040 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20638), .A(
        n12165), .ZN(n12075) );
  NAND2_X1 U15041 ( .A1(n12161), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12074) );
  OAI211_X1 U15042 ( .C1(n12077), .C2(n12076), .A(n12075), .B(n12074), .ZN(
        n12078) );
  OAI21_X1 U15043 ( .B1(n12079), .B2(n14629), .A(n12078), .ZN(n14397) );
  NOR2_X1 U15044 ( .A1(n12081), .A2(n12080), .ZN(n12108) );
  OAI22_X1 U15045 ( .A1(n12085), .A2(n12084), .B1(n9592), .B2(n12082), .ZN(
        n12091) );
  INV_X1 U15046 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12088) );
  INV_X1 U15047 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12086) );
  OAI22_X1 U15048 ( .A1(n12089), .A2(n12088), .B1(n12087), .B2(n12086), .ZN(
        n12090) );
  AOI211_X1 U15049 ( .C1(n11860), .C2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12091), .B(n12090), .ZN(n12094) );
  AOI22_X1 U15050 ( .A1(n11944), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12092), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12093) );
  OAI211_X1 U15051 ( .C1(n9617), .C2(n12095), .A(n12094), .B(n12093), .ZN(
        n12106) );
  AOI22_X1 U15052 ( .A1(n9624), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12096), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15053 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15054 ( .A1(n12099), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9601), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15055 ( .A1(n9636), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12100), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15056 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12105) );
  NOR2_X1 U15057 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  XNOR2_X1 U15058 ( .A(n12108), .B(n12107), .ZN(n12110) );
  NAND2_X1 U15059 ( .A1(n12110), .A2(n12109), .ZN(n12115) );
  INV_X1 U15060 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12169) );
  AOI21_X1 U15061 ( .B1(n12169), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12111) );
  AOI21_X1 U15062 ( .B1(n12161), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12111), .ZN(
        n12114) );
  XNOR2_X1 U15063 ( .A(n12170), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14384) );
  AND2_X1 U15064 ( .A1(n14384), .A2(n12112), .ZN(n12113) );
  AOI21_X1 U15065 ( .B1(n12115), .B2(n12114), .A(n12113), .ZN(n12162) );
  AND2_X1 U15066 ( .A1(n20635), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U15067 ( .A1(n12166), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16145) );
  NOR2_X2 U15068 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20499) );
  INV_X1 U15069 ( .A(n14384), .ZN(n12122) );
  OR2_X1 U15070 ( .A1(n12119), .A2(n20499), .ZN(n20740) );
  AND2_X1 U15071 ( .A1(n20740), .A2(n20635), .ZN(n12116) );
  NAND2_X1 U15072 ( .A1(n20635), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15875) );
  INV_X1 U15073 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20496) );
  NAND2_X1 U15074 ( .A1(n20496), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12117) );
  AND2_X1 U15075 ( .A1(n15875), .A2(n12117), .ZN(n13332) );
  INV_X1 U15076 ( .A(n13332), .ZN(n12118) );
  NAND2_X1 U15077 ( .A1(n19973), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14764) );
  OAI21_X1 U15078 ( .B1(n14741), .B2(n12169), .A(n14764), .ZN(n12120) );
  INV_X1 U15079 ( .A(n12120), .ZN(n12121) );
  OAI21_X1 U15080 ( .B1(n12122), .B2(n19985), .A(n12121), .ZN(n12123) );
  INV_X1 U15081 ( .A(n12123), .ZN(n12124) );
  AND2_X1 U15082 ( .A1(n19203), .A2(n19721), .ZN(n12125) );
  NAND2_X1 U15083 ( .A1(n12126), .A2(n12125), .ZN(n13110) );
  INV_X1 U15084 ( .A(n13110), .ZN(n12127) );
  NAND2_X1 U15085 ( .A1(n12127), .A2(n19849), .ZN(n19194) );
  NOR2_X2 U15086 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19800) );
  OR2_X1 U15087 ( .A1(n19800), .A2(n19799), .ZN(n19815) );
  NAND2_X1 U15088 ( .A1(n19815), .A2(n19716), .ZN(n12129) );
  AND2_X1 U15089 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19816) );
  NAND2_X1 U15090 ( .A1(n19716), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12387) );
  INV_X1 U15091 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19847) );
  NAND2_X1 U15092 ( .A1(n19847), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12130) );
  NAND2_X1 U15093 ( .A1(n12387), .A2(n12130), .ZN(n13310) );
  INV_X1 U15094 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16235) );
  NAND2_X1 U15095 ( .A1(n12334), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12332) );
  NAND2_X1 U15096 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n12331), .ZN(
        n12343) );
  INV_X1 U15097 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15307) );
  INV_X1 U15098 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15290) );
  AND2_X1 U15099 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12132) );
  INV_X1 U15100 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15262) );
  INV_X1 U15101 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15231) );
  INV_X1 U15102 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15237) );
  NOR2_X1 U15103 ( .A1(n15231), .A2(n15237), .ZN(n12133) );
  AND2_X1 U15104 ( .A1(n12133), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12134) );
  AND2_X1 U15105 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12135) );
  INV_X1 U15106 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15192) );
  INV_X1 U15107 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12310) );
  XNOR2_X1 U15108 ( .A(n12312), .B(n12310), .ZN(n14260) );
  NAND2_X1 U15109 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12136) );
  OAI211_X1 U15110 ( .C1(n19191), .C2(n14260), .A(n12137), .B(n12136), .ZN(
        n12138) );
  AOI21_X1 U15111 ( .B1(n12673), .B2(n19198), .A(n12138), .ZN(n12139) );
  INV_X1 U15112 ( .A(n12139), .ZN(n12140) );
  NOR2_X1 U15113 ( .A1(n9869), .A2(n12140), .ZN(n12141) );
  OAI21_X1 U15114 ( .B1(n12142), .B2(n19194), .A(n12141), .ZN(P2_U2984) );
  INV_X1 U15115 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20675) );
  INV_X1 U15116 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20661) );
  OR3_X1 U15117 ( .A1(n12146), .A2(n12145), .A3(n12144), .ZN(n12147) );
  NOR2_X1 U15118 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  NOR2_X1 U15119 ( .A1(n12150), .A2(n12149), .ZN(n13496) );
  INV_X1 U15120 ( .A(n13496), .ZN(n12151) );
  NOR2_X1 U15121 ( .A1(n12143), .A2(n12151), .ZN(n13252) );
  NAND2_X1 U15122 ( .A1(n13252), .A2(n13501), .ZN(n13227) );
  INV_X1 U15123 ( .A(n12152), .ZN(n13348) );
  NOR2_X1 U15124 ( .A1(n13817), .A2(n11136), .ZN(n12153) );
  NAND2_X1 U15125 ( .A1(n14311), .A2(n12154), .ZN(n12155) );
  INV_X1 U15126 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20650) );
  NAND2_X1 U15127 ( .A1(n12157), .A2(n20650), .ZN(n15900) );
  INV_X1 U15128 ( .A(n15900), .ZN(n13459) );
  OR2_X1 U15129 ( .A1(n20054), .A2(n13459), .ZN(n13503) );
  NAND2_X1 U15130 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20741) );
  AND2_X1 U15131 ( .A1(n20741), .A2(n20496), .ZN(n12289) );
  NAND2_X1 U15132 ( .A1(n13503), .A2(n12289), .ZN(n15877) );
  INV_X1 U15133 ( .A(n15877), .ZN(n12158) );
  INV_X1 U15134 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20659) );
  NAND3_X1 U15135 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19954) );
  NOR2_X1 U15136 ( .A1(n20659), .A2(n19954), .ZN(n12296) );
  NAND2_X1 U15137 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19927), .ZN(n19917) );
  NAND2_X1 U15138 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n12159) );
  NAND3_X1 U15139 ( .A1(n19899), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16020) );
  INV_X1 U15140 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20669) );
  INV_X1 U15141 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20678) );
  NAND2_X1 U15142 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15960) );
  NOR2_X2 U15143 ( .A1(n15975), .A2(n15960), .ZN(n15956) );
  NAND2_X1 U15144 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n12299) );
  INV_X1 U15145 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20694) );
  AND2_X1 U15146 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n12300) );
  NAND2_X1 U15147 ( .A1(n15925), .A2(n12300), .ZN(n14414) );
  INV_X1 U15148 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20700) );
  INV_X1 U15149 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20704) );
  OR3_X2 U15150 ( .A1(n14414), .A2(n20700), .A3(n20704), .ZN(n14408) );
  INV_X1 U15151 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14383) );
  INV_X1 U15152 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20702) );
  AOI22_X1 U15153 ( .A1(n12161), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12160), .ZN(n12164) );
  NAND2_X1 U15154 ( .A1(n14396), .A2(n12162), .ZN(n12163) );
  XOR2_X1 U15155 ( .A(n12164), .B(n12163), .Z(n14315) );
  NAND2_X1 U15156 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  NAND2_X1 U15157 ( .A1(n20638), .A2(n20634), .ZN(n16149) );
  INV_X1 U15158 ( .A(n16149), .ZN(n20745) );
  NAND3_X1 U15159 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_3__SCAN_IN), .A3(n20745), .ZN(n15887) );
  NAND2_X1 U15160 ( .A1(n12167), .A2(n15887), .ZN(n12168) );
  NOR2_X1 U15161 ( .A1(n12170), .A2(n12169), .ZN(n12171) );
  XNOR2_X1 U15162 ( .A(n12171), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14304) );
  NOR2_X1 U15163 ( .A1(n14304), .A2(n20634), .ZN(n12172) );
  OR2_X1 U15164 ( .A1(n12279), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12180) );
  INV_X1 U15165 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U15166 ( .A1(n9633), .A2(n13730), .ZN(n12178) );
  INV_X1 U15167 ( .A(n20064), .ZN(n12175) );
  INV_X1 U15168 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U15169 ( .A1(n12189), .A2(n20012), .ZN(n12177) );
  NAND3_X1 U15170 ( .A1(n12178), .A2(n12177), .A3(n14380), .ZN(n12179) );
  NAND2_X1 U15171 ( .A1(n12189), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12182) );
  INV_X1 U15172 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13738) );
  NAND2_X1 U15173 ( .A1(n14380), .A2(n13738), .ZN(n12181) );
  NAND2_X1 U15174 ( .A1(n12182), .A2(n12181), .ZN(n13517) );
  OR2_X1 U15175 ( .A1(n12279), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12186) );
  INV_X1 U15176 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13866) );
  NAND2_X1 U15177 ( .A1(n9633), .A2(n13866), .ZN(n12184) );
  NAND2_X1 U15178 ( .A1(n12189), .A2(n20026), .ZN(n12183) );
  NAND3_X1 U15179 ( .A1(n12184), .A2(n12183), .A3(n14380), .ZN(n12185) );
  NAND2_X1 U15180 ( .A1(n12186), .A2(n12185), .ZN(n13862) );
  MUX2_X1 U15181 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12188) );
  OR2_X1 U15182 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12187) );
  OR2_X1 U15183 ( .A1(n12279), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U15184 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12190) );
  NAND2_X1 U15185 ( .A1(n12190), .A2(n12189), .ZN(n12193) );
  INV_X1 U15186 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15187 ( .A1(n9633), .A2(n12191), .ZN(n12192) );
  NAND2_X1 U15188 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  INV_X1 U15189 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13874) );
  NAND2_X1 U15190 ( .A1(n9633), .A2(n13874), .ZN(n12199) );
  NAND2_X1 U15191 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12198) );
  NAND3_X1 U15192 ( .A1(n12199), .A2(n12189), .A3(n12198), .ZN(n12200) );
  OAI21_X1 U15193 ( .B1(n12276), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12200), .ZN(
        n13869) );
  OR2_X1 U15194 ( .A1(n12279), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U15195 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12201) );
  NAND2_X1 U15196 ( .A1(n12201), .A2(n12189), .ZN(n12204) );
  INV_X1 U15197 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n12202) );
  NAND2_X1 U15198 ( .A1(n9633), .A2(n12202), .ZN(n12203) );
  NAND2_X1 U15199 ( .A1(n12204), .A2(n12203), .ZN(n12205) );
  NAND2_X1 U15200 ( .A1(n12206), .A2(n12205), .ZN(n13796) );
  OR2_X1 U15201 ( .A1(n12276), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12210) );
  INV_X1 U15202 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13891) );
  NAND2_X1 U15203 ( .A1(n9633), .A2(n13891), .ZN(n12208) );
  NAND2_X1 U15204 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12207) );
  NAND3_X1 U15205 ( .A1(n12208), .A2(n12189), .A3(n12207), .ZN(n12209) );
  OR2_X1 U15206 ( .A1(n12279), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U15207 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U15208 ( .A1(n12211), .A2(n12189), .ZN(n12214) );
  INV_X1 U15209 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U15210 ( .A1(n9633), .A2(n12212), .ZN(n12213) );
  NAND2_X1 U15211 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  INV_X1 U15212 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19972) );
  NAND2_X1 U15213 ( .A1(n9633), .A2(n19972), .ZN(n12218) );
  NAND2_X1 U15214 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12217) );
  NAND3_X1 U15215 ( .A1(n12218), .A2(n12189), .A3(n12217), .ZN(n12219) );
  OAI21_X1 U15216 ( .B1(n12276), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12219), .ZN(
        n16105) );
  OR2_X1 U15217 ( .A1(n12279), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12223) );
  INV_X1 U15218 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U15219 ( .A1(n9633), .A2(n14044), .ZN(n12221) );
  NAND2_X1 U15220 ( .A1(n12189), .A2(n14747), .ZN(n12220) );
  NAND3_X1 U15221 ( .A1(n12221), .A2(n12220), .A3(n14380), .ZN(n12222) );
  MUX2_X1 U15222 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12224) );
  MUX2_X1 U15223 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12226) );
  OR2_X1 U15224 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U15225 ( .A1(n12226), .A2(n12225), .ZN(n14544) );
  INV_X1 U15226 ( .A(n14544), .ZN(n12233) );
  OR2_X1 U15227 ( .A1(n12279), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n12232) );
  NAND2_X1 U15228 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12227) );
  NAND2_X1 U15229 ( .A1(n12227), .A2(n12189), .ZN(n12230) );
  INV_X1 U15230 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U15231 ( .A1(n9633), .A2(n12228), .ZN(n12229) );
  NAND2_X1 U15232 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U15233 ( .A1(n12232), .A2(n12231), .ZN(n14543) );
  NAND2_X1 U15234 ( .A1(n12233), .A2(n14543), .ZN(n12234) );
  OR2_X1 U15235 ( .A1(n12279), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n12238) );
  INV_X1 U15236 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14536) );
  NAND2_X1 U15237 ( .A1(n9633), .A2(n14536), .ZN(n12236) );
  NAND2_X1 U15238 ( .A1(n12189), .A2(n14926), .ZN(n12235) );
  NAND3_X1 U15239 ( .A1(n12236), .A2(n12235), .A3(n14380), .ZN(n12237) );
  MUX2_X1 U15240 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12240) );
  OR2_X1 U15241 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12239) );
  AND2_X1 U15242 ( .A1(n12240), .A2(n12239), .ZN(n14527) );
  OR2_X1 U15243 ( .A1(n12279), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12244) );
  INV_X1 U15244 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U15245 ( .A1(n9633), .A2(n14524), .ZN(n12242) );
  INV_X1 U15246 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14883) );
  NAND2_X1 U15247 ( .A1(n12189), .A2(n14883), .ZN(n12241) );
  NAND3_X1 U15248 ( .A1(n12242), .A2(n12241), .A3(n14380), .ZN(n12243) );
  NAND2_X1 U15249 ( .A1(n12244), .A2(n12243), .ZN(n14449) );
  MUX2_X1 U15250 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12245) );
  OAI21_X1 U15251 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13516), .A(
        n12245), .ZN(n14519) );
  OR2_X1 U15252 ( .A1(n12279), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12249) );
  INV_X1 U15253 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U15254 ( .A1(n9633), .A2(n14512), .ZN(n12247) );
  NAND2_X1 U15255 ( .A1(n12189), .A2(n14699), .ZN(n12246) );
  NAND3_X1 U15256 ( .A1(n12247), .A2(n12246), .A3(n14380), .ZN(n12248) );
  AND2_X1 U15257 ( .A1(n12249), .A2(n12248), .ZN(n14158) );
  MUX2_X1 U15258 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12250) );
  OAI21_X1 U15259 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13516), .A(
        n12250), .ZN(n14510) );
  OR2_X1 U15260 ( .A1(n12279), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U15261 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12251) );
  NAND2_X1 U15262 ( .A1(n12251), .A2(n12189), .ZN(n12254) );
  INV_X1 U15263 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n12252) );
  NAND2_X1 U15264 ( .A1(n9633), .A2(n12252), .ZN(n12253) );
  NAND2_X1 U15265 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NAND2_X1 U15266 ( .A1(n12256), .A2(n12255), .ZN(n14502) );
  MUX2_X1 U15267 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12257) );
  OAI21_X1 U15268 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13516), .A(
        n12257), .ZN(n14494) );
  OR2_X1 U15269 ( .A1(n12279), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12261) );
  INV_X1 U15270 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U15271 ( .A1(n9633), .A2(n14491), .ZN(n12259) );
  NAND2_X1 U15272 ( .A1(n12189), .A2(n11462), .ZN(n12258) );
  NAND3_X1 U15273 ( .A1(n12259), .A2(n12258), .A3(n14380), .ZN(n12260) );
  AND2_X1 U15274 ( .A1(n12261), .A2(n12260), .ZN(n14436) );
  INV_X1 U15275 ( .A(n12276), .ZN(n12262) );
  INV_X1 U15276 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n20759) );
  NAND2_X1 U15277 ( .A1(n12262), .A2(n20759), .ZN(n12266) );
  NAND2_X1 U15278 ( .A1(n9633), .A2(n20759), .ZN(n12264) );
  NAND2_X1 U15279 ( .A1(n14380), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12263) );
  NAND3_X1 U15280 ( .A1(n12264), .A2(n12189), .A3(n12263), .ZN(n12265) );
  AND2_X1 U15281 ( .A1(n12266), .A2(n12265), .ZN(n14830) );
  OR2_X1 U15282 ( .A1(n12279), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12270) );
  INV_X1 U15283 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14488) );
  NAND2_X1 U15284 ( .A1(n9633), .A2(n14488), .ZN(n12268) );
  NAND2_X1 U15285 ( .A1(n12189), .A2(n11468), .ZN(n12267) );
  NAND3_X1 U15286 ( .A1(n12268), .A2(n12267), .A3(n14380), .ZN(n12269) );
  NAND2_X1 U15287 ( .A1(n12270), .A2(n12269), .ZN(n14423) );
  MUX2_X1 U15288 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12271) );
  NAND2_X1 U15289 ( .A1(n9888), .A2(n12271), .ZN(n14486) );
  OR2_X1 U15290 ( .A1(n12279), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12275) );
  INV_X1 U15291 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U15292 ( .A1(n9633), .A2(n14477), .ZN(n12273) );
  INV_X1 U15293 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14803) );
  NAND2_X1 U15294 ( .A1(n12189), .A2(n14803), .ZN(n12272) );
  NAND3_X1 U15295 ( .A1(n12273), .A2(n12272), .A3(n14380), .ZN(n12274) );
  AND2_X1 U15296 ( .A1(n12275), .A2(n12274), .ZN(n14474) );
  MUX2_X1 U15297 ( .A(n12276), .B(n14380), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12278) );
  OR2_X1 U15298 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12277) );
  AND2_X1 U15299 ( .A1(n12278), .A2(n12277), .ZN(n14213) );
  OR2_X1 U15300 ( .A1(n12279), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12283) );
  INV_X1 U15301 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U15302 ( .A1(n9633), .A2(n14468), .ZN(n12281) );
  INV_X1 U15303 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14784) );
  NAND2_X1 U15304 ( .A1(n12189), .A2(n14784), .ZN(n12280) );
  NAND3_X1 U15305 ( .A1(n12281), .A2(n12280), .A3(n14380), .ZN(n12282) );
  NAND2_X1 U15306 ( .A1(n12283), .A2(n12282), .ZN(n14410) );
  INV_X1 U15307 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14467) );
  NAND2_X1 U15308 ( .A1(n9633), .A2(n14467), .ZN(n12285) );
  OR2_X1 U15309 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12284) );
  NAND2_X1 U15310 ( .A1(n12284), .A2(n12285), .ZN(n14379) );
  MUX2_X1 U15311 ( .A(n12285), .B(n14379), .S(n14380), .Z(n14399) );
  INV_X1 U15312 ( .A(n9633), .ZN(n13729) );
  NAND2_X1 U15313 ( .A1(n13729), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12287) );
  NAND2_X1 U15314 ( .A1(n13516), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U15315 ( .A1(n12287), .A2(n12286), .ZN(n14381) );
  AOI22_X1 U15316 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13729), .B1(
        n13516), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U15317 ( .A1(n20054), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12291) );
  NOR2_X1 U15318 ( .A1(n12291), .A2(n12289), .ZN(n12290) );
  AND2_X1 U15319 ( .A1(n15877), .A2(n12291), .ZN(n12292) );
  AND2_X2 U15320 ( .A1(n12293), .A2(n12292), .ZN(n19955) );
  AOI22_X1 U15321 ( .A1(n19955), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19953), .ZN(n12294) );
  OAI21_X1 U15322 ( .B1(n14466), .B2(n19948), .A(n12294), .ZN(n12295) );
  NAND2_X1 U15323 ( .A1(n14363), .A2(n14357), .ZN(n19932) );
  INV_X1 U15324 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20692) );
  INV_X1 U15325 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20677) );
  NAND2_X1 U15326 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n12297) );
  INV_X1 U15327 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20663) );
  NAND2_X1 U15328 ( .A1(n12296), .A2(n14357), .ZN(n19931) );
  NOR3_X1 U15329 ( .A1(n20663), .A2(n20661), .A3(n19931), .ZN(n19904) );
  NAND3_X1 U15330 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n19904), .ZN(n13977) );
  NOR2_X1 U15331 ( .A1(n12297), .A2(n13977), .ZN(n14058) );
  NAND3_X1 U15332 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n14058), .ZN(n15995) );
  NOR3_X1 U15333 ( .A1(n20677), .A2(n20675), .A3(n15995), .ZN(n14127) );
  NAND4_X1 U15334 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n14127), .ZN(n15961) );
  NOR2_X1 U15335 ( .A1(n15960), .A2(n15961), .ZN(n12298) );
  INV_X1 U15336 ( .A(n19932), .ZN(n19905) );
  AOI221_X1 U15337 ( .B1(n12299), .B2(n19932), .C1(n20692), .C2(n19932), .A(
        n15957), .ZN(n14425) );
  NAND2_X1 U15338 ( .A1(n12300), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n12301) );
  NAND2_X1 U15339 ( .A1(n19932), .A2(n12301), .ZN(n12302) );
  NAND2_X1 U15340 ( .A1(n14425), .A2(n12302), .ZN(n15913) );
  NAND2_X1 U15341 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n12303) );
  AND2_X1 U15342 ( .A1(n19932), .A2(n12303), .ZN(n12304) );
  NAND2_X1 U15343 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12305) );
  AND2_X1 U15344 ( .A1(n19932), .A2(n12305), .ZN(n12306) );
  NAND4_X1 U15345 ( .A1(n9657), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        P1_U2809) );
  INV_X1 U15346 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14341) );
  INV_X1 U15347 ( .A(n12312), .ZN(n12313) );
  AOI21_X1 U15348 ( .B1(n12311), .B2(n15192), .A(n12313), .ZN(n16154) );
  AND2_X1 U15349 ( .A1(n12314), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12315) );
  OAI21_X1 U15350 ( .B1(n12315), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12311), .ZN(n15208) );
  INV_X1 U15351 ( .A(n15208), .ZN(n14975) );
  INV_X1 U15352 ( .A(n12314), .ZN(n12318) );
  AOI21_X1 U15353 ( .B1(n15216), .B2(n12318), .A(n12315), .ZN(n16166) );
  NAND2_X1 U15354 ( .A1(n12316), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12321) );
  OR2_X1 U15355 ( .A1(n12321), .A2(n15237), .ZN(n12319) );
  NAND2_X1 U15356 ( .A1(n12319), .A2(n15231), .ZN(n12317) );
  AND2_X1 U15357 ( .A1(n12318), .A2(n12317), .ZN(n15229) );
  INV_X1 U15358 ( .A(n12319), .ZN(n12320) );
  AOI21_X1 U15359 ( .B1(n15237), .B2(n12321), .A(n12320), .ZN(n15235) );
  OAI21_X1 U15360 ( .B1(n12316), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12321), .ZN(n12322) );
  INV_X1 U15361 ( .A(n12322), .ZN(n15256) );
  AOI21_X1 U15362 ( .B1(n15262), .B2(n12323), .A(n12316), .ZN(n15260) );
  NAND2_X1 U15363 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12324), .ZN(
        n12327) );
  INV_X1 U15364 ( .A(n12327), .ZN(n12325) );
  AND2_X1 U15365 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12325), .ZN(
        n12326) );
  OAI21_X1 U15366 ( .B1(n12326), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12323), .ZN(n15282) );
  INV_X1 U15367 ( .A(n15282), .ZN(n15033) );
  AOI21_X1 U15368 ( .B1(n12327), .B2(n14189), .A(n12326), .ZN(n14192) );
  OAI21_X1 U15369 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12324), .A(
        n12327), .ZN(n14233) );
  INV_X1 U15370 ( .A(n14233), .ZN(n15051) );
  AOI21_X1 U15371 ( .B1(n15290), .B2(n9671), .A(n12324), .ZN(n18916) );
  OR2_X1 U15372 ( .A1(n12344), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12328) );
  NAND2_X1 U15373 ( .A1(n9671), .A2(n12328), .ZN(n18936) );
  AOI21_X1 U15374 ( .B1(n10801), .B2(n12330), .A(n12331), .ZN(n18971) );
  AOI21_X1 U15375 ( .B1(n10795), .B2(n12340), .A(n12342), .ZN(n13084) );
  NOR2_X1 U15376 ( .A1(n10778), .A2(n12332), .ZN(n12341) );
  AOI21_X1 U15377 ( .B1(n10778), .B2(n12332), .A(n12341), .ZN(n18987) );
  AOI21_X1 U15378 ( .B1(n16235), .B2(n12333), .A(n12334), .ZN(n18998) );
  AOI21_X1 U15379 ( .B1(n15350), .B2(n12335), .A(n9677), .ZN(n19008) );
  AOI21_X1 U15380 ( .B1(n16256), .B2(n12336), .A(n12337), .ZN(n19039) );
  NOR2_X1 U15381 ( .A1(n10080), .A2(n12338), .ZN(n12339) );
  AOI21_X1 U15382 ( .B1(n10080), .B2(n12338), .A(n12339), .ZN(n16257) );
  INV_X1 U15383 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19059) );
  AOI22_X1 U15384 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13790), .B1(n19059), 
        .B2(n19716), .ZN(n19047) );
  INV_X1 U15385 ( .A(n19047), .ZN(n13791) );
  INV_X1 U15386 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13547) );
  OAI22_X1 U15387 ( .A1(n19716), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13547), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13553) );
  AND2_X1 U15388 ( .A1(n13791), .A2(n13553), .ZN(n13432) );
  OAI21_X1 U15389 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12338), .ZN(n19190) );
  NAND2_X1 U15390 ( .A1(n13432), .A2(n19190), .ZN(n13446) );
  NOR2_X1 U15391 ( .A1(n16257), .A2(n13446), .ZN(n13419) );
  OAI21_X1 U15392 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12339), .A(
        n12336), .ZN(n19189) );
  NAND2_X1 U15393 ( .A1(n13419), .A2(n19189), .ZN(n19037) );
  NOR2_X1 U15394 ( .A1(n19039), .A2(n19037), .ZN(n19022) );
  OAI21_X1 U15395 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12337), .A(
        n12335), .ZN(n19024) );
  NAND2_X1 U15396 ( .A1(n19022), .A2(n19024), .ZN(n19007) );
  NOR2_X1 U15397 ( .A1(n19008), .A2(n19007), .ZN(n13407) );
  OAI21_X1 U15398 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9677), .A(
        n12333), .ZN(n16250) );
  NAND2_X1 U15399 ( .A1(n13407), .A2(n16250), .ZN(n18997) );
  NOR2_X1 U15400 ( .A1(n18998), .A2(n18997), .ZN(n13616) );
  OAI21_X1 U15401 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12334), .A(
        n12332), .ZN(n16228) );
  NAND2_X1 U15402 ( .A1(n13616), .A2(n16228), .ZN(n18986) );
  NOR2_X1 U15403 ( .A1(n18987), .A2(n18986), .ZN(n18979) );
  OAI21_X1 U15404 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12341), .A(
        n12340), .ZN(n18980) );
  NAND2_X1 U15405 ( .A1(n18979), .A2(n18980), .ZN(n13083) );
  NOR2_X1 U15406 ( .A1(n13084), .A2(n13083), .ZN(n13955) );
  OAI21_X1 U15407 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12342), .A(
        n12330), .ZN(n16205) );
  NAND2_X1 U15408 ( .A1(n13955), .A2(n16205), .ZN(n18969) );
  NOR2_X1 U15409 ( .A1(n18971), .A2(n18969), .ZN(n18955) );
  OAI21_X1 U15410 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12331), .A(
        n12343), .ZN(n18956) );
  AND2_X1 U15411 ( .A1(n18955), .A2(n18956), .ZN(n18951) );
  AOI21_X1 U15412 ( .B1(n15307), .B2(n12343), .A(n12344), .ZN(n12345) );
  INV_X1 U15413 ( .A(n12345), .ZN(n18950) );
  NAND2_X1 U15414 ( .A1(n18951), .A2(n18950), .ZN(n12346) );
  NOR2_X1 U15415 ( .A1(n18916), .A2(n18917), .ZN(n18915) );
  NOR2_X1 U15416 ( .A1(n12329), .A2(n18915), .ZN(n15050) );
  NOR2_X1 U15417 ( .A1(n15051), .A2(n15050), .ZN(n15049) );
  NOR2_X1 U15418 ( .A1(n12329), .A2(n15049), .ZN(n13055) );
  NOR2_X1 U15419 ( .A1(n15260), .A2(n13068), .ZN(n13067) );
  NOR2_X1 U15420 ( .A1(n12329), .A2(n13067), .ZN(n15016) );
  NOR2_X1 U15421 ( .A1(n15229), .A2(n14987), .ZN(n14986) );
  NOR2_X1 U15422 ( .A1(n12329), .A2(n14986), .ZN(n16167) );
  NOR2_X1 U15423 ( .A1(n16154), .A2(n16155), .ZN(n14259) );
  NOR2_X1 U15424 ( .A1(n12329), .A2(n14259), .ZN(n12348) );
  XNOR2_X1 U15425 ( .A(n12348), .B(n14260), .ZN(n12349) );
  NOR3_X1 U15426 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15904) );
  NAND2_X1 U15427 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15904), .ZN(n19724) );
  NAND2_X1 U15428 ( .A1(n12349), .A2(n19042), .ZN(n12372) );
  NAND2_X1 U15429 ( .A1(n16341), .A2(n13099), .ZN(n12366) );
  INV_X1 U15430 ( .A(n12366), .ZN(n19858) );
  NOR2_X1 U15431 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19853), .ZN(n12356) );
  INV_X1 U15432 ( .A(n12356), .ZN(n12363) );
  NOR2_X1 U15433 ( .A1(n12350), .A2(n12363), .ZN(n12351) );
  INV_X1 U15434 ( .A(n12352), .ZN(n16368) );
  AND2_X1 U15435 ( .A1(n16368), .A2(n13099), .ZN(n13112) );
  INV_X1 U15436 ( .A(n13108), .ZN(n13178) );
  NOR2_X1 U15437 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13178), .ZN(n16367) );
  NAND2_X1 U15438 ( .A1(n19852), .A2(n13789), .ZN(n15903) );
  NOR3_X1 U15439 ( .A1(n19716), .A2(n19240), .A3(n15903), .ZN(n16366) );
  NOR2_X1 U15440 ( .A1(n19042), .A2(n16366), .ZN(n12353) );
  AND2_X1 U15441 ( .A1(n18941), .A2(n12353), .ZN(n12354) );
  INV_X1 U15442 ( .A(n19030), .ZN(n19048) );
  AOI22_X1 U15443 ( .A1(n19036), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        n19048), .B2(P2_REIP_REG_30__SCAN_IN), .ZN(n12360) );
  INV_X1 U15444 ( .A(n16367), .ZN(n12355) );
  NAND2_X1 U15445 ( .A1(n13161), .A2(n12355), .ZN(n14267) );
  NOR2_X1 U15446 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12356), .ZN(n12357) );
  NAND2_X1 U15447 ( .A1(n13112), .A2(n12357), .ZN(n12358) );
  NAND2_X1 U15448 ( .A1(n14267), .A2(n12358), .ZN(n19049) );
  NAND2_X1 U15449 ( .A1(n19049), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12359) );
  OAI211_X1 U15450 ( .C1(n14352), .C2(n19046), .A(n12360), .B(n12359), .ZN(
        n12361) );
  AOI21_X1 U15451 ( .B1(n12673), .B2(n19041), .A(n12361), .ZN(n12370) );
  INV_X1 U15452 ( .A(n12362), .ZN(n12368) );
  NAND3_X1 U15453 ( .A1(n12364), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12363), 
        .ZN(n12365) );
  NAND2_X1 U15454 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  NAND2_X1 U15455 ( .A1(n12372), .A2(n12371), .ZN(P2_U2825) );
  NAND2_X1 U15456 ( .A1(n19224), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15457 ( .A1(n12403), .A2(n19240), .ZN(n12397) );
  NAND2_X1 U15458 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19300) );
  INV_X1 U15459 ( .A(n19300), .ZN(n19529) );
  INV_X1 U15460 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19807) );
  NAND2_X1 U15461 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19807), .ZN(
        n19396) );
  INV_X1 U15462 ( .A(n19396), .ZN(n12373) );
  NAND2_X1 U15463 ( .A1(n19529), .A2(n12373), .ZN(n15714) );
  NOR2_X1 U15464 ( .A1(n12395), .A2(n19824), .ZN(n15721) );
  NAND2_X1 U15465 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15721), .ZN(
        n15688) );
  NAND2_X1 U15466 ( .A1(n15688), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12374) );
  NAND2_X1 U15467 ( .A1(n15714), .A2(n12374), .ZN(n12375) );
  AND2_X1 U15468 ( .A1(n12375), .A2(n19800), .ZN(n19558) );
  AOI21_X1 U15469 ( .B1(n12397), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19558), .ZN(n12382) );
  INV_X1 U15470 ( .A(n12382), .ZN(n12378) );
  NAND2_X1 U15471 ( .A1(n12378), .A2(n12380), .ZN(n12406) );
  INV_X1 U15472 ( .A(n12387), .ZN(n12394) );
  NAND2_X1 U15473 ( .A1(n12379), .A2(n12394), .ZN(n12384) );
  INV_X1 U15474 ( .A(n12380), .ZN(n12381) );
  AND2_X1 U15475 ( .A1(n12382), .A2(n12381), .ZN(n12383) );
  NAND2_X1 U15476 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  AOI22_X1 U15477 ( .A1(n12397), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19800), .B2(n19833), .ZN(n12386) );
  XNOR2_X1 U15478 ( .A(n13219), .B(n12390), .ZN(n13248) );
  NAND2_X1 U15479 ( .A1(n12397), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12388) );
  NAND2_X1 U15480 ( .A1(n19824), .A2(n19833), .ZN(n19441) );
  AND2_X1 U15481 ( .A1(n19300), .A2(n19441), .ZN(n19331) );
  NAND2_X1 U15482 ( .A1(n19331), .A2(n19800), .ZN(n19500) );
  NAND2_X1 U15483 ( .A1(n12388), .A2(n19500), .ZN(n12389) );
  INV_X1 U15484 ( .A(n12390), .ZN(n12391) );
  NOR2_X1 U15485 ( .A1(n13219), .A2(n12391), .ZN(n12392) );
  NAND2_X1 U15486 ( .A1(n19300), .A2(n12395), .ZN(n12396) );
  AND2_X1 U15487 ( .A1(n12396), .A2(n15688), .ZN(n19332) );
  AOI22_X1 U15488 ( .A1(n12397), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19800), .B2(n19332), .ZN(n12398) );
  NAND2_X1 U15489 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  INV_X1 U15490 ( .A(n12403), .ZN(n12404) );
  NAND2_X1 U15491 ( .A1(n12404), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12405) );
  AOI22_X1 U15492 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15493 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15494 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15495 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15496 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12417) );
  AOI22_X1 U15497 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15498 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15499 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15500 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15501 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  NOR2_X1 U15502 ( .A1(n12417), .A2(n12416), .ZN(n14016) );
  INV_X1 U15503 ( .A(n14016), .ZN(n12445) );
  AOI22_X1 U15504 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15505 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15506 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15507 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10604), .B1(
        n9593), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U15508 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12427) );
  AOI22_X1 U15509 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10300), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15511 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12513), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15512 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12422) );
  NAND4_X1 U15513 ( .A1(n12425), .A2(n12424), .A3(n12423), .A4(n12422), .ZN(
        n12426) );
  NOR2_X1 U15514 ( .A1(n12427), .A2(n12426), .ZN(n13992) );
  INV_X1 U15515 ( .A(n13992), .ZN(n12444) );
  AOI22_X1 U15516 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10211), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15517 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15518 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15519 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10604), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12428) );
  NAND4_X1 U15520 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12437) );
  AOI22_X1 U15521 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10300), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15522 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12512), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15523 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12513), .B1(
        n10159), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12432) );
  NAND4_X1 U15525 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12436) );
  OR2_X1 U15526 ( .A1(n12437), .A2(n12436), .ZN(n13846) );
  OR2_X1 U15527 ( .A1(n13663), .A2(n13601), .ZN(n13661) );
  OR2_X1 U15528 ( .A1(n12438), .A2(n13661), .ZN(n13832) );
  OR2_X1 U15529 ( .A1(n12439), .A2(n13832), .ZN(n12440) );
  NOR2_X1 U15530 ( .A1(n12440), .A2(n13532), .ZN(n13844) );
  AND2_X1 U15531 ( .A1(n13846), .A2(n13844), .ZN(n12443) );
  AND4_X1 U15532 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__7__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12441) );
  NAND4_X1 U15533 ( .A1(n13722), .A2(n13777), .A3(n13774), .A4(n12441), .ZN(
        n12442) );
  NOR2_X1 U15534 ( .A1(n13397), .A2(n12442), .ZN(n13531) );
  AOI22_X1 U15535 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15536 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15537 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15538 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10604), .B1(
        n9593), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U15539 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12456) );
  AOI22_X1 U15540 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15541 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10259), .B1(
        n12512), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15542 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15543 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10160), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12451) );
  NAND4_X1 U15544 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12455) );
  OR2_X1 U15545 ( .A1(n12456), .A2(n12455), .ZN(n14048) );
  AOI22_X1 U15546 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15547 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15548 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15549 ( .A1(n9593), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15550 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12466) );
  AOI22_X1 U15551 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15552 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15553 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15554 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15555 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12465) );
  OR2_X1 U15556 ( .A1(n12466), .A2(n12465), .ZN(n15116) );
  AOI22_X1 U15557 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15558 ( .A1(n9628), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15559 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U15560 ( .A1(n9594), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12467) );
  NAND4_X1 U15561 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12476) );
  AOI22_X1 U15562 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15563 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15564 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15565 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12471) );
  NAND4_X1 U15566 ( .A1(n12474), .A2(n12473), .A3(n12472), .A4(n12471), .ZN(
        n12475) );
  NOR2_X1 U15567 ( .A1(n12476), .A2(n12475), .ZN(n14068) );
  AOI22_X1 U15568 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10154), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15569 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15570 ( .A1(n12478), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15571 ( .A1(n9593), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12479) );
  NAND4_X1 U15572 ( .A1(n12482), .A2(n12481), .A3(n12480), .A4(n12479), .ZN(
        n12489) );
  AOI22_X1 U15573 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15682), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15574 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15575 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15576 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15577 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12488) );
  NOR2_X1 U15578 ( .A1(n12489), .A2(n12488), .ZN(n15112) );
  AOI22_X1 U15579 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15580 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15581 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12496) );
  NAND2_X1 U15582 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U15583 ( .A1(n12649), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12493) );
  AND2_X1 U15584 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12492) );
  OR2_X1 U15585 ( .A1(n12492), .A2(n12491), .ZN(n12661) );
  AND3_X1 U15586 ( .A1(n12494), .A2(n12493), .A3(n12661), .ZN(n12495) );
  NAND4_X1 U15587 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12506) );
  AOI22_X1 U15588 ( .A1(n12658), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15589 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15590 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12502) );
  INV_X1 U15591 ( .A(n12661), .ZN(n12635) );
  NAND2_X1 U15592 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12500) );
  NAND2_X1 U15593 ( .A1(n12649), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12499) );
  AND3_X1 U15594 ( .A1(n12635), .A2(n12500), .A3(n12499), .ZN(n12501) );
  NAND4_X1 U15595 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12505) );
  NAND2_X1 U15596 ( .A1(n12506), .A2(n12505), .ZN(n12545) );
  NOR2_X1 U15597 ( .A1(n10566), .A2(n12545), .ZN(n12522) );
  AOI22_X1 U15598 ( .A1(n9630), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12478), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15599 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10168), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15600 ( .A1(n10154), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10153), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15601 ( .A1(n15682), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9594), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12508) );
  NAND4_X1 U15602 ( .A1(n12511), .A2(n12510), .A3(n12509), .A4(n12508), .ZN(
        n12521) );
  AOI22_X1 U15603 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15604 ( .A1(n12512), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10259), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15605 ( .A1(n10159), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12513), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15606 ( .A1(n10160), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12514), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12516) );
  NAND4_X1 U15607 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12520) );
  NOR2_X1 U15608 ( .A1(n12521), .A2(n12520), .ZN(n12539) );
  XNOR2_X1 U15609 ( .A(n12522), .B(n12539), .ZN(n12543) );
  XNOR2_X1 U15610 ( .A(n15111), .B(n12543), .ZN(n15107) );
  INV_X1 U15611 ( .A(n12545), .ZN(n12540) );
  NAND2_X1 U15612 ( .A1(n10566), .A2(n12540), .ZN(n15106) );
  AOI22_X1 U15613 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15614 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9583), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15615 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9930), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15616 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U15617 ( .A1(n12649), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12525) );
  AND3_X1 U15618 ( .A1(n12526), .A2(n12525), .A3(n12661), .ZN(n12527) );
  NAND4_X1 U15619 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n12538) );
  AOI22_X1 U15620 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15621 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15622 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12531) );
  AND3_X1 U15623 ( .A1(n12635), .A2(n12532), .A3(n12531), .ZN(n12535) );
  AOI22_X1 U15624 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15625 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12533) );
  NAND4_X1 U15626 ( .A1(n12536), .A2(n12535), .A3(n12534), .A4(n12533), .ZN(
        n12537) );
  NAND2_X1 U15627 ( .A1(n12538), .A2(n12537), .ZN(n12548) );
  INV_X1 U15628 ( .A(n12539), .ZN(n12541) );
  NAND2_X1 U15629 ( .A1(n12541), .A2(n12540), .ZN(n12549) );
  XOR2_X1 U15630 ( .A(n12548), .B(n12549), .Z(n12542) );
  NAND2_X1 U15631 ( .A1(n12542), .A2(n12606), .ZN(n15099) );
  INV_X1 U15632 ( .A(n12543), .ZN(n12546) );
  INV_X1 U15633 ( .A(n12548), .ZN(n12544) );
  NAND2_X1 U15634 ( .A1(n10566), .A2(n12544), .ZN(n15102) );
  NOR3_X1 U15635 ( .A1(n12546), .A2(n12545), .A3(n15102), .ZN(n12547) );
  NOR2_X1 U15636 ( .A1(n12549), .A2(n12548), .ZN(n12564) );
  AOI22_X1 U15637 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15638 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15639 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12553) );
  NAND2_X1 U15640 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U15641 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12550) );
  AND3_X1 U15642 ( .A1(n12551), .A2(n12550), .A3(n12661), .ZN(n12552) );
  NAND4_X1 U15643 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12563) );
  AOI22_X1 U15644 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15645 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12632), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U15646 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12557) );
  NAND2_X1 U15647 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12556) );
  AND3_X1 U15648 ( .A1(n12635), .A2(n12557), .A3(n12556), .ZN(n12559) );
  AOI22_X1 U15649 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12558) );
  NAND4_X1 U15650 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12562) );
  AND2_X1 U15651 ( .A1(n12563), .A2(n12562), .ZN(n12565) );
  NAND2_X1 U15652 ( .A1(n12564), .A2(n12565), .ZN(n12603) );
  OAI211_X1 U15653 ( .C1(n12564), .C2(n12565), .A(n12606), .B(n12603), .ZN(
        n12567) );
  INV_X1 U15654 ( .A(n12565), .ZN(n12566) );
  NOR2_X1 U15655 ( .A1(n19849), .A2(n12566), .ZN(n15093) );
  NAND2_X1 U15656 ( .A1(n15094), .A2(n15093), .ZN(n15092) );
  NAND2_X1 U15657 ( .A1(n15092), .A2(n12569), .ZN(n12586) );
  AOI22_X1 U15658 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U15659 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U15660 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12571) );
  AND3_X1 U15661 ( .A1(n12635), .A2(n12572), .A3(n12571), .ZN(n12575) );
  AOI22_X1 U15662 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15663 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12636), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U15664 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12584) );
  AOI22_X1 U15665 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15666 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15667 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15668 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12578) );
  NAND2_X1 U15669 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12577) );
  AND3_X1 U15670 ( .A1(n12578), .A2(n12577), .A3(n12661), .ZN(n12579) );
  NAND4_X1 U15671 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12583) );
  AND2_X1 U15672 ( .A1(n12584), .A2(n12583), .ZN(n12601) );
  XNOR2_X1 U15673 ( .A(n12603), .B(n12601), .ZN(n12585) );
  NAND2_X1 U15674 ( .A1(n10566), .A2(n12601), .ZN(n15087) );
  AOI22_X1 U15675 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15676 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9583), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15677 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U15678 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U15679 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12587) );
  AND3_X1 U15680 ( .A1(n12588), .A2(n12587), .A3(n12661), .ZN(n12589) );
  NAND4_X1 U15681 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12600) );
  AOI22_X1 U15682 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U15683 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12594) );
  NAND2_X1 U15684 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12593) );
  AND3_X1 U15685 ( .A1(n12635), .A2(n12594), .A3(n12593), .ZN(n12597) );
  AOI22_X1 U15686 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15687 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U15688 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12599) );
  NAND2_X1 U15689 ( .A1(n12600), .A2(n12599), .ZN(n12604) );
  INV_X1 U15690 ( .A(n12604), .ZN(n12609) );
  INV_X1 U15691 ( .A(n12601), .ZN(n12602) );
  OR2_X1 U15692 ( .A1(n12603), .A2(n12602), .ZN(n12605) );
  INV_X1 U15693 ( .A(n12605), .ZN(n12607) );
  OR2_X1 U15694 ( .A1(n12605), .A2(n12604), .ZN(n15071) );
  OAI211_X1 U15695 ( .C1(n12609), .C2(n12607), .A(n15071), .B(n12606), .ZN(
        n12608) );
  NAND2_X1 U15696 ( .A1(n10566), .A2(n12609), .ZN(n15082) );
  AOI22_X1 U15697 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U15698 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U15699 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12610) );
  AND3_X1 U15700 ( .A1(n12635), .A2(n12611), .A3(n12610), .ZN(n12614) );
  AOI22_X1 U15701 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15702 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9930), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12612) );
  NAND4_X1 U15703 ( .A1(n12615), .A2(n12614), .A3(n12613), .A4(n12612), .ZN(
        n12623) );
  AOI22_X1 U15704 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15705 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15706 ( .A1(n10001), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12636), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U15707 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U15708 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12616) );
  AND3_X1 U15709 ( .A1(n12617), .A2(n12616), .A3(n12661), .ZN(n12618) );
  NAND4_X1 U15710 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12622) );
  AND2_X1 U15711 ( .A1(n12623), .A2(n12622), .ZN(n15073) );
  OAI21_X1 U15712 ( .B1(n15081), .B2(n12624), .A(n15073), .ZN(n15068) );
  NAND2_X1 U15713 ( .A1(n19849), .A2(n15073), .ZN(n12625) );
  NOR2_X1 U15714 ( .A1(n15071), .A2(n12625), .ZN(n12644) );
  AOI22_X1 U15715 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15716 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9618), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12630) );
  INV_X1 U15717 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U15718 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12655), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12629) );
  NAND2_X1 U15719 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12627) );
  NAND2_X1 U15720 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12626) );
  AND3_X1 U15721 ( .A1(n12627), .A2(n12626), .A3(n12661), .ZN(n12628) );
  NAND4_X1 U15722 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12642) );
  AOI22_X1 U15723 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9970), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15724 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9618), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U15725 ( .A1(n20914), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12634) );
  NAND2_X1 U15726 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12633) );
  AND3_X1 U15727 ( .A1(n12635), .A2(n12634), .A3(n12633), .ZN(n12638) );
  INV_X1 U15728 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U15729 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9583), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12637) );
  NAND4_X1 U15730 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12641) );
  AND2_X1 U15731 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U15732 ( .A1(n12644), .A2(n12643), .ZN(n12645) );
  OAI21_X1 U15733 ( .B1(n12644), .B2(n12643), .A(n12645), .ZN(n15067) );
  NOR2_X1 U15734 ( .A1(n15068), .A2(n15067), .ZN(n15066) );
  INV_X1 U15735 ( .A(n12645), .ZN(n12646) );
  NOR2_X1 U15736 ( .A1(n15066), .A2(n12646), .ZN(n12670) );
  AOI22_X1 U15737 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10001), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15738 ( .A1(n9623), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9583), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15739 ( .A1(n12648), .A2(n12647), .ZN(n12668) );
  INV_X1 U15740 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15741 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12651) );
  AOI21_X1 U15742 ( .B1(n12649), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n12661), .ZN(n12650) );
  OAI211_X1 U15743 ( .C1(n12653), .C2(n12652), .A(n12651), .B(n12650), .ZN(
        n12667) );
  AOI22_X1 U15744 ( .A1(n12654), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9623), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U15745 ( .A1(n9618), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9584), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12656) );
  NAND2_X1 U15746 ( .A1(n12657), .A2(n12656), .ZN(n12666) );
  AOI22_X1 U15747 ( .A1(n10146), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20914), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U15748 ( .A1(n12659), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12663) );
  NAND2_X1 U15749 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12662) );
  NAND4_X1 U15750 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12665) );
  OAI22_X1 U15751 ( .A1(n12668), .A2(n12667), .B1(n12666), .B2(n12665), .ZN(
        n12669) );
  XNOR2_X1 U15752 ( .A(n12670), .B(n12669), .ZN(n14355) );
  INV_X1 U15753 ( .A(n16345), .ZN(n12671) );
  INV_X1 U15754 ( .A(n13782), .ZN(n16342) );
  NAND2_X1 U15755 ( .A1(n12671), .A2(n16342), .ZN(n13185) );
  NAND2_X1 U15756 ( .A1(n13185), .A2(n13784), .ZN(n12672) );
  NAND2_X1 U15757 ( .A1(n12673), .A2(n15123), .ZN(n12675) );
  NAND2_X1 U15758 ( .A1(n13579), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12674) );
  OAI21_X1 U15759 ( .B1(n14355), .B2(n15130), .A(n12676), .ZN(P2_U2857) );
  INV_X2 U15760 ( .A(n18663), .ZN(n17334) );
  NOR2_X1 U15761 ( .A1(n12685), .A2(n12683), .ZN(n12678) );
  INV_X2 U15762 ( .A(n12893), .ZN(n17185) );
  AOI22_X1 U15763 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12682) );
  NOR2_X2 U15764 ( .A1(n18675), .A2(n12683), .ZN(n12904) );
  AOI22_X1 U15765 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12681) );
  INV_X4 U15766 ( .A(n12718), .ZN(n17339) );
  AOI22_X1 U15767 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12680) );
  OR3_X2 U15768 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15834), .A3(
        n18849), .ZN(n12760) );
  AOI22_X1 U15769 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12679) );
  NAND4_X1 U15770 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12695) );
  INV_X4 U15771 ( .A(n17022), .ZN(n17332) );
  AOI22_X1 U15772 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12693) );
  NOR2_X1 U15773 ( .A1(n12683), .A2(n16932), .ZN(n12735) );
  AOI22_X1 U15774 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12692) );
  NOR2_X2 U15775 ( .A1(n18675), .A2(n12687), .ZN(n12686) );
  AOI22_X1 U15776 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15777 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U15778 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12694) );
  AOI22_X1 U15779 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15780 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U15781 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15782 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12696) );
  NAND4_X1 U15783 ( .A1(n12699), .A2(n12698), .A3(n12697), .A4(n12696), .ZN(
        n12705) );
  AOI22_X1 U15784 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15785 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12702) );
  INV_X1 U15786 ( .A(n12882), .ZN(n16973) );
  AOI22_X1 U15787 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15788 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15789 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12704) );
  AOI22_X1 U15790 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15791 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12708) );
  INV_X2 U15792 ( .A(n12848), .ZN(n17146) );
  AOI22_X1 U15793 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12707) );
  INV_X2 U15794 ( .A(n12893), .ZN(n17328) );
  AOI22_X1 U15795 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12706) );
  NAND4_X1 U15796 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12715) );
  AOI22_X1 U15797 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15798 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15799 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15800 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12710) );
  NAND4_X1 U15801 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n12710), .ZN(
        n12714) );
  AOI22_X1 U15802 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12725) );
  INV_X2 U15803 ( .A(n15797), .ZN(n15786) );
  AOI22_X1 U15804 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15805 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12684), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12717) );
  OAI21_X1 U15806 ( .B1(n17022), .B2(n20851), .A(n12717), .ZN(n12723) );
  AOI22_X1 U15807 ( .A1(n12905), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15808 ( .A1(n12686), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12678), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15809 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15810 ( .A1(n12871), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15811 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12726), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15812 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17201), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n12905), .ZN(n12729) );
  AOI22_X1 U15813 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15814 ( .A1(n12871), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15815 ( .A1(n12686), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9596), .ZN(n12734) );
  AOI22_X1 U15816 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17331), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12684), .ZN(n12733) );
  INV_X2 U15817 ( .A(n18663), .ZN(n17058) );
  NAND2_X1 U15818 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12732) );
  AOI22_X1 U15819 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17185), .B1(
        n12735), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12736) );
  OAI21_X1 U15820 ( .B1(n20805), .B2(n17188), .A(n12736), .ZN(n12737) );
  INV_X1 U15821 ( .A(n12737), .ZN(n12738) );
  NAND3_X1 U15822 ( .A1(n9873), .A2(n9876), .A3(n12738), .ZN(n12980) );
  NAND2_X1 U15823 ( .A1(n17421), .A2(n12980), .ZN(n12775) );
  AOI22_X1 U15824 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15825 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15826 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17201), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12739) );
  OAI21_X1 U15827 ( .B1(n12848), .B2(n20867), .A(n12739), .ZN(n12745) );
  AOI22_X1 U15828 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15829 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15830 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15831 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12740) );
  NAND4_X1 U15832 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n12740), .ZN(
        n12744) );
  AOI211_X1 U15833 ( .C1(n17058), .C2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n12745), .B(n12744), .ZN(n12746) );
  NAND3_X1 U15834 ( .A1(n12748), .A2(n12747), .A3(n12746), .ZN(n12968) );
  NAND2_X1 U15835 ( .A1(n12778), .A2(n12968), .ZN(n12780) );
  AOI22_X1 U15836 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15837 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12757) );
  INV_X2 U15838 ( .A(n15797), .ZN(n17218) );
  INV_X1 U15839 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U15840 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12749) );
  OAI21_X1 U15841 ( .B1(n18663), .B2(n17238), .A(n12749), .ZN(n12755) );
  AOI22_X1 U15842 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U15843 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15844 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15845 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U15846 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12754) );
  AOI211_X1 U15847 ( .C1(n17218), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12755), .B(n12754), .ZN(n12756) );
  NAND3_X1 U15848 ( .A1(n12758), .A2(n12757), .A3(n12756), .ZN(n12969) );
  NOR2_X4 U15849 ( .A1(n17402), .A2(n12788), .ZN(n17811) );
  NAND2_X1 U15850 ( .A1(n17432), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12771) );
  AOI22_X1 U15851 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12684), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15852 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12763) );
  INV_X2 U15853 ( .A(n12760), .ZN(n17333) );
  AOI22_X1 U15854 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15855 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12761) );
  NAND4_X1 U15856 ( .A1(n12764), .A2(n12763), .A3(n12762), .A4(n12761), .ZN(
        n12770) );
  AOI22_X1 U15857 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12686), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15858 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15859 ( .A1(n12871), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15860 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U15861 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12769) );
  INV_X1 U15862 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18222) );
  NOR2_X1 U15863 ( .A1(n17900), .A2(n18222), .ZN(n17899) );
  NAND2_X1 U15864 ( .A1(n17891), .A2(n17899), .ZN(n17890) );
  NAND2_X1 U15865 ( .A1(n12771), .A2(n17890), .ZN(n17882) );
  NAND2_X1 U15866 ( .A1(n17883), .A2(n17882), .ZN(n17881) );
  NAND2_X1 U15867 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12772), .ZN(
        n12773) );
  XOR2_X1 U15868 ( .A(n17417), .B(n12775), .Z(n17871) );
  NAND2_X1 U15869 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12776), .ZN(
        n12777) );
  INV_X1 U15870 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18178) );
  INV_X1 U15871 ( .A(n12968), .ZN(n17413) );
  XNOR2_X1 U15872 ( .A(n17413), .B(n12778), .ZN(n12779) );
  XNOR2_X1 U15873 ( .A(n18178), .B(n12779), .ZN(n17862) );
  XOR2_X1 U15874 ( .A(n17409), .B(n12780), .Z(n12783) );
  NAND2_X1 U15875 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17848), .ZN(
        n17847) );
  NAND2_X1 U15876 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  NAND2_X1 U15877 ( .A1(n17847), .A2(n12784), .ZN(n17833) );
  INV_X1 U15878 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18129) );
  INV_X1 U15879 ( .A(n12969), .ZN(n17406) );
  XNOR2_X1 U15880 ( .A(n17406), .B(n12785), .ZN(n12786) );
  XNOR2_X1 U15881 ( .A(n18129), .B(n12786), .ZN(n17834) );
  NAND2_X1 U15882 ( .A1(n17833), .A2(n17834), .ZN(n17832) );
  NAND2_X1 U15883 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12786), .ZN(
        n12787) );
  NAND2_X1 U15884 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  INV_X1 U15885 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18122) );
  INV_X1 U15886 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18108) );
  NAND2_X1 U15887 ( .A1(n17762), .A2(n18108), .ZN(n17755) );
  INV_X1 U15888 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17734) );
  NAND2_X1 U15889 ( .A1(n17731), .A2(n17734), .ZN(n17705) );
  INV_X1 U15890 ( .A(n17705), .ZN(n12794) );
  INV_X1 U15891 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18060) );
  INV_X1 U15892 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18058) );
  NAND2_X1 U15893 ( .A1(n18060), .A2(n18058), .ZN(n12795) );
  INV_X1 U15894 ( .A(n12807), .ZN(n12799) );
  NAND2_X1 U15895 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18107) );
  NOR2_X1 U15896 ( .A1(n18107), .A2(n18108), .ZN(n17758) );
  NAND3_X1 U15897 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17706) );
  OR2_X1 U15898 ( .A1(n12793), .A2(n17706), .ZN(n18059) );
  NOR2_X1 U15899 ( .A1(n18058), .A2(n18059), .ZN(n18013) );
  INV_X1 U15900 ( .A(n18013), .ZN(n16412) );
  NAND2_X2 U15901 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12796), .ZN(
        n18096) );
  NOR2_X2 U15902 ( .A1(n16410), .A2(n12797), .ZN(n18143) );
  INV_X1 U15903 ( .A(n12797), .ZN(n12798) );
  INV_X1 U15904 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17958) );
  NAND2_X1 U15905 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17631) );
  INV_X1 U15906 ( .A(n17631), .ZN(n18022) );
  INV_X1 U15907 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17671) );
  INV_X1 U15908 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17986) );
  INV_X1 U15909 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18006) );
  INV_X1 U15910 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17968) );
  NOR2_X1 U15911 ( .A1(n18006), .A2(n17968), .ZN(n17963) );
  INV_X1 U15912 ( .A(n17963), .ZN(n17985) );
  NOR3_X1 U15913 ( .A1(n17671), .A2(n17986), .A3(n17985), .ZN(n12811) );
  AND2_X1 U15914 ( .A1(n18022), .A2(n12811), .ZN(n17970) );
  NAND2_X1 U15915 ( .A1(n17970), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16413) );
  NOR2_X1 U15916 ( .A1(n17958), .A2(n16413), .ZN(n12997) );
  INV_X1 U15917 ( .A(n12997), .ZN(n12802) );
  NAND2_X1 U15918 ( .A1(n17671), .A2(n12810), .ZN(n17670) );
  NOR2_X1 U15919 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17670), .ZN(
        n12800) );
  NAND2_X1 U15920 ( .A1(n12800), .A2(n17968), .ZN(n17637) );
  INV_X1 U15921 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17973) );
  NAND3_X1 U15922 ( .A1(n17627), .A2(n17958), .A3(n17973), .ZN(n12801) );
  OAI21_X1 U15923 ( .B1(n17689), .B2(n12802), .A(n12801), .ZN(n12803) );
  INV_X1 U15924 ( .A(n12803), .ZN(n12808) );
  INV_X1 U15925 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17703) );
  INV_X1 U15926 ( .A(n12805), .ZN(n12806) );
  INV_X1 U15927 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17603) );
  INV_X1 U15928 ( .A(n17598), .ZN(n17590) );
  INV_X1 U15929 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17930) );
  NOR2_X2 U15930 ( .A1(n17605), .A2(n17636), .ZN(n17672) );
  NAND2_X1 U15931 ( .A1(n12811), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13001) );
  NAND3_X1 U15932 ( .A1(n17604), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17598), .ZN(n12814) );
  NAND2_X1 U15933 ( .A1(n12814), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12812) );
  INV_X1 U15934 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20800) );
  NAND2_X1 U15935 ( .A1(n17811), .A2(n12814), .ZN(n17589) );
  NOR2_X1 U15936 ( .A1(n20800), .A2(n17930), .ZN(n17912) );
  INV_X1 U15937 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16415) );
  INV_X1 U15938 ( .A(n16426), .ZN(n17564) );
  NOR2_X1 U15939 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17811), .ZN(
        n16416) );
  NAND2_X1 U15940 ( .A1(n17564), .A2(n16416), .ZN(n15839) );
  NOR2_X2 U15941 ( .A1(n15839), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15889) );
  NOR2_X1 U15942 ( .A1(n17811), .A2(n15889), .ZN(n12822) );
  INV_X1 U15943 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15893) );
  INV_X1 U15944 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16396) );
  INV_X1 U15945 ( .A(n15890), .ZN(n12817) );
  OAI21_X1 U15946 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15893), .A(
        n12817), .ZN(n12818) );
  NAND2_X1 U15947 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17811), .ZN(
        n12820) );
  OAI22_X1 U15948 ( .A1(n12822), .A2(n12818), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12820), .ZN(n12819) );
  INV_X1 U15949 ( .A(n12819), .ZN(n12827) );
  OAI21_X1 U15950 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17811), .A(
        n12820), .ZN(n12821) );
  INV_X1 U15951 ( .A(n12821), .ZN(n12826) );
  OAI22_X1 U15952 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15890), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12822), .ZN(n12823) );
  INV_X1 U15953 ( .A(n12823), .ZN(n12824) );
  NAND2_X1 U15954 ( .A1(n12824), .A2(n12826), .ZN(n12825) );
  OAI21_X1 U15955 ( .B1(n12827), .B2(n12826), .A(n12825), .ZN(n13014) );
  AOI22_X1 U15956 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U15957 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U15958 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U15959 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12828) );
  NAND4_X1 U15960 ( .A1(n12831), .A2(n12830), .A3(n12829), .A4(n12828), .ZN(
        n12837) );
  INV_X2 U15961 ( .A(n12870), .ZN(n17219) );
  AOI22_X1 U15962 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15963 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15964 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12726), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15965 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U15966 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  AOI22_X1 U15967 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15968 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12905), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15969 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12838) );
  OAI21_X1 U15970 ( .B1(n12760), .B2(n20851), .A(n12838), .ZN(n12844) );
  AOI22_X1 U15971 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15972 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U15973 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U15974 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12839) );
  NAND4_X1 U15975 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n12843) );
  AOI211_X1 U15976 ( .C1(n17340), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n12844), .B(n12843), .ZN(n12845) );
  NAND3_X1 U15977 ( .A1(n12847), .A2(n12846), .A3(n12845), .ZN(n18251) );
  NOR2_X1 U15978 ( .A1(n18877), .A2(n18251), .ZN(n12954) );
  AOI22_X1 U15979 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15980 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12857) );
  INV_X1 U15981 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17251) );
  INV_X2 U15982 ( .A(n12848), .ZN(n17342) );
  AOI22_X1 U15983 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12849) );
  OAI21_X1 U15984 ( .B1(n15808), .B2(n17251), .A(n12849), .ZN(n12855) );
  AOI22_X1 U15985 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U15986 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15987 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15988 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12850) );
  NAND4_X1 U15989 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12854) );
  AOI211_X1 U15990 ( .C1(n16971), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n12855), .B(n12854), .ZN(n12856) );
  NAND3_X1 U15991 ( .A1(n12858), .A2(n12857), .A3(n12856), .ZN(n18255) );
  INV_X1 U15992 ( .A(n18255), .ZN(n12923) );
  AOI22_X1 U15993 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U15994 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U15995 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U15996 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17201), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12859) );
  NAND4_X1 U15997 ( .A1(n12862), .A2(n12861), .A3(n12860), .A4(n12859), .ZN(
        n12868) );
  AOI22_X1 U15998 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U15999 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16000 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16001 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12863) );
  NAND4_X1 U16002 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  AOI22_X1 U16003 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U16004 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16005 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U16006 ( .B1(n12870), .B2(n20794), .A(n12869), .ZN(n12877) );
  AOI22_X1 U16007 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U16008 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U16009 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U16010 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12872) );
  NAND4_X1 U16011 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12872), .ZN(
        n12876) );
  INV_X1 U16012 ( .A(n12932), .ZN(n12915) );
  AOI22_X1 U16013 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16014 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16015 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17201), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12881) );
  OAI21_X1 U16016 ( .B1(n12882), .B2(n20867), .A(n12881), .ZN(n12888) );
  AOI22_X1 U16017 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U16018 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U16019 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U16020 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12883) );
  NAND4_X1 U16021 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12887) );
  AOI211_X1 U16022 ( .C1(n17332), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n12888), .B(n12887), .ZN(n12889) );
  NAND3_X1 U16023 ( .A1(n12891), .A2(n12890), .A3(n12889), .ZN(n18260) );
  AOI22_X1 U16024 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16025 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12901) );
  INV_X1 U16026 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U16027 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12892) );
  OAI21_X1 U16028 ( .B1(n12893), .B2(n20791), .A(n12892), .ZN(n12899) );
  AOI22_X1 U16029 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U16030 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16031 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16032 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12894) );
  NAND4_X1 U16033 ( .A1(n12897), .A2(n12896), .A3(n12895), .A4(n12894), .ZN(
        n12898) );
  AOI22_X1 U16034 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16035 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17218), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U16036 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12903) );
  OAI21_X1 U16037 ( .B1(n15808), .B2(n17238), .A(n12903), .ZN(n12911) );
  AOI22_X1 U16038 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U16039 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16040 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12905), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16041 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12906) );
  NAND4_X1 U16042 ( .A1(n12909), .A2(n12908), .A3(n12907), .A4(n12906), .ZN(
        n12910) );
  AOI211_X1 U16043 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12911), .B(n12910), .ZN(n12912) );
  NAND3_X1 U16044 ( .A1(n12914), .A2(n12913), .A3(n12912), .ZN(n18269) );
  NAND2_X1 U16045 ( .A1(n18264), .A2(n18269), .ZN(n12963) );
  NOR2_X1 U16046 ( .A1(n18260), .A2(n12963), .ZN(n12918) );
  NOR2_X1 U16047 ( .A1(n18269), .A2(n18260), .ZN(n12921) );
  NAND2_X1 U16048 ( .A1(n12966), .A2(n17433), .ZN(n12917) );
  INV_X1 U16049 ( .A(n12963), .ZN(n12916) );
  NOR2_X1 U16050 ( .A1(n12927), .A2(n12916), .ZN(n12919) );
  AOI22_X1 U16051 ( .A1(n12966), .A2(n12919), .B1(n12918), .B2(n12917), .ZN(
        n12920) );
  AOI21_X1 U16052 ( .B1(n12921), .B2(n12922), .A(n12920), .ZN(n12949) );
  NAND2_X1 U16053 ( .A1(n12949), .A2(n18274), .ZN(n12930) );
  OAI211_X1 U16054 ( .C1(n12921), .C2(n18264), .A(n12966), .B(n18255), .ZN(
        n12931) );
  INV_X1 U16055 ( .A(n18269), .ZN(n12928) );
  NAND2_X1 U16056 ( .A1(n12966), .A2(n12923), .ZN(n18661) );
  NOR3_X1 U16057 ( .A1(n12928), .A2(n18264), .A3(n18661), .ZN(n15739) );
  NAND3_X1 U16058 ( .A1(n18877), .A2(n12924), .A3(n15739), .ZN(n12925) );
  NAND2_X1 U16059 ( .A1(n12928), .A2(n18260), .ZN(n18662) );
  NOR2_X1 U16060 ( .A1(n17433), .A2(n18248), .ZN(n12929) );
  NOR2_X1 U16061 ( .A1(n12927), .A2(n12929), .ZN(n18888) );
  NAND2_X1 U16062 ( .A1(n12928), .A2(n18264), .ZN(n18694) );
  INV_X1 U16063 ( .A(n18694), .ZN(n15909) );
  AOI211_X1 U16064 ( .C1(n12932), .C2(n12931), .A(n12951), .B(n12930), .ZN(
        n18660) );
  INV_X1 U16065 ( .A(n18260), .ZN(n15738) );
  AOI22_X1 U16066 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20892), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18849), .ZN(n12957) );
  OAI22_X1 U16067 ( .A1(n9714), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18240), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12940) );
  INV_X1 U16068 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18706) );
  OAI22_X1 U16069 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18706), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12937), .ZN(n12944) );
  NOR2_X1 U16070 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18706), .ZN(
        n12938) );
  NAND2_X1 U16071 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12937), .ZN(
        n12943) );
  AOI22_X1 U16072 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12944), .B1(
        n12938), .B2(n12943), .ZN(n12946) );
  NAND2_X1 U16073 ( .A1(n12941), .A2(n12940), .ZN(n12939) );
  OAI211_X1 U16074 ( .C1(n12941), .C2(n12940), .A(n12946), .B(n12939), .ZN(
        n12942) );
  INV_X1 U16075 ( .A(n12942), .ZN(n12962) );
  INV_X1 U16076 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18716) );
  AND2_X1 U16077 ( .A1(n12943), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12945) );
  OAI22_X1 U16078 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18716), .B1(
        n12945), .B2(n12944), .ZN(n12958) );
  NOR2_X1 U16079 ( .A1(n12962), .A2(n12958), .ZN(n12948) );
  AOI21_X1 U16080 ( .B1(n12933), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12956), .ZN(n12961) );
  NAND3_X1 U16081 ( .A1(n12957), .A2(n12946), .A3(n12961), .ZN(n12947) );
  NAND2_X1 U16082 ( .A1(n12950), .A2(n12949), .ZN(n12953) );
  AOI21_X1 U16083 ( .B1(n12953), .B2(n12952), .A(n12951), .ZN(n15829) );
  NAND2_X1 U16084 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18878) );
  INV_X1 U16085 ( .A(n18878), .ZN(n18750) );
  NAND2_X1 U16086 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18741), .ZN(n18885) );
  INV_X2 U16087 ( .A(n18885), .ZN(n18822) );
  NAND2_X1 U16088 ( .A1(n18822), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18816) );
  NOR2_X1 U16089 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16541) );
  INV_X1 U16090 ( .A(n16541), .ZN(n18740) );
  NAND3_X1 U16091 ( .A1(n18741), .A2(n18810), .A3(n18740), .ZN(n18875) );
  INV_X1 U16092 ( .A(n18875), .ZN(n16564) );
  AOI211_X1 U16093 ( .C1(n18877), .C2(n18251), .A(n12954), .B(n16564), .ZN(
        n12955) );
  NOR2_X1 U16094 ( .A1(n18750), .A2(n12955), .ZN(n16543) );
  XOR2_X1 U16095 ( .A(n12957), .B(n12956), .Z(n12959) );
  OAI211_X1 U16096 ( .C1(n17272), .C2(n18251), .A(n16543), .B(n18682), .ZN(
        n12960) );
  OAI211_X1 U16097 ( .C1(n15738), .C2(n18688), .A(n15829), .B(n12960), .ZN(
        n12967) );
  INV_X1 U16098 ( .A(n18682), .ZN(n15824) );
  AOI21_X1 U16099 ( .B1(n12962), .B2(n12961), .A(n15824), .ZN(n18685) );
  INV_X1 U16100 ( .A(n18685), .ZN(n13013) );
  NAND2_X1 U16101 ( .A1(n18248), .A2(n18269), .ZN(n12964) );
  OAI22_X1 U16102 ( .A1(n13013), .A2(n12964), .B1(n12963), .B2(n18688), .ZN(
        n12965) );
  INV_X1 U16103 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n16561) );
  NOR2_X1 U16104 ( .A1(n16561), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18731) );
  NAND2_X1 U16105 ( .A1(n18731), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18725) );
  NOR3_X4 U16106 ( .A1(n17402), .A2(n18684), .A3(n18182), .ZN(n18141) );
  NAND2_X1 U16107 ( .A1(n13014), .A2(n18141), .ZN(n13012) );
  NAND2_X1 U16108 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18086) );
  NOR2_X1 U16109 ( .A1(n12976), .A2(n17421), .ZN(n12974) );
  NOR2_X1 U16110 ( .A1(n12974), .A2(n17417), .ZN(n12972) );
  NAND2_X1 U16111 ( .A1(n12972), .A2(n12968), .ZN(n12985) );
  NOR2_X1 U16112 ( .A1(n17409), .A2(n12985), .ZN(n12971) );
  NAND2_X1 U16113 ( .A1(n12971), .A2(n12969), .ZN(n12970) );
  NOR2_X1 U16114 ( .A1(n17402), .A2(n12970), .ZN(n12994) );
  INV_X1 U16115 ( .A(n17402), .ZN(n16419) );
  XNOR2_X1 U16116 ( .A(n12970), .B(n16419), .ZN(n17825) );
  XNOR2_X1 U16117 ( .A(n12971), .B(n17406), .ZN(n12987) );
  XNOR2_X1 U16118 ( .A(n12972), .B(n17413), .ZN(n12973) );
  NAND2_X1 U16119 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12973), .ZN(
        n12983) );
  XNOR2_X1 U16120 ( .A(n18178), .B(n12973), .ZN(n17856) );
  XOR2_X1 U16121 ( .A(n17417), .B(n12974), .Z(n12975) );
  NAND2_X1 U16122 ( .A1(n12975), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12982) );
  XNOR2_X1 U16123 ( .A(n12774), .B(n12975), .ZN(n17869) );
  XNOR2_X1 U16124 ( .A(n17421), .B(n12976), .ZN(n12977) );
  NAND2_X1 U16125 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12977), .ZN(
        n12981) );
  XOR2_X1 U16126 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12977), .Z(
        n17880) );
  INV_X1 U16127 ( .A(n17900), .ZN(n15910) );
  AOI21_X1 U16128 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12980), .A(
        n15910), .ZN(n12979) );
  NOR2_X1 U16129 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12980), .ZN(
        n12978) );
  AOI221_X1 U16130 ( .B1(n15910), .B2(n12980), .C1(n12979), .C2(n18222), .A(
        n12978), .ZN(n17879) );
  NAND2_X1 U16131 ( .A1(n17880), .A2(n17879), .ZN(n17878) );
  NAND2_X1 U16132 ( .A1(n12981), .A2(n17878), .ZN(n17868) );
  NAND2_X1 U16133 ( .A1(n17869), .A2(n17868), .ZN(n17867) );
  NAND2_X1 U16134 ( .A1(n12982), .A2(n17867), .ZN(n17855) );
  NAND2_X1 U16135 ( .A1(n17856), .A2(n17855), .ZN(n17854) );
  NAND2_X1 U16136 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12984), .ZN(
        n12986) );
  XOR2_X1 U16137 ( .A(n12985), .B(n17409), .Z(n17842) );
  NAND2_X1 U16138 ( .A1(n17843), .A2(n17842), .ZN(n17841) );
  NAND2_X1 U16139 ( .A1(n12986), .A2(n17841), .ZN(n12988) );
  NAND2_X1 U16140 ( .A1(n12987), .A2(n12988), .ZN(n12989) );
  INV_X1 U16141 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18130) );
  NAND2_X1 U16142 ( .A1(n12994), .A2(n12990), .ZN(n12995) );
  INV_X1 U16143 ( .A(n12990), .ZN(n12993) );
  NAND2_X1 U16144 ( .A1(n17825), .A2(n17824), .ZN(n12992) );
  NAND2_X1 U16145 ( .A1(n12994), .A2(n12993), .ZN(n12991) );
  NAND2_X1 U16146 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17801), .ZN(
        n17800) );
  NOR2_X2 U16147 ( .A1(n17941), .A2(n17603), .ZN(n17588) );
  INV_X1 U16148 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16425) );
  NOR2_X1 U16149 ( .A1(n16415), .A2(n16425), .ZN(n16393) );
  NAND2_X1 U16150 ( .A1(n16393), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15892) );
  NAND2_X1 U16151 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n9602), .ZN(
        n12996) );
  XNOR2_X1 U16152 ( .A(n12996), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13026) );
  NOR2_X1 U16153 ( .A1(n18201), .A2(n18182), .ZN(n18225) );
  NAND2_X1 U16154 ( .A1(n12997), .A2(n18045), .ZN(n17940) );
  NAND2_X1 U16155 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16394), .ZN(
        n12998) );
  XOR2_X1 U16156 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12998), .Z(
        n13024) );
  NOR2_X1 U16157 ( .A1(n18684), .A2(n18182), .ZN(n18227) );
  NAND2_X1 U16158 ( .A1(n17402), .A2(n18227), .ZN(n18139) );
  INV_X1 U16159 ( .A(n18135), .ZN(n17972) );
  NAND2_X1 U16160 ( .A1(n18218), .A2(n17972), .ZN(n18173) );
  NOR2_X1 U16161 ( .A1(n17958), .A2(n17603), .ZN(n17907) );
  NAND2_X1 U16162 ( .A1(n17912), .A2(n17907), .ZN(n16414) );
  INV_X1 U16163 ( .A(n16413), .ZN(n17955) );
  NOR3_X1 U16164 ( .A1(n18130), .A2(n18129), .A3(n9811), .ZN(n18011) );
  NAND3_X1 U16165 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18010) );
  NAND2_X1 U16166 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18008) );
  NOR2_X1 U16167 ( .A1(n18010), .A2(n18008), .ZN(n18131) );
  NAND2_X1 U16168 ( .A1(n18011), .A2(n18131), .ZN(n12999) );
  NOR2_X1 U16169 ( .A1(n16412), .A2(n12999), .ZN(n18017) );
  NAND2_X1 U16170 ( .A1(n17955), .A2(n18017), .ZN(n17906) );
  NOR2_X1 U16171 ( .A1(n16414), .A2(n17906), .ZN(n13003) );
  INV_X1 U16172 ( .A(n16414), .ZN(n17914) );
  INV_X1 U16173 ( .A(n12999), .ZN(n18099) );
  NAND2_X1 U16174 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18099), .ZN(
        n18101) );
  NOR2_X1 U16175 ( .A1(n16412), .A2(n18101), .ZN(n18033) );
  NAND3_X1 U16176 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17914), .A3(
        n18033), .ZN(n13000) );
  OAI21_X1 U16177 ( .B1(n16413), .B2(n13000), .A(n18668), .ZN(n13002) );
  AOI21_X1 U16178 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18198) );
  NOR2_X1 U16179 ( .A1(n18198), .A2(n18010), .ZN(n18132) );
  NAND2_X1 U16180 ( .A1(n18132), .A2(n18011), .ZN(n18034) );
  NOR2_X1 U16181 ( .A1(n16412), .A2(n18034), .ZN(n17926) );
  NAND2_X1 U16182 ( .A1(n18022), .A2(n17926), .ZN(n18020) );
  NOR2_X1 U16183 ( .A1(n13001), .A2(n18020), .ZN(n17944) );
  NAND2_X1 U16184 ( .A1(n17944), .A2(n17914), .ZN(n13005) );
  NAND2_X1 U16185 ( .A1(n18689), .A2(n13005), .ZN(n17910) );
  OAI211_X1 U16186 ( .C1(n18100), .C2(n13003), .A(n13002), .B(n17910), .ZN(
        n15842) );
  INV_X1 U16187 ( .A(n18173), .ZN(n18210) );
  AOI22_X1 U16188 ( .A1(n18218), .A2(n15842), .B1(n18210), .B2(n15892), .ZN(
        n15895) );
  INV_X1 U16189 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18853) );
  NAND2_X1 U16190 ( .A1(n18853), .A2(n18830), .ZN(n18852) );
  NOR2_X1 U16191 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18852), .ZN(n18887) );
  AND2_X2 U16192 ( .A1(n18887), .A2(n16561), .ZN(n18209) );
  INV_X2 U16193 ( .A(n18209), .ZN(n18175) );
  OAI211_X1 U16194 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18173), .A(
        n15895), .B(n18221), .ZN(n13008) );
  INV_X1 U16195 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18813) );
  NOR2_X1 U16196 ( .A1(n18813), .A2(n18175), .ZN(n13022) );
  INV_X1 U16197 ( .A(n13003), .ZN(n13004) );
  INV_X1 U16198 ( .A(n18100), .ZN(n18699) );
  AOI21_X1 U16199 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18668), .A(
        n18699), .ZN(n18194) );
  OAI22_X1 U16200 ( .A1(n18670), .A2(n13005), .B1(n13004), .B2(n18194), .ZN(
        n13006) );
  NAND2_X1 U16201 ( .A1(n18218), .A2(n13006), .ZN(n15847) );
  NOR4_X1 U16202 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15892), .A3(
        n15893), .A4(n15847), .ZN(n13007) );
  AOI211_X1 U16203 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13008), .A(
        n13022), .B(n13007), .ZN(n13009) );
  NAND2_X1 U16204 ( .A1(n13012), .A2(n13011), .ZN(P3_U2831) );
  NAND2_X1 U16205 ( .A1(n13014), .A2(n17812), .ZN(n13028) );
  NOR2_X2 U16206 ( .A1(n18248), .A2(n16544), .ZN(n17893) );
  NAND2_X1 U16207 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17858) );
  NAND2_X1 U16208 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18229) );
  NAND2_X1 U16209 ( .A1(n18830), .A2(n18229), .ZN(n18872) );
  INV_X1 U16210 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20809) );
  INV_X1 U16211 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17680) );
  INV_X1 U16212 ( .A(n16883), .ZN(n17859) );
  NAND2_X1 U16213 ( .A1(n17859), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17845) );
  NAND2_X1 U16214 ( .A1(n17819), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17804) );
  NAND3_X1 U16215 ( .A1(n17802), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16798) );
  NOR2_X2 U16216 ( .A1(n17804), .A2(n16798), .ZN(n17775) );
  NAND2_X1 U16217 ( .A1(n17775), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17720) );
  INV_X1 U16218 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17750) );
  NAND2_X1 U16219 ( .A1(n17736), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17695) );
  NAND3_X1 U16220 ( .A1(n17691), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17681) );
  NOR2_X2 U16221 ( .A1(n17680), .A2(n17681), .ZN(n17665) );
  NAND3_X1 U16222 ( .A1(n17665), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17643) );
  NOR2_X2 U16223 ( .A1(n20809), .A2(n17643), .ZN(n17619) );
  NAND3_X1 U16224 ( .A1(n17619), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17610) );
  INV_X1 U16225 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17609) );
  NOR2_X2 U16226 ( .A1(n17610), .A2(n17609), .ZN(n17583) );
  NAND2_X1 U16227 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17584) );
  NAND2_X1 U16228 ( .A1(n17548), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16574) );
  INV_X1 U16229 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17546) );
  INV_X1 U16230 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16610) );
  NOR2_X2 U16231 ( .A1(n16572), .A2(n16610), .ZN(n16397) );
  NAND2_X1 U16232 ( .A1(n16397), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13016) );
  XOR2_X2 U16233 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13016), .Z(
        n16874) );
  INV_X1 U16234 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17573) );
  NAND3_X1 U16235 ( .A1(n17583), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17572) );
  NOR2_X1 U16236 ( .A1(n17573), .A2(n17572), .ZN(n17547) );
  NAND3_X1 U16237 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n17547), .ZN(n16392) );
  NOR2_X1 U16238 ( .A1(n16610), .A2(n16392), .ZN(n13017) );
  INV_X1 U16239 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17894) );
  INV_X1 U16240 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16562) );
  NOR2_X1 U16241 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n16562), .ZN(n13097) );
  NOR2_X1 U16242 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18830), .ZN(
        n18847) );
  NOR2_X1 U16243 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18880) );
  AOI21_X1 U16244 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18880), .ZN(n18735) );
  NOR2_X1 U16245 ( .A1(n18847), .A2(n18735), .ZN(n18238) );
  INV_X1 U16246 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18876) );
  NOR3_X1 U16247 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18876), .ZN(n18243) );
  NAND2_X1 U16248 ( .A1(n18579), .A2(n18243), .ZN(n18278) );
  NAND2_X1 U16249 ( .A1(n13017), .A2(n17694), .ZN(n16385) );
  INV_X1 U16250 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16583) );
  XOR2_X1 U16251 ( .A(n16583), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13020) );
  NOR2_X1 U16252 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17678), .ZN(
        n16398) );
  INV_X1 U16253 ( .A(n13017), .ZN(n13018) );
  AOI22_X1 U16254 ( .A1(n18607), .A2(n13018), .B1(n13097), .B2(n16572), .ZN(
        n13019) );
  NAND2_X1 U16255 ( .A1(n13019), .A2(n17901), .ZN(n16403) );
  NOR2_X1 U16256 ( .A1(n16398), .A2(n16403), .ZN(n16383) );
  OAI22_X1 U16257 ( .A1(n16385), .A2(n13020), .B1(n16383), .B2(n16583), .ZN(
        n13021) );
  AOI211_X1 U16258 ( .C1(n17754), .C2(n16903), .A(n13022), .B(n13021), .ZN(
        n13023) );
  NAND2_X1 U16259 ( .A1(n13028), .A2(n13027), .ZN(P3_U2799) );
  NOR4_X1 U16260 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13032) );
  NOR4_X1 U16261 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13031) );
  NOR4_X1 U16262 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13030) );
  NOR4_X1 U16263 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13029) );
  AND4_X1 U16264 ( .A1(n13032), .A2(n13031), .A3(n13030), .A4(n13029), .ZN(
        n13037) );
  NOR4_X1 U16265 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13035) );
  NOR4_X1 U16266 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13034) );
  NOR4_X1 U16267 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13033) );
  INV_X1 U16268 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20657) );
  AND4_X1 U16269 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n20657), .ZN(
        n13036) );
  NAND2_X1 U16270 ( .A1(n13037), .A2(n13036), .ZN(n13038) );
  AND2_X2 U16271 ( .A1(n13038), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20032)
         );
  INV_X1 U16272 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20738) );
  NOR3_X1 U16273 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20738), .ZN(n13040) );
  NOR4_X1 U16274 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13039) );
  NAND4_X1 U16275 ( .A1(n20032), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13040), .A4(
        n13039), .ZN(U214) );
  NOR4_X1 U16276 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13044) );
  NOR4_X1 U16277 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n13043) );
  NOR4_X1 U16278 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13042) );
  NOR4_X1 U16279 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13041) );
  NAND4_X1 U16280 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13049) );
  NOR4_X1 U16281 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n13047) );
  NOR4_X1 U16282 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n13046) );
  NOR4_X1 U16283 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13045) );
  INV_X1 U16284 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19745) );
  NAND4_X1 U16285 ( .A1(n13047), .A2(n13046), .A3(n13045), .A4(n19745), .ZN(
        n13048) );
  OAI21_X1 U16286 ( .B1(n13049), .B2(n13048), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13050) );
  NOR2_X1 U16287 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13052) );
  NOR4_X1 U16288 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13051) );
  NAND4_X1 U16289 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13052), .A4(n13051), .ZN(n13053) );
  NOR2_X1 U16290 ( .A1(n15696), .A2(n13053), .ZN(n16433) );
  NAND2_X1 U16291 ( .A1(n16433), .A2(U214), .ZN(U212) );
  NOR2_X1 U16292 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13053), .ZN(n16521)
         );
  AOI211_X1 U16293 ( .C1(n14192), .C2(n13055), .A(n13054), .B(n19724), .ZN(
        n13066) );
  INV_X1 U16294 ( .A(n19036), .ZN(n19060) );
  OAI22_X1 U16295 ( .A1(n19765), .A2(n19030), .B1(n14189), .B2(n19060), .ZN(
        n13065) );
  INV_X1 U16296 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n13056) );
  INV_X1 U16297 ( .A(n19049), .ZN(n19032) );
  OAI22_X1 U16298 ( .A1(n13057), .A2(n19052), .B1(n13056), .B2(n19032), .ZN(
        n13064) );
  OAI21_X1 U16299 ( .B1(n13058), .B2(n13059), .A(n15036), .ZN(n14203) );
  NOR2_X1 U16300 ( .A1(n14239), .A2(n13061), .ZN(n13062) );
  OR2_X1 U16301 ( .A1(n13060), .A2(n13062), .ZN(n14198) );
  OAI22_X1 U16302 ( .A1(n14203), .A2(n19057), .B1(n14198), .B2(n19046), .ZN(
        n13063) );
  OR4_X1 U16303 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        P2_U2834) );
  AOI211_X1 U16304 ( .C1(n15260), .C2(n13068), .A(n13067), .B(n19724), .ZN(
        n13080) );
  INV_X1 U16305 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19768) );
  OAI22_X1 U16306 ( .A1(n15262), .A2(n19060), .B1(n19768), .B2(n19030), .ZN(
        n13079) );
  INV_X1 U16307 ( .A(n13069), .ZN(n13070) );
  OAI22_X1 U16308 ( .A1(n13070), .A2(n19052), .B1(n19032), .B2(n10830), .ZN(
        n13078) );
  AND2_X1 U16309 ( .A1(n15038), .A2(n13071), .ZN(n13072) );
  NOR2_X1 U16310 ( .A1(n15020), .A2(n13072), .ZN(n15451) );
  INV_X1 U16311 ( .A(n15451), .ZN(n13076) );
  NAND2_X1 U16312 ( .A1(n13073), .A2(n13074), .ZN(n13075) );
  NAND2_X1 U16313 ( .A1(n15023), .A2(n13075), .ZN(n15447) );
  OAI22_X1 U16314 ( .A1(n13076), .A2(n19057), .B1(n19046), .B2(n15447), .ZN(
        n13077) );
  OR4_X1 U16315 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        P2_U2832) );
  NAND2_X1 U16316 ( .A1(n19042), .A2(n12347), .ZN(n13082) );
  AOI211_X1 U16317 ( .C1(n13084), .C2(n13083), .A(n13955), .B(n13082), .ZN(
        n13096) );
  INV_X1 U16318 ( .A(n13084), .ZN(n15338) );
  NAND2_X1 U16319 ( .A1(n19042), .A2(n12329), .ZN(n18942) );
  AOI22_X1 U16320 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19036), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19048), .ZN(n13085) );
  OAI211_X1 U16321 ( .C1(n15338), .C2(n18942), .A(n13085), .B(n10856), .ZN(
        n13095) );
  INV_X1 U16322 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13660) );
  OAI22_X1 U16323 ( .A1(n13086), .A2(n19052), .B1(n19032), .B2(n13660), .ZN(
        n13094) );
  AOI21_X1 U16324 ( .B1(n13088), .B2(n13599), .A(n13087), .ZN(n15528) );
  INV_X1 U16325 ( .A(n15528), .ZN(n13092) );
  OAI21_X1 U16326 ( .B1(n13091), .B2(n13090), .A(n13089), .ZN(n19086) );
  OAI22_X1 U16327 ( .A1(n13092), .A2(n19057), .B1(n19046), .B2(n19086), .ZN(
        n13093) );
  OR4_X1 U16328 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        P2_U2842) );
  INV_X1 U16329 ( .A(n13097), .ZN(n18739) );
  OR2_X1 U16330 ( .A1(n18853), .A2(n18739), .ZN(n17457) );
  NAND2_X1 U16331 ( .A1(n18873), .A2(n18682), .ZN(n17493) );
  INV_X1 U16332 ( .A(n17493), .ZN(n17492) );
  OAI21_X1 U16333 ( .B1(n17494), .B2(n18248), .A(n16560), .ZN(n13098) );
  AND2_X1 U16334 ( .A1(n17488), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U16335 ( .A(n13099), .ZN(n13100) );
  NOR2_X1 U16336 ( .A1(n10511), .A2(n13100), .ZN(n19064) );
  INV_X1 U16337 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19866) );
  INV_X1 U16338 ( .A(n13101), .ZN(n13102) );
  NOR2_X1 U16339 ( .A1(n13112), .A2(n13102), .ZN(n13106) );
  OAI21_X1 U16340 ( .B1(n19064), .B2(n19866), .A(n13106), .ZN(P2_U2814) );
  INV_X1 U16341 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18896) );
  INV_X1 U16342 ( .A(n19800), .ZN(n19795) );
  OAI22_X1 U16343 ( .A1(n19858), .A2(n18896), .B1(n13103), .B2(n19795), .ZN(
        P2_U2816) );
  NOR2_X1 U16344 ( .A1(n19064), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13105)
         );
  AOI22_X1 U16345 ( .A1(n13106), .A2(n13105), .B1(n13104), .B2(n19858), .ZN(
        P2_U3612) );
  NAND2_X1 U16346 ( .A1(n16341), .A2(n16340), .ZN(n13181) );
  NAND2_X1 U16347 ( .A1(n13107), .A2(n19861), .ZN(n13180) );
  INV_X1 U16348 ( .A(n13180), .ZN(n13109) );
  NOR3_X1 U16349 ( .A1(n13181), .A2(n13109), .A3(n13108), .ZN(n16335) );
  INV_X1 U16350 ( .A(n19721), .ZN(n13188) );
  NOR2_X1 U16351 ( .A1(n16335), .A2(n13188), .ZN(n19836) );
  OAI21_X1 U16352 ( .B1(n13111), .B2(n19836), .A(n13110), .ZN(P2_U2819) );
  OAI21_X1 U16353 ( .B1(n10566), .B2(n19861), .A(n13112), .ZN(n13138) );
  INV_X1 U16354 ( .A(n13138), .ZN(n13141) );
  AOI22_X1 U16355 ( .A1(n13161), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13138), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13113) );
  NAND3_X1 U16356 ( .A1(n13112), .A2(n19861), .A3(n19849), .ZN(n13156) );
  INV_X1 U16357 ( .A(n13156), .ZN(n13166) );
  AOI22_X1 U16358 ( .A1(n15698), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15696), .ZN(n19121) );
  INV_X1 U16359 ( .A(n19121), .ZN(n14053) );
  NAND2_X1 U16360 ( .A1(n13166), .A2(n14053), .ZN(n13168) );
  NAND2_X1 U16361 ( .A1(n13113), .A2(n13168), .ZN(P2_U2955) );
  AOI22_X1 U16362 ( .A1(n13161), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13138), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16363 ( .A1(n15698), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15696), .ZN(n19209) );
  INV_X1 U16364 ( .A(n19209), .ZN(n14007) );
  NAND2_X1 U16365 ( .A1(n13166), .A2(n14007), .ZN(n13154) );
  NAND2_X1 U16366 ( .A1(n13114), .A2(n13154), .ZN(P2_U2953) );
  AOI22_X1 U16367 ( .A1(n13161), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13196), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16368 ( .A1(n15698), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15696), .ZN(n19232) );
  INV_X1 U16369 ( .A(n19232), .ZN(n13115) );
  NAND2_X1 U16370 ( .A1(n13166), .A2(n13115), .ZN(n13162) );
  NAND2_X1 U16371 ( .A1(n13116), .A2(n13162), .ZN(P2_U2959) );
  AOI22_X1 U16372 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n13161), .B1(n13196), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13117) );
  OAI22_X1 U16373 ( .A1(n15696), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15698), .ZN(n19225) );
  INV_X1 U16374 ( .A(n19225), .ZN(n16182) );
  NAND2_X1 U16375 ( .A1(n13166), .A2(n16182), .ZN(n13170) );
  NAND2_X1 U16376 ( .A1(n13117), .A2(n13170), .ZN(P2_U2958) );
  INV_X1 U16377 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U16378 ( .A1(n15696), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13120) );
  INV_X1 U16379 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13118) );
  OR2_X1 U16380 ( .A1(n15696), .A2(n13118), .ZN(n13119) );
  NAND2_X1 U16381 ( .A1(n13120), .A2(n13119), .ZN(n19082) );
  NAND2_X1 U16382 ( .A1(n13166), .A2(n19082), .ZN(n13143) );
  NAND2_X1 U16383 ( .A1(n13138), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U16384 ( .C1(n13201), .C2(n19143), .A(n13143), .B(n13121), .ZN(
        P2_U2981) );
  INV_X1 U16385 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19153) );
  NAND2_X1 U16386 ( .A1(n15696), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13123) );
  INV_X1 U16387 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16475) );
  OR2_X1 U16388 ( .A1(n15696), .A2(n16475), .ZN(n13122) );
  NAND2_X1 U16389 ( .A1(n13123), .A2(n13122), .ZN(n19095) );
  NAND2_X1 U16390 ( .A1(n13166), .A2(n19095), .ZN(n13147) );
  NAND2_X1 U16391 ( .A1(n13138), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13124) );
  OAI211_X1 U16392 ( .C1(n13201), .C2(n19153), .A(n13147), .B(n13124), .ZN(
        P2_U2976) );
  INV_X1 U16393 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16394 ( .A1(n15696), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13126) );
  INV_X1 U16395 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16473) );
  OR2_X1 U16396 ( .A1(n15696), .A2(n16473), .ZN(n13125) );
  NAND2_X1 U16397 ( .A1(n13126), .A2(n13125), .ZN(n19092) );
  NAND2_X1 U16398 ( .A1(n13166), .A2(n19092), .ZN(n13140) );
  NAND2_X1 U16399 ( .A1(n13138), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13127) );
  OAI211_X1 U16400 ( .C1(n13201), .C2(n13206), .A(n13140), .B(n13127), .ZN(
        P2_U2962) );
  INV_X1 U16401 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19147) );
  NAND2_X1 U16402 ( .A1(n15696), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13129) );
  INV_X1 U16403 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16470) );
  OR2_X1 U16404 ( .A1(n15696), .A2(n16470), .ZN(n13128) );
  NAND2_X1 U16405 ( .A1(n13129), .A2(n13128), .ZN(n19087) );
  NAND2_X1 U16406 ( .A1(n13166), .A2(n19087), .ZN(n13132) );
  NAND2_X1 U16407 ( .A1(n13138), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13130) );
  OAI211_X1 U16408 ( .C1(n13201), .C2(n19147), .A(n13132), .B(n13130), .ZN(
        P2_U2979) );
  INV_X1 U16409 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13216) );
  NAND2_X1 U16410 ( .A1(n13138), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13131) );
  OAI211_X1 U16411 ( .C1(n13201), .C2(n13216), .A(n13132), .B(n13131), .ZN(
        P2_U2964) );
  INV_X1 U16412 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19155) );
  NAND2_X1 U16413 ( .A1(n15696), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13134) );
  INV_X1 U16414 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16476) );
  OR2_X1 U16415 ( .A1(n15696), .A2(n16476), .ZN(n13133) );
  NAND2_X1 U16416 ( .A1(n13134), .A2(n13133), .ZN(n19099) );
  NAND2_X1 U16417 ( .A1(n13166), .A2(n19099), .ZN(n13137) );
  NAND2_X1 U16418 ( .A1(n13138), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13135) );
  OAI211_X1 U16419 ( .C1(n13201), .C2(n19155), .A(n13137), .B(n13135), .ZN(
        P2_U2975) );
  INV_X1 U16420 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U16421 ( .A1(n13138), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13136) );
  OAI211_X1 U16422 ( .C1(n13201), .C2(n13210), .A(n13137), .B(n13136), .ZN(
        P2_U2960) );
  INV_X1 U16423 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19151) );
  NAND2_X1 U16424 ( .A1(n13138), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13139) );
  OAI211_X1 U16425 ( .C1(n13201), .C2(n19151), .A(n13140), .B(n13139), .ZN(
        P2_U2977) );
  AOI22_X1 U16426 ( .A1(n15698), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15696), .ZN(n19079) );
  INV_X1 U16427 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19141) );
  INV_X1 U16428 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n20861) );
  OAI222_X1 U16429 ( .A1(n13156), .A2(n19079), .B1(n13201), .B2(n19141), .C1(
        n20861), .C2(n13141), .ZN(P2_U2982) );
  INV_X1 U16430 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13208) );
  NAND2_X1 U16431 ( .A1(n13196), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13142) );
  OAI211_X1 U16432 ( .C1(n13201), .C2(n13208), .A(n13143), .B(n13142), .ZN(
        P2_U2966) );
  AOI22_X1 U16433 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13161), .B1(n13196), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13146) );
  INV_X1 U16434 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16468) );
  OR2_X1 U16435 ( .A1(n15696), .A2(n16468), .ZN(n13145) );
  NAND2_X1 U16436 ( .A1(n15696), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13144) );
  AND2_X1 U16437 ( .A1(n13145), .A2(n13144), .ZN(n19085) );
  INV_X1 U16438 ( .A(n19085), .ZN(n15134) );
  NAND2_X1 U16439 ( .A1(n13166), .A2(n15134), .ZN(n13159) );
  NAND2_X1 U16440 ( .A1(n13146), .A2(n13159), .ZN(P2_U2965) );
  AOI22_X1 U16441 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n13161), .B1(n13196), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U16442 ( .A1(n13148), .A2(n13147), .ZN(P2_U2961) );
  AOI22_X1 U16443 ( .A1(n13161), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13196), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13149) );
  INV_X1 U16444 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16492) );
  INV_X1 U16445 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U16446 ( .A1(n15698), .A2(n16492), .B1(n18241), .B2(n15696), .ZN(
        n19070) );
  INV_X1 U16447 ( .A(n19070), .ZN(n19204) );
  OR2_X1 U16448 ( .A1(n13156), .A2(n19204), .ZN(n13174) );
  NAND2_X1 U16449 ( .A1(n13149), .A2(n13174), .ZN(P2_U2952) );
  AOI22_X1 U16450 ( .A1(n13161), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13196), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13153) );
  INV_X1 U16451 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13150) );
  OR2_X1 U16452 ( .A1(n15696), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U16453 ( .A1(n15696), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13151) );
  AND2_X1 U16454 ( .A1(n13152), .A2(n13151), .ZN(n19090) );
  INV_X1 U16455 ( .A(n19090), .ZN(n15148) );
  NAND2_X1 U16456 ( .A1(n13166), .A2(n15148), .ZN(n13197) );
  NAND2_X1 U16457 ( .A1(n13153), .A2(n13197), .ZN(P2_U2978) );
  AOI22_X1 U16458 ( .A1(n13161), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16459 ( .A1(n13155), .A2(n13154), .ZN(P2_U2968) );
  AOI22_X1 U16460 ( .A1(n13161), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13157) );
  INV_X1 U16461 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16482) );
  INV_X1 U16462 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U16463 ( .A1(n15698), .A2(n16482), .B1(n18261), .B2(n15696), .ZN(
        n16189) );
  INV_X1 U16464 ( .A(n16189), .ZN(n19216) );
  OR2_X1 U16465 ( .A1(n13156), .A2(n19216), .ZN(n13176) );
  NAND2_X1 U16466 ( .A1(n13157), .A2(n13176), .ZN(P2_U2971) );
  AOI22_X1 U16467 ( .A1(n13161), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16468 ( .A1(n15698), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15696), .ZN(n19221) );
  INV_X1 U16469 ( .A(n19221), .ZN(n19106) );
  NAND2_X1 U16470 ( .A1(n13166), .A2(n19106), .ZN(n13164) );
  NAND2_X1 U16471 ( .A1(n13158), .A2(n13164), .ZN(P2_U2972) );
  AOI22_X1 U16472 ( .A1(n13161), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13196), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U16473 ( .A1(n13160), .A2(n13159), .ZN(P2_U2980) );
  AOI22_X1 U16474 ( .A1(n13161), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13163) );
  NAND2_X1 U16475 ( .A1(n13163), .A2(n13162), .ZN(P2_U2974) );
  AOI22_X1 U16476 ( .A1(n13161), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13196), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13165) );
  NAND2_X1 U16477 ( .A1(n13165), .A2(n13164), .ZN(P2_U2957) );
  AOI22_X1 U16478 ( .A1(n13161), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13196), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U16479 ( .A1(n15698), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15696), .ZN(n19128) );
  INV_X1 U16480 ( .A(n19128), .ZN(n14028) );
  NAND2_X1 U16481 ( .A1(n13166), .A2(n14028), .ZN(n13172) );
  NAND2_X1 U16482 ( .A1(n13167), .A2(n13172), .ZN(P2_U2954) );
  AOI22_X1 U16483 ( .A1(n13161), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U16484 ( .A1(n13169), .A2(n13168), .ZN(P2_U2970) );
  AOI22_X1 U16485 ( .A1(n13161), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U16486 ( .A1(n13171), .A2(n13170), .ZN(P2_U2973) );
  AOI22_X1 U16487 ( .A1(n13161), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16488 ( .A1(n13173), .A2(n13172), .ZN(P2_U2969) );
  AOI22_X1 U16489 ( .A1(n13161), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13196), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U16490 ( .A1(n13175), .A2(n13174), .ZN(P2_U2967) );
  AOI22_X1 U16491 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n13161), .B1(n13196), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13177) );
  NAND2_X1 U16492 ( .A1(n13177), .A2(n13176), .ZN(P2_U2956) );
  NOR2_X1 U16493 ( .A1(n10511), .A2(n13178), .ZN(n13179) );
  NAND2_X1 U16494 ( .A1(n13200), .A2(n13179), .ZN(n13187) );
  NOR2_X1 U16495 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  AOI21_X1 U16496 ( .B1(n16345), .B2(n13183), .A(n13182), .ZN(n13230) );
  INV_X1 U16497 ( .A(n13184), .ZN(n13186) );
  AND4_X1 U16498 ( .A1(n13187), .A2(n13230), .A3(n13186), .A4(n13185), .ZN(
        n16357) );
  OR2_X1 U16499 ( .A1(n16357), .A2(n13188), .ZN(n13190) );
  NOR2_X1 U16500 ( .A1(n19852), .A2(n13789), .ZN(n19830) );
  NAND2_X1 U16501 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19830), .ZN(n16378) );
  INV_X1 U16502 ( .A(n16378), .ZN(n16379) );
  AOI22_X1 U16503 ( .A1(n16379), .A2(P2_FLUSH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(n19716), .ZN(n13189) );
  NAND2_X1 U16504 ( .A1(n13190), .A2(n13189), .ZN(n15685) );
  AND3_X1 U16505 ( .A1(n13193), .A2(n13192), .A3(n13191), .ZN(n16336) );
  NAND3_X1 U16506 ( .A1(n15685), .A2(n19799), .A3(n16336), .ZN(n13194) );
  OAI21_X1 U16507 ( .B1(n15685), .B2(n13195), .A(n13194), .ZN(P2_U3595) );
  AOI22_X1 U16508 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13161), .B1(n13196), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16509 ( .A1(n13198), .A2(n13197), .ZN(P2_U2963) );
  INV_X1 U16510 ( .A(n10511), .ZN(n13199) );
  NAND3_X1 U16511 ( .A1(n13200), .A2(n13199), .A3(n19721), .ZN(n13202) );
  NAND2_X1 U16512 ( .A1(n13202), .A2(n13201), .ZN(n13204) );
  INV_X1 U16513 ( .A(n19848), .ZN(n13203) );
  NAND2_X1 U16514 ( .A1(n19139), .A2(n19846), .ZN(n13327) );
  INV_X1 U16515 ( .A(n19830), .ZN(n15690) );
  NOR2_X1 U16516 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15690), .ZN(n19165) );
  AOI22_X1 U16517 ( .A1(n19860), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13205) );
  OAI21_X1 U16518 ( .B1(n13206), .B2(n13327), .A(n13205), .ZN(P2_U2925) );
  AOI22_X1 U16519 ( .A1(n19860), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13207) );
  OAI21_X1 U16520 ( .B1(n13208), .B2(n13327), .A(n13207), .ZN(P2_U2921) );
  AOI22_X1 U16521 ( .A1(n19860), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13209) );
  OAI21_X1 U16522 ( .B1(n13210), .B2(n13327), .A(n13209), .ZN(P2_U2927) );
  INV_X1 U16523 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U16524 ( .A1(n19860), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13211) );
  OAI21_X1 U16525 ( .B1(n13212), .B2(n13327), .A(n13211), .ZN(P2_U2922) );
  INV_X1 U16526 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16527 ( .A1(n19860), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13213) );
  OAI21_X1 U16528 ( .B1(n13214), .B2(n13327), .A(n13213), .ZN(P2_U2926) );
  AOI22_X1 U16529 ( .A1(n19860), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13215) );
  OAI21_X1 U16530 ( .B1(n13216), .B2(n13327), .A(n13215), .ZN(P2_U2923) );
  INV_X1 U16531 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U16532 ( .A1(n19860), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13217) );
  OAI21_X1 U16533 ( .B1(n13218), .B2(n13327), .A(n13217), .ZN(P2_U2924) );
  INV_X1 U16534 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19208) );
  NAND2_X1 U16535 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19240), .ZN(n13220) );
  NOR2_X1 U16536 ( .A1(n19224), .A2(n13220), .ZN(n13221) );
  OAI21_X1 U16537 ( .B1(n10566), .B2(n19208), .A(n13221), .ZN(n13222) );
  INV_X1 U16538 ( .A(n13222), .ZN(n13223) );
  NOR2_X1 U16539 ( .A1(n19058), .A2(n13579), .ZN(n13224) );
  AOI21_X1 U16540 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n13579), .A(n13224), .ZN(
        n13225) );
  OAI21_X1 U16541 ( .B1(n19827), .B2(n15130), .A(n13225), .ZN(P2_U2887) );
  AND2_X1 U16542 ( .A1(n20499), .A2(n20634), .ZN(n13242) );
  NAND2_X1 U16543 ( .A1(n13507), .A2(n13251), .ZN(n13893) );
  INV_X1 U16544 ( .A(n13893), .ZN(n13226) );
  AOI211_X1 U16545 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13227), .A(n13242), 
        .B(n13226), .ZN(n13228) );
  INV_X1 U16546 ( .A(n13228), .ZN(P1_U2801) );
  NAND2_X1 U16547 ( .A1(n13230), .A2(n13229), .ZN(n13231) );
  NAND2_X1 U16548 ( .A1(n19103), .A2(n13232), .ZN(n19134) );
  NAND2_X1 U16549 ( .A1(n19103), .A2(n10509), .ZN(n16191) );
  AOI21_X1 U16550 ( .B1(n19827), .B2(n19108), .A(n19130), .ZN(n13241) );
  INV_X1 U16551 ( .A(n13233), .ZN(n13234) );
  XNOR2_X1 U16552 ( .A(n13235), .B(n13234), .ZN(n19054) );
  INV_X1 U16553 ( .A(n19054), .ZN(n16317) );
  NOR2_X1 U16554 ( .A1(n19134), .A2(n19054), .ZN(n13236) );
  AOI22_X1 U16555 ( .A1(n19063), .A2(n13236), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19129), .ZN(n13240) );
  AND2_X1 U16556 ( .A1(n19103), .A2(n13238), .ZN(n14006) );
  NAND2_X1 U16557 ( .A1(n19105), .A2(n19070), .ZN(n13239) );
  OAI211_X1 U16558 ( .C1(n13241), .C2(n16317), .A(n13240), .B(n13239), .ZN(
        P2_U2919) );
  NOR2_X1 U16559 ( .A1(n13242), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13246)
         );
  OAI21_X1 U16560 ( .B1(n13815), .B2(n13244), .A(n20739), .ZN(n13245) );
  OAI21_X1 U16561 ( .B1(n13246), .B2(n20739), .A(n13245), .ZN(P1_U3487) );
  INV_X1 U16562 ( .A(n13247), .ZN(n13249) );
  MUX2_X1 U16563 ( .A(n13548), .B(n15641), .S(n15123), .Z(n13250) );
  OAI21_X1 U16564 ( .B1(n19817), .B2(n15130), .A(n13250), .ZN(P2_U2886) );
  OR2_X1 U16565 ( .A1(n13252), .A2(n13251), .ZN(n13254) );
  OR2_X1 U16566 ( .A1(n13499), .A2(n13815), .ZN(n13253) );
  NAND2_X1 U16567 ( .A1(n13254), .A2(n13253), .ZN(n19871) );
  OR2_X1 U16568 ( .A1(n13255), .A2(n13459), .ZN(n13256) );
  AND2_X1 U16569 ( .A1(n13256), .A2(n20741), .ZN(n20743) );
  NOR2_X1 U16570 ( .A1(n19871), .A2(n20743), .ZN(n15866) );
  INV_X1 U16571 ( .A(n13501), .ZN(n19870) );
  OR2_X1 U16572 ( .A1(n15866), .A2(n19870), .ZN(n13270) );
  INV_X1 U16573 ( .A(n13270), .ZN(n19879) );
  INV_X1 U16574 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16575 ( .A1(n13353), .A2(n11136), .ZN(n13257) );
  NAND2_X1 U16576 ( .A1(n13363), .A2(n13257), .ZN(n13510) );
  NAND3_X1 U16577 ( .A1(n13259), .A2(n13258), .A3(n20037), .ZN(n13260) );
  NAND2_X1 U16578 ( .A1(n13510), .A2(n13260), .ZN(n13267) );
  NAND2_X1 U16579 ( .A1(n13516), .A2(n13261), .ZN(n13264) );
  INV_X1 U16580 ( .A(n13817), .ZN(n13262) );
  NAND2_X1 U16581 ( .A1(n13262), .A2(n11136), .ZN(n13263) );
  NAND2_X1 U16582 ( .A1(n13266), .A2(n13265), .ZN(n13500) );
  INV_X1 U16583 ( .A(n13384), .ZN(n13519) );
  MUX2_X1 U16584 ( .A(n13267), .B(n13519), .S(n13499), .Z(n13269) );
  NOR2_X1 U16585 ( .A1(n12143), .A2(n13496), .ZN(n13268) );
  OAI21_X1 U16586 ( .B1(n13269), .B2(n13268), .A(n9635), .ZN(n15868) );
  OR2_X1 U16587 ( .A1(n13270), .A2(n15868), .ZN(n13271) );
  OAI21_X1 U16588 ( .B1(n19879), .B2(n13272), .A(n13271), .ZN(P1_U3484) );
  NAND2_X1 U16589 ( .A1(n13275), .A2(n13274), .ZN(n13277) );
  AND2_X1 U16590 ( .A1(n13277), .A2(n9857), .ZN(n15179) );
  INV_X1 U16591 ( .A(n15179), .ZN(n19809) );
  AOI22_X1 U16592 ( .A1(n19809), .A2(n16307), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13278), .ZN(n13295) );
  INV_X1 U16593 ( .A(n13279), .ZN(n13292) );
  INV_X1 U16594 ( .A(n13280), .ZN(n13283) );
  OR2_X1 U16595 ( .A1(n10856), .A2(n13281), .ZN(n19199) );
  OAI211_X1 U16596 ( .C1(n15490), .C2(n13283), .A(n13282), .B(n19199), .ZN(
        n13291) );
  NAND2_X1 U16597 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  NAND2_X1 U16598 ( .A1(n13287), .A2(n13286), .ZN(n19195) );
  XNOR2_X1 U16599 ( .A(n13289), .B(n13288), .ZN(n19193) );
  OAI22_X1 U16600 ( .A1(n16299), .A2(n19195), .B1(n19193), .B2(n16330), .ZN(
        n13290) );
  AOI211_X1 U16601 ( .C1(n13293), .C2(n13292), .A(n13291), .B(n13290), .ZN(
        n13294) );
  OAI211_X1 U16602 ( .C1(n13273), .C2(n16319), .A(n13295), .B(n13294), .ZN(
        P2_U3044) );
  INV_X1 U16603 ( .A(n19194), .ZN(n19180) );
  OAI21_X1 U16604 ( .B1(n13544), .B2(n13305), .A(n13296), .ZN(n13297) );
  XNOR2_X1 U16605 ( .A(n13297), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15645) );
  AOI22_X1 U16606 ( .A1(n19180), .A2(n15645), .B1(n19177), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13301) );
  AOI21_X1 U16607 ( .B1(n15642), .B2(n13299), .A(n13298), .ZN(n15646) );
  AOI22_X1 U16608 ( .A1(n9578), .A2(n15646), .B1(P2_REIP_REG_1__SCAN_IN), .B2(
        n19176), .ZN(n13300) );
  NAND2_X1 U16609 ( .A1(n13301), .A2(n13300), .ZN(n13302) );
  AOI21_X1 U16610 ( .B1(n16258), .B2(n13547), .A(n13302), .ZN(n13303) );
  OAI21_X1 U16611 ( .B1(n15641), .B2(n19185), .A(n13303), .ZN(P2_U3013) );
  NAND2_X1 U16612 ( .A1(n19051), .A2(n13790), .ZN(n13304) );
  AND2_X1 U16613 ( .A1(n13305), .A2(n13304), .ZN(n16325) );
  OR2_X1 U16614 ( .A1(n13306), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13307) );
  NAND2_X1 U16615 ( .A1(n13308), .A2(n13307), .ZN(n16329) );
  OR2_X1 U16616 ( .A1(n10856), .A2(n10052), .ZN(n16327) );
  OAI21_X1 U16617 ( .B1(n19192), .B2(n16329), .A(n16327), .ZN(n13309) );
  AOI21_X1 U16618 ( .B1(n19180), .B2(n16325), .A(n13309), .ZN(n13312) );
  OAI21_X1 U16619 ( .B1(n19177), .B2(n13310), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13311) );
  OAI211_X1 U16620 ( .C1(n19185), .C2(n19058), .A(n13312), .B(n13311), .ZN(
        P2_U3014) );
  INV_X1 U16621 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U16622 ( .A1(n19860), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13313) );
  OAI21_X1 U16623 ( .B1(n13314), .B2(n13327), .A(n13313), .ZN(P2_U2929) );
  INV_X1 U16624 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U16625 ( .A1(n19860), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13315) );
  OAI21_X1 U16626 ( .B1(n15171), .B2(n13327), .A(n13315), .ZN(P2_U2928) );
  INV_X1 U16627 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16628 ( .A1(n19860), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13316) );
  OAI21_X1 U16629 ( .B1(n13317), .B2(n13327), .A(n13316), .ZN(P2_U2933) );
  INV_X1 U16630 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U16631 ( .A1(n19860), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13318) );
  OAI21_X1 U16632 ( .B1(n13319), .B2(n13327), .A(n13318), .ZN(P2_U2932) );
  INV_X1 U16633 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16634 ( .A1(n19860), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13320) );
  OAI21_X1 U16635 ( .B1(n13321), .B2(n13327), .A(n13320), .ZN(P2_U2930) );
  INV_X1 U16636 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16637 ( .A1(n19860), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13322) );
  OAI21_X1 U16638 ( .B1(n13323), .B2(n13327), .A(n13322), .ZN(P2_U2934) );
  INV_X1 U16639 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U16640 ( .A1(n19860), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U16641 ( .B1(n13325), .B2(n13327), .A(n13324), .ZN(P2_U2935) );
  INV_X1 U16642 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U16643 ( .A1(n19860), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U16644 ( .B1(n13328), .B2(n13327), .A(n13326), .ZN(P2_U2931) );
  OAI21_X1 U16645 ( .B1(n13331), .B2(n13330), .A(n13329), .ZN(n14464) );
  NAND2_X1 U16646 ( .A1(n13332), .A2(n14741), .ZN(n13336) );
  AND2_X1 U16647 ( .A1(n19973), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13527) );
  OAI21_X1 U16648 ( .B1(n13334), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13333), .ZN(n13529) );
  NOR2_X1 U16649 ( .A1(n13529), .A2(n19877), .ZN(n13335) );
  AOI211_X1 U16650 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13336), .A(
        n13527), .B(n13335), .ZN(n13337) );
  OAI21_X1 U16651 ( .B1(n20031), .B2(n14464), .A(n13337), .ZN(P1_U2999) );
  INV_X1 U16652 ( .A(n13339), .ZN(n13340) );
  INV_X1 U16653 ( .A(n19810), .ZN(n15178) );
  MUX2_X1 U16654 ( .A(n13434), .B(n13273), .S(n15123), .Z(n13342) );
  OAI21_X1 U16655 ( .B1(n15178), .B2(n15130), .A(n13342), .ZN(P2_U2885) );
  NAND2_X1 U16656 ( .A1(n9633), .A2(n20741), .ZN(n13344) );
  NAND2_X1 U16657 ( .A1(n13363), .A2(n13815), .ZN(n13385) );
  OAI21_X1 U16658 ( .B1(n13343), .B2(n13344), .A(n13385), .ZN(n13345) );
  NAND2_X1 U16659 ( .A1(n13345), .A2(n13499), .ZN(n13350) );
  NAND2_X1 U16660 ( .A1(n13815), .A2(n13346), .ZN(n13347) );
  NOR2_X1 U16661 ( .A1(n13348), .A2(n13347), .ZN(n13697) );
  NAND3_X1 U16662 ( .A1(n13697), .A2(n13496), .A3(n20741), .ZN(n13349) );
  NOR2_X1 U16663 ( .A1(n20073), .A2(n19870), .ZN(n13352) );
  NOR2_X1 U16664 ( .A1(n9634), .A2(n11115), .ZN(n13351) );
  NAND4_X1 U16665 ( .A1(n13371), .A2(n13352), .A3(n13351), .A4(n20078), .ZN(
        n13726) );
  OR2_X1 U16666 ( .A1(n13726), .A2(n13353), .ZN(n13354) );
  NAND2_X1 U16667 ( .A1(n13360), .A2(n9635), .ZN(n13356) );
  NAND2_X2 U16668 ( .A1(n14614), .A2(n13356), .ZN(n14622) );
  NAND2_X1 U16669 ( .A1(n20030), .A2(DATAI_0_), .ZN(n13358) );
  NAND2_X1 U16670 ( .A1(n20032), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13357) );
  AND2_X1 U16671 ( .A1(n13358), .A2(n13357), .ZN(n20048) );
  INV_X1 U16672 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13762) );
  OAI222_X1 U16673 ( .A1(n14464), .A2(n14622), .B1(n14617), .B2(n20048), .C1(
        n14614), .C2(n13762), .ZN(P1_U2904) );
  INV_X1 U16674 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20451) );
  AND2_X1 U16675 ( .A1(n14311), .A2(n13343), .ZN(n13369) );
  NAND3_X1 U16676 ( .A1(n13499), .A2(n13459), .A3(n20741), .ZN(n13368) );
  INV_X1 U16677 ( .A(n13359), .ZN(n13367) );
  OAI21_X1 U16678 ( .B1(n13360), .B2(n11495), .A(n20037), .ZN(n13361) );
  INV_X1 U16679 ( .A(n13361), .ZN(n13362) );
  NAND2_X1 U16680 ( .A1(n11149), .A2(n13362), .ZN(n13377) );
  NAND2_X1 U16681 ( .A1(n13363), .A2(n13377), .ZN(n13364) );
  NAND2_X1 U16682 ( .A1(n13364), .A2(n12143), .ZN(n13498) );
  OAI211_X1 U16683 ( .C1(n13817), .C2(n20059), .A(n13498), .B(n13728), .ZN(
        n13365) );
  INV_X1 U16684 ( .A(n13365), .ZN(n13366) );
  NOR2_X1 U16685 ( .A1(n20638), .A2(n20634), .ZN(n16147) );
  INV_X1 U16686 ( .A(n16147), .ZN(n16152) );
  NOR2_X1 U16687 ( .A1(n20635), .A2(n16152), .ZN(n13701) );
  AOI22_X1 U16688 ( .A1(n13501), .A2(n15854), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13701), .ZN(n16143) );
  OAI21_X1 U16689 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20451), .A(n16143), 
        .ZN(n20727) );
  INV_X1 U16690 ( .A(n20727), .ZN(n13395) );
  INV_X1 U16691 ( .A(n20448), .ZN(n20043) );
  INV_X1 U16692 ( .A(n13371), .ZN(n13372) );
  NAND2_X1 U16693 ( .A1(n13373), .A2(n13372), .ZN(n13375) );
  AOI21_X1 U16694 ( .B1(n20054), .B2(n13375), .A(n13374), .ZN(n13379) );
  NAND2_X1 U16695 ( .A1(n13376), .A2(n13815), .ZN(n13378) );
  AND3_X1 U16696 ( .A1(n13379), .A2(n13378), .A3(n13377), .ZN(n13521) );
  NAND2_X1 U16697 ( .A1(n13522), .A2(n20073), .ZN(n13380) );
  NOR2_X1 U16698 ( .A1(n13697), .A2(n13380), .ZN(n13381) );
  NAND2_X1 U16699 ( .A1(n13521), .A2(n13381), .ZN(n14965) );
  NOR2_X1 U16700 ( .A1(n14311), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14964) );
  NOR2_X1 U16701 ( .A1(n14311), .A2(n9701), .ZN(n13382) );
  MUX2_X1 U16702 ( .A(n14964), .B(n13382), .S(n11166), .Z(n13389) );
  NOR2_X1 U16703 ( .A1(n13383), .A2(n14962), .ZN(n13683) );
  NAND2_X1 U16704 ( .A1(n13385), .A2(n13384), .ZN(n13678) );
  INV_X1 U16705 ( .A(n13682), .ZN(n13387) );
  INV_X1 U16706 ( .A(n10968), .ZN(n13386) );
  NAND2_X1 U16707 ( .A1(n13386), .A2(n11166), .ZN(n13676) );
  NAND2_X1 U16708 ( .A1(n13387), .A2(n13676), .ZN(n13391) );
  MUX2_X1 U16709 ( .A(n13683), .B(n13678), .S(n13391), .Z(n13388) );
  AOI211_X1 U16710 ( .C1(n20043), .C2(n14965), .A(n13389), .B(n13388), .ZN(
        n13390) );
  INV_X1 U16711 ( .A(n13390), .ZN(n13675) );
  INV_X1 U16712 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14309) );
  NOR2_X1 U16713 ( .A1(n20634), .A2(n14309), .ZN(n14968) );
  AOI22_X1 U16714 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20012), .B2(n14279), .ZN(
        n14966) );
  INV_X1 U16715 ( .A(n15880), .ZN(n20722) );
  INV_X1 U16716 ( .A(n13391), .ZN(n13392) );
  AOI222_X1 U16717 ( .A1(n13675), .A2(n20724), .B1(n14968), .B2(n14966), .C1(
        n20722), .C2(n13392), .ZN(n13394) );
  NAND2_X1 U16718 ( .A1(n13395), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13393) );
  OAI21_X1 U16719 ( .B1(n13395), .B2(n13394), .A(n13393), .ZN(P1_U3472) );
  INV_X1 U16720 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19219) );
  NOR2_X1 U16721 ( .A1(n13397), .A2(n19219), .ZN(n13398) );
  NAND2_X1 U16722 ( .A1(n13396), .A2(n13398), .ZN(n13581) );
  OAI21_X1 U16723 ( .B1(n13396), .B2(n13398), .A(n13581), .ZN(n19107) );
  NAND2_X1 U16724 ( .A1(n13401), .A2(n13400), .ZN(n13402) );
  NAND2_X1 U16725 ( .A1(n13399), .A2(n13402), .ZN(n19184) );
  MUX2_X1 U16726 ( .A(n19184), .B(n13403), .S(n13579), .Z(n13404) );
  OAI21_X1 U16727 ( .B1(n19107), .B2(n15130), .A(n13404), .ZN(P2_U2883) );
  NOR2_X1 U16728 ( .A1(n13574), .A2(n13405), .ZN(n13406) );
  OR2_X1 U16729 ( .A1(n13670), .A2(n13406), .ZN(n16309) );
  NOR2_X1 U16730 ( .A1(n12329), .A2(n13407), .ZN(n13408) );
  XNOR2_X1 U16731 ( .A(n13408), .B(n16250), .ZN(n13409) );
  NAND2_X1 U16732 ( .A1(n13409), .A2(n19042), .ZN(n13418) );
  INV_X1 U16733 ( .A(n19046), .ZN(n19055) );
  AOI21_X1 U16734 ( .B1(n13411), .B2(n13410), .A(n15582), .ZN(n19098) );
  AOI22_X1 U16735 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19049), .ZN(n13412) );
  OAI211_X1 U16736 ( .C1(n19030), .C2(n13413), .A(n13412), .B(n18941), .ZN(
        n13416) );
  NOR2_X1 U16737 ( .A1(n13414), .A2(n19052), .ZN(n13415) );
  AOI211_X1 U16738 ( .C1(n19055), .C2(n19098), .A(n13416), .B(n13415), .ZN(
        n13417) );
  OAI211_X1 U16739 ( .C1(n16309), .C2(n19057), .A(n13418), .B(n13417), .ZN(
        P2_U2847) );
  INV_X1 U16740 ( .A(n19064), .ZN(n13458) );
  INV_X1 U16741 ( .A(n19189), .ZN(n13422) );
  NOR2_X1 U16742 ( .A1(n12329), .A2(n13419), .ZN(n13421) );
  AOI21_X1 U16743 ( .B1(n13422), .B2(n13421), .A(n19724), .ZN(n13420) );
  OAI21_X1 U16744 ( .B1(n13422), .B2(n13421), .A(n13420), .ZN(n13431) );
  INV_X1 U16745 ( .A(n19184), .ZN(n13949) );
  XNOR2_X1 U16746 ( .A(n13424), .B(n13423), .ZN(n15181) );
  AOI22_X1 U16747 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19036), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19048), .ZN(n13425) );
  OAI211_X1 U16748 ( .C1(n19046), .C2(n15181), .A(n13425), .B(n18941), .ZN(
        n13426) );
  AOI21_X1 U16749 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n19049), .A(n13426), .ZN(
        n13427) );
  OAI21_X1 U16750 ( .B1(n13428), .B2(n19052), .A(n13427), .ZN(n13429) );
  AOI21_X1 U16751 ( .B1(n13949), .B2(n19041), .A(n13429), .ZN(n13430) );
  OAI211_X1 U16752 ( .C1(n19107), .C2(n13458), .A(n13431), .B(n13430), .ZN(
        P2_U2851) );
  NOR2_X1 U16753 ( .A1(n12329), .A2(n13432), .ZN(n13552) );
  XNOR2_X1 U16754 ( .A(n13552), .B(n19190), .ZN(n13433) );
  NAND2_X1 U16755 ( .A1(n13433), .A2(n19042), .ZN(n13441) );
  OAI22_X1 U16756 ( .A1(n19032), .A2(n13434), .B1(n15179), .B2(n19046), .ZN(
        n13436) );
  NOR2_X1 U16757 ( .A1(n19030), .A2(n13281), .ZN(n13435) );
  AOI211_X1 U16758 ( .C1(n19036), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13436), .B(n13435), .ZN(n13437) );
  OAI21_X1 U16759 ( .B1(n13438), .B2(n19052), .A(n13437), .ZN(n13439) );
  AOI21_X1 U16760 ( .B1(n9595), .B2(n19041), .A(n13439), .ZN(n13440) );
  OAI211_X1 U16761 ( .C1(n13458), .C2(n15178), .A(n13441), .B(n13440), .ZN(
        P2_U2853) );
  NAND2_X1 U16762 ( .A1(n12347), .A2(n13446), .ZN(n13447) );
  XNOR2_X1 U16763 ( .A(n16257), .B(n13447), .ZN(n13448) );
  NAND2_X1 U16764 ( .A1(n13448), .A2(n19042), .ZN(n13457) );
  XNOR2_X1 U16765 ( .A(n13449), .B(n9648), .ZN(n19805) );
  CLKBUF_X1 U16766 ( .A(n13450), .Z(n16261) );
  NOR2_X1 U16767 ( .A1(n13451), .A2(n19052), .ZN(n13453) );
  OAI22_X1 U16768 ( .A1(n10080), .A2(n19060), .B1(n10081), .B2(n19030), .ZN(
        n13452) );
  AOI211_X1 U16769 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19049), .A(n13453), .B(
        n13452), .ZN(n13454) );
  OAI21_X1 U16770 ( .B1(n16261), .B2(n19057), .A(n13454), .ZN(n13455) );
  AOI21_X1 U16771 ( .B1(n19805), .B2(n19055), .A(n13455), .ZN(n13456) );
  OAI211_X1 U16772 ( .C1(n13458), .C2(n19801), .A(n13457), .B(n13456), .ZN(
        P2_U2852) );
  NAND2_X1 U16773 ( .A1(n14311), .A2(n20054), .ZN(n13460) );
  NAND2_X1 U16774 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  NOR2_X1 U16775 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16152), .ZN(n20742) );
  INV_X1 U16776 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13465) );
  INV_X1 U16777 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14086) );
  INV_X1 U16778 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13464) );
  OAI222_X1 U16779 ( .A1(n13739), .A2(n13465), .B1(n13769), .B2(n14086), .C1(
        n13464), .C2(n13766), .ZN(P1_U2906) );
  INV_X1 U16780 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n13467) );
  INV_X1 U16781 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n13466) );
  OAI222_X1 U16782 ( .A1(n13467), .A2(n13739), .B1(n13772), .B2(n11582), .C1(
        n13766), .C2(n13466), .ZN(P1_U2929) );
  INV_X1 U16783 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n13469) );
  INV_X1 U16784 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n13468) );
  OAI222_X1 U16785 ( .A1(n13469), .A2(n13739), .B1(n13772), .B2(n11575), .C1(
        n13766), .C2(n13468), .ZN(P1_U2930) );
  INV_X1 U16786 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13471) );
  INV_X1 U16787 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14083) );
  INV_X1 U16788 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n13470) );
  OAI222_X1 U16789 ( .A1(n13471), .A2(n13739), .B1(n13769), .B2(n14083), .C1(
        n13470), .C2(n13766), .ZN(P1_U2907) );
  INV_X1 U16790 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n13473) );
  INV_X1 U16791 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n13472) );
  OAI222_X1 U16792 ( .A1(n13473), .A2(n13739), .B1(n13772), .B2(n11532), .C1(
        n13766), .C2(n13472), .ZN(P1_U2935) );
  INV_X1 U16793 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n13475) );
  INV_X1 U16794 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13635) );
  INV_X1 U16795 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n13474) );
  OAI222_X1 U16796 ( .A1(n13475), .A2(n13739), .B1(n13772), .B2(n13635), .C1(
        n13766), .C2(n13474), .ZN(P1_U2931) );
  INV_X1 U16797 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n13477) );
  INV_X1 U16798 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13596) );
  INV_X1 U16799 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n13476) );
  OAI222_X1 U16800 ( .A1(n13477), .A2(n13739), .B1(n13772), .B2(n13596), .C1(
        n13766), .C2(n13476), .ZN(P1_U2932) );
  INV_X1 U16801 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n13479) );
  INV_X1 U16802 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13591) );
  INV_X1 U16803 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n13478) );
  OAI222_X1 U16804 ( .A1(n13479), .A2(n13739), .B1(n13772), .B2(n13591), .C1(
        n13766), .C2(n13478), .ZN(P1_U2933) );
  XOR2_X1 U16805 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13581), .Z(n13485)
         );
  NAND2_X1 U16806 ( .A1(n13399), .A2(n13481), .ZN(n13482) );
  AND2_X1 U16807 ( .A1(n13480), .A2(n13482), .ZN(n19040) );
  NOR2_X1 U16808 ( .A1(n15123), .A2(n19031), .ZN(n13483) );
  AOI21_X1 U16809 ( .B1(n19040), .B2(n15123), .A(n13483), .ZN(n13484) );
  OAI21_X1 U16810 ( .B1(n13485), .B2(n15130), .A(n13484), .ZN(P2_U2882) );
  MUX2_X1 U16811 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n12379), .S(n15123), .Z(
        n13486) );
  AOI21_X1 U16812 ( .B1(n15727), .B2(n15118), .A(n13486), .ZN(n13487) );
  INV_X1 U16813 ( .A(n13487), .ZN(P2_U2884) );
  OAI21_X1 U16814 ( .B1(n13489), .B2(n13488), .A(n13560), .ZN(n13861) );
  NAND2_X1 U16815 ( .A1(n19952), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14951) );
  OAI21_X1 U16816 ( .B1(n14741), .B2(n13853), .A(n14951), .ZN(n13490) );
  AOI21_X1 U16817 ( .B1(n16048), .B2(n13853), .A(n13490), .ZN(n13494) );
  OR2_X1 U16818 ( .A1(n13491), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14949) );
  NAND3_X1 U16819 ( .A1(n14949), .A2(n13492), .A3(n19981), .ZN(n13493) );
  OAI211_X1 U16820 ( .C1(n13861), .C2(n20031), .A(n13494), .B(n13493), .ZN(
        P1_U2998) );
  NAND2_X1 U16821 ( .A1(n20054), .A2(n15900), .ZN(n13495) );
  NAND4_X1 U16822 ( .A1(n13496), .A2(n20059), .A3(n20741), .A4(n13495), .ZN(
        n13497) );
  OAI211_X1 U16823 ( .C1(n13500), .C2(n13499), .A(n13498), .B(n13497), .ZN(
        n13502) );
  NAND2_X1 U16824 ( .A1(n13502), .A2(n13501), .ZN(n13509) );
  NAND2_X1 U16825 ( .A1(n13503), .A2(n20741), .ZN(n13504) );
  OAI211_X1 U16826 ( .C1(n13343), .C2(n13504), .A(n20037), .B(n14316), .ZN(
        n13505) );
  NAND3_X1 U16827 ( .A1(n13507), .A2(n13506), .A3(n13505), .ZN(n13508) );
  OAI211_X1 U16828 ( .C1(n13512), .C2(n13514), .A(n13511), .B(n13510), .ZN(
        n13513) );
  OR2_X1 U16829 ( .A1(n13343), .A2(n20744), .ZN(n15878) );
  OAI21_X1 U16830 ( .B1(n13514), .B2(n11115), .A(n15878), .ZN(n13515) );
  OR2_X1 U16831 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13518) );
  AND2_X1 U16832 ( .A1(n13518), .A2(n13517), .ZN(n13737) );
  OAI211_X1 U16833 ( .C1(n13522), .C2(n20037), .A(n13521), .B(n13520), .ZN(
        n13523) );
  NAND2_X1 U16834 ( .A1(n13524), .A2(n13523), .ZN(n14916) );
  NAND2_X1 U16835 ( .A1(n20018), .A2(n14916), .ZN(n14291) );
  INV_X1 U16836 ( .A(n14291), .ZN(n13525) );
  NOR2_X1 U16837 ( .A1(n13524), .A2(n19952), .ZN(n14920) );
  AOI21_X1 U16838 ( .B1(n14309), .B2(n14291), .A(n14920), .ZN(n14952) );
  INV_X1 U16839 ( .A(n14311), .ZN(n13685) );
  AOI22_X1 U16840 ( .A1(n13525), .A2(n14309), .B1(n14952), .B2(n14914), .ZN(
        n13526) );
  AOI211_X1 U16841 ( .C1(n20021), .C2(n13737), .A(n13527), .B(n13526), .ZN(
        n13528) );
  OAI21_X1 U16842 ( .B1(n13529), .B2(n16120), .A(n13528), .ZN(P1_U3031) );
  INV_X1 U16843 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16488) );
  NAND2_X1 U16844 ( .A1(n20032), .A2(n16488), .ZN(n13530) );
  OAI21_X1 U16845 ( .B1(n20032), .B2(DATAI_1_), .A(n13530), .ZN(n20056) );
  OAI222_X1 U16846 ( .A1(n14617), .A2(n20056), .B1(n14614), .B2(n11532), .C1(
        n14622), .C2(n13861), .ZN(P1_U2903) );
  NAND2_X1 U16847 ( .A1(n13396), .A2(n13531), .ZN(n13776) );
  INV_X1 U16848 ( .A(n13776), .ZN(n13845) );
  INV_X1 U16849 ( .A(n13532), .ZN(n13533) );
  OAI211_X1 U16850 ( .C1(n13845), .C2(n13533), .A(n15118), .B(n13833), .ZN(
        n13540) );
  INV_X1 U16851 ( .A(n13534), .ZN(n13536) );
  NAND2_X1 U16852 ( .A1(n13535), .A2(n13670), .ZN(n13622) );
  NAND2_X1 U16853 ( .A1(n13536), .A2(n13622), .ZN(n13538) );
  INV_X1 U16854 ( .A(n13597), .ZN(n13537) );
  AND2_X1 U16855 ( .A1(n13538), .A2(n13537), .ZN(n18991) );
  NAND2_X1 U16856 ( .A1(n15123), .A2(n18991), .ZN(n13539) );
  OAI211_X1 U16857 ( .C1(n15123), .C2(n13541), .A(n13540), .B(n13539), .ZN(
        P2_U2876) );
  XNOR2_X1 U16858 ( .A(n13543), .B(n13542), .ZN(n19822) );
  INV_X1 U16859 ( .A(n13544), .ZN(n13545) );
  AOI22_X1 U16860 ( .A1(n19048), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n12367), 
        .B2(n13545), .ZN(n13546) );
  OAI21_X1 U16861 ( .B1(n19060), .B2(n13547), .A(n13546), .ZN(n13550) );
  NOR2_X1 U16862 ( .A1(n19032), .A2(n13548), .ZN(n13549) );
  AOI211_X1 U16863 ( .C1(n19822), .C2(n19055), .A(n13550), .B(n13549), .ZN(
        n13551) );
  OAI21_X1 U16864 ( .B1(n15641), .B2(n19057), .A(n13551), .ZN(n13555) );
  OAI21_X1 U16865 ( .B1(n13791), .B2(n13553), .A(n13552), .ZN(n13792) );
  OAI22_X1 U16866 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18942), .B1(
        n13792), .B2(n19724), .ZN(n13554) );
  AOI211_X1 U16867 ( .C1(n19820), .C2(n19064), .A(n13555), .B(n13554), .ZN(
        n13556) );
  INV_X1 U16868 ( .A(n13556), .ZN(P2_U2854) );
  INV_X1 U16869 ( .A(n13558), .ZN(n13559) );
  AOI21_X1 U16870 ( .B1(n13557), .B2(n13560), .A(n13559), .ZN(n14356) );
  INV_X1 U16871 ( .A(n20031), .ZN(n19980) );
  AOI22_X1 U16872 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13561) );
  OAI21_X1 U16873 ( .B1(n14361), .B2(n19985), .A(n13561), .ZN(n13562) );
  AOI21_X1 U16874 ( .B1(n14356), .B2(n19980), .A(n13562), .ZN(n13567) );
  OR2_X1 U16875 ( .A1(n13564), .A2(n13563), .ZN(n20014) );
  NAND3_X1 U16876 ( .A1(n20014), .A2(n13565), .A3(n19981), .ZN(n13566) );
  NAND2_X1 U16877 ( .A1(n13567), .A2(n13566), .ZN(P1_U2997) );
  INV_X1 U16878 ( .A(n14356), .ZN(n13570) );
  NAND2_X1 U16879 ( .A1(n20030), .A2(DATAI_2_), .ZN(n13569) );
  NAND2_X1 U16880 ( .A1(n20032), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13568) );
  AND2_X1 U16881 ( .A1(n13569), .A2(n13568), .ZN(n20061) );
  INV_X1 U16882 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13650) );
  OAI222_X1 U16883 ( .A1(n13570), .A2(n14622), .B1(n14617), .B2(n20061), .C1(
        n14614), .C2(n13650), .ZN(P1_U2902) );
  INV_X1 U16884 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13580) );
  NOR3_X1 U16885 ( .A1(n13581), .A2(n13580), .A3(n19228), .ZN(n13667) );
  XNOR2_X1 U16886 ( .A(n13667), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13576) );
  NOR2_X1 U16887 ( .A1(n13571), .A2(n13572), .ZN(n13573) );
  OR2_X1 U16888 ( .A1(n13574), .A2(n13573), .ZN(n19013) );
  MUX2_X1 U16889 ( .A(n19013), .B(n10352), .S(n13579), .Z(n13575) );
  OAI21_X1 U16890 ( .B1(n13576), .B2(n15130), .A(n13575), .ZN(P2_U2880) );
  AND2_X1 U16891 ( .A1(n13480), .A2(n13577), .ZN(n13578) );
  NOR2_X1 U16892 ( .A1(n13571), .A2(n13578), .ZN(n15609) );
  INV_X1 U16893 ( .A(n15609), .ZN(n19025) );
  NOR2_X1 U16894 ( .A1(n13581), .A2(n13580), .ZN(n13583) );
  INV_X1 U16895 ( .A(n13667), .ZN(n13582) );
  OAI211_X1 U16896 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13583), .A(
        n13582), .B(n15118), .ZN(n13585) );
  NAND2_X1 U16897 ( .A1(n13579), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13584) );
  OAI211_X1 U16898 ( .C1(n19025), .C2(n13579), .A(n13585), .B(n13584), .ZN(
        P2_U2881) );
  OAI21_X1 U16899 ( .B1(n13588), .B2(n13587), .A(n13586), .ZN(n13831) );
  NAND2_X1 U16900 ( .A1(n20030), .A2(DATAI_3_), .ZN(n13590) );
  NAND2_X1 U16901 ( .A1(n20032), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13589) );
  AND2_X1 U16902 ( .A1(n13590), .A2(n13589), .ZN(n20066) );
  OAI222_X1 U16903 ( .A1(n13831), .A2(n14622), .B1(n14617), .B2(n20066), .C1(
        n14614), .C2(n13591), .ZN(P1_U2901) );
  INV_X1 U16904 ( .A(n13592), .ZN(n13593) );
  XNOR2_X1 U16905 ( .A(n13586), .B(n13593), .ZN(n19979) );
  INV_X1 U16906 ( .A(n19979), .ZN(n13735) );
  NAND2_X1 U16907 ( .A1(n20030), .A2(DATAI_4_), .ZN(n13595) );
  NAND2_X1 U16908 ( .A1(n20032), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13594) );
  AND2_X1 U16909 ( .A1(n13595), .A2(n13594), .ZN(n20070) );
  OAI222_X1 U16910 ( .A1(n14622), .A2(n13735), .B1(n14617), .B2(n20070), .C1(
        n14614), .C2(n13596), .ZN(P1_U2900) );
  OR2_X1 U16911 ( .A1(n13598), .A2(n13597), .ZN(n13600) );
  AND2_X1 U16912 ( .A1(n13600), .A2(n13599), .ZN(n18982) );
  INV_X1 U16913 ( .A(n18982), .ZN(n13606) );
  INV_X1 U16914 ( .A(n13833), .ZN(n13603) );
  INV_X1 U16915 ( .A(n13601), .ZN(n13602) );
  OR2_X1 U16916 ( .A1(n13833), .A2(n13601), .ZN(n13662) );
  OAI211_X1 U16917 ( .C1(n13603), .C2(n13602), .A(n15118), .B(n13662), .ZN(
        n13605) );
  NAND2_X1 U16918 ( .A1(n13579), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13604) );
  OAI211_X1 U16919 ( .C1(n13606), .C2(n13579), .A(n13605), .B(n13604), .ZN(
        P2_U2875) );
  OAI21_X1 U16920 ( .B1(n13609), .B2(n13608), .A(n13607), .ZN(n13610) );
  INV_X1 U16921 ( .A(n13610), .ZN(n20004) );
  NAND2_X1 U16922 ( .A1(n20004), .A2(n19981), .ZN(n13613) );
  AND2_X1 U16923 ( .A1(n19973), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20001) );
  NOR2_X1 U16924 ( .A1(n19985), .A2(n13821), .ZN(n13611) );
  AOI211_X1 U16925 ( .C1(n19974), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20001), .B(n13611), .ZN(n13612) );
  OAI211_X1 U16926 ( .C1(n20031), .C2(n13831), .A(n13613), .B(n13612), .ZN(
        P1_U2996) );
  AOI21_X1 U16927 ( .B1(n13614), .B2(n13615), .A(n15567), .ZN(n16292) );
  INV_X1 U16928 ( .A(n16292), .ZN(n19094) );
  NOR2_X1 U16929 ( .A1(n12329), .A2(n13616), .ZN(n13617) );
  XNOR2_X1 U16930 ( .A(n13617), .B(n16228), .ZN(n13618) );
  NAND2_X1 U16931 ( .A1(n13618), .A2(n19042), .ZN(n13628) );
  AOI22_X1 U16932 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n19049), .ZN(n13619) );
  OAI211_X1 U16933 ( .C1(n19030), .C2(n13620), .A(n13619), .B(n18941), .ZN(
        n13625) );
  AND2_X1 U16934 ( .A1(n13670), .A2(n13669), .ZN(n13672) );
  OR2_X1 U16935 ( .A1(n13672), .A2(n13621), .ZN(n13623) );
  NAND2_X1 U16936 ( .A1(n13623), .A2(n13622), .ZN(n16224) );
  NOR2_X1 U16937 ( .A1(n16224), .A2(n19057), .ZN(n13624) );
  AOI211_X1 U16938 ( .C1(n12367), .C2(n13626), .A(n13625), .B(n13624), .ZN(
        n13627) );
  OAI211_X1 U16939 ( .C1(n19046), .C2(n19094), .A(n13628), .B(n13627), .ZN(
        P2_U2845) );
  OR2_X1 U16940 ( .A1(n13631), .A2(n13630), .ZN(n13632) );
  AND2_X1 U16941 ( .A1(n13629), .A2(n13632), .ZN(n19942) );
  INV_X1 U16942 ( .A(n19942), .ZN(n13636) );
  NAND2_X1 U16943 ( .A1(n20030), .A2(DATAI_5_), .ZN(n13634) );
  NAND2_X1 U16944 ( .A1(n20032), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13633) );
  AND2_X1 U16945 ( .A1(n13634), .A2(n13633), .ZN(n20075) );
  OAI222_X1 U16946 ( .A1(n13636), .A2(n14622), .B1(n14617), .B2(n20075), .C1(
        n14614), .C2(n13635), .ZN(P1_U2899) );
  INV_X1 U16947 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13639) );
  INV_X1 U16948 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13638) );
  INV_X1 U16949 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n13637) );
  OAI222_X1 U16950 ( .A1(n13639), .A2(n13739), .B1(n13769), .B2(n13638), .C1(
        n13637), .C2(n13766), .ZN(P1_U2914) );
  INV_X1 U16951 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13642) );
  INV_X1 U16952 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13641) );
  INV_X1 U16953 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n13640) );
  OAI222_X1 U16954 ( .A1(n13642), .A2(n13739), .B1(n13769), .B2(n13641), .C1(
        n13640), .C2(n13766), .ZN(P1_U2913) );
  INV_X1 U16955 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13644) );
  INV_X1 U16956 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14096) );
  INV_X1 U16957 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n13643) );
  OAI222_X1 U16958 ( .A1(n13644), .A2(n13739), .B1(n13769), .B2(n14096), .C1(
        n13643), .C2(n13766), .ZN(P1_U2912) );
  INV_X1 U16959 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13646) );
  INV_X1 U16960 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14093) );
  INV_X1 U16961 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n13645) );
  OAI222_X1 U16962 ( .A1(n13646), .A2(n13739), .B1(n13769), .B2(n14093), .C1(
        n13645), .C2(n13766), .ZN(P1_U2911) );
  INV_X1 U16963 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13648) );
  INV_X1 U16964 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14089) );
  INV_X1 U16965 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n13647) );
  OAI222_X1 U16966 ( .A1(n13648), .A2(n13739), .B1(n13769), .B2(n14089), .C1(
        n13647), .C2(n13766), .ZN(P1_U2908) );
  INV_X1 U16967 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13651) );
  INV_X1 U16968 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n13649) );
  OAI222_X1 U16969 ( .A1(n13651), .A2(n13739), .B1(n13772), .B2(n13650), .C1(
        n13766), .C2(n13649), .ZN(P1_U2934) );
  INV_X1 U16970 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13653) );
  INV_X1 U16971 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14100) );
  INV_X1 U16972 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n13652) );
  OAI222_X1 U16973 ( .A1(n13653), .A2(n13739), .B1(n13769), .B2(n14100), .C1(
        n13652), .C2(n13766), .ZN(P1_U2909) );
  INV_X1 U16974 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13655) );
  INV_X1 U16975 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14107) );
  INV_X1 U16976 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n13654) );
  OAI222_X1 U16977 ( .A1(n13655), .A2(n13739), .B1(n13772), .B2(n14107), .C1(
        n13654), .C2(n13766), .ZN(P1_U2926) );
  INV_X1 U16978 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13657) );
  INV_X1 U16979 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14102) );
  INV_X1 U16980 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n13656) );
  OAI222_X1 U16981 ( .A1(n13657), .A2(n13739), .B1(n13769), .B2(n14102), .C1(
        n13656), .C2(n13766), .ZN(P1_U2910) );
  INV_X1 U16982 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13659) );
  INV_X1 U16983 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14610) );
  INV_X1 U16984 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13658) );
  OAI222_X1 U16985 ( .A1(n13659), .A2(n13766), .B1(n13772), .B2(n14610), .C1(
        n13658), .C2(n13739), .ZN(P1_U2921) );
  NOR2_X1 U16986 ( .A1(n15123), .A2(n13660), .ZN(n13665) );
  NOR2_X1 U16987 ( .A1(n13833), .A2(n13661), .ZN(n13836) );
  AOI211_X1 U16988 ( .C1(n13663), .C2(n13662), .A(n15130), .B(n13836), .ZN(
        n13664) );
  AOI211_X1 U16989 ( .C1(n15528), .C2(n15123), .A(n13665), .B(n13664), .ZN(
        n13666) );
  INV_X1 U16990 ( .A(n13666), .ZN(P2_U2874) );
  NAND2_X1 U16991 ( .A1(n13667), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13720) );
  NOR2_X1 U16992 ( .A1(n13720), .A2(n13668), .ZN(n13775) );
  XNOR2_X1 U16993 ( .A(n13775), .B(n13774), .ZN(n13674) );
  NOR2_X1 U16994 ( .A1(n13670), .A2(n13669), .ZN(n13671) );
  OR2_X1 U16995 ( .A1(n13672), .A2(n13671), .ZN(n19002) );
  MUX2_X1 U16996 ( .A(n19002), .B(n10367), .S(n13579), .Z(n13673) );
  OAI21_X1 U16997 ( .B1(n13674), .B2(n15130), .A(n13673), .ZN(P2_U2878) );
  NOR2_X1 U16998 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20634), .ZN(n13700) );
  MUX2_X1 U16999 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13675), .S(
        n15854), .Z(n15859) );
  AOI22_X1 U17000 ( .A1(n13700), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15859), .B2(n20634), .ZN(n13693) );
  NAND2_X1 U17001 ( .A1(n20319), .A2(n14965), .ZN(n13689) );
  XNOR2_X1 U17002 ( .A(n13676), .B(n9759), .ZN(n13677) );
  NAND2_X1 U17003 ( .A1(n13678), .A2(n13677), .ZN(n13687) );
  NAND2_X1 U17004 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U17005 ( .A1(n13680), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n9759), .B2(n13679), .ZN(n13684) );
  OAI21_X1 U17006 ( .B1(n13682), .B2(n9759), .A(n9617), .ZN(n20723) );
  AOI22_X1 U17007 ( .A1(n13685), .A2(n13684), .B1(n13683), .B2(n20723), .ZN(
        n13686) );
  AND2_X1 U17008 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  NAND2_X1 U17009 ( .A1(n13689), .A2(n13688), .ZN(n20725) );
  NAND2_X1 U17010 ( .A1(n20725), .A2(n15854), .ZN(n13691) );
  OR2_X1 U17011 ( .A1(n15854), .A2(n9759), .ZN(n13690) );
  NAND2_X1 U17012 ( .A1(n13691), .A2(n13690), .ZN(n15860) );
  AOI22_X1 U17013 ( .A1(n15860), .A2(n20634), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13700), .ZN(n13692) );
  INV_X1 U17014 ( .A(n20197), .ZN(n20447) );
  NOR2_X1 U17015 ( .A1(n13695), .A2(n20447), .ZN(n13696) );
  XNOR2_X1 U17016 ( .A(n13696), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19950) );
  INV_X1 U17017 ( .A(n13697), .ZN(n13698) );
  NOR2_X1 U17018 ( .A1(n19950), .A2(n13698), .ZN(n16140) );
  MUX2_X1 U17019 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n16140), .S(
        n15854), .Z(n13699) );
  AOI22_X1 U17020 ( .A1(n13700), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n13699), .B2(n20634), .ZN(n15870) );
  OAI21_X1 U17021 ( .B1(n15864), .B2(n13694), .A(n15870), .ZN(n13716) );
  OAI21_X1 U17022 ( .B1(n13716), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13701), .ZN(
        n13702) );
  AND2_X1 U17023 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20451), .ZN(n14960) );
  NOR2_X1 U17024 ( .A1(n20448), .A2(n14960), .ZN(n13706) );
  AOI21_X1 U17025 ( .B1(n9631), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20574), 
        .ZN(n20415) );
  NOR3_X1 U17026 ( .A1(n20318), .A2(n20496), .A3(n20574), .ZN(n20579) );
  MUX2_X1 U17027 ( .A(n20415), .B(n20579), .S(n20034), .Z(n13705) );
  OAI21_X1 U17028 ( .B1(n13706), .B2(n13705), .A(n20028), .ZN(n13707) );
  OAI21_X1 U17029 ( .B1(n20028), .B2(n20320), .A(n13707), .ZN(P1_U3476) );
  INV_X1 U17030 ( .A(n20034), .ZN(n13708) );
  INV_X1 U17031 ( .A(n13709), .ZN(n13710) );
  NOR4_X1 U17032 ( .A1(n20413), .A2(n20492), .A3(n20287), .A4(n20496), .ZN(
        n13711) );
  AOI211_X1 U17033 ( .C1(n20035), .C2(n20496), .A(n20574), .B(n13711), .ZN(
        n13714) );
  INV_X1 U17034 ( .A(n20319), .ZN(n13712) );
  NOR2_X1 U17035 ( .A1(n13712), .A2(n14960), .ZN(n13713) );
  OAI21_X1 U17036 ( .B1(n13714), .B2(n13713), .A(n20028), .ZN(n13715) );
  OAI21_X1 U17037 ( .B1(n20125), .B2(n20028), .A(n13715), .ZN(P1_U3475) );
  NOR2_X1 U17038 ( .A1(n13716), .A2(n16152), .ZN(n15882) );
  INV_X1 U17039 ( .A(n20160), .ZN(n13717) );
  OAI22_X1 U17040 ( .A1(n9632), .A2(n20574), .B1(n13717), .B2(n14960), .ZN(
        n13718) );
  OAI21_X1 U17041 ( .B1(n15882), .B2(n13718), .A(n20028), .ZN(n13719) );
  OAI21_X1 U17042 ( .B1(n20028), .B2(n20493), .A(n13719), .ZN(P1_U3478) );
  INV_X1 U17043 ( .A(n13720), .ZN(n13723) );
  INV_X1 U17044 ( .A(n13775), .ZN(n13721) );
  OAI211_X1 U17045 ( .C1(n13723), .C2(n13722), .A(n13721), .B(n15118), .ZN(
        n13725) );
  NAND2_X1 U17046 ( .A1(n13579), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13724) );
  OAI211_X1 U17047 ( .C1(n16309), .C2(n13579), .A(n13725), .B(n13724), .ZN(
        P2_U2879) );
  OAI21_X4 U17048 ( .B1(n13728), .B2(n19870), .A(n13727), .ZN(n14535) );
  NAND2_X2 U17049 ( .A1(n14535), .A2(n14389), .ZN(n19967) );
  XNOR2_X1 U17050 ( .A(n13852), .B(n13729), .ZN(n14950) );
  OAI22_X1 U17051 ( .A1(n19967), .A2(n14950), .B1(n13730), .B2(n14535), .ZN(
        n13731) );
  INV_X1 U17052 ( .A(n13731), .ZN(n13732) );
  OAI21_X1 U17053 ( .B1(n13861), .B2(n14550), .A(n13732), .ZN(P1_U2871) );
  NAND2_X1 U17054 ( .A1(n13736), .A2(n13733), .ZN(n13734) );
  NAND2_X1 U17055 ( .A1(n13870), .A2(n13734), .ZN(n19994) );
  OAI222_X1 U17056 ( .A1(n19994), .A2(n19967), .B1(n14535), .B2(n12191), .C1(
        n14550), .C2(n13735), .ZN(P1_U2868) );
  OAI21_X1 U17057 ( .B1(n13865), .B2(n9654), .A(n13736), .ZN(n20000) );
  INV_X1 U17058 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13825) );
  OAI222_X1 U17059 ( .A1(n20000), .A2(n19967), .B1(n14535), .B2(n13825), .C1(
        n14550), .C2(n13831), .ZN(P1_U2869) );
  INV_X1 U17060 ( .A(n13737), .ZN(n14459) );
  OAI222_X1 U17061 ( .A1(n14459), .A2(n19967), .B1(n14535), .B2(n13738), .C1(
        n14464), .C2(n14550), .ZN(P1_U2872) );
  INV_X1 U17062 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13741) );
  INV_X1 U17063 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13740) );
  INV_X1 U17064 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n13929) );
  OAI222_X1 U17065 ( .A1(n13741), .A2(n13739), .B1(n13769), .B2(n13740), .C1(
        n13929), .C2(n13766), .ZN(P1_U2920) );
  INV_X1 U17066 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n13743) );
  INV_X1 U17067 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14110) );
  INV_X1 U17068 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n13742) );
  OAI222_X1 U17069 ( .A1(n13743), .A2(n13739), .B1(n13772), .B2(n14110), .C1(
        n13742), .C2(n13766), .ZN(P1_U2925) );
  INV_X1 U17070 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13745) );
  INV_X1 U17071 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n13744) );
  OAI222_X1 U17072 ( .A1(n13745), .A2(n13739), .B1(n13772), .B2(n14147), .C1(
        n13744), .C2(n13766), .ZN(P1_U2924) );
  INV_X1 U17073 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13748) );
  INV_X1 U17074 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13747) );
  INV_X1 U17075 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n13746) );
  OAI222_X1 U17076 ( .A1(n13748), .A2(n13739), .B1(n13769), .B2(n13747), .C1(
        n13746), .C2(n13766), .ZN(P1_U2915) );
  INV_X1 U17077 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n13750) );
  INV_X1 U17078 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n13749) );
  OAI222_X1 U17079 ( .A1(n13750), .A2(n13739), .B1(n13772), .B2(n14615), .C1(
        n13749), .C2(n13766), .ZN(P1_U2923) );
  INV_X1 U17080 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n13752) );
  INV_X1 U17081 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14077) );
  INV_X1 U17082 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n13751) );
  OAI222_X1 U17083 ( .A1(n13752), .A2(n13739), .B1(n13772), .B2(n14077), .C1(
        n13751), .C2(n13766), .ZN(P1_U2922) );
  INV_X1 U17084 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13755) );
  INV_X1 U17085 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13754) );
  INV_X1 U17086 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n13753) );
  OAI222_X1 U17087 ( .A1(n13755), .A2(n13739), .B1(n13769), .B2(n13754), .C1(
        n13753), .C2(n13766), .ZN(P1_U2916) );
  INV_X1 U17088 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13757) );
  INV_X1 U17089 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n13756) );
  OAI222_X1 U17090 ( .A1(n13757), .A2(n13739), .B1(n13769), .B2(n11959), .C1(
        n13756), .C2(n13766), .ZN(P1_U2918) );
  INV_X1 U17091 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13760) );
  INV_X1 U17092 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13759) );
  INV_X1 U17093 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n13758) );
  OAI222_X1 U17094 ( .A1(n13760), .A2(n13739), .B1(n13769), .B2(n13759), .C1(
        n13758), .C2(n13766), .ZN(P1_U2917) );
  INV_X1 U17095 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13763) );
  INV_X1 U17096 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n13761) );
  OAI222_X1 U17097 ( .A1(n13763), .A2(n13739), .B1(n13772), .B2(n13762), .C1(
        n13766), .C2(n13761), .ZN(P1_U2936) );
  INV_X1 U17098 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13765) );
  INV_X1 U17099 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14091) );
  INV_X1 U17100 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n13764) );
  OAI222_X1 U17101 ( .A1(n13765), .A2(n13739), .B1(n13772), .B2(n14091), .C1(
        n13764), .C2(n13766), .ZN(P1_U2928) );
  INV_X1 U17102 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13770) );
  INV_X1 U17103 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13768) );
  INV_X1 U17104 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n13767) );
  OAI222_X1 U17105 ( .A1(n13770), .A2(n13739), .B1(n13769), .B2(n13768), .C1(
        n13767), .C2(n13766), .ZN(P1_U2919) );
  INV_X1 U17106 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n13773) );
  INV_X1 U17107 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n13771) );
  OAI222_X1 U17108 ( .A1(n13773), .A2(n13739), .B1(n13772), .B2(n14024), .C1(
        n13771), .C2(n13766), .ZN(P1_U2927) );
  INV_X1 U17109 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13781) );
  AND2_X1 U17110 ( .A1(n13775), .A2(n13774), .ZN(n13778) );
  OAI211_X1 U17111 ( .C1(n13778), .C2(n13777), .A(n15118), .B(n13776), .ZN(
        n13780) );
  INV_X1 U17112 ( .A(n16224), .ZN(n16293) );
  NAND2_X1 U17113 ( .A1(n16293), .A2(n15123), .ZN(n13779) );
  OAI211_X1 U17114 ( .C1(n15123), .C2(n13781), .A(n13780), .B(n13779), .ZN(
        P2_U2877) );
  AND2_X1 U17115 ( .A1(n16344), .A2(n13782), .ZN(n15671) );
  NOR2_X1 U17116 ( .A1(n10143), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15674) );
  NOR2_X1 U17117 ( .A1(n15674), .A2(n20914), .ZN(n13788) );
  INV_X1 U17118 ( .A(n15651), .ZN(n15683) );
  NAND2_X1 U17119 ( .A1(n9595), .A2(n15683), .ZN(n13787) );
  NAND2_X1 U17120 ( .A1(n13784), .A2(n13783), .ZN(n15673) );
  AOI22_X1 U17121 ( .A1(n15673), .A2(n13788), .B1(n13785), .B2(n15676), .ZN(
        n13786) );
  OAI211_X1 U17122 ( .C1(n15671), .C2(n13788), .A(n13787), .B(n13786), .ZN(
        n16333) );
  AOI221_X1 U17123 ( .B1(n13791), .B2(n12347), .C1(n13790), .C2(n12329), .A(
        n13789), .ZN(n15660) );
  OAI21_X1 U17124 ( .B1(n12347), .B2(n15642), .A(n13792), .ZN(n15666) );
  AOI222_X1 U17125 ( .A1(n16333), .A2(n19799), .B1(n15660), .B2(n15666), .C1(
        n16371), .C2(n19810), .ZN(n13793) );
  MUX2_X1 U17126 ( .A(n13794), .B(n13793), .S(n15685), .Z(n13795) );
  INV_X1 U17127 ( .A(n13795), .ZN(P2_U3599) );
  NOR2_X1 U17128 ( .A1(n9679), .A2(n13796), .ZN(n13797) );
  OR2_X1 U17129 ( .A1(n9680), .A2(n13797), .ZN(n19920) );
  AOI21_X1 U17130 ( .B1(n13799), .B2(n13629), .A(n11586), .ZN(n13925) );
  INV_X1 U17131 ( .A(n13925), .ZN(n19925) );
  OAI222_X1 U17132 ( .A1(n19920), .A2(n19967), .B1(n14535), .B2(n12202), .C1(
        n14550), .C2(n19925), .ZN(P1_U2866) );
  INV_X1 U17133 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16479) );
  NAND2_X1 U17134 ( .A1(n20032), .A2(n16479), .ZN(n13800) );
  OAI21_X1 U17135 ( .B1(n20032), .B2(DATAI_6_), .A(n13800), .ZN(n20080) );
  OAI222_X1 U17136 ( .A1(n14617), .A2(n20080), .B1(n14614), .B2(n11575), .C1(
        n14622), .C2(n19925), .ZN(P1_U2898) );
  XNOR2_X1 U17137 ( .A(n13801), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13802) );
  XNOR2_X1 U17138 ( .A(n13803), .B(n13802), .ZN(n16263) );
  INV_X1 U17139 ( .A(n16263), .ZN(n13814) );
  OAI22_X1 U17140 ( .A1(n16261), .A2(n16319), .B1(n10081), .B2(n18941), .ZN(
        n13808) );
  NAND2_X1 U17141 ( .A1(n13806), .A2(n16322), .ZN(n13804) );
  OAI22_X1 U17142 ( .A1(n13945), .A2(n13806), .B1(n13805), .B2(n13804), .ZN(
        n13807) );
  AOI211_X1 U17143 ( .C1(n16307), .C2(n19805), .A(n13808), .B(n13807), .ZN(
        n13813) );
  OR2_X1 U17144 ( .A1(n13810), .A2(n13809), .ZN(n16259) );
  NAND3_X1 U17145 ( .A1(n16259), .A2(n16295), .A3(n13811), .ZN(n13812) );
  OAI211_X1 U17146 ( .C1(n13814), .C2(n16299), .A(n13813), .B(n13812), .ZN(
        P2_U3043) );
  NAND2_X1 U17147 ( .A1(n20739), .A2(n13815), .ZN(n13816) );
  NAND2_X1 U17148 ( .A1(n19924), .A2(n13816), .ZN(n19958) );
  INV_X1 U17149 ( .A(n19958), .ZN(n14463) );
  NOR2_X1 U17150 ( .A1(n13818), .A2(n13817), .ZN(n14461) );
  INV_X1 U17151 ( .A(n19955), .ZN(n15986) );
  OAI221_X1 U17152 ( .B1(n14363), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n14363), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14357), .ZN(n13819) );
  AOI22_X1 U17153 ( .A1(n19953), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13819), .ZN(n13824) );
  AND2_X1 U17154 ( .A1(n14304), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13820) );
  AND2_X1 U17155 ( .A1(n14357), .A2(n13820), .ZN(n19909) );
  INV_X1 U17156 ( .A(n13821), .ZN(n13822) );
  NAND2_X1 U17157 ( .A1(n19909), .A2(n13822), .ZN(n13823) );
  OAI211_X1 U17158 ( .C1(n15986), .C2(n13825), .A(n13824), .B(n13823), .ZN(
        n13829) );
  INV_X1 U17159 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13826) );
  NAND4_X1 U17160 ( .A1(n19957), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n13826), .ZN(n13827) );
  OAI21_X1 U17161 ( .B1(n19948), .B2(n20000), .A(n13827), .ZN(n13828) );
  AOI211_X1 U17162 ( .C1(n20319), .C2(n14461), .A(n13829), .B(n13828), .ZN(
        n13830) );
  OAI21_X1 U17163 ( .B1(n13831), .B2(n14463), .A(n13830), .ZN(P1_U2837) );
  NOR2_X1 U17164 ( .A1(n13833), .A2(n13832), .ZN(n13878) );
  INV_X1 U17165 ( .A(n13878), .ZN(n13834) );
  OAI211_X1 U17166 ( .C1(n13836), .C2(n13835), .A(n13834), .B(n15118), .ZN(
        n13841) );
  INV_X1 U17167 ( .A(n13837), .ZN(n13839) );
  INV_X1 U17168 ( .A(n13087), .ZN(n13838) );
  AOI21_X1 U17169 ( .B1(n13839), .B2(n13838), .A(n13880), .ZN(n16277) );
  NAND2_X1 U17170 ( .A1(n16277), .A2(n15123), .ZN(n13840) );
  OAI211_X1 U17171 ( .C1(n15123), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        P2_U2873) );
  OAI21_X1 U17172 ( .B1(n13882), .B2(n13843), .A(n13987), .ZN(n15514) );
  AND2_X1 U17173 ( .A1(n13845), .A2(n13844), .ZN(n13875) );
  OR2_X1 U17174 ( .A1(n13875), .A2(n13846), .ZN(n13848) );
  NAND2_X1 U17175 ( .A1(n13396), .A2(n13847), .ZN(n13991) );
  AND2_X1 U17176 ( .A1(n13848), .A2(n13991), .ZN(n19075) );
  NAND2_X1 U17177 ( .A1(n19075), .A2(n15118), .ZN(n13850) );
  NAND2_X1 U17178 ( .A1(n13579), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13849) );
  OAI211_X1 U17179 ( .C1(n15514), .C2(n13579), .A(n13850), .B(n13849), .ZN(
        P2_U2871) );
  INV_X1 U17180 ( .A(n14461), .ZN(n19949) );
  INV_X1 U17181 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20729) );
  AOI22_X1 U17182 ( .A1(n19957), .A2(n20729), .B1(n19936), .B2(n13852), .ZN(
        n13858) );
  NAND2_X1 U17183 ( .A1(n19909), .A2(n13853), .ZN(n13855) );
  NAND2_X1 U17184 ( .A1(n19953), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13854) );
  OAI211_X1 U17185 ( .C1(n20729), .C2(n14357), .A(n13855), .B(n13854), .ZN(
        n13856) );
  AOI21_X1 U17186 ( .B1(n19955), .B2(P1_EBX_REG_1__SCAN_IN), .A(n13856), .ZN(
        n13857) );
  OAI211_X1 U17187 ( .C1(n20449), .C2(n19949), .A(n13858), .B(n13857), .ZN(
        n13859) );
  INV_X1 U17188 ( .A(n13859), .ZN(n13860) );
  OAI21_X1 U17189 ( .B1(n13861), .B2(n14463), .A(n13860), .ZN(P1_U2839) );
  INV_X1 U17190 ( .A(n14550), .ZN(n16023) );
  NOR2_X1 U17191 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  OR2_X1 U17192 ( .A1(n13865), .A2(n13864), .ZN(n14362) );
  OAI22_X1 U17193 ( .A1(n14362), .A2(n19967), .B1(n13866), .B2(n14535), .ZN(
        n13867) );
  AOI21_X1 U17194 ( .B1(n14356), .B2(n16023), .A(n13867), .ZN(n13868) );
  INV_X1 U17195 ( .A(n13868), .ZN(P1_U2870) );
  NAND2_X1 U17196 ( .A1(n19942), .A2(n16023), .ZN(n13873) );
  AND2_X1 U17197 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  NOR2_X1 U17198 ( .A1(n9679), .A2(n13871), .ZN(n19937) );
  NAND2_X1 U17199 ( .A1(n19937), .A2(n16021), .ZN(n13872) );
  OAI211_X1 U17200 ( .C1(n13874), .C2(n14535), .A(n13873), .B(n13872), .ZN(
        P1_U2867) );
  INV_X1 U17201 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18965) );
  INV_X1 U17202 ( .A(n13875), .ZN(n13876) );
  OAI211_X1 U17203 ( .C1(n13878), .C2(n13877), .A(n13876), .B(n15118), .ZN(
        n13884) );
  NOR2_X1 U17204 ( .A1(n13880), .A2(n13879), .ZN(n13881) );
  OR2_X1 U17205 ( .A1(n13882), .A2(n13881), .ZN(n15327) );
  NAND2_X1 U17206 ( .A1(n18972), .A2(n15123), .ZN(n13883) );
  OAI211_X1 U17207 ( .C1(n15123), .C2(n18965), .A(n13884), .B(n13883), .ZN(
        P2_U2872) );
  NAND2_X1 U17208 ( .A1(n13798), .A2(n13885), .ZN(n13886) );
  AND2_X1 U17209 ( .A1(n13968), .A2(n13886), .ZN(n19903) );
  INV_X1 U17210 ( .A(n19903), .ZN(n13890) );
  NAND2_X1 U17211 ( .A1(n20030), .A2(DATAI_7_), .ZN(n13888) );
  NAND2_X1 U17212 ( .A1(n20032), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13887) );
  AND2_X1 U17213 ( .A1(n13888), .A2(n13887), .ZN(n20087) );
  OAI222_X1 U17214 ( .A1(n13890), .A2(n14622), .B1(n14617), .B2(n20087), .C1(
        n14614), .C2(n11582), .ZN(P1_U2897) );
  OAI21_X1 U17215 ( .B1(n9680), .B2(n13889), .A(n13975), .ZN(n16127) );
  OAI222_X1 U17216 ( .A1(n16127), .A2(n19967), .B1(n13891), .B2(n14535), .C1(
        n14550), .C2(n13890), .ZN(P1_U2865) );
  INV_X1 U17217 ( .A(n20741), .ZN(n15899) );
  AND2_X1 U17218 ( .A1(n20744), .A2(n15899), .ZN(n13892) );
  OR2_X2 U17219 ( .A1(n13893), .A2(n13892), .ZN(n13894) );
  NOR2_X2 U17220 ( .A1(n13894), .A2(n20054), .ZN(n14071) );
  AOI22_X1 U17221 ( .A1(n14071), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n13894), .ZN(n13895) );
  NOR2_X2 U17222 ( .A1(n13894), .A2(n11495), .ZN(n14111) );
  INV_X1 U17223 ( .A(n20075), .ZN(n14586) );
  NAND2_X1 U17224 ( .A1(n14111), .A2(n14586), .ZN(n13905) );
  NAND2_X1 U17225 ( .A1(n13895), .A2(n13905), .ZN(P1_U2942) );
  AOI22_X1 U17226 ( .A1(n14071), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n13894), .ZN(n13896) );
  INV_X1 U17227 ( .A(n20066), .ZN(n14592) );
  NAND2_X1 U17228 ( .A1(n14111), .A2(n14592), .ZN(n13902) );
  NAND2_X1 U17229 ( .A1(n13896), .A2(n13902), .ZN(P1_U2940) );
  AOI22_X1 U17230 ( .A1(n14071), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n13894), .ZN(n13898) );
  INV_X1 U17231 ( .A(n20087), .ZN(n13897) );
  NAND2_X1 U17232 ( .A1(n14111), .A2(n13897), .ZN(n13908) );
  NAND2_X1 U17233 ( .A1(n13898), .A2(n13908), .ZN(P1_U2944) );
  AOI22_X1 U17234 ( .A1(n14071), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n13894), .ZN(n13899) );
  INV_X1 U17235 ( .A(n20048), .ZN(n14605) );
  NAND2_X1 U17236 ( .A1(n14111), .A2(n14605), .ZN(n13928) );
  NAND2_X1 U17237 ( .A1(n13899), .A2(n13928), .ZN(P1_U2952) );
  AOI22_X1 U17238 ( .A1(n14071), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13894), .ZN(n13900) );
  INV_X1 U17239 ( .A(n20056), .ZN(n14599) );
  NAND2_X1 U17240 ( .A1(n14111), .A2(n14599), .ZN(n13912) );
  NAND2_X1 U17241 ( .A1(n13900), .A2(n13912), .ZN(P1_U2953) );
  AOI22_X1 U17242 ( .A1(n14071), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n13894), .ZN(n13901) );
  INV_X1 U17243 ( .A(n20061), .ZN(n14596) );
  NAND2_X1 U17244 ( .A1(n14111), .A2(n14596), .ZN(n13914) );
  NAND2_X1 U17245 ( .A1(n13901), .A2(n13914), .ZN(P1_U2954) );
  AOI22_X1 U17246 ( .A1(n14071), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n13894), .ZN(n13903) );
  NAND2_X1 U17247 ( .A1(n13903), .A2(n13902), .ZN(P1_U2955) );
  AOI22_X1 U17248 ( .A1(n14071), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n13894), .ZN(n13904) );
  INV_X1 U17249 ( .A(n20070), .ZN(n14589) );
  NAND2_X1 U17250 ( .A1(n14111), .A2(n14589), .ZN(n13910) );
  NAND2_X1 U17251 ( .A1(n13904), .A2(n13910), .ZN(P1_U2956) );
  AOI22_X1 U17252 ( .A1(n14071), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13894), .ZN(n13906) );
  NAND2_X1 U17253 ( .A1(n13906), .A2(n13905), .ZN(P1_U2957) );
  AOI22_X1 U17254 ( .A1(n14071), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n13894), .ZN(n13907) );
  INV_X1 U17255 ( .A(n20080), .ZN(n14582) );
  NAND2_X1 U17256 ( .A1(n14111), .A2(n14582), .ZN(n13916) );
  NAND2_X1 U17257 ( .A1(n13907), .A2(n13916), .ZN(P1_U2958) );
  AOI22_X1 U17258 ( .A1(n14071), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n13894), .ZN(n13909) );
  NAND2_X1 U17259 ( .A1(n13909), .A2(n13908), .ZN(P1_U2959) );
  AOI22_X1 U17260 ( .A1(n14071), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13894), .ZN(n13911) );
  NAND2_X1 U17261 ( .A1(n13911), .A2(n13910), .ZN(P1_U2941) );
  AOI22_X1 U17262 ( .A1(n14071), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n13894), .ZN(n13913) );
  NAND2_X1 U17263 ( .A1(n13913), .A2(n13912), .ZN(P1_U2938) );
  AOI22_X1 U17264 ( .A1(n14071), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n13894), .ZN(n13915) );
  NAND2_X1 U17265 ( .A1(n13915), .A2(n13914), .ZN(P1_U2939) );
  AOI22_X1 U17266 ( .A1(n14071), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n13894), .ZN(n13917) );
  NAND2_X1 U17267 ( .A1(n13917), .A2(n13916), .ZN(P1_U2943) );
  NAND2_X1 U17268 ( .A1(n13918), .A2(n16069), .ZN(n16068) );
  NAND2_X1 U17269 ( .A1(n16068), .A2(n13919), .ZN(n13922) );
  XOR2_X1 U17270 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13920), .Z(
        n13921) );
  XNOR2_X1 U17271 ( .A(n13922), .B(n13921), .ZN(n13940) );
  NAND2_X1 U17272 ( .A1(n19952), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n13930) );
  NAND2_X1 U17273 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13923) );
  OAI211_X1 U17274 ( .C1(n19985), .C2(n19923), .A(n13930), .B(n13923), .ZN(
        n13924) );
  AOI21_X1 U17275 ( .B1(n13925), .B2(n19980), .A(n13924), .ZN(n13926) );
  OAI21_X1 U17276 ( .B1(n13940), .B2(n19877), .A(n13926), .ZN(P1_U2993) );
  NAND2_X1 U17277 ( .A1(n14071), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n13927) );
  OAI211_X1 U17278 ( .C1(n14114), .C2(n13929), .A(n13928), .B(n13927), .ZN(
        P1_U2937) );
  NAND2_X1 U17279 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19991) );
  NOR2_X1 U17280 ( .A1(n16138), .A2(n19991), .ZN(n14935) );
  NOR2_X1 U17281 ( .A1(n20026), .A2(n20012), .ZN(n19987) );
  NAND2_X1 U17282 ( .A1(n14916), .A2(n14914), .ZN(n20011) );
  NAND2_X1 U17283 ( .A1(n14914), .A2(n14309), .ZN(n14955) );
  AOI21_X1 U17284 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20015) );
  INV_X1 U17285 ( .A(n16123), .ZN(n13933) );
  INV_X1 U17286 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13932) );
  OAI21_X1 U17287 ( .B1(n19920), .B2(n19993), .A(n13930), .ZN(n13931) );
  AOI21_X1 U17288 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(n13939) );
  NOR2_X1 U17289 ( .A1(n19991), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16134) );
  INV_X1 U17290 ( .A(n16134), .ZN(n13937) );
  INV_X1 U17291 ( .A(n20011), .ZN(n19988) );
  NOR2_X1 U17292 ( .A1(n14916), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13934) );
  INV_X1 U17293 ( .A(n20010), .ZN(n19986) );
  INV_X1 U17294 ( .A(n20018), .ZN(n19990) );
  INV_X1 U17295 ( .A(n20015), .ZN(n13935) );
  NAND2_X1 U17296 ( .A1(n14935), .A2(n13935), .ZN(n16098) );
  NAND2_X1 U17297 ( .A1(n19990), .A2(n16098), .ZN(n13936) );
  OAI211_X1 U17298 ( .C1(n19988), .C2(n19987), .A(n19986), .B(n13936), .ZN(
        n16097) );
  AOI21_X1 U17299 ( .B1(n20011), .B2(n19991), .A(n16097), .ZN(n16139) );
  OAI21_X1 U17300 ( .B1(n14936), .B2(n13937), .A(n16139), .ZN(n16117) );
  NAND2_X1 U17301 ( .A1(n16117), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13938) );
  OAI211_X1 U17302 ( .C1(n13940), .C2(n16120), .A(n13939), .B(n13938), .ZN(
        P1_U3025) );
  XNOR2_X1 U17303 ( .A(n13941), .B(n15630), .ZN(n19179) );
  INV_X1 U17304 ( .A(n19179), .ZN(n13953) );
  INV_X1 U17305 ( .A(n13943), .ZN(n13944) );
  XNOR2_X1 U17306 ( .A(n13942), .B(n13944), .ZN(n19181) );
  NAND2_X1 U17307 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15602), .ZN(
        n15629) );
  OAI21_X1 U17308 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14342), .A(
        n13945), .ZN(n15634) );
  NOR2_X1 U17309 ( .A1(n10755), .A2(n10856), .ZN(n13946) );
  AOI21_X1 U17310 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15634), .A(
        n13946), .ZN(n13947) );
  OAI21_X1 U17311 ( .B1(n16318), .B2(n15181), .A(n13947), .ZN(n13948) );
  AOI21_X1 U17312 ( .B1(n13949), .B2(n16294), .A(n13948), .ZN(n13950) );
  OAI21_X1 U17313 ( .B1(n15629), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13950), .ZN(n13951) );
  AOI21_X1 U17314 ( .B1(n19181), .B2(n16326), .A(n13951), .ZN(n13952) );
  OAI21_X1 U17315 ( .B1(n13953), .B2(n16330), .A(n13952), .ZN(P2_U3042) );
  INV_X1 U17316 ( .A(n13954), .ZN(n13966) );
  NOR2_X1 U17317 ( .A1(n12329), .A2(n13955), .ZN(n13956) );
  XNOR2_X1 U17318 ( .A(n13956), .B(n16205), .ZN(n13957) );
  NAND2_X1 U17319 ( .A1(n13957), .A2(n19042), .ZN(n13965) );
  AOI21_X1 U17320 ( .B1(n13958), .B2(n13089), .A(n9643), .ZN(n19081) );
  AOI22_X1 U17321 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19049), .ZN(n13959) );
  OAI211_X1 U17322 ( .C1(n19030), .C2(n13960), .A(n13959), .B(n18941), .ZN(
        n13963) );
  INV_X1 U17323 ( .A(n16277), .ZN(n13961) );
  NOR2_X1 U17324 ( .A1(n13961), .A2(n19057), .ZN(n13962) );
  AOI211_X1 U17325 ( .C1(n19055), .C2(n19081), .A(n13963), .B(n13962), .ZN(
        n13964) );
  OAI211_X1 U17326 ( .C1(n19052), .C2(n13966), .A(n13965), .B(n13964), .ZN(
        P2_U2841) );
  AOI21_X1 U17327 ( .B1(n13969), .B2(n13968), .A(n13967), .ZN(n14002) );
  INV_X1 U17328 ( .A(n14002), .ZN(n13984) );
  INV_X1 U17329 ( .A(n14617), .ZN(n14620) );
  INV_X1 U17330 ( .A(DATAI_8_), .ZN(n13971) );
  NAND2_X1 U17331 ( .A1(n20032), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13970) );
  OAI21_X1 U17332 ( .B1(n20032), .B2(n13971), .A(n13970), .ZN(n14571) );
  AOI22_X1 U17333 ( .A1(n14620), .A2(n14571), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14618), .ZN(n13972) );
  OAI21_X1 U17334 ( .B1(n13984), .B2(n14622), .A(n13972), .ZN(P1_U2896) );
  INV_X1 U17335 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13973) );
  OAI22_X1 U17336 ( .A1(n14000), .A2(n19965), .B1(n19919), .B2(n13973), .ZN(
        n13980) );
  INV_X1 U17337 ( .A(n19973), .ZN(n19933) );
  INV_X1 U17338 ( .A(n19933), .ZN(n19952) );
  NAND2_X1 U17339 ( .A1(n13975), .A2(n13974), .ZN(n13976) );
  NAND2_X1 U17340 ( .A1(n16106), .A2(n13976), .ZN(n16121) );
  AND2_X1 U17341 ( .A1(n19932), .A2(n13977), .ZN(n19898) );
  AOI22_X1 U17342 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(n19955), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n19898), .ZN(n13978) );
  OAI21_X1 U17343 ( .B1(n19948), .B2(n16121), .A(n13978), .ZN(n13979) );
  NOR3_X1 U17344 ( .A1(n13980), .A2(n19952), .A3(n13979), .ZN(n13983) );
  NOR2_X1 U17345 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19917), .ZN(n13981) );
  NAND2_X1 U17346 ( .A1(n13981), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n13982) );
  OAI211_X1 U17347 ( .C1(n13984), .C2(n19924), .A(n13983), .B(n13982), .ZN(
        P1_U2832) );
  OAI222_X1 U17348 ( .A1(n16121), .A2(n19967), .B1(n14535), .B2(n12212), .C1(
        n14550), .C2(n13984), .ZN(P1_U2864) );
  INV_X1 U17349 ( .A(n13985), .ZN(n13986) );
  AOI21_X1 U17350 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n18945) );
  INV_X1 U17351 ( .A(n18945), .ZN(n13995) );
  NAND2_X1 U17352 ( .A1(n13396), .A2(n13989), .ZN(n14015) );
  INV_X1 U17353 ( .A(n14015), .ZN(n13990) );
  AOI21_X1 U17354 ( .B1(n13992), .B2(n13991), .A(n13990), .ZN(n14011) );
  NAND2_X1 U17355 ( .A1(n14011), .A2(n15118), .ZN(n13994) );
  NAND2_X1 U17356 ( .A1(n13579), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13993) );
  OAI211_X1 U17357 ( .C1(n13995), .C2(n13579), .A(n13994), .B(n13993), .ZN(
        P2_U2870) );
  XNOR2_X1 U17358 ( .A(n13996), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13997) );
  XNOR2_X1 U17359 ( .A(n9612), .B(n13997), .ZN(n16119) );
  AOI22_X1 U17360 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U17361 ( .B1(n14000), .B2(n19985), .A(n13999), .ZN(n14001) );
  AOI21_X1 U17362 ( .B1(n14002), .B2(n19980), .A(n14001), .ZN(n14003) );
  OAI21_X1 U17363 ( .B1(n16119), .B2(n19877), .A(n14003), .ZN(P1_U2991) );
  OR2_X1 U17364 ( .A1(n15512), .A2(n14004), .ZN(n14005) );
  NAND2_X1 U17365 ( .A1(n14027), .A2(n14005), .ZN(n18954) );
  AOI22_X1 U17366 ( .A1(n19073), .A2(BUF1_REG_17__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17367 ( .A1(n19071), .A2(n14007), .B1(n19129), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14008) );
  OAI211_X1 U17368 ( .C1(n16191), .C2(n18954), .A(n14009), .B(n14008), .ZN(
        n14010) );
  AOI21_X1 U17369 ( .B1(n14011), .B2(n19108), .A(n14010), .ZN(n14012) );
  INV_X1 U17370 ( .A(n14012), .ZN(P2_U2902) );
  OR2_X1 U17371 ( .A1(n13985), .A2(n14013), .ZN(n15125) );
  NAND2_X1 U17372 ( .A1(n13985), .A2(n14013), .ZN(n14014) );
  NAND2_X1 U17373 ( .A1(n15125), .A2(n14014), .ZN(n18934) );
  AOI21_X1 U17374 ( .B1(n14016), .B2(n14015), .A(n14049), .ZN(n14032) );
  NAND2_X1 U17375 ( .A1(n14032), .A2(n15118), .ZN(n14018) );
  NAND2_X1 U17376 ( .A1(n13579), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14017) );
  OAI211_X1 U17377 ( .C1(n18934), .C2(n13579), .A(n14018), .B(n14017), .ZN(
        P2_U2869) );
  AND2_X1 U17378 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  OR2_X1 U17379 ( .A1(n14021), .A2(n14035), .ZN(n19969) );
  INV_X1 U17380 ( .A(DATAI_9_), .ZN(n14023) );
  NAND2_X1 U17381 ( .A1(n20032), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14022) );
  OAI21_X1 U17382 ( .B1(n20032), .B2(n14023), .A(n14022), .ZN(n14567) );
  INV_X1 U17383 ( .A(n14567), .ZN(n14025) );
  OAI222_X1 U17384 ( .A1(n19969), .A2(n14622), .B1(n14617), .B2(n14025), .C1(
        n14024), .C2(n14614), .ZN(P1_U2895) );
  XNOR2_X1 U17385 ( .A(n14027), .B(n14026), .ZN(n18939) );
  AOI22_X1 U17386 ( .A1(n19073), .A2(BUF1_REG_18__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17387 ( .A1(n19071), .A2(n14028), .B1(n19129), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n14029) );
  OAI211_X1 U17388 ( .C1(n18939), .C2(n16191), .A(n14030), .B(n14029), .ZN(
        n14031) );
  AOI21_X1 U17389 ( .B1(n14032), .B2(n19108), .A(n14031), .ZN(n14033) );
  INV_X1 U17390 ( .A(n14033), .ZN(P2_U2901) );
  INV_X1 U17391 ( .A(n14034), .ZN(n14037) );
  INV_X1 U17392 ( .A(n14035), .ZN(n14036) );
  AOI21_X1 U17393 ( .B1(n14037), .B2(n14036), .A(n9656), .ZN(n14757) );
  INV_X1 U17394 ( .A(n14757), .ZN(n14041) );
  INV_X1 U17395 ( .A(DATAI_10_), .ZN(n14039) );
  NAND2_X1 U17396 ( .A1(n20032), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14038) );
  OAI21_X1 U17397 ( .B1(n20032), .B2(n14039), .A(n14038), .ZN(n14564) );
  AOI22_X1 U17398 ( .A1(n14620), .A2(n14564), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14618), .ZN(n14040) );
  OAI21_X1 U17399 ( .B1(n14041), .B2(n14622), .A(n14040), .ZN(P1_U2894) );
  AND2_X1 U17400 ( .A1(n16108), .A2(n14042), .ZN(n14043) );
  OR2_X1 U17401 ( .A1(n14043), .A2(n14552), .ZN(n16099) );
  OAI22_X1 U17402 ( .A1(n16099), .A2(n19967), .B1(n14044), .B2(n14535), .ZN(
        n14045) );
  AOI21_X1 U17403 ( .B1(n14757), .B2(n16023), .A(n14045), .ZN(n14046) );
  INV_X1 U17404 ( .A(n14046), .ZN(P1_U2862) );
  INV_X1 U17405 ( .A(n9686), .ZN(n14047) );
  OAI21_X1 U17406 ( .B1(n14049), .B2(n14048), .A(n14047), .ZN(n15131) );
  OR2_X1 U17407 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U17408 ( .A1(n14052), .A2(n9639), .ZN(n18926) );
  AOI22_X1 U17409 ( .A1(n19073), .A2(BUF1_REG_19__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17410 ( .A1(n19071), .A2(n14053), .B1(n19129), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14054) );
  OAI211_X1 U17411 ( .C1(n16191), .C2(n18926), .A(n14055), .B(n14054), .ZN(
        n14056) );
  INV_X1 U17412 ( .A(n14056), .ZN(n14057) );
  OAI21_X1 U17413 ( .B1(n15131), .B2(n19134), .A(n14057), .ZN(P2_U2900) );
  AOI21_X1 U17414 ( .B1(n19953), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19952), .ZN(n14060) );
  NOR2_X1 U17415 ( .A1(n19905), .A2(n14058), .ZN(n16013) );
  AOI22_X1 U17416 ( .A1(n16013), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n19955), 
        .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n14059) );
  OAI211_X1 U17417 ( .C1(n19948), .C2(n16099), .A(n14060), .B(n14059), .ZN(
        n14063) );
  INV_X1 U17418 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20671) );
  NAND3_X1 U17419 ( .A1(n19899), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n20671), 
        .ZN(n14061) );
  OAI21_X1 U17420 ( .B1(n14755), .B2(n19965), .A(n14061), .ZN(n14062) );
  AOI211_X1 U17421 ( .C1(n14757), .C2(n19902), .A(n14063), .B(n14062), .ZN(
        n14064) );
  INV_X1 U17422 ( .A(n14064), .ZN(P1_U2830) );
  INV_X1 U17423 ( .A(n14066), .ZN(n14067) );
  AOI21_X1 U17424 ( .B1(n14068), .B2(n14065), .A(n14067), .ZN(n14145) );
  NAND2_X1 U17425 ( .A1(n14145), .A2(n15118), .ZN(n14070) );
  NAND2_X1 U17426 ( .A1(n13579), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14069) );
  OAI211_X1 U17427 ( .C1(n14203), .C2(n13579), .A(n14070), .B(n14069), .ZN(
        P2_U2866) );
  NAND2_X1 U17428 ( .A1(n13894), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14073) );
  INV_X1 U17429 ( .A(DATAI_13_), .ZN(n20834) );
  NAND2_X1 U17430 ( .A1(n20032), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14072) );
  OAI21_X1 U17431 ( .B1(n20032), .B2(n20834), .A(n14072), .ZN(n14613) );
  NAND2_X1 U17432 ( .A1(n14111), .A2(n14613), .ZN(n14081) );
  OAI211_X1 U17433 ( .C1(n14116), .C2(n14615), .A(n14073), .B(n14081), .ZN(
        P1_U2965) );
  NAND2_X1 U17434 ( .A1(n13894), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14076) );
  INV_X1 U17435 ( .A(DATAI_14_), .ZN(n14075) );
  NAND2_X1 U17436 ( .A1(n20032), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14074) );
  OAI21_X1 U17437 ( .B1(n20032), .B2(n14075), .A(n14074), .ZN(n14390) );
  NAND2_X1 U17438 ( .A1(n14111), .A2(n14390), .ZN(n14084) );
  OAI211_X1 U17439 ( .C1(n14116), .C2(n14077), .A(n14076), .B(n14084), .ZN(
        P1_U2966) );
  NAND2_X1 U17440 ( .A1(n13894), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14080) );
  INV_X1 U17441 ( .A(DATAI_12_), .ZN(n14079) );
  NAND2_X1 U17442 ( .A1(n20032), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14078) );
  OAI21_X1 U17443 ( .B1(n20032), .B2(n14079), .A(n14078), .ZN(n14559) );
  NAND2_X1 U17444 ( .A1(n14111), .A2(n14559), .ZN(n14087) );
  OAI211_X1 U17445 ( .C1(n14116), .C2(n14147), .A(n14080), .B(n14087), .ZN(
        P1_U2964) );
  NAND2_X1 U17446 ( .A1(n13894), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U17447 ( .C1(n14116), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        P1_U2950) );
  NAND2_X1 U17448 ( .A1(n13894), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14085) );
  OAI211_X1 U17449 ( .C1(n14116), .C2(n14086), .A(n14085), .B(n14084), .ZN(
        P1_U2951) );
  NAND2_X1 U17450 ( .A1(n13894), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14088) );
  OAI211_X1 U17451 ( .C1(n14116), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        P1_U2949) );
  NAND2_X1 U17452 ( .A1(n13894), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U17453 ( .A1(n14111), .A2(n14571), .ZN(n14094) );
  OAI211_X1 U17454 ( .C1(n14116), .C2(n14091), .A(n14090), .B(n14094), .ZN(
        P1_U2960) );
  NAND2_X1 U17455 ( .A1(n13894), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U17456 ( .A1(n14111), .A2(n14567), .ZN(n14103) );
  OAI211_X1 U17457 ( .C1(n14116), .C2(n14093), .A(n14092), .B(n14103), .ZN(
        P1_U2946) );
  NAND2_X1 U17458 ( .A1(n13894), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14095) );
  OAI211_X1 U17459 ( .C1(n14116), .C2(n14096), .A(n14095), .B(n14094), .ZN(
        P1_U2945) );
  NAND2_X1 U17460 ( .A1(n13894), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14099) );
  INV_X1 U17461 ( .A(DATAI_11_), .ZN(n14098) );
  NAND2_X1 U17462 ( .A1(n20032), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14097) );
  OAI21_X1 U17463 ( .B1(n20032), .B2(n14098), .A(n14097), .ZN(n14619) );
  NAND2_X1 U17464 ( .A1(n14111), .A2(n14619), .ZN(n14108) );
  OAI211_X1 U17465 ( .C1(n14116), .C2(n14100), .A(n14099), .B(n14108), .ZN(
        P1_U2948) );
  NAND2_X1 U17466 ( .A1(n13894), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14101) );
  NAND2_X1 U17467 ( .A1(n14111), .A2(n14564), .ZN(n14105) );
  OAI211_X1 U17468 ( .C1(n14116), .C2(n14102), .A(n14101), .B(n14105), .ZN(
        P1_U2947) );
  NAND2_X1 U17469 ( .A1(n13894), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14104) );
  OAI211_X1 U17470 ( .C1(n14116), .C2(n14024), .A(n14104), .B(n14103), .ZN(
        P1_U2961) );
  NAND2_X1 U17471 ( .A1(n13894), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14106) );
  OAI211_X1 U17472 ( .C1(n14116), .C2(n14107), .A(n14106), .B(n14105), .ZN(
        P1_U2962) );
  NAND2_X1 U17473 ( .A1(n13894), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14109) );
  OAI211_X1 U17474 ( .C1(n14116), .C2(n14110), .A(n14109), .B(n14108), .ZN(
        P1_U2963) );
  INV_X1 U17475 ( .A(n14111), .ZN(n14115) );
  INV_X1 U17476 ( .A(DATAI_15_), .ZN(n14113) );
  INV_X1 U17477 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14112) );
  MUX2_X1 U17478 ( .A(n14113), .B(n14112), .S(n20032), .Z(n14611) );
  OAI222_X1 U17479 ( .A1(n14116), .A2(n14610), .B1(n14115), .B2(n14611), .C1(
        n14114), .C2(n13659), .ZN(P1_U2967) );
  XNOR2_X1 U17480 ( .A(n14751), .B(n16115), .ZN(n14117) );
  XNOR2_X1 U17481 ( .A(n9611), .B(n14117), .ZN(n16112) );
  NAND2_X1 U17482 ( .A1(n16112), .A2(n19981), .ZN(n14123) );
  INV_X1 U17483 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U17484 ( .A1(n19973), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16109) );
  OAI21_X1 U17485 ( .B1(n14741), .B2(n14119), .A(n16109), .ZN(n14120) );
  AOI21_X1 U17486 ( .B1(n16048), .B2(n14121), .A(n14120), .ZN(n14122) );
  OAI211_X1 U17487 ( .C1(n20031), .C2(n19969), .A(n14123), .B(n14122), .ZN(
        P1_U2990) );
  OAI21_X1 U17488 ( .B1(n14540), .B2(n14125), .A(n14124), .ZN(n14534) );
  AOI22_X1 U17489 ( .A1(n14620), .A2(n14390), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14618), .ZN(n14126) );
  OAI21_X1 U17490 ( .B1(n14534), .B2(n14622), .A(n14126), .ZN(P1_U2890) );
  NOR2_X1 U17491 ( .A1(n19905), .A2(n14127), .ZN(n15984) );
  OAI21_X1 U17492 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14128), .A(n15984), 
        .ZN(n14135) );
  INV_X1 U17493 ( .A(n14727), .ZN(n14133) );
  AND2_X1 U17494 ( .A1(n14546), .A2(n14129), .ZN(n14130) );
  OR2_X1 U17495 ( .A1(n14130), .A2(n14528), .ZN(n14924) );
  AOI22_X1 U17496 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19953), .B1(
        n19955), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n14131) );
  OAI211_X1 U17497 ( .C1(n14924), .C2(n19948), .A(n14131), .B(n19933), .ZN(
        n14132) );
  AOI21_X1 U17498 ( .B1(n14133), .B2(n19909), .A(n14132), .ZN(n14134) );
  OAI211_X1 U17499 ( .C1(n14534), .C2(n19924), .A(n14135), .B(n14134), .ZN(
        P1_U2826) );
  OAI21_X1 U17500 ( .B1(n9656), .B2(n11659), .A(n14137), .ZN(n14553) );
  OAI21_X1 U17501 ( .B1(n14553), .B2(n14554), .A(n14137), .ZN(n14139) );
  NAND2_X1 U17502 ( .A1(n14139), .A2(n14138), .ZN(n14542) );
  OAI21_X1 U17503 ( .B1(n14139), .B2(n14138), .A(n14542), .ZN(n16004) );
  XNOR2_X1 U17504 ( .A(n14140), .B(n14543), .ZN(n16003) );
  AOI22_X1 U17505 ( .A1(n16003), .A2(n16021), .B1(n14548), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14141) );
  OAI21_X1 U17506 ( .B1(n16004), .B2(n19968), .A(n14141), .ZN(P1_U2860) );
  AOI22_X1 U17507 ( .A1(n19073), .A2(BUF1_REG_21__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17508 ( .A1(n19071), .A2(n19106), .B1(n19129), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14142) );
  OAI211_X1 U17509 ( .C1(n16191), .C2(n14198), .A(n14143), .B(n14142), .ZN(
        n14144) );
  AOI21_X1 U17510 ( .B1(n14145), .B2(n19108), .A(n14144), .ZN(n14146) );
  INV_X1 U17511 ( .A(n14146), .ZN(P2_U2898) );
  INV_X1 U17512 ( .A(n14559), .ZN(n14148) );
  OAI222_X1 U17513 ( .A1(n16004), .A2(n14622), .B1(n14617), .B2(n14148), .C1(
        n14147), .C2(n14614), .ZN(P1_U2892) );
  OAI211_X1 U17514 ( .C1(n18849), .C2(n15834), .A(n17022), .B(n18716), .ZN(
        n18230) );
  NOR2_X1 U17515 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18230), .ZN(n14149) );
  NAND3_X1 U17516 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18829)
         );
  OAI21_X1 U17517 ( .B1(n14149), .B2(n18829), .A(n18285), .ZN(n18236) );
  INV_X1 U17518 ( .A(n18236), .ZN(n14150) );
  INV_X1 U17519 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18482) );
  NOR2_X1 U17520 ( .A1(n18482), .A2(n18830), .ZN(n18244) );
  INV_X1 U17521 ( .A(n17858), .ZN(n17805) );
  NOR2_X1 U17522 ( .A1(n17805), .A2(n18872), .ZN(n15821) );
  NOR2_X1 U17523 ( .A1(n18244), .A2(n15821), .ZN(n15822) );
  NOR2_X1 U17524 ( .A1(n14150), .A2(n15822), .ZN(n14152) );
  NOR2_X1 U17525 ( .A1(n18830), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18284) );
  OR2_X1 U17526 ( .A1(n18284), .A2(n14150), .ZN(n15820) );
  OR2_X1 U17527 ( .A1(n18243), .A2(n15820), .ZN(n14151) );
  MUX2_X1 U17528 ( .A(n14152), .B(n14151), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17529 ( .A(n14914), .ZN(n14848) );
  INV_X1 U17530 ( .A(n16118), .ZN(n14894) );
  INV_X1 U17531 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14887) );
  NOR4_X1 U17532 ( .A1(n14926), .A2(n11457), .A3(n14883), .A4(n14887), .ZN(
        n14281) );
  NAND3_X1 U17533 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16102) );
  NOR3_X1 U17534 ( .A1(n14747), .A2(n16115), .A3(n16102), .ZN(n14937) );
  NAND2_X1 U17535 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14937), .ZN(
        n14934) );
  INV_X1 U17536 ( .A(n14934), .ZN(n14942) );
  NAND2_X1 U17537 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14942), .ZN(
        n14284) );
  OR2_X1 U17538 ( .A1(n16088), .A2(n14284), .ZN(n14157) );
  NAND2_X1 U17539 ( .A1(n19987), .A2(n14935), .ZN(n14939) );
  NOR2_X1 U17540 ( .A1(n14939), .A2(n14157), .ZN(n14915) );
  AOI21_X1 U17541 ( .B1(n19990), .B2(n16098), .A(n20010), .ZN(n14941) );
  OAI21_X1 U17542 ( .B1(n19988), .B2(n14915), .A(n14941), .ZN(n14153) );
  AOI21_X1 U17543 ( .B1(n19990), .B2(n14157), .A(n14153), .ZN(n14893) );
  OAI21_X1 U17544 ( .B1(n14894), .B2(n14281), .A(n14893), .ZN(n14891) );
  INV_X1 U17545 ( .A(n14891), .ZN(n14164) );
  OR2_X1 U17546 ( .A1(n14155), .A2(n14154), .ZN(n14165) );
  NAND3_X1 U17547 ( .A1(n14165), .A2(n14156), .A3(n20013), .ZN(n14163) );
  AND2_X1 U17548 ( .A1(n14699), .A2(n14281), .ZN(n14161) );
  NAND2_X1 U17549 ( .A1(n14522), .A2(n14158), .ZN(n14159) );
  NAND2_X1 U17550 ( .A1(n14509), .A2(n14159), .ZN(n15969) );
  NAND2_X1 U17551 ( .A1(n19952), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14166) );
  OAI21_X1 U17552 ( .B1(n15969), .B2(n19993), .A(n14166), .ZN(n14160) );
  AOI21_X1 U17553 ( .B1(n14927), .B2(n14161), .A(n14160), .ZN(n14162) );
  OAI211_X1 U17554 ( .C1(n14164), .C2(n14699), .A(n14163), .B(n14162), .ZN(
        P1_U3013) );
  OAI21_X1 U17555 ( .B1(n14516), .B2(n14432), .A(n14506), .ZN(n15970) );
  NAND3_X1 U17556 ( .A1(n14165), .A2(n14156), .A3(n19981), .ZN(n14169) );
  OAI21_X1 U17557 ( .B1(n14741), .B2(n15968), .A(n14166), .ZN(n14167) );
  AOI21_X1 U17558 ( .B1(n15973), .B2(n16048), .A(n14167), .ZN(n14168) );
  OAI211_X1 U17559 ( .C1(n20031), .C2(n15970), .A(n14169), .B(n14168), .ZN(
        P1_U2981) );
  NAND2_X1 U17560 ( .A1(n15557), .A2(n14170), .ZN(n14172) );
  INV_X1 U17561 ( .A(n15331), .ZN(n14173) );
  INV_X1 U17562 ( .A(n16199), .ZN(n14174) );
  INV_X1 U17563 ( .A(n15321), .ZN(n14175) );
  OAI21_X1 U17564 ( .B1(n15323), .B2(n14175), .A(n15322), .ZN(n15314) );
  NAND2_X1 U17565 ( .A1(n14179), .A2(n14178), .ZN(n15306) );
  INV_X1 U17566 ( .A(n14222), .ZN(n14183) );
  INV_X1 U17567 ( .A(n14184), .ZN(n14186) );
  NAND2_X1 U17568 ( .A1(n14186), .A2(n14185), .ZN(n14187) );
  XNOR2_X1 U17569 ( .A(n14188), .B(n14187), .ZN(n14210) );
  OR2_X1 U17570 ( .A1(n10856), .A2(n19765), .ZN(n14202) );
  OAI21_X1 U17571 ( .B1(n19202), .B2(n14189), .A(n14202), .ZN(n14191) );
  NOR2_X1 U17572 ( .A1(n14203), .A2(n19185), .ZN(n14190) );
  AOI211_X1 U17573 ( .C1(n16258), .C2(n14192), .A(n14191), .B(n14190), .ZN(
        n14197) );
  OR2_X1 U17574 ( .A1(n14193), .A2(n14194), .ZN(n15280) );
  OR2_X1 U17575 ( .A1(n14193), .A2(n14195), .ZN(n14225) );
  NAND2_X1 U17576 ( .A1(n14225), .A2(n14199), .ZN(n14207) );
  NAND3_X1 U17577 ( .A1(n15280), .A2(n9578), .A3(n14207), .ZN(n14196) );
  OAI211_X1 U17578 ( .C1(n14210), .C2(n19194), .A(n14197), .B(n14196), .ZN(
        P2_U2993) );
  NOR2_X1 U17579 ( .A1(n16318), .A2(n14198), .ZN(n14205) );
  NAND2_X1 U17580 ( .A1(n14200), .A2(n14199), .ZN(n14201) );
  OAI211_X1 U17581 ( .C1(n14203), .C2(n16319), .A(n14202), .B(n14201), .ZN(
        n14204) );
  AOI211_X1 U17582 ( .C1(n14206), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14205), .B(n14204), .ZN(n14209) );
  NAND3_X1 U17583 ( .A1(n15280), .A2(n16295), .A3(n14207), .ZN(n14208) );
  OAI211_X1 U17584 ( .C1(n14210), .C2(n16299), .A(n14209), .B(n14208), .ZN(
        P2_U3025) );
  AOI21_X1 U17585 ( .B1(n14212), .B2(n14472), .A(n14211), .ZN(n14469) );
  NAND2_X1 U17586 ( .A1(n14469), .A2(n19902), .ZN(n14220) );
  NOR2_X1 U17587 ( .A1(n14475), .A2(n14213), .ZN(n14214) );
  OR2_X1 U17588 ( .A1(n14411), .A2(n14214), .ZN(n14792) );
  INV_X1 U17589 ( .A(n14643), .ZN(n14215) );
  AOI22_X1 U17590 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19953), .B1(
        n19909), .B2(n14215), .ZN(n14217) );
  NAND2_X1 U17591 ( .A1(n19955), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14216) );
  OAI211_X1 U17592 ( .C1(n14792), .C2(n19948), .A(n14217), .B(n14216), .ZN(
        n14218) );
  AOI21_X1 U17593 ( .B1(n15913), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14218), 
        .ZN(n14219) );
  OAI211_X1 U17594 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14414), .A(n14220), 
        .B(n14219), .ZN(P1_U2813) );
  NAND2_X1 U17595 ( .A1(n14222), .A2(n14221), .ZN(n14224) );
  XOR2_X1 U17596 ( .A(n14224), .B(n14223), .Z(n14251) );
  INV_X1 U17597 ( .A(n14225), .ZN(n14229) );
  OR2_X2 U17598 ( .A1(n14193), .A2(n14226), .ZN(n15317) );
  NOR2_X2 U17599 ( .A1(n15317), .A2(n15502), .ZN(n15492) );
  AND2_X2 U17600 ( .A1(n15492), .A2(n14227), .ZN(n15299) );
  AOI21_X1 U17601 ( .B1(n15299), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14228) );
  NOR2_X1 U17602 ( .A1(n14229), .A2(n14228), .ZN(n14248) );
  NOR2_X1 U17603 ( .A1(n13985), .A2(n14230), .ZN(n15126) );
  NOR2_X1 U17604 ( .A1(n15126), .A2(n14231), .ZN(n14232) );
  OR2_X1 U17605 ( .A1(n13058), .A2(n14232), .ZN(n15053) );
  NOR2_X1 U17606 ( .A1(n10856), .A2(n19763), .ZN(n14241) );
  NOR2_X1 U17607 ( .A1(n19191), .A2(n14233), .ZN(n14234) );
  AOI211_X1 U17608 ( .C1(n19177), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14241), .B(n14234), .ZN(n14235) );
  OAI21_X1 U17609 ( .B1(n15053), .B2(n19185), .A(n14235), .ZN(n14236) );
  AOI21_X1 U17610 ( .B1(n14248), .B2(n9578), .A(n14236), .ZN(n14237) );
  OAI21_X1 U17611 ( .B1(n14251), .B2(n19194), .A(n14237), .ZN(P2_U2994) );
  AND2_X1 U17612 ( .A1(n9639), .A2(n14238), .ZN(n14240) );
  OR2_X1 U17613 ( .A1(n14240), .A2(n14239), .ZN(n16190) );
  NOR2_X1 U17614 ( .A1(n16318), .A2(n16190), .ZN(n14247) );
  INV_X1 U17615 ( .A(n14241), .ZN(n14245) );
  INV_X1 U17616 ( .A(n14242), .ZN(n15472) );
  OAI211_X1 U17617 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15472), .B(n14243), .ZN(
        n14244) );
  OAI211_X1 U17618 ( .C1(n15053), .C2(n16319), .A(n14245), .B(n14244), .ZN(
        n14246) );
  AOI211_X1 U17619 ( .C1(n15479), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14247), .B(n14246), .ZN(n14250) );
  NAND2_X1 U17620 ( .A1(n14248), .A2(n16295), .ZN(n14249) );
  OAI211_X1 U17621 ( .C1(n14251), .C2(n16299), .A(n14250), .B(n14249), .ZN(
        P2_U3026) );
  INV_X1 U17622 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17623 ( .A1(n14252), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14253) );
  OAI21_X1 U17624 ( .B1(n14254), .B2(n14268), .A(n14253), .ZN(n14255) );
  AOI21_X1 U17625 ( .B1(n14256), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14255), .ZN(n14257) );
  XNOR2_X2 U17626 ( .A(n14258), .B(n14257), .ZN(n15061) );
  NAND4_X1 U17627 ( .A1(n14259), .A2(n19042), .A3(n13081), .A4(n14260), .ZN(
        n14273) );
  INV_X1 U17628 ( .A(n14261), .ZN(n14264) );
  NOR2_X1 U17629 ( .A1(n14262), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14263) );
  MUX2_X1 U17630 ( .A(n14264), .B(n14263), .S(n10477), .Z(n14321) );
  AOI222_X1 U17631 ( .A1(n10712), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10725), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10577), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14265) );
  OAI22_X1 U17632 ( .A1(n9742), .A2(n19060), .B1(n14268), .B2(n14267), .ZN(
        n14269) );
  AOI21_X1 U17633 ( .B1(n19048), .B2(P2_REIP_REG_31__SCAN_IN), .A(n14269), 
        .ZN(n14270) );
  OAI21_X1 U17634 ( .B1(n19066), .B2(n19046), .A(n14270), .ZN(n14271) );
  AOI21_X1 U17635 ( .B1(n14321), .B2(n12367), .A(n14271), .ZN(n14272) );
  OAI211_X1 U17636 ( .C1(n15061), .C2(n19057), .A(n14273), .B(n14272), .ZN(
        P2_U2824) );
  NOR2_X1 U17637 ( .A1(n14625), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14278) );
  INV_X1 U17638 ( .A(n14276), .ZN(n14277) );
  AOI22_X1 U17639 ( .A1(n14626), .A2(n14278), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14277), .ZN(n14280) );
  XNOR2_X1 U17640 ( .A(n14280), .B(n14279), .ZN(n14307) );
  AND2_X1 U17641 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14281), .ZN(
        n14814) );
  AND2_X1 U17642 ( .A1(n14817), .A2(n14814), .ZN(n14282) );
  NAND2_X1 U17643 ( .A1(n14927), .A2(n14282), .ZN(n14822) );
  NAND2_X1 U17644 ( .A1(n11471), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14283) );
  NOR2_X1 U17645 ( .A1(n14798), .A2(n14780), .ZN(n14772) );
  NAND4_X1 U17646 ( .A1(n14772), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n14279), .ZN(n14298) );
  NAND2_X1 U17647 ( .A1(n19973), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14303) );
  NOR2_X1 U17648 ( .A1(n14939), .A2(n14284), .ZN(n16082) );
  NAND2_X1 U17649 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14814), .ZN(
        n14847) );
  INV_X1 U17650 ( .A(n14847), .ZN(n14285) );
  NAND2_X1 U17651 ( .A1(n16082), .A2(n14285), .ZN(n14842) );
  AND2_X1 U17652 ( .A1(n20011), .A2(n14842), .ZN(n14288) );
  NOR2_X1 U17653 ( .A1(n14284), .A2(n16098), .ZN(n14918) );
  AND2_X1 U17654 ( .A1(n14918), .A2(n14285), .ZN(n14286) );
  NOR2_X1 U17655 ( .A1(n20018), .A2(n14286), .ZN(n14287) );
  OAI22_X1 U17656 ( .A1(n16073), .A2(n14850), .B1(n16118), .B2(n20010), .ZN(
        n14861) );
  NAND2_X1 U17657 ( .A1(n16118), .A2(n14856), .ZN(n14289) );
  NAND2_X1 U17658 ( .A1(n14861), .A2(n14289), .ZN(n14835) );
  NOR2_X1 U17659 ( .A1(n20018), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14290) );
  NOR2_X1 U17660 ( .A1(n14835), .A2(n14290), .ZN(n14818) );
  AND2_X1 U17661 ( .A1(n14291), .A2(n11468), .ZN(n14293) );
  OAI22_X1 U17662 ( .A1(n11471), .A2(n14914), .B1(n14916), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14292) );
  NOR2_X1 U17663 ( .A1(n14293), .A2(n14292), .ZN(n14294) );
  NAND2_X1 U17664 ( .A1(n14809), .A2(n14894), .ZN(n14769) );
  NAND3_X1 U17665 ( .A1(n14809), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U17666 ( .A1(n14769), .A2(n14295), .ZN(n14791) );
  NAND2_X1 U17667 ( .A1(n14791), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14770) );
  OAI21_X1 U17668 ( .B1(n14770), .B2(n14780), .A(n14769), .ZN(n14296) );
  NAND2_X1 U17669 ( .A1(n14296), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14761) );
  NAND3_X1 U17670 ( .A1(n14761), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14769), .ZN(n14297) );
  NAND3_X1 U17671 ( .A1(n14298), .A2(n14303), .A3(n14297), .ZN(n14299) );
  OAI21_X1 U17672 ( .B1(n14307), .B2(n16120), .A(n14301), .ZN(P1_U3000) );
  NAND2_X1 U17673 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14302) );
  OAI211_X1 U17674 ( .C1(n19985), .C2(n14304), .A(n14303), .B(n14302), .ZN(
        n14305) );
  AOI21_X1 U17675 ( .B1(n14315), .B2(n19980), .A(n14305), .ZN(n14306) );
  OAI21_X1 U17676 ( .B1(n14307), .B2(n19877), .A(n14306), .ZN(P1_U2968) );
  INV_X1 U17677 ( .A(n14962), .ZN(n14308) );
  AOI22_X1 U17678 ( .A1(n20160), .A2(n14965), .B1(n14308), .B2(n9848), .ZN(
        n15850) );
  INV_X1 U17679 ( .A(n20724), .ZN(n14971) );
  AOI22_X1 U17680 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n14309), .B1(n9848), 
        .B2(n20722), .ZN(n14310) );
  OAI21_X1 U17681 ( .B1(n15850), .B2(n14971), .A(n14310), .ZN(n14312) );
  NOR2_X1 U17682 ( .A1(n14311), .A2(n9848), .ZN(n15851) );
  AOI22_X1 U17683 ( .A1(n20727), .A2(n14312), .B1(n20724), .B2(n15851), .ZN(
        n14313) );
  OAI21_X1 U17684 ( .B1(n20727), .B2(n9848), .A(n14313), .ZN(P1_U3474) );
  NOR2_X1 U17685 ( .A1(n14316), .A2(n20030), .ZN(n14314) );
  NAND2_X1 U17686 ( .A1(n14614), .A2(n14314), .ZN(n14577) );
  INV_X1 U17687 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16434) );
  NAND3_X1 U17688 ( .A1(n14315), .A2(n14389), .A3(n14614), .ZN(n14319) );
  NOR3_X1 U17689 ( .A1(n14618), .A2(n20032), .A3(n14316), .ZN(n14317) );
  AOI22_X1 U17690 ( .A1(n14604), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14618), .ZN(n14318) );
  OAI211_X1 U17691 ( .C1(n14577), .C2(n16434), .A(n14319), .B(n14318), .ZN(
        P1_U2873) );
  INV_X1 U17692 ( .A(n14327), .ZN(n14323) );
  NAND2_X1 U17693 ( .A1(n14321), .A2(n14320), .ZN(n14326) );
  INV_X1 U17694 ( .A(n14326), .ZN(n14322) );
  AOI21_X1 U17695 ( .B1(n14323), .B2(n14341), .A(n14322), .ZN(n14336) );
  AND2_X1 U17696 ( .A1(n14324), .A2(n15186), .ZN(n14331) );
  INV_X1 U17697 ( .A(n14331), .ZN(n14325) );
  AOI21_X1 U17698 ( .B1(n14341), .B2(n14325), .A(n14326), .ZN(n14335) );
  XNOR2_X1 U17699 ( .A(n14326), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14329) );
  NAND3_X1 U17700 ( .A1(n14328), .A2(n14329), .A3(n14327), .ZN(n14334) );
  INV_X1 U17701 ( .A(n14329), .ZN(n14330) );
  NAND3_X1 U17702 ( .A1(n14332), .A2(n14331), .A3(n14330), .ZN(n14333) );
  OAI211_X1 U17703 ( .C1(n14336), .C2(n14335), .A(n14334), .B(n14333), .ZN(
        n14378) );
  NAND2_X1 U17704 ( .A1(n19176), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14371) );
  NAND3_X1 U17705 ( .A1(n14337), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14341), .ZN(n14338) );
  OAI211_X1 U17706 ( .C1(n19066), .C2(n16318), .A(n14371), .B(n14338), .ZN(
        n14339) );
  INV_X1 U17707 ( .A(n14339), .ZN(n14345) );
  AOI211_X1 U17708 ( .C1(n16316), .C2(n14342), .A(n14341), .B(n14340), .ZN(
        n14343) );
  INV_X1 U17709 ( .A(n14343), .ZN(n14344) );
  INV_X1 U17710 ( .A(n14346), .ZN(n14349) );
  NAND2_X1 U17711 ( .A1(n15194), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14347) );
  XNOR2_X1 U17712 ( .A(n14347), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14376) );
  NAND2_X1 U17713 ( .A1(n14376), .A2(n16295), .ZN(n14348) );
  OAI211_X1 U17714 ( .C1(n14378), .C2(n16299), .A(n14349), .B(n14348), .ZN(
        P2_U3015) );
  AOI22_X1 U17715 ( .A1(n19071), .A2(n19082), .B1(n19129), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U17716 ( .A1(n19073), .A2(BUF1_REG_30__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14350) );
  OAI211_X1 U17717 ( .C1(n14352), .C2(n16191), .A(n14351), .B(n14350), .ZN(
        n14353) );
  INV_X1 U17718 ( .A(n14353), .ZN(n14354) );
  OAI21_X1 U17719 ( .B1(n14355), .B2(n19134), .A(n14354), .ZN(P2_U2889) );
  NAND2_X1 U17720 ( .A1(n14356), .A2(n19958), .ZN(n14369) );
  NAND2_X1 U17721 ( .A1(n19955), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14360) );
  OAI21_X1 U17722 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n14363), .A(n14357), .ZN(
        n14358) );
  AOI22_X1 U17723 ( .A1(n19953), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n14358), .ZN(n14359) );
  OAI211_X1 U17724 ( .C1(n19965), .C2(n14361), .A(n14360), .B(n14359), .ZN(
        n14367) );
  INV_X1 U17725 ( .A(n14362), .ZN(n20020) );
  NAND2_X1 U17726 ( .A1(n19936), .A2(n20020), .ZN(n14365) );
  OR3_X1 U17727 ( .A1(n14363), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n20729), .ZN(
        n14364) );
  NAND2_X1 U17728 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  NOR2_X1 U17729 ( .A1(n14367), .A2(n14366), .ZN(n14368) );
  OAI211_X1 U17730 ( .C1(n19949), .C2(n20448), .A(n14369), .B(n14368), .ZN(
        P1_U2838) );
  NAND2_X1 U17731 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14370) );
  OAI211_X1 U17732 ( .C1(n19191), .C2(n14372), .A(n14371), .B(n14370), .ZN(
        n14373) );
  INV_X1 U17733 ( .A(n14373), .ZN(n14374) );
  AOI21_X1 U17734 ( .B1(n14376), .B2(n9578), .A(n14375), .ZN(n14377) );
  OAI21_X1 U17735 ( .B1(n14378), .B2(n19194), .A(n14377), .ZN(P2_U2983) );
  OAI22_X1 U17736 ( .A1(n14401), .A2(n14380), .B1(n14379), .B2(n14398), .ZN(
        n14382) );
  XNOR2_X1 U17737 ( .A(n14382), .B(n14381), .ZN(n14765) );
  AOI22_X1 U17738 ( .A1(n14384), .A2(n19909), .B1(n19953), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U17739 ( .A1(n19955), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14385) );
  NAND2_X1 U17740 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  OAI21_X1 U17741 ( .B1(n14394), .B2(n19924), .A(n14388), .ZN(P1_U2810) );
  AOI22_X1 U17742 ( .A1(n14603), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14618), .ZN(n14392) );
  NOR3_X4 U17743 ( .A1(n14618), .A2(n14389), .A3(n20073), .ZN(n14606) );
  AOI22_X1 U17744 ( .A1(n14606), .A2(n14390), .B1(n14604), .B2(DATAI_30_), 
        .ZN(n14391) );
  OAI211_X1 U17745 ( .C1(n14394), .C2(n14622), .A(n14392), .B(n14391), .ZN(
        P1_U2874) );
  INV_X1 U17746 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14393) );
  OAI222_X1 U17747 ( .A1(n14550), .A2(n14394), .B1(n14535), .B2(n14393), .C1(
        n14765), .C2(n19967), .ZN(P1_U2842) );
  AOI21_X1 U17748 ( .B1(n14397), .B2(n14395), .A(n14396), .ZN(n14631) );
  NAND2_X1 U17749 ( .A1(n14631), .A2(n19902), .ZN(n14407) );
  AND2_X1 U17750 ( .A1(n14398), .A2(n14399), .ZN(n14400) );
  OR2_X1 U17751 ( .A1(n14401), .A2(n14400), .ZN(n14775) );
  INV_X1 U17752 ( .A(n14629), .ZN(n14402) );
  AOI22_X1 U17753 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19953), .B1(
        n19909), .B2(n14402), .ZN(n14404) );
  NAND2_X1 U17754 ( .A1(n19955), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14403) );
  OAI211_X1 U17755 ( .C1(n14775), .C2(n19948), .A(n14404), .B(n14403), .ZN(
        n14405) );
  AOI21_X1 U17756 ( .B1(n14417), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14405), 
        .ZN(n14406) );
  OAI211_X1 U17757 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14408), .A(n14407), 
        .B(n14406), .ZN(P1_U2811) );
  OAI21_X1 U17758 ( .B1(n14211), .B2(n14409), .A(n14395), .ZN(n14638) );
  OAI21_X1 U17759 ( .B1(n14411), .B2(n14410), .A(n14398), .ZN(n14779) );
  AOI22_X1 U17760 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19953), .B1(
        n19909), .B2(n14641), .ZN(n14413) );
  NAND2_X1 U17761 ( .A1(n19955), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14412) );
  OAI211_X1 U17762 ( .C1(n14779), .C2(n19948), .A(n14413), .B(n14412), .ZN(
        n14416) );
  NOR3_X1 U17763 ( .A1(n14414), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n20700), 
        .ZN(n14415) );
  OAI21_X1 U17764 ( .B1(n14638), .B2(n19924), .A(n14418), .ZN(P1_U2812) );
  NAND2_X1 U17765 ( .A1(n14516), .A2(n14419), .ZN(n14481) );
  NAND2_X1 U17766 ( .A1(n14516), .A2(n14420), .ZN(n14574) );
  NAND2_X1 U17767 ( .A1(n14574), .A2(n14421), .ZN(n14422) );
  NAND2_X1 U17768 ( .A1(n14481), .A2(n14422), .ZN(n14673) );
  OR2_X1 U17769 ( .A1(n14833), .A2(n14423), .ZN(n14424) );
  NAND2_X1 U17770 ( .A1(n14485), .A2(n14424), .ZN(n14825) );
  INV_X1 U17771 ( .A(n14425), .ZN(n15937) );
  AOI22_X1 U17772 ( .A1(n15937), .A2(P1_REIP_REG_24__SCAN_IN), .B1(n19955), 
        .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17773 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19953), .B1(
        n14670), .B2(n19909), .ZN(n14426) );
  OAI211_X1 U17774 ( .C1(n14825), .C2(n19948), .A(n14427), .B(n14426), .ZN(
        n14429) );
  NOR2_X1 U17775 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14428), .ZN(n15927) );
  NOR2_X1 U17776 ( .A1(n14429), .A2(n15927), .ZN(n14430) );
  OAI21_X1 U17777 ( .B1(n14673), .B2(n19924), .A(n14430), .ZN(P1_U2816) );
  AND2_X1 U17778 ( .A1(n14516), .A2(n14432), .ZN(n14434) );
  INV_X1 U17779 ( .A(n14691), .ZN(n14585) );
  NOR2_X1 U17780 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n14439), .ZN(n15948) );
  OAI21_X1 U17781 ( .B1(n15957), .B2(n15948), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14443) );
  AND2_X1 U17782 ( .A1(n14495), .A2(n14436), .ZN(n14437) );
  OR2_X1 U17783 ( .A1(n14437), .A2(n14831), .ZN(n14853) );
  AOI22_X1 U17784 ( .A1(n14687), .A2(n19909), .B1(n19955), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n14438) );
  OAI21_X1 U17785 ( .B1(n19948), .B2(n14853), .A(n14438), .ZN(n14441) );
  INV_X1 U17786 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20689) );
  NOR3_X1 U17787 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14439), .A3(n20689), 
        .ZN(n14440) );
  AOI211_X1 U17788 ( .C1(n19953), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14441), .B(n14440), .ZN(n14442) );
  OAI211_X1 U17789 ( .C1(n14585), .C2(n19924), .A(n14443), .B(n14442), .ZN(
        P1_U2818) );
  AOI21_X1 U17790 ( .B1(n14445), .B2(n14533), .A(n14444), .ZN(n14719) );
  INV_X1 U17791 ( .A(n14719), .ZN(n14609) );
  INV_X1 U17792 ( .A(n15979), .ZN(n14448) );
  NOR2_X1 U17793 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14446), .ZN(n15992) );
  NOR2_X1 U17794 ( .A1(n15984), .A2(n15992), .ZN(n14447) );
  MUX2_X1 U17795 ( .A(n14448), .B(n14447), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14455) );
  OR2_X1 U17796 ( .A1(n14530), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U17797 ( .A1(n14520), .A2(n14450), .ZN(n14897) );
  INV_X1 U17798 ( .A(n14717), .ZN(n14451) );
  AOI22_X1 U17799 ( .A1(n19955), .A2(P1_EBX_REG_16__SCAN_IN), .B1(n14451), 
        .B2(n19909), .ZN(n14452) );
  OAI21_X1 U17800 ( .B1(n19948), .B2(n14897), .A(n14452), .ZN(n14453) );
  AOI211_X1 U17801 ( .C1(n19953), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14453), .B(n19952), .ZN(n14454) );
  OAI211_X1 U17802 ( .C1(n14609), .C2(n19924), .A(n14455), .B(n14454), .ZN(
        P1_U2824) );
  NAND2_X1 U17803 ( .A1(n19919), .A2(n19965), .ZN(n14456) );
  AOI22_X1 U17804 ( .A1(n19955), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n14456), .B2(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U17805 ( .A1(n19932), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14457) );
  OAI211_X1 U17806 ( .C1(n19948), .C2(n14459), .A(n14458), .B(n14457), .ZN(
        n14460) );
  AOI21_X1 U17807 ( .B1(n20160), .B2(n14461), .A(n14460), .ZN(n14462) );
  OAI21_X1 U17808 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(P1_U2840) );
  INV_X1 U17809 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14465) );
  OAI22_X1 U17810 ( .A1(n14466), .A2(n19967), .B1(n14465), .B2(n14535), .ZN(
        P1_U2841) );
  INV_X1 U17811 ( .A(n14631), .ZN(n14558) );
  OAI222_X1 U17812 ( .A1(n14467), .A2(n14535), .B1(n19967), .B2(n14775), .C1(
        n14558), .C2(n14550), .ZN(P1_U2843) );
  OAI222_X1 U17813 ( .A1(n14468), .A2(n14535), .B1(n19967), .B2(n14779), .C1(
        n14638), .C2(n19968), .ZN(P1_U2844) );
  INV_X1 U17814 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14470) );
  INV_X1 U17815 ( .A(n14469), .ZN(n14650) );
  OAI222_X1 U17816 ( .A1(n14470), .A2(n14535), .B1(n19967), .B2(n14792), .C1(
        n14650), .C2(n14550), .ZN(P1_U2845) );
  OAI21_X1 U17817 ( .B1(n14471), .B2(n14473), .A(n14472), .ZN(n15914) );
  AND2_X1 U17818 ( .A1(n14483), .A2(n14474), .ZN(n14476) );
  OR2_X1 U17819 ( .A1(n14476), .A2(n14475), .ZN(n15915) );
  OAI22_X1 U17820 ( .A1(n15915), .A2(n19967), .B1(n14477), .B2(n14535), .ZN(
        n14478) );
  INV_X1 U17821 ( .A(n14478), .ZN(n14479) );
  OAI21_X1 U17822 ( .B1(n15914), .B2(n19968), .A(n14479), .ZN(P1_U2846) );
  AND2_X1 U17823 ( .A1(n14481), .A2(n14480), .ZN(n14482) );
  NOR2_X1 U17824 ( .A1(n14471), .A2(n14482), .ZN(n15926) );
  INV_X1 U17825 ( .A(n15926), .ZN(n14570) );
  INV_X1 U17826 ( .A(n14483), .ZN(n14484) );
  AOI21_X1 U17827 ( .B1(n14486), .B2(n14485), .A(n14484), .ZN(n15923) );
  AOI22_X1 U17828 ( .A1(n15923), .A2(n16021), .B1(n14548), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14487) );
  OAI21_X1 U17829 ( .B1(n14570), .B2(n14550), .A(n14487), .ZN(P1_U2847) );
  OAI22_X1 U17830 ( .A1(n14825), .A2(n19967), .B1(n14488), .B2(n14535), .ZN(
        n14489) );
  INV_X1 U17831 ( .A(n14489), .ZN(n14490) );
  OAI21_X1 U17832 ( .B1(n14673), .B2(n14550), .A(n14490), .ZN(P1_U2848) );
  OAI22_X1 U17833 ( .A1(n14853), .A2(n19967), .B1(n14491), .B2(n14535), .ZN(
        n14492) );
  AOI21_X1 U17834 ( .B1(n14691), .B2(n16023), .A(n14492), .ZN(n14493) );
  INV_X1 U17835 ( .A(n14493), .ZN(P1_U2850) );
  INV_X1 U17836 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14500) );
  INV_X1 U17837 ( .A(n14494), .ZN(n14496) );
  OAI21_X1 U17838 ( .B1(n9672), .B2(n14496), .A(n14495), .ZN(n15945) );
  OAI21_X1 U17839 ( .B1(n14504), .B2(n14501), .A(n14497), .ZN(n14499) );
  NAND2_X1 U17840 ( .A1(n14499), .A2(n14498), .ZN(n15944) );
  OAI222_X1 U17841 ( .A1(n14500), .A2(n14535), .B1(n19967), .B2(n15945), .C1(
        n15944), .C2(n14550), .ZN(P1_U2851) );
  INV_X1 U17842 ( .A(n14508), .ZN(n14503) );
  AOI21_X1 U17843 ( .B1(n9829), .B2(n14503), .A(n9672), .ZN(n14876) );
  INV_X1 U17844 ( .A(n14876), .ZN(n15954) );
  OAI222_X1 U17845 ( .A1(n14550), .A2(n15955), .B1(n14535), .B2(n12252), .C1(
        n15954), .C2(n19967), .ZN(P1_U2852) );
  INV_X1 U17846 ( .A(n14504), .ZN(n14505) );
  AOI21_X1 U17847 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n16032) );
  INV_X1 U17848 ( .A(n16032), .ZN(n14595) );
  AOI21_X1 U17849 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n16074) );
  AOI22_X1 U17850 ( .A1(n16074), .A2(n16021), .B1(n14548), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14511) );
  OAI21_X1 U17851 ( .B1(n14595), .B2(n14550), .A(n14511), .ZN(P1_U2853) );
  OAI22_X1 U17852 ( .A1(n15969), .A2(n19967), .B1(n14512), .B2(n14535), .ZN(
        n14513) );
  INV_X1 U17853 ( .A(n14513), .ZN(n14514) );
  OAI21_X1 U17854 ( .B1(n15970), .B2(n19968), .A(n14514), .ZN(P1_U2854) );
  INV_X1 U17855 ( .A(n14515), .ZN(n14518) );
  INV_X1 U17856 ( .A(n14444), .ZN(n14517) );
  AOI21_X1 U17857 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n16037) );
  INV_X1 U17858 ( .A(n16037), .ZN(n14602) );
  NAND2_X1 U17859 ( .A1(n14520), .A2(n14519), .ZN(n14521) );
  NAND2_X1 U17860 ( .A1(n14522), .A2(n14521), .ZN(n15976) );
  INV_X1 U17861 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14523) );
  OAI222_X1 U17862 ( .A1(n14602), .A2(n14550), .B1(n19967), .B2(n15976), .C1(
        n14535), .C2(n14523), .ZN(P1_U2855) );
  OAI22_X1 U17863 ( .A1(n14897), .A2(n19967), .B1(n14524), .B2(n14535), .ZN(
        n14525) );
  AOI21_X1 U17864 ( .B1(n14719), .B2(n16023), .A(n14525), .ZN(n14526) );
  INV_X1 U17865 ( .A(n14526), .ZN(P1_U2856) );
  NOR2_X1 U17866 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  OR2_X1 U17867 ( .A1(n14530), .A2(n14529), .ZN(n15987) );
  INV_X1 U17868 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U17869 ( .A1(n14124), .A2(n14531), .ZN(n14532) );
  OAI222_X1 U17870 ( .A1(n15987), .A2(n19967), .B1(n15985), .B2(n14535), .C1(
        n14612), .C2(n14550), .ZN(P1_U2857) );
  INV_X1 U17871 ( .A(n14534), .ZN(n14731) );
  OAI22_X1 U17872 ( .A1(n14924), .A2(n19967), .B1(n14536), .B2(n14535), .ZN(
        n14537) );
  AOI21_X1 U17873 ( .B1(n14731), .B2(n16023), .A(n14537), .ZN(n14538) );
  INV_X1 U17874 ( .A(n14538), .ZN(P1_U2858) );
  INV_X1 U17875 ( .A(n14539), .ZN(n14541) );
  AOI21_X1 U17876 ( .B1(n14542), .B2(n14541), .A(n14540), .ZN(n14743) );
  INV_X1 U17877 ( .A(n14743), .ZN(n15998) );
  INV_X1 U17878 ( .A(n14543), .ZN(n14545) );
  OAI21_X1 U17879 ( .B1(n14140), .B2(n14545), .A(n14544), .ZN(n14547) );
  AND2_X1 U17880 ( .A1(n14547), .A2(n14546), .ZN(n16084) );
  AOI22_X1 U17881 ( .A1(n16084), .A2(n16021), .B1(n14548), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14549) );
  OAI21_X1 U17882 ( .B1(n15998), .B2(n14550), .A(n14549), .ZN(P1_U2859) );
  OAI21_X1 U17883 ( .B1(n14552), .B2(n14551), .A(n14140), .ZN(n16012) );
  INV_X1 U17884 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14555) );
  XOR2_X1 U17885 ( .A(n14554), .B(n14553), .Z(n16057) );
  INV_X1 U17886 ( .A(n16057), .ZN(n14623) );
  OAI222_X1 U17887 ( .A1(n16012), .A2(n19967), .B1(n14555), .B2(n14535), .C1(
        n19968), .C2(n14623), .ZN(P1_U2861) );
  AOI22_X1 U17888 ( .A1(n14603), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14618), .ZN(n14557) );
  AOI22_X1 U17889 ( .A1(n14606), .A2(n14613), .B1(n14604), .B2(DATAI_29_), 
        .ZN(n14556) );
  OAI211_X1 U17890 ( .C1(n14558), .C2(n14622), .A(n14557), .B(n14556), .ZN(
        P1_U2875) );
  AOI22_X1 U17891 ( .A1(n14603), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14618), .ZN(n14561) );
  AOI22_X1 U17892 ( .A1(n14606), .A2(n14559), .B1(n14604), .B2(DATAI_28_), 
        .ZN(n14560) );
  OAI211_X1 U17893 ( .C1(n14638), .C2(n14622), .A(n14561), .B(n14560), .ZN(
        P1_U2876) );
  AOI22_X1 U17894 ( .A1(n14603), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14618), .ZN(n14563) );
  AOI22_X1 U17895 ( .A1(n14606), .A2(n14619), .B1(n14604), .B2(DATAI_27_), 
        .ZN(n14562) );
  OAI211_X1 U17896 ( .C1(n14650), .C2(n14622), .A(n14563), .B(n14562), .ZN(
        P1_U2877) );
  AOI22_X1 U17897 ( .A1(n14603), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14618), .ZN(n14566) );
  AOI22_X1 U17898 ( .A1(n14606), .A2(n14564), .B1(n14604), .B2(DATAI_26_), 
        .ZN(n14565) );
  OAI211_X1 U17899 ( .C1(n15914), .C2(n14622), .A(n14566), .B(n14565), .ZN(
        P1_U2878) );
  AOI22_X1 U17900 ( .A1(n14603), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14618), .ZN(n14569) );
  AOI22_X1 U17901 ( .A1(n14606), .A2(n14567), .B1(n14604), .B2(DATAI_25_), 
        .ZN(n14568) );
  OAI211_X1 U17902 ( .C1(n14570), .C2(n14622), .A(n14569), .B(n14568), .ZN(
        P1_U2879) );
  AOI22_X1 U17903 ( .A1(n14603), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14618), .ZN(n14573) );
  AOI22_X1 U17904 ( .A1(n14606), .A2(n14571), .B1(n14604), .B2(DATAI_24_), 
        .ZN(n14572) );
  OAI211_X1 U17905 ( .C1(n14673), .C2(n14622), .A(n14573), .B(n14572), .ZN(
        P1_U2880) );
  OAI21_X1 U17906 ( .B1(n14576), .B2(n14575), .A(n14574), .ZN(n15935) );
  INV_X1 U17907 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16450) );
  OAI22_X1 U17908 ( .A1(n14577), .A2(n16450), .B1(n13641), .B2(n14614), .ZN(
        n14580) );
  INV_X1 U17909 ( .A(n14606), .ZN(n14578) );
  NOR2_X1 U17910 ( .A1(n14578), .A2(n20087), .ZN(n14579) );
  AOI211_X1 U17911 ( .C1(n14604), .C2(DATAI_23_), .A(n14580), .B(n14579), .ZN(
        n14581) );
  OAI21_X1 U17912 ( .B1(n15935), .B2(n14622), .A(n14581), .ZN(P1_U2881) );
  AOI22_X1 U17913 ( .A1(n14603), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14618), .ZN(n14584) );
  AOI22_X1 U17914 ( .A1(n14606), .A2(n14582), .B1(n14604), .B2(DATAI_22_), 
        .ZN(n14583) );
  OAI211_X1 U17915 ( .C1(n14585), .C2(n14622), .A(n14584), .B(n14583), .ZN(
        P1_U2882) );
  AOI22_X1 U17916 ( .A1(n14603), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14618), .ZN(n14588) );
  AOI22_X1 U17917 ( .A1(n14606), .A2(n14586), .B1(n14604), .B2(DATAI_21_), 
        .ZN(n14587) );
  OAI211_X1 U17918 ( .C1(n15944), .C2(n14622), .A(n14588), .B(n14587), .ZN(
        P1_U2883) );
  AOI22_X1 U17919 ( .A1(n14603), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14618), .ZN(n14591) );
  AOI22_X1 U17920 ( .A1(n14606), .A2(n14589), .B1(n14604), .B2(DATAI_20_), 
        .ZN(n14590) );
  OAI211_X1 U17921 ( .C1(n15955), .C2(n14622), .A(n14591), .B(n14590), .ZN(
        P1_U2884) );
  AOI22_X1 U17922 ( .A1(n14603), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14618), .ZN(n14594) );
  AOI22_X1 U17923 ( .A1(n14606), .A2(n14592), .B1(n14604), .B2(DATAI_19_), 
        .ZN(n14593) );
  OAI211_X1 U17924 ( .C1(n14595), .C2(n14622), .A(n14594), .B(n14593), .ZN(
        P1_U2885) );
  AOI22_X1 U17925 ( .A1(n14603), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14618), .ZN(n14598) );
  AOI22_X1 U17926 ( .A1(n14606), .A2(n14596), .B1(n14604), .B2(DATAI_18_), 
        .ZN(n14597) );
  OAI211_X1 U17927 ( .C1(n15970), .C2(n14622), .A(n14598), .B(n14597), .ZN(
        P1_U2886) );
  AOI22_X1 U17928 ( .A1(n14603), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14618), .ZN(n14601) );
  AOI22_X1 U17929 ( .A1(n14606), .A2(n14599), .B1(n14604), .B2(DATAI_17_), 
        .ZN(n14600) );
  OAI211_X1 U17930 ( .C1(n14602), .C2(n14622), .A(n14601), .B(n14600), .ZN(
        P1_U2887) );
  AOI22_X1 U17931 ( .A1(n14603), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14618), .ZN(n14608) );
  AOI22_X1 U17932 ( .A1(n14606), .A2(n14605), .B1(n14604), .B2(DATAI_16_), 
        .ZN(n14607) );
  OAI211_X1 U17933 ( .C1(n14609), .C2(n14622), .A(n14608), .B(n14607), .ZN(
        P1_U2888) );
  OAI222_X1 U17934 ( .A1(n14612), .A2(n14622), .B1(n14617), .B2(n14611), .C1(
        n14614), .C2(n14610), .ZN(P1_U2889) );
  INV_X1 U17935 ( .A(n14613), .ZN(n14616) );
  OAI222_X1 U17936 ( .A1(n14622), .A2(n15998), .B1(n14617), .B2(n14616), .C1(
        n14615), .C2(n14614), .ZN(P1_U2891) );
  AOI22_X1 U17937 ( .A1(n14620), .A2(n14619), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14618), .ZN(n14621) );
  OAI21_X1 U17938 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(P1_U2893) );
  NAND2_X1 U17939 ( .A1(n14625), .A2(n14624), .ZN(n14627) );
  XOR2_X1 U17940 ( .A(n14627), .B(n14626), .Z(n14778) );
  NAND2_X1 U17941 ( .A1(n19973), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14774) );
  NAND2_X1 U17942 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14628) );
  OAI211_X1 U17943 ( .C1(n19985), .C2(n14629), .A(n14774), .B(n14628), .ZN(
        n14630) );
  AOI21_X1 U17944 ( .B1(n14631), .B2(n19980), .A(n14630), .ZN(n14632) );
  OAI21_X1 U17945 ( .B1(n19877), .B2(n14778), .A(n14632), .ZN(P1_U2970) );
  NAND2_X1 U17946 ( .A1(n14653), .A2(n14803), .ZN(n14645) );
  NAND2_X1 U17947 ( .A1(n14748), .A2(n14633), .ZN(n14651) );
  NAND3_X1 U17948 ( .A1(n14677), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14651), .ZN(n14635) );
  MUX2_X1 U17949 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14803), .S(
        n14748), .Z(n14634) );
  AOI21_X1 U17950 ( .B1(n14645), .B2(n14635), .A(n14634), .ZN(n14636) );
  XNOR2_X1 U17951 ( .A(n14636), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14789) );
  NAND2_X1 U17952 ( .A1(n19973), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14783) );
  OAI21_X1 U17953 ( .B1(n14741), .B2(n14637), .A(n14783), .ZN(n14640) );
  NOR2_X1 U17954 ( .A1(n14638), .A2(n20031), .ZN(n14639) );
  AOI211_X1 U17955 ( .C1(n16048), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14642) );
  OAI21_X1 U17956 ( .B1(n19877), .B2(n14789), .A(n14642), .ZN(P1_U2971) );
  NOR2_X1 U17957 ( .A1(n19933), .A2(n20700), .ZN(n14794) );
  NOR2_X1 U17958 ( .A1(n19985), .A2(n14643), .ZN(n14644) );
  AOI211_X1 U17959 ( .C1(n19974), .C2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14794), .B(n14644), .ZN(n14649) );
  NAND2_X1 U17960 ( .A1(n14790), .A2(n19981), .ZN(n14648) );
  OAI211_X1 U17961 ( .C1(n14650), .C2(n20031), .A(n14649), .B(n14648), .ZN(
        P1_U2972) );
  NOR2_X1 U17962 ( .A1(n14666), .A2(n16052), .ZN(n14652) );
  OAI21_X1 U17963 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14654) );
  XNOR2_X1 U17964 ( .A(n14654), .B(n14803), .ZN(n14807) );
  NAND2_X1 U17965 ( .A1(n19973), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U17966 ( .B1(n14741), .B2(n14655), .A(n14800), .ZN(n14657) );
  NOR2_X1 U17967 ( .A1(n15914), .A2(n20031), .ZN(n14656) );
  AOI211_X1 U17968 ( .C1(n16048), .C2(n15912), .A(n14657), .B(n14656), .ZN(
        n14658) );
  OAI21_X1 U17969 ( .B1(n19877), .B2(n14807), .A(n14658), .ZN(P1_U2973) );
  NAND2_X1 U17970 ( .A1(n14659), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14667) );
  INV_X1 U17971 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20806) );
  NAND2_X1 U17972 ( .A1(n14666), .A2(n20806), .ZN(n14660) );
  MUX2_X1 U17973 ( .A(n14660), .B(n11468), .S(n14748), .Z(n14661) );
  XNOR2_X1 U17974 ( .A(n14662), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14813) );
  NAND2_X1 U17975 ( .A1(n19952), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U17976 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14663) );
  OAI211_X1 U17977 ( .C1(n19985), .C2(n15922), .A(n14808), .B(n14663), .ZN(
        n14664) );
  AOI21_X1 U17978 ( .B1(n15926), .B2(n19980), .A(n14664), .ZN(n14665) );
  OAI21_X1 U17979 ( .B1(n14813), .B2(n19877), .A(n14665), .ZN(P1_U2974) );
  NAND2_X1 U17980 ( .A1(n14666), .A2(n14667), .ZN(n14668) );
  MUX2_X1 U17981 ( .A(n14668), .B(n14667), .S(n14748), .Z(n14669) );
  XNOR2_X1 U17982 ( .A(n14669), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14827) );
  AND2_X1 U17983 ( .A1(n19952), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14820) );
  AOI21_X1 U17984 ( .B1(n19974), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14820), .ZN(n14672) );
  NAND2_X1 U17985 ( .A1(n16048), .A2(n14670), .ZN(n14671) );
  OAI211_X1 U17986 ( .C1(n14673), .C2(n20031), .A(n14672), .B(n14671), .ZN(
        n14674) );
  AOI21_X1 U17987 ( .B1(n14827), .B2(n19981), .A(n14674), .ZN(n14675) );
  INV_X1 U17988 ( .A(n14675), .ZN(P1_U2975) );
  XNOR2_X1 U17989 ( .A(n14751), .B(n20806), .ZN(n14676) );
  XNOR2_X1 U17990 ( .A(n14677), .B(n14676), .ZN(n14829) );
  NAND2_X1 U17991 ( .A1(n14829), .A2(n19981), .ZN(n14680) );
  AND2_X1 U17992 ( .A1(n19973), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14834) );
  NOR2_X1 U17993 ( .A1(n19985), .A2(n15932), .ZN(n14678) );
  AOI211_X1 U17994 ( .C1(n19974), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14834), .B(n14678), .ZN(n14679) );
  OAI211_X1 U17995 ( .C1(n20031), .C2(n15935), .A(n14680), .B(n14679), .ZN(
        P1_U2976) );
  INV_X1 U17996 ( .A(n14850), .ZN(n14681) );
  NAND2_X1 U17997 ( .A1(n14681), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14682) );
  OR2_X1 U17998 ( .A1(n14156), .A2(n14682), .ZN(n14683) );
  NAND2_X1 U17999 ( .A1(n14683), .A2(n14751), .ZN(n14684) );
  NAND2_X1 U18000 ( .A1(n14685), .A2(n14684), .ZN(n14686) );
  XNOR2_X1 U18001 ( .A(n14686), .B(n11462), .ZN(n14859) );
  INV_X1 U18002 ( .A(n14687), .ZN(n14689) );
  NAND2_X1 U18003 ( .A1(n19952), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U18004 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14688) );
  OAI211_X1 U18005 ( .C1(n19985), .C2(n14689), .A(n14852), .B(n14688), .ZN(
        n14690) );
  AOI21_X1 U18006 ( .B1(n14691), .B2(n19980), .A(n14690), .ZN(n14692) );
  OAI21_X1 U18007 ( .B1(n19877), .B2(n14859), .A(n14692), .ZN(P1_U2977) );
  NAND2_X1 U18008 ( .A1(n14751), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16030) );
  NOR2_X1 U18009 ( .A1(n14156), .A2(n16030), .ZN(n14698) );
  NAND2_X1 U18010 ( .A1(n14698), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14702) );
  OAI21_X1 U18011 ( .B1(n14693), .B2(n14751), .A(n14702), .ZN(n14694) );
  XOR2_X1 U18012 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14694), .Z(
        n14860) );
  NAND2_X1 U18013 ( .A1(n14860), .A2(n19981), .ZN(n14697) );
  NOR2_X1 U18014 ( .A1(n19933), .A2(n20689), .ZN(n14863) );
  NOR2_X1 U18015 ( .A1(n19985), .A2(n15942), .ZN(n14695) );
  AOI211_X1 U18016 ( .C1(n19974), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14863), .B(n14695), .ZN(n14696) );
  OAI211_X1 U18017 ( .C1(n20031), .C2(n15944), .A(n14697), .B(n14696), .ZN(
        P1_U2978) );
  OR2_X1 U18018 ( .A1(n14698), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14701) );
  OAI21_X1 U18019 ( .B1(n14748), .B2(n14699), .A(n14156), .ZN(n16031) );
  NAND2_X1 U18020 ( .A1(n16052), .A2(n14700), .ZN(n16027) );
  NOR2_X1 U18021 ( .A1(n16031), .A2(n16027), .ZN(n16026) );
  MUX2_X1 U18022 ( .A(n14701), .B(n14868), .S(n16026), .Z(n14703) );
  NAND2_X1 U18023 ( .A1(n14703), .A2(n14702), .ZN(n14878) );
  NAND2_X1 U18024 ( .A1(n16048), .A2(n15953), .ZN(n14704) );
  NAND2_X1 U18025 ( .A1(n19952), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14872) );
  OAI211_X1 U18026 ( .C1(n14741), .C2(n15959), .A(n14704), .B(n14872), .ZN(
        n14705) );
  AOI21_X1 U18027 ( .B1(n14706), .B2(n19980), .A(n14705), .ZN(n14707) );
  OAI21_X1 U18028 ( .B1(n14878), .B2(n19877), .A(n14707), .ZN(P1_U2979) );
  INV_X1 U18029 ( .A(n16053), .ZN(n14736) );
  INV_X1 U18030 ( .A(n14709), .ZN(n14711) );
  AOI21_X1 U18031 ( .B1(n14736), .B2(n14711), .A(n14710), .ZN(n14905) );
  AND2_X1 U18032 ( .A1(n14712), .A2(n14713), .ZN(n14904) );
  NAND2_X1 U18033 ( .A1(n14905), .A2(n14904), .ZN(n14903) );
  NAND2_X1 U18034 ( .A1(n14903), .A2(n14713), .ZN(n14714) );
  XOR2_X1 U18035 ( .A(n14715), .B(n14714), .Z(n14902) );
  NAND2_X1 U18036 ( .A1(n19952), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U18037 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14716) );
  OAI211_X1 U18038 ( .C1(n14717), .C2(n19985), .A(n14896), .B(n14716), .ZN(
        n14718) );
  AOI21_X1 U18039 ( .B1(n14719), .B2(n19980), .A(n14718), .ZN(n14720) );
  OAI21_X1 U18040 ( .B1(n14902), .B2(n19877), .A(n14720), .ZN(P1_U2983) );
  NAND2_X1 U18041 ( .A1(n16053), .A2(n14721), .ZN(n14882) );
  NAND3_X1 U18042 ( .A1(n14882), .A2(n14722), .A3(n14735), .ZN(n14724) );
  NAND2_X1 U18043 ( .A1(n14724), .A2(n14723), .ZN(n14726) );
  XNOR2_X1 U18044 ( .A(n14751), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14725) );
  XNOR2_X1 U18045 ( .A(n14726), .B(n14725), .ZN(n14929) );
  NOR2_X1 U18046 ( .A1(n14727), .A2(n19985), .ZN(n14730) );
  INV_X1 U18047 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14728) );
  OAI22_X1 U18048 ( .A1(n14741), .A2(n14728), .B1(n19933), .B2(n20677), .ZN(
        n14729) );
  AOI211_X1 U18049 ( .C1(n14731), .C2(n19980), .A(n14730), .B(n14729), .ZN(
        n14732) );
  OAI21_X1 U18050 ( .B1(n14929), .B2(n19877), .A(n14732), .ZN(P1_U2985) );
  AOI21_X1 U18051 ( .B1(n14747), .B2(n14733), .A(n14751), .ZN(n14734) );
  AOI21_X1 U18052 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14931) );
  AOI21_X1 U18053 ( .B1(n16052), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14737), .ZN(n14930) );
  AND2_X1 U18054 ( .A1(n14931), .A2(n14930), .ZN(n14932) );
  NOR2_X1 U18055 ( .A1(n14932), .A2(n14737), .ZN(n14738) );
  XOR2_X1 U18056 ( .A(n14739), .B(n14738), .Z(n16083) );
  OAI22_X1 U18057 ( .A1(n14741), .A2(n14740), .B1(n19933), .B2(n20675), .ZN(
        n14742) );
  AOI21_X1 U18058 ( .B1(n16048), .B2(n16001), .A(n14742), .ZN(n14745) );
  NAND2_X1 U18059 ( .A1(n14743), .A2(n19980), .ZN(n14744) );
  OAI211_X1 U18060 ( .C1(n16083), .C2(n19877), .A(n14745), .B(n14744), .ZN(
        P1_U2986) );
  NAND2_X1 U18061 ( .A1(n14746), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14750) );
  XNOR2_X1 U18062 ( .A(n16053), .B(n14747), .ZN(n14749) );
  MUX2_X1 U18063 ( .A(n14750), .B(n14749), .S(n14748), .Z(n14753) );
  NOR3_X1 U18064 ( .A1(n14746), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14751), .ZN(n16054) );
  INV_X1 U18065 ( .A(n16054), .ZN(n14752) );
  NAND2_X1 U18066 ( .A1(n14753), .A2(n14752), .ZN(n16101) );
  INV_X1 U18067 ( .A(n16101), .ZN(n14759) );
  AOI22_X1 U18068 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14754) );
  OAI21_X1 U18069 ( .B1(n14755), .B2(n19985), .A(n14754), .ZN(n14756) );
  AOI21_X1 U18070 ( .B1(n14757), .B2(n19980), .A(n14756), .ZN(n14758) );
  OAI21_X1 U18071 ( .B1(n14759), .B2(n19877), .A(n14758), .ZN(P1_U2989) );
  NOR3_X1 U18072 ( .A1(n14798), .A2(n14780), .A3(n14760), .ZN(n14762) );
  OAI21_X1 U18073 ( .B1(n14762), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14761), .ZN(n14763) );
  OAI211_X1 U18074 ( .C1(n14765), .C2(n19993), .A(n14764), .B(n14763), .ZN(
        n14766) );
  INV_X1 U18075 ( .A(n14766), .ZN(n14767) );
  OAI21_X1 U18076 ( .B1(n14768), .B2(n16120), .A(n14767), .ZN(P1_U3001) );
  AND2_X1 U18077 ( .A1(n14769), .A2(n14780), .ZN(n14771) );
  OAI22_X1 U18078 ( .A1(n14772), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n14771), .B2(n14770), .ZN(n14773) );
  OAI211_X1 U18079 ( .C1(n14775), .C2(n19993), .A(n14774), .B(n14773), .ZN(
        n14776) );
  INV_X1 U18080 ( .A(n14776), .ZN(n14777) );
  OAI21_X1 U18081 ( .B1(n14778), .B2(n16120), .A(n14777), .ZN(P1_U3002) );
  INV_X1 U18082 ( .A(n14779), .ZN(n14787) );
  INV_X1 U18083 ( .A(n14780), .ZN(n14782) );
  NOR3_X1 U18084 ( .A1(n14798), .A2(n14782), .A3(n14781), .ZN(n14786) );
  OAI21_X1 U18085 ( .B1(n14791), .B2(n14784), .A(n14783), .ZN(n14785) );
  AOI211_X1 U18086 ( .C1(n14787), .C2(n20021), .A(n14786), .B(n14785), .ZN(
        n14788) );
  OAI21_X1 U18087 ( .B1(n14789), .B2(n16120), .A(n14788), .ZN(P1_U3003) );
  NAND2_X1 U18088 ( .A1(n14790), .A2(n20013), .ZN(n14797) );
  INV_X1 U18089 ( .A(n14791), .ZN(n14795) );
  NOR2_X1 U18090 ( .A1(n14792), .A2(n19993), .ZN(n14793) );
  AOI211_X1 U18091 ( .C1(n14795), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14794), .B(n14793), .ZN(n14796) );
  OAI211_X1 U18092 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14798), .A(
        n14797), .B(n14796), .ZN(P1_U3004) );
  INV_X1 U18093 ( .A(n14822), .ZN(n14802) );
  NAND3_X1 U18094 ( .A1(n14802), .A2(n11471), .A3(n14803), .ZN(n14799) );
  OAI211_X1 U18095 ( .C1(n15915), .C2(n19993), .A(n14800), .B(n14799), .ZN(
        n14805) );
  NAND3_X1 U18096 ( .A1(n14802), .A2(n14801), .A3(n11467), .ZN(n14811) );
  AOI21_X1 U18097 ( .B1(n14811), .B2(n14809), .A(n14803), .ZN(n14804) );
  NOR2_X1 U18098 ( .A1(n14805), .A2(n14804), .ZN(n14806) );
  OAI21_X1 U18099 ( .B1(n14807), .B2(n16120), .A(n14806), .ZN(P1_U3005) );
  OAI21_X1 U18100 ( .B1(n14809), .B2(n11467), .A(n14808), .ZN(n14810) );
  AOI21_X1 U18101 ( .B1(n15923), .B2(n20021), .A(n14810), .ZN(n14812) );
  OAI211_X1 U18102 ( .C1(n14813), .C2(n16120), .A(n14812), .B(n14811), .ZN(
        P1_U3006) );
  INV_X1 U18103 ( .A(n14814), .ZN(n14815) );
  NOR2_X1 U18104 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14815), .ZN(
        n14816) );
  NAND2_X1 U18105 ( .A1(n14817), .A2(n14816), .ZN(n14841) );
  INV_X1 U18106 ( .A(n20009), .ZN(n14819) );
  OAI21_X1 U18107 ( .B1(n14841), .B2(n14819), .A(n14818), .ZN(n14821) );
  AOI21_X1 U18108 ( .B1(n14821), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14820), .ZN(n14824) );
  OR3_X1 U18109 ( .A1(n14822), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n20806), .ZN(n14823) );
  OAI211_X1 U18110 ( .C1(n14825), .C2(n19993), .A(n14824), .B(n14823), .ZN(
        n14826) );
  AOI21_X1 U18111 ( .B1(n14827), .B2(n20013), .A(n14826), .ZN(n14828) );
  INV_X1 U18112 ( .A(n14828), .ZN(P1_U3007) );
  INV_X1 U18113 ( .A(n14927), .ZN(n14840) );
  NAND2_X1 U18114 ( .A1(n14829), .A2(n20013), .ZN(n14839) );
  NOR2_X1 U18115 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  OR2_X1 U18116 ( .A1(n14833), .A2(n14832), .ZN(n15936) );
  AOI21_X1 U18117 ( .B1(n14835), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14834), .ZN(n14836) );
  OAI21_X1 U18118 ( .B1(n15936), .B2(n19993), .A(n14836), .ZN(n14837) );
  INV_X1 U18119 ( .A(n14837), .ZN(n14838) );
  OAI211_X1 U18120 ( .C1(n14841), .C2(n14840), .A(n14839), .B(n14838), .ZN(
        P1_U3008) );
  INV_X1 U18121 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14864) );
  INV_X1 U18122 ( .A(n14842), .ZN(n14849) );
  AND2_X1 U18123 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16082), .ZN(
        n14917) );
  INV_X1 U18124 ( .A(n14917), .ZN(n14843) );
  OR2_X1 U18125 ( .A1(n14916), .A2(n14843), .ZN(n14846) );
  INV_X1 U18126 ( .A(n14918), .ZN(n14844) );
  OR2_X1 U18127 ( .A1(n20018), .A2(n14844), .ZN(n14845) );
  AND2_X1 U18128 ( .A1(n14846), .A2(n14845), .ZN(n14913) );
  NOR2_X1 U18129 ( .A1(n14913), .A2(n14847), .ZN(n14869) );
  AOI21_X1 U18130 ( .B1(n14849), .B2(n14848), .A(n14869), .ZN(n16078) );
  NOR2_X1 U18131 ( .A1(n16078), .A2(n14850), .ZN(n14865) );
  INV_X1 U18132 ( .A(n14865), .ZN(n14851) );
  AOI21_X1 U18133 ( .B1(n14864), .B2(n11462), .A(n14851), .ZN(n14857) );
  OAI21_X1 U18134 ( .B1(n14861), .B2(n11462), .A(n14852), .ZN(n14855) );
  NOR2_X1 U18135 ( .A1(n14853), .A2(n19993), .ZN(n14854) );
  AOI211_X1 U18136 ( .C1(n14857), .C2(n14856), .A(n14855), .B(n14854), .ZN(
        n14858) );
  OAI21_X1 U18137 ( .B1(n14859), .B2(n16120), .A(n14858), .ZN(P1_U3009) );
  NAND2_X1 U18138 ( .A1(n14860), .A2(n20013), .ZN(n14867) );
  NOR2_X1 U18139 ( .A1(n14861), .A2(n14864), .ZN(n14862) );
  AOI211_X1 U18140 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14866) );
  OAI211_X1 U18141 ( .C1(n19993), .C2(n15945), .A(n14867), .B(n14866), .ZN(
        P1_U3010) );
  NAND2_X1 U18142 ( .A1(n14868), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14874) );
  INV_X1 U18143 ( .A(n14869), .ZN(n14870) );
  AOI21_X1 U18144 ( .B1(n14870), .B2(n14914), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14871) );
  OAI21_X1 U18145 ( .B1(n14871), .B2(n16073), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14873) );
  OAI211_X1 U18146 ( .C1(n16078), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14875) );
  AOI21_X1 U18147 ( .B1(n14876), .B2(n20021), .A(n14875), .ZN(n14877) );
  OAI21_X1 U18148 ( .B1(n14878), .B2(n16120), .A(n14877), .ZN(P1_U3011) );
  INV_X1 U18149 ( .A(n14879), .ZN(n14881) );
  OAI21_X1 U18150 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14885) );
  NAND2_X1 U18151 ( .A1(n14885), .A2(n14883), .ZN(n14884) );
  MUX2_X1 U18152 ( .A(n14885), .B(n14884), .S(n16052), .Z(n14886) );
  XOR2_X1 U18153 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n14886), .Z(
        n16040) );
  NAND2_X1 U18154 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14899) );
  NAND2_X1 U18155 ( .A1(n14927), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14907) );
  OAI21_X1 U18156 ( .B1(n14899), .B2(n14907), .A(n14887), .ZN(n14890) );
  INV_X1 U18157 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14888) );
  OAI22_X1 U18158 ( .A1(n15976), .A2(n19993), .B1(n19933), .B2(n14888), .ZN(
        n14889) );
  AOI21_X1 U18159 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14892) );
  OAI21_X1 U18160 ( .B1(n16040), .B2(n16120), .A(n14892), .ZN(P1_U3014) );
  AOI21_X1 U18161 ( .B1(n11457), .B2(n14883), .A(n14907), .ZN(n14900) );
  OAI21_X1 U18162 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14894), .A(
        n14893), .ZN(n14908) );
  NAND2_X1 U18163 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14908), .ZN(
        n14895) );
  OAI211_X1 U18164 ( .C1(n14897), .C2(n19993), .A(n14896), .B(n14895), .ZN(
        n14898) );
  AOI21_X1 U18165 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14901) );
  OAI21_X1 U18166 ( .B1(n14902), .B2(n16120), .A(n14901), .ZN(P1_U3015) );
  OAI21_X1 U18167 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(n14906) );
  INV_X1 U18168 ( .A(n14906), .ZN(n16045) );
  INV_X1 U18169 ( .A(n14907), .ZN(n14911) );
  AOI22_X1 U18170 ( .A1(n19952), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14908), .ZN(n14909) );
  OAI21_X1 U18171 ( .B1(n15987), .B2(n19993), .A(n14909), .ZN(n14910) );
  AOI21_X1 U18172 ( .B1(n14911), .B2(n11457), .A(n14910), .ZN(n14912) );
  OAI21_X1 U18173 ( .B1(n16045), .B2(n16120), .A(n14912), .ZN(P1_U3016) );
  NOR2_X1 U18174 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14913), .ZN(
        n16079) );
  NOR2_X1 U18175 ( .A1(n14915), .A2(n14914), .ZN(n16081) );
  OAI22_X1 U18176 ( .A1(n14918), .A2(n20018), .B1(n14917), .B2(n14916), .ZN(
        n14919) );
  NOR3_X1 U18177 ( .A1(n14920), .A2(n16081), .A3(n14919), .ZN(n16089) );
  INV_X1 U18178 ( .A(n16089), .ZN(n14922) );
  NOR2_X1 U18179 ( .A1(n19933), .A2(n20677), .ZN(n14921) );
  AOI221_X1 U18180 ( .B1(n16079), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n14922), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n14921), .ZN(
        n14923) );
  OAI21_X1 U18181 ( .B1(n19993), .B2(n14924), .A(n14923), .ZN(n14925) );
  AOI21_X1 U18182 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  OAI21_X1 U18183 ( .B1(n14929), .B2(n16120), .A(n14928), .ZN(P1_U3017) );
  NOR2_X1 U18184 ( .A1(n14931), .A2(n14930), .ZN(n14933) );
  NOR2_X1 U18185 ( .A1(n14933), .A2(n14932), .ZN(n16051) );
  NOR3_X1 U18186 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14934), .A3(
        n16123), .ZN(n14947) );
  NAND3_X1 U18187 ( .A1(n14935), .A2(n14937), .A3(n14733), .ZN(n16095) );
  NOR2_X1 U18188 ( .A1(n16095), .A2(n14936), .ZN(n14943) );
  INV_X1 U18189 ( .A(n14937), .ZN(n14938) );
  OAI21_X1 U18190 ( .B1(n14939), .B2(n14938), .A(n20011), .ZN(n14940) );
  OAI211_X1 U18191 ( .C1(n14942), .C2(n20018), .A(n14941), .B(n14940), .ZN(
        n16091) );
  OAI21_X1 U18192 ( .B1(n14943), .B2(n16091), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U18193 ( .A1(n16003), .A2(n20021), .B1(n19973), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U18194 ( .A1(n14945), .A2(n14944), .ZN(n14946) );
  NOR2_X1 U18195 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  OAI21_X1 U18196 ( .B1(n16051), .B2(n16120), .A(n14948), .ZN(P1_U3019) );
  NAND3_X1 U18197 ( .A1(n14949), .A2(n13492), .A3(n20013), .ZN(n14958) );
  INV_X1 U18198 ( .A(n14950), .ZN(n14954) );
  OAI21_X1 U18199 ( .B1(n14952), .B2(n20012), .A(n14951), .ZN(n14953) );
  AOI21_X1 U18200 ( .B1(n20021), .B2(n14954), .A(n14953), .ZN(n14957) );
  NAND3_X1 U18201 ( .A1(n16118), .A2(n20012), .A3(n14955), .ZN(n14956) );
  NAND3_X1 U18202 ( .A1(n14958), .A2(n14957), .A3(n14956), .ZN(P1_U3030) );
  OAI21_X1 U18203 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9631), .A(n20415), 
        .ZN(n14959) );
  OAI21_X1 U18204 ( .B1(n14960), .B2(n20449), .A(n14959), .ZN(n14961) );
  MUX2_X1 U18205 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14961), .S(
        n20028), .Z(P1_U3477) );
  INV_X1 U18206 ( .A(n20449), .ZN(n20520) );
  NOR3_X1 U18207 ( .A1(n14962), .A2(n13694), .A3(n10968), .ZN(n14963) );
  AOI211_X1 U18208 ( .C1(n20520), .C2(n14965), .A(n14964), .B(n14963), .ZN(
        n15853) );
  INV_X1 U18209 ( .A(n14966), .ZN(n14969) );
  NOR3_X1 U18210 ( .A1(n13694), .A2(n10968), .A3(n15880), .ZN(n14967) );
  AOI21_X1 U18211 ( .B1(n14969), .B2(n14968), .A(n14967), .ZN(n14970) );
  OAI21_X1 U18212 ( .B1(n15853), .B2(n14971), .A(n14970), .ZN(n14972) );
  MUX2_X1 U18213 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14972), .S(
        n20727), .Z(P1_U3473) );
  OAI21_X1 U18214 ( .B1(n15080), .B2(n14973), .A(n15064), .ZN(n15380) );
  AOI21_X1 U18215 ( .B1(n9676), .B2(n14975), .A(n14974), .ZN(n14976) );
  NAND2_X1 U18216 ( .A1(n14976), .A2(n19042), .ZN(n14985) );
  AOI21_X1 U18217 ( .B1(n14978), .B2(n9674), .A(n14977), .ZN(n15378) );
  NAND2_X1 U18218 ( .A1(n15378), .A2(n19055), .ZN(n14980) );
  AOI22_X1 U18219 ( .A1(n19036), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n19048), .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n14979) );
  OAI211_X1 U18220 ( .C1(n19032), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n14982) );
  AOI21_X1 U18221 ( .B1(n14983), .B2(n12367), .A(n14982), .ZN(n14984) );
  OAI211_X1 U18222 ( .C1(n19057), .C2(n15380), .A(n14985), .B(n14984), .ZN(
        P2_U2827) );
  AOI21_X1 U18223 ( .B1(n14987), .B2(n15229), .A(n14986), .ZN(n15000) );
  OR2_X1 U18224 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  NAND2_X1 U18225 ( .A1(n14988), .A2(n14991), .ZN(n15404) );
  INV_X1 U18226 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U18227 ( .A1(n14992), .A2(n12367), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19036), .ZN(n14993) );
  OAI21_X1 U18228 ( .B1(n19773), .B2(n19030), .A(n14993), .ZN(n14994) );
  AOI21_X1 U18229 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n19049), .A(n14994), .ZN(
        n14998) );
  AND2_X1 U18230 ( .A1(n15009), .A2(n14995), .ZN(n14996) );
  NOR2_X1 U18231 ( .A1(n15078), .A2(n14996), .ZN(n15403) );
  NAND2_X1 U18232 ( .A1(n15403), .A2(n19041), .ZN(n14997) );
  OAI211_X1 U18233 ( .C1(n15404), .C2(n19046), .A(n14998), .B(n14997), .ZN(
        n14999) );
  AOI21_X1 U18234 ( .B1(n15000), .B2(n19042), .A(n14999), .ZN(n15001) );
  INV_X1 U18235 ( .A(n15001), .ZN(P2_U2829) );
  AOI211_X1 U18236 ( .C1(n15235), .C2(n15003), .A(n15002), .B(n19724), .ZN(
        n15015) );
  INV_X1 U18237 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U18238 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19049), .ZN(n15007) );
  OAI211_X1 U18239 ( .C1(n15018), .C2(n15005), .A(n15004), .B(n12367), .ZN(
        n15006) );
  OAI211_X1 U18240 ( .C1(n19030), .C2(n19771), .A(n15007), .B(n15006), .ZN(
        n15014) );
  INV_X1 U18241 ( .A(n15009), .ZN(n15010) );
  AOI21_X1 U18242 ( .B1(n15011), .B2(n15008), .A(n15010), .ZN(n15424) );
  INV_X1 U18243 ( .A(n15424), .ZN(n15095) );
  XNOR2_X1 U18244 ( .A(n15025), .B(n15012), .ZN(n15419) );
  OAI22_X1 U18245 ( .A1(n15095), .A2(n19057), .B1(n15419), .B2(n19046), .ZN(
        n15013) );
  OR3_X1 U18246 ( .A1(n15015), .A2(n15014), .A3(n15013), .ZN(P2_U2830) );
  AOI211_X1 U18247 ( .C1(n15256), .C2(n15016), .A(n15017), .B(n19724), .ZN(
        n15031) );
  AOI211_X1 U18248 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n10466), .A(n19052), .B(
        n15018), .ZN(n15030) );
  OR2_X1 U18249 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  NAND2_X1 U18250 ( .A1(n15008), .A2(n15021), .ZN(n15438) );
  NAND2_X1 U18251 ( .A1(n15023), .A2(n15022), .ZN(n15024) );
  AND2_X1 U18252 ( .A1(n15025), .A2(n15024), .ZN(n15435) );
  AOI22_X1 U18253 ( .A1(n15435), .A2(n19055), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19049), .ZN(n15028) );
  OAI22_X1 U18254 ( .A1(n15253), .A2(n19030), .B1(n15254), .B2(n19060), .ZN(
        n15026) );
  INV_X1 U18255 ( .A(n15026), .ZN(n15027) );
  OAI211_X1 U18256 ( .C1(n15438), .C2(n19057), .A(n15028), .B(n15027), .ZN(
        n15029) );
  OR3_X1 U18257 ( .A1(n15031), .A2(n15030), .A3(n15029), .ZN(P2_U2831) );
  AOI211_X1 U18258 ( .C1(n15033), .C2(n15032), .A(n9748), .B(n19724), .ZN(
        n15034) );
  INV_X1 U18259 ( .A(n15034), .ZN(n15047) );
  NAND2_X1 U18260 ( .A1(n15036), .A2(n15035), .ZN(n15037) );
  AND2_X1 U18261 ( .A1(n15038), .A2(n15037), .ZN(n15465) );
  OR2_X1 U18262 ( .A1(n13060), .A2(n15039), .ZN(n15040) );
  NAND2_X1 U18263 ( .A1(n13073), .A2(n15040), .ZN(n16183) );
  INV_X1 U18264 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U18265 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19049), .ZN(n15041) );
  OAI21_X1 U18266 ( .B1(n19030), .B2(n15042), .A(n15041), .ZN(n15043) );
  AOI21_X1 U18267 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19036), .A(
        n15043), .ZN(n15044) );
  OAI21_X1 U18268 ( .B1(n16183), .B2(n19046), .A(n15044), .ZN(n15045) );
  AOI21_X1 U18269 ( .B1(n15465), .B2(n19041), .A(n15045), .ZN(n15046) );
  OAI211_X1 U18270 ( .C1(n19052), .C2(n15048), .A(n15047), .B(n15046), .ZN(
        P2_U2833) );
  AOI211_X1 U18271 ( .C1(n15051), .C2(n15050), .A(n15049), .B(n19724), .ZN(
        n15052) );
  INV_X1 U18272 ( .A(n15052), .ZN(n15059) );
  INV_X1 U18273 ( .A(n15053), .ZN(n15119) );
  AOI22_X1 U18274 ( .A1(n19049), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19048), .ZN(n15054) );
  INV_X1 U18275 ( .A(n15054), .ZN(n15055) );
  AOI21_X1 U18276 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19036), .A(
        n15055), .ZN(n15056) );
  OAI21_X1 U18277 ( .B1(n19046), .B2(n16190), .A(n15056), .ZN(n15057) );
  AOI21_X1 U18278 ( .B1(n15119), .B2(n19041), .A(n15057), .ZN(n15058) );
  OAI211_X1 U18279 ( .C1(n19052), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        P2_U2835) );
  INV_X1 U18280 ( .A(n15061), .ZN(n15062) );
  MUX2_X1 U18281 ( .A(n15062), .B(P2_EBX_REG_31__SCAN_IN), .S(n13579), .Z(
        P2_U2856) );
  AOI21_X1 U18282 ( .B1(n15065), .B2(n15064), .A(n15063), .ZN(n16158) );
  INV_X1 U18283 ( .A(n16158), .ZN(n15368) );
  INV_X1 U18284 ( .A(n15066), .ZN(n15133) );
  NAND2_X1 U18285 ( .A1(n15068), .A2(n15067), .ZN(n15132) );
  NAND3_X1 U18286 ( .A1(n15133), .A2(n15118), .A3(n15132), .ZN(n15070) );
  NAND2_X1 U18287 ( .A1(n13579), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15069) );
  OAI211_X1 U18288 ( .C1(n15368), .C2(n13579), .A(n15070), .B(n15069), .ZN(
        P2_U2858) );
  NAND2_X1 U18289 ( .A1(n15072), .A2(n15071), .ZN(n15074) );
  XNOR2_X1 U18290 ( .A(n15074), .B(n15073), .ZN(n15146) );
  NOR2_X1 U18291 ( .A1(n15380), .A2(n13579), .ZN(n15075) );
  AOI21_X1 U18292 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13579), .A(n15075), .ZN(
        n15076) );
  OAI21_X1 U18293 ( .B1(n15146), .B2(n15130), .A(n15076), .ZN(P2_U2859) );
  NOR2_X1 U18294 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  OR2_X1 U18295 ( .A1(n15080), .A2(n15079), .ZN(n16177) );
  AOI21_X1 U18296 ( .B1(n15083), .B2(n15082), .A(n15081), .ZN(n15147) );
  NAND2_X1 U18297 ( .A1(n15147), .A2(n15118), .ZN(n15085) );
  NAND2_X1 U18298 ( .A1(n13579), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15084) );
  OAI211_X1 U18299 ( .C1(n16177), .C2(n13579), .A(n15085), .B(n15084), .ZN(
        P2_U2860) );
  AOI21_X1 U18300 ( .B1(n15088), .B2(n15087), .A(n15086), .ZN(n15159) );
  NAND2_X1 U18301 ( .A1(n15159), .A2(n15118), .ZN(n15090) );
  NAND2_X1 U18302 ( .A1(n15403), .A2(n15123), .ZN(n15089) );
  OAI211_X1 U18303 ( .C1(n15123), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        P2_U2861) );
  OAI21_X1 U18304 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15165) );
  NOR2_X1 U18305 ( .A1(n15095), .A2(n13579), .ZN(n15096) );
  AOI21_X1 U18306 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n13579), .A(n15096), .ZN(
        n15097) );
  OAI21_X1 U18307 ( .B1(n15165), .B2(n15130), .A(n15097), .ZN(P2_U2862) );
  AOI21_X1 U18308 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15101) );
  XOR2_X1 U18309 ( .A(n15102), .B(n15101), .Z(n15170) );
  NOR2_X1 U18310 ( .A1(n15438), .A2(n13579), .ZN(n15103) );
  AOI21_X1 U18311 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n13579), .A(n15103), .ZN(
        n15104) );
  OAI21_X1 U18312 ( .B1(n15170), .B2(n15130), .A(n15104), .ZN(P2_U2863) );
  AOI21_X1 U18313 ( .B1(n15107), .B2(n15106), .A(n15105), .ZN(n15108) );
  INV_X1 U18314 ( .A(n15108), .ZN(n15177) );
  NAND2_X1 U18315 ( .A1(n13579), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15110) );
  NAND2_X1 U18316 ( .A1(n15451), .A2(n15123), .ZN(n15109) );
  OAI211_X1 U18317 ( .C1(n15177), .C2(n15130), .A(n15110), .B(n15109), .ZN(
        P2_U2864) );
  AOI21_X1 U18318 ( .B1(n15112), .B2(n14066), .A(n15111), .ZN(n16185) );
  NAND2_X1 U18319 ( .A1(n16185), .A2(n15118), .ZN(n15114) );
  NAND2_X1 U18320 ( .A1(n15465), .A2(n15123), .ZN(n15113) );
  OAI211_X1 U18321 ( .C1(n15123), .C2(n15115), .A(n15114), .B(n15113), .ZN(
        P2_U2865) );
  OR2_X1 U18322 ( .A1(n9686), .A2(n15116), .ZN(n15117) );
  AND2_X1 U18323 ( .A1(n14065), .A2(n15117), .ZN(n16193) );
  NAND2_X1 U18324 ( .A1(n16193), .A2(n15118), .ZN(n15121) );
  NAND2_X1 U18325 ( .A1(n15119), .A2(n15123), .ZN(n15120) );
  OAI211_X1 U18326 ( .C1(n15123), .C2(n15122), .A(n15121), .B(n15120), .ZN(
        P2_U2867) );
  AND2_X1 U18327 ( .A1(n15125), .A2(n15124), .ZN(n15127) );
  NOR2_X1 U18328 ( .A1(n18919), .A2(n13579), .ZN(n15128) );
  AOI21_X1 U18329 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n13579), .A(n15128), .ZN(
        n15129) );
  OAI21_X1 U18330 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(P2_U2868) );
  NAND3_X1 U18331 ( .A1(n15133), .A2(n19108), .A3(n15132), .ZN(n15141) );
  AOI22_X1 U18332 ( .A1(n19071), .A2(n15134), .B1(n19129), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15140) );
  AOI22_X1 U18333 ( .A1(n19073), .A2(BUF1_REG_29__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15139) );
  NOR2_X1 U18334 ( .A1(n14977), .A2(n15135), .ZN(n15136) );
  INV_X1 U18335 ( .A(n16164), .ZN(n15137) );
  NAND2_X1 U18336 ( .A1(n15137), .A2(n19130), .ZN(n15138) );
  NAND4_X1 U18337 ( .A1(n15141), .A2(n15140), .A3(n15139), .A4(n15138), .ZN(
        P2_U2890) );
  INV_X1 U18338 ( .A(n19071), .ZN(n15172) );
  INV_X1 U18339 ( .A(n19087), .ZN(n15142) );
  OAI22_X1 U18340 ( .A1(n15172), .A2(n15142), .B1(n19103), .B2(n13216), .ZN(
        n15143) );
  AOI21_X1 U18341 ( .B1(n15378), .B2(n19130), .A(n15143), .ZN(n15145) );
  AOI22_X1 U18342 ( .A1(n19073), .A2(BUF1_REG_28__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15144) );
  OAI211_X1 U18343 ( .C1(n15146), .C2(n19134), .A(n15145), .B(n15144), .ZN(
        P2_U2891) );
  NAND2_X1 U18344 ( .A1(n15147), .A2(n19108), .ZN(n15155) );
  AOI22_X1 U18345 ( .A1(n19071), .A2(n15148), .B1(n19129), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U18346 ( .A1(n19073), .A2(BUF1_REG_27__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U18347 ( .A1(n14988), .A2(n15149), .ZN(n15150) );
  NAND2_X1 U18348 ( .A1(n9674), .A2(n15150), .ZN(n16181) );
  INV_X1 U18349 ( .A(n16181), .ZN(n15151) );
  NAND2_X1 U18350 ( .A1(n15151), .A2(n19130), .ZN(n15152) );
  NAND4_X1 U18351 ( .A1(n15155), .A2(n15154), .A3(n15153), .A4(n15152), .ZN(
        P2_U2892) );
  AOI22_X1 U18352 ( .A1(n19073), .A2(BUF1_REG_26__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U18353 ( .A1(n19071), .A2(n19092), .B1(n19129), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15156) );
  OAI211_X1 U18354 ( .C1(n16191), .C2(n15404), .A(n15157), .B(n15156), .ZN(
        n15158) );
  AOI21_X1 U18355 ( .B1(n15159), .B2(n19108), .A(n15158), .ZN(n15160) );
  INV_X1 U18356 ( .A(n15160), .ZN(P2_U2893) );
  AOI22_X1 U18357 ( .A1(n19073), .A2(BUF1_REG_25__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U18358 ( .A1(n19071), .A2(n19095), .B1(n19129), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15161) );
  OAI211_X1 U18359 ( .C1(n15419), .C2(n16191), .A(n15162), .B(n15161), .ZN(
        n15163) );
  INV_X1 U18360 ( .A(n15163), .ZN(n15164) );
  OAI21_X1 U18361 ( .B1(n15165), .B2(n19134), .A(n15164), .ZN(P2_U2894) );
  INV_X1 U18362 ( .A(n19099), .ZN(n15166) );
  OAI22_X1 U18363 ( .A1(n15172), .A2(n15166), .B1(n19103), .B2(n13210), .ZN(
        n15167) );
  AOI21_X1 U18364 ( .B1(n19130), .B2(n15435), .A(n15167), .ZN(n15169) );
  AOI22_X1 U18365 ( .A1(n19073), .A2(BUF1_REG_24__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15168) );
  OAI211_X1 U18366 ( .C1(n15170), .C2(n19134), .A(n15169), .B(n15168), .ZN(
        P2_U2895) );
  INV_X1 U18367 ( .A(n15447), .ZN(n15174) );
  OAI22_X1 U18368 ( .A1(n15172), .A2(n19232), .B1(n15171), .B2(n19103), .ZN(
        n15173) );
  AOI21_X1 U18369 ( .B1(n19130), .B2(n15174), .A(n15173), .ZN(n15176) );
  AOI22_X1 U18370 ( .A1(n19073), .A2(BUF1_REG_23__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15175) );
  OAI211_X1 U18371 ( .C1(n15177), .C2(n19134), .A(n15176), .B(n15175), .ZN(
        P2_U2896) );
  INV_X1 U18372 ( .A(n19822), .ZN(n15640) );
  XNOR2_X1 U18373 ( .A(n19820), .B(n19822), .ZN(n19132) );
  NOR2_X1 U18374 ( .A1(n19827), .A2(n16317), .ZN(n19133) );
  NOR2_X1 U18375 ( .A1(n19132), .A2(n19133), .ZN(n19131) );
  AOI21_X1 U18376 ( .B1(n19817), .B2(n15640), .A(n19131), .ZN(n19123) );
  XNOR2_X1 U18377 ( .A(n15178), .B(n15179), .ZN(n19124) );
  NOR2_X1 U18378 ( .A1(n19123), .A2(n19124), .ZN(n19122) );
  AOI21_X1 U18379 ( .B1(n15179), .B2(n15178), .A(n19122), .ZN(n19116) );
  XNOR2_X1 U18380 ( .A(n15727), .B(n19805), .ZN(n19117) );
  NOR2_X1 U18381 ( .A1(n19116), .A2(n19117), .ZN(n19115) );
  NOR2_X1 U18382 ( .A1(n15727), .A2(n19805), .ZN(n15180) );
  OAI21_X1 U18383 ( .B1(n19115), .B2(n15180), .A(n15181), .ZN(n19110) );
  XOR2_X1 U18384 ( .A(n19107), .B(n19110), .Z(n15185) );
  INV_X1 U18385 ( .A(n15181), .ZN(n15182) );
  AOI22_X1 U18386 ( .A1(n19130), .A2(n15182), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19129), .ZN(n15184) );
  NAND2_X1 U18387 ( .A1(n19105), .A2(n16189), .ZN(n15183) );
  OAI211_X1 U18388 ( .C1(n15185), .C2(n19134), .A(n15184), .B(n15183), .ZN(
        P2_U2915) );
  INV_X1 U18389 ( .A(n15186), .ZN(n15187) );
  NOR2_X1 U18390 ( .A1(n15188), .A2(n15187), .ZN(n15190) );
  XOR2_X1 U18391 ( .A(n15190), .B(n15189), .Z(n15374) );
  NAND2_X1 U18392 ( .A1(n16258), .A2(n16154), .ZN(n15191) );
  NAND2_X1 U18393 ( .A1(n19176), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15367) );
  OAI211_X1 U18394 ( .C1(n15192), .C2(n19202), .A(n15191), .B(n15367), .ZN(
        n15193) );
  AOI21_X1 U18395 ( .B1(n16158), .B2(n19198), .A(n15193), .ZN(n15196) );
  AOI21_X1 U18396 ( .B1(n15210), .B2(n15364), .A(n15194), .ZN(n15371) );
  NAND2_X1 U18397 ( .A1(n15371), .A2(n9578), .ZN(n15195) );
  OAI211_X1 U18398 ( .C1(n15374), .C2(n19194), .A(n15196), .B(n15195), .ZN(
        P2_U2985) );
  NOR2_X1 U18399 ( .A1(n15197), .A2(n15198), .ZN(n15203) );
  INV_X1 U18400 ( .A(n15198), .ZN(n15200) );
  NAND2_X1 U18401 ( .A1(n10472), .A2(n15202), .ZN(n15199) );
  AND2_X1 U18402 ( .A1(n15200), .A2(n15199), .ZN(n15201) );
  AND2_X1 U18403 ( .A1(n15201), .A2(n9890), .ZN(n15215) );
  NAND2_X1 U18404 ( .A1(n15215), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15389) );
  OAI21_X1 U18405 ( .B1(n15203), .B2(n15202), .A(n15389), .ZN(n15206) );
  XNOR2_X1 U18406 ( .A(n15204), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15205) );
  XNOR2_X1 U18407 ( .A(n15206), .B(n15205), .ZN(n15387) );
  INV_X1 U18408 ( .A(n15380), .ZN(n15213) );
  NOR2_X1 U18409 ( .A1(n10856), .A2(n19776), .ZN(n15377) );
  AOI21_X1 U18410 ( .B1(n19177), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15377), .ZN(n15207) );
  OAI21_X1 U18411 ( .B1(n19191), .B2(n15208), .A(n15207), .ZN(n15212) );
  NOR2_X1 U18412 ( .A1(n15209), .A2(n15391), .ZN(n15401) );
  OAI21_X1 U18413 ( .B1(n15401), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15210), .ZN(n15381) );
  NOR2_X1 U18414 ( .A1(n15381), .A2(n19192), .ZN(n15211) );
  OAI21_X1 U18415 ( .B1(n15387), .B2(n19194), .A(n15214), .ZN(P2_U2986) );
  NAND2_X1 U18416 ( .A1(n15209), .A2(n15391), .ZN(n15388) );
  NAND2_X1 U18417 ( .A1(n15388), .A2(n9578), .ZN(n15221) );
  OR2_X1 U18418 ( .A1(n15215), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15390) );
  NAND3_X1 U18419 ( .A1(n15390), .A2(n19180), .A3(n15389), .ZN(n15220) );
  NAND2_X1 U18420 ( .A1(n19176), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15394) );
  OAI21_X1 U18421 ( .B1(n19202), .B2(n15216), .A(n15394), .ZN(n15218) );
  NOR2_X1 U18422 ( .A1(n16177), .A2(n19185), .ZN(n15217) );
  AOI211_X1 U18423 ( .C1(n16258), .C2(n16166), .A(n15218), .B(n15217), .ZN(
        n15219) );
  OAI211_X1 U18424 ( .C1(n15401), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        P2_U2987) );
  INV_X1 U18425 ( .A(n15222), .ZN(n15239) );
  NOR2_X1 U18426 ( .A1(n15223), .A2(n15239), .ZN(n15224) );
  XOR2_X1 U18427 ( .A(n15225), .B(n15224), .Z(n15417) );
  INV_X1 U18428 ( .A(n15209), .ZN(n15228) );
  AOI21_X1 U18429 ( .B1(n15226), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15227) );
  NOR2_X1 U18430 ( .A1(n15228), .A2(n15227), .ZN(n15415) );
  NAND2_X1 U18431 ( .A1(n15415), .A2(n9578), .ZN(n15234) );
  NAND2_X1 U18432 ( .A1(n16258), .A2(n15229), .ZN(n15230) );
  OR2_X1 U18433 ( .A1(n10856), .A2(n19773), .ZN(n15407) );
  OAI211_X1 U18434 ( .C1(n19202), .C2(n15231), .A(n15230), .B(n15407), .ZN(
        n15232) );
  AOI21_X1 U18435 ( .B1(n15403), .B2(n19198), .A(n15232), .ZN(n15233) );
  OAI211_X1 U18436 ( .C1(n15417), .C2(n19194), .A(n15234), .B(n15233), .ZN(
        P2_U2988) );
  XNOR2_X1 U18437 ( .A(n15226), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15431) );
  NAND2_X1 U18438 ( .A1(n16258), .A2(n15235), .ZN(n15236) );
  NAND2_X1 U18439 ( .A1(n19176), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18440 ( .C1(n19202), .C2(n15237), .A(n15236), .B(n15420), .ZN(
        n15245) );
  NOR2_X1 U18441 ( .A1(n15239), .A2(n15238), .ZN(n15243) );
  NAND2_X1 U18442 ( .A1(n15241), .A2(n15240), .ZN(n15242) );
  XOR2_X1 U18443 ( .A(n15243), .B(n15242), .Z(n15418) );
  NOR2_X1 U18444 ( .A1(n15418), .A2(n19194), .ZN(n15244) );
  AOI211_X1 U18445 ( .C1(n19198), .C2(n15424), .A(n15245), .B(n15244), .ZN(
        n15246) );
  OAI21_X1 U18446 ( .B1(n19192), .B2(n15431), .A(n15246), .ZN(P2_U2989) );
  INV_X1 U18447 ( .A(n15247), .ZN(n15248) );
  NAND2_X1 U18448 ( .A1(n15249), .A2(n15248), .ZN(n15252) );
  XNOR2_X1 U18449 ( .A(n15250), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15251) );
  XNOR2_X1 U18450 ( .A(n15252), .B(n15251), .ZN(n15443) );
  AOI21_X1 U18451 ( .B1(n15402), .B2(n9655), .A(n15226), .ZN(n15432) );
  NOR2_X1 U18452 ( .A1(n10856), .A2(n15253), .ZN(n15433) );
  NOR2_X1 U18453 ( .A1(n19202), .A2(n15254), .ZN(n15255) );
  AOI211_X1 U18454 ( .C1(n15256), .C2(n16258), .A(n15433), .B(n15255), .ZN(
        n15257) );
  OAI21_X1 U18455 ( .B1(n15438), .B2(n19185), .A(n15257), .ZN(n15258) );
  AOI21_X1 U18456 ( .B1(n15432), .B2(n9578), .A(n15258), .ZN(n15259) );
  OAI21_X1 U18457 ( .B1(n15443), .B2(n19194), .A(n15259), .ZN(P2_U2990) );
  NOR2_X1 U18458 ( .A1(n15280), .A2(n15461), .ZN(n15279) );
  OAI21_X1 U18459 ( .B1(n15279), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9655), .ZN(n15455) );
  NAND2_X1 U18460 ( .A1(n16258), .A2(n15260), .ZN(n15261) );
  NAND2_X1 U18461 ( .A1(n19176), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15446) );
  OAI211_X1 U18462 ( .C1(n19202), .C2(n15262), .A(n15261), .B(n15446), .ZN(
        n15270) );
  OR2_X1 U18463 ( .A1(n15334), .A2(n15264), .ZN(n15266) );
  NAND2_X1 U18464 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  XNOR2_X1 U18465 ( .A(n15268), .B(n15267), .ZN(n15452) );
  NOR2_X1 U18466 ( .A1(n15452), .A2(n19194), .ZN(n15269) );
  AOI211_X1 U18467 ( .C1(n19198), .C2(n15451), .A(n15270), .B(n15269), .ZN(
        n15271) );
  OAI21_X1 U18468 ( .B1(n15455), .B2(n19192), .A(n15271), .ZN(P2_U2991) );
  NAND2_X1 U18469 ( .A1(n15273), .A2(n15272), .ZN(n15278) );
  OR2_X1 U18470 ( .A1(n15334), .A2(n15274), .ZN(n15276) );
  NAND2_X1 U18471 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  XOR2_X1 U18472 ( .A(n15278), .B(n15277), .Z(n15468) );
  INV_X1 U18473 ( .A(n15279), .ZN(n15457) );
  NAND2_X1 U18474 ( .A1(n15280), .A2(n15461), .ZN(n15456) );
  NAND3_X1 U18475 ( .A1(n15457), .A2(n9578), .A3(n15456), .ZN(n15285) );
  NAND2_X1 U18476 ( .A1(n19176), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15460) );
  NAND2_X1 U18477 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15281) );
  OAI211_X1 U18478 ( .C1(n19191), .C2(n15282), .A(n15460), .B(n15281), .ZN(
        n15283) );
  AOI21_X1 U18479 ( .B1(n15465), .B2(n19198), .A(n15283), .ZN(n15284) );
  OAI211_X1 U18480 ( .C1(n15468), .C2(n19194), .A(n15285), .B(n15284), .ZN(
        P2_U2992) );
  NAND2_X1 U18481 ( .A1(n15287), .A2(n15286), .ZN(n15289) );
  AOI21_X1 U18482 ( .B1(n15298), .B2(n15296), .A(n15295), .ZN(n15288) );
  XOR2_X1 U18483 ( .A(n15289), .B(n15288), .Z(n15478) );
  XNOR2_X1 U18484 ( .A(n15299), .B(n15471), .ZN(n15476) );
  INV_X1 U18485 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19761) );
  NOR2_X1 U18486 ( .A1(n10856), .A2(n19761), .ZN(n15470) );
  NOR2_X1 U18487 ( .A1(n19202), .A2(n15290), .ZN(n15291) );
  AOI211_X1 U18488 ( .C1(n18916), .C2(n16258), .A(n15470), .B(n15291), .ZN(
        n15292) );
  OAI21_X1 U18489 ( .B1(n19185), .B2(n18919), .A(n15292), .ZN(n15293) );
  AOI21_X1 U18490 ( .B1(n15476), .B2(n9578), .A(n15293), .ZN(n15294) );
  OAI21_X1 U18491 ( .B1(n15478), .B2(n19194), .A(n15294), .ZN(P2_U2995) );
  NAND2_X1 U18492 ( .A1(n14180), .A2(n15296), .ZN(n15297) );
  XNOR2_X1 U18493 ( .A(n15298), .B(n15297), .ZN(n15489) );
  AOI21_X1 U18494 ( .B1(n15492), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15300) );
  NOR2_X1 U18495 ( .A1(n15300), .A2(n15299), .ZN(n15487) );
  INV_X1 U18496 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19759) );
  NOR2_X1 U18497 ( .A1(n10856), .A2(n19759), .ZN(n15482) );
  NOR2_X1 U18498 ( .A1(n19191), .A2(n18936), .ZN(n15301) );
  AOI211_X1 U18499 ( .C1(n19177), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15482), .B(n15301), .ZN(n15302) );
  OAI21_X1 U18500 ( .B1(n19185), .B2(n18934), .A(n15302), .ZN(n15303) );
  AOI21_X1 U18501 ( .B1(n15487), .B2(n9578), .A(n15303), .ZN(n15304) );
  OAI21_X1 U18502 ( .B1(n15489), .B2(n19194), .A(n15304), .ZN(P2_U2996) );
  XNOR2_X1 U18503 ( .A(n15492), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15312) );
  XNOR2_X1 U18504 ( .A(n15305), .B(n15306), .ZN(n15499) );
  NAND2_X1 U18505 ( .A1(n15499), .A2(n19180), .ZN(n15311) );
  INV_X1 U18506 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19757) );
  NOR2_X1 U18507 ( .A1(n19757), .A2(n18941), .ZN(n15309) );
  OAI22_X1 U18508 ( .A1(n19202), .A2(n15307), .B1(n19191), .B2(n18950), .ZN(
        n15308) );
  AOI211_X1 U18509 ( .C1(n18945), .C2(n19198), .A(n15309), .B(n15308), .ZN(
        n15310) );
  OAI211_X1 U18510 ( .C1(n19192), .C2(n15312), .A(n15311), .B(n15310), .ZN(
        P2_U2997) );
  XNOR2_X1 U18511 ( .A(n15314), .B(n15313), .ZN(n15521) );
  INV_X1 U18512 ( .A(n15514), .ZN(n18961) );
  NOR2_X1 U18513 ( .A1(n15513), .A2(n18941), .ZN(n15316) );
  OAI22_X1 U18514 ( .A1(n19202), .A2(n10804), .B1(n19191), .B2(n18956), .ZN(
        n15315) );
  AOI211_X1 U18515 ( .C1(n19198), .C2(n18961), .A(n15316), .B(n15315), .ZN(
        n15320) );
  INV_X1 U18516 ( .A(n15317), .ZN(n15501) );
  INV_X1 U18517 ( .A(n15492), .ZN(n15318) );
  OAI211_X1 U18518 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15501), .A(
        n15318), .B(n9578), .ZN(n15319) );
  OAI211_X1 U18519 ( .C1(n15521), .C2(n19194), .A(n15320), .B(n15319), .ZN(
        P2_U2998) );
  NAND2_X1 U18520 ( .A1(n15322), .A2(n15321), .ZN(n15324) );
  XOR2_X1 U18521 ( .A(n15324), .B(n15323), .Z(n16275) );
  XNOR2_X1 U18522 ( .A(n14193), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16272) );
  INV_X1 U18523 ( .A(n18971), .ZN(n15325) );
  OAI22_X1 U18524 ( .A1(n19202), .A2(n10801), .B1(n19191), .B2(n15325), .ZN(
        n15329) );
  OAI22_X1 U18525 ( .A1(n19185), .A2(n15327), .B1(n10856), .B2(n15326), .ZN(
        n15328) );
  AOI211_X1 U18526 ( .C1(n16272), .C2(n9578), .A(n15329), .B(n15328), .ZN(
        n15330) );
  OAI21_X1 U18527 ( .B1(n16275), .B2(n19194), .A(n15330), .ZN(P2_U2999) );
  NAND2_X1 U18528 ( .A1(n15332), .A2(n15331), .ZN(n15333) );
  XNOR2_X1 U18529 ( .A(n15334), .B(n15333), .ZN(n15535) );
  NAND2_X1 U18530 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15335), .ZN(
        n15536) );
  INV_X1 U18531 ( .A(n16282), .ZN(n15523) );
  OR2_X1 U18532 ( .A1(n10856), .A2(n15336), .ZN(n15526) );
  OAI21_X1 U18533 ( .B1(n19192), .B2(n15337), .A(n15526), .ZN(n15340) );
  OAI22_X1 U18534 ( .A1(n19202), .A2(n10795), .B1(n19191), .B2(n15338), .ZN(
        n15339) );
  OAI21_X1 U18535 ( .B1(n15535), .B2(n19194), .A(n15341), .ZN(P2_U3001) );
  NAND2_X1 U18536 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15343) );
  NAND2_X1 U18537 ( .A1(n15343), .A2(n15342), .ZN(n16243) );
  AND2_X1 U18538 ( .A1(n15345), .A2(n15344), .ZN(n15346) );
  NAND2_X1 U18539 ( .A1(n16243), .A2(n15346), .ZN(n15347) );
  XNOR2_X1 U18540 ( .A(n15347), .B(n16304), .ZN(n15599) );
  NAND2_X1 U18541 ( .A1(n10361), .A2(n16237), .ZN(n15349) );
  XNOR2_X1 U18542 ( .A(n15348), .B(n15349), .ZN(n15597) );
  OAI22_X1 U18543 ( .A1(n19202), .A2(n15350), .B1(n10771), .B2(n10856), .ZN(
        n15351) );
  AOI21_X1 U18544 ( .B1(n16258), .B2(n19008), .A(n15351), .ZN(n15352) );
  OAI21_X1 U18545 ( .B1(n19013), .B2(n19185), .A(n15352), .ZN(n15353) );
  AOI21_X1 U18546 ( .B1(n15597), .B2(n19180), .A(n15353), .ZN(n15354) );
  OAI21_X1 U18547 ( .B1(n15599), .B2(n19192), .A(n15354), .ZN(P2_U3007) );
  XNOR2_X1 U18548 ( .A(n15355), .B(n15356), .ZN(n15601) );
  XNOR2_X1 U18549 ( .A(n15358), .B(n15357), .ZN(n15600) );
  NAND2_X1 U18550 ( .A1(n15600), .A2(n9578), .ZN(n15362) );
  OAI22_X1 U18551 ( .A1(n10767), .A2(n10856), .B1(n19191), .B2(n19024), .ZN(
        n15360) );
  NOR2_X1 U18552 ( .A1(n19202), .A2(n9739), .ZN(n15359) );
  AOI211_X1 U18553 ( .C1(n15609), .C2(n19198), .A(n15360), .B(n15359), .ZN(
        n15361) );
  OAI211_X1 U18554 ( .C1(n19194), .C2(n15601), .A(n15362), .B(n15361), .ZN(
        P2_U3008) );
  OAI21_X1 U18555 ( .B1(n15365), .B2(n15376), .A(n15363), .ZN(n15385) );
  INV_X1 U18556 ( .A(n15376), .ZN(n15392) );
  NAND3_X1 U18557 ( .A1(n15392), .A2(n15365), .A3(n15364), .ZN(n15366) );
  OAI211_X1 U18558 ( .C1(n16164), .C2(n16318), .A(n15367), .B(n15366), .ZN(
        n15370) );
  NOR2_X1 U18559 ( .A1(n15368), .A2(n16319), .ZN(n15369) );
  NAND2_X1 U18560 ( .A1(n15371), .A2(n16295), .ZN(n15372) );
  OAI211_X1 U18561 ( .C1(n15374), .C2(n16299), .A(n15373), .B(n15372), .ZN(
        P2_U3017) );
  OAI21_X1 U18562 ( .B1(n15376), .B2(n15391), .A(n15375), .ZN(n15384) );
  AOI21_X1 U18563 ( .B1(n15378), .B2(n16307), .A(n15377), .ZN(n15379) );
  OAI21_X1 U18564 ( .B1(n15380), .B2(n16319), .A(n15379), .ZN(n15383) );
  NOR2_X1 U18565 ( .A1(n15381), .A2(n16330), .ZN(n15382) );
  OAI21_X1 U18566 ( .B1(n15387), .B2(n16299), .A(n15386), .ZN(P2_U3018) );
  NAND2_X1 U18567 ( .A1(n15388), .A2(n16295), .ZN(n15400) );
  NAND3_X1 U18568 ( .A1(n15390), .A2(n16326), .A3(n15389), .ZN(n15399) );
  NAND2_X1 U18569 ( .A1(n15392), .A2(n15391), .ZN(n15393) );
  OAI211_X1 U18570 ( .C1(n16181), .C2(n16318), .A(n15394), .B(n15393), .ZN(
        n15396) );
  NOR2_X1 U18571 ( .A1(n16177), .A2(n16319), .ZN(n15395) );
  AOI211_X1 U18572 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15397), .A(
        n15396), .B(n15395), .ZN(n15398) );
  OAI211_X1 U18573 ( .C1(n15401), .C2(n15400), .A(n15399), .B(n15398), .ZN(
        P2_U3019) );
  AND2_X1 U18574 ( .A1(n15405), .A2(n15402), .ZN(n15434) );
  NOR2_X1 U18575 ( .A1(n15440), .A2(n15434), .ZN(n15427) );
  NAND2_X1 U18576 ( .A1(n15403), .A2(n16294), .ZN(n15412) );
  INV_X1 U18577 ( .A(n15404), .ZN(n15410) );
  NAND2_X1 U18578 ( .A1(n15405), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15421) );
  OAI21_X1 U18579 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15406), .ZN(n15408) );
  OAI21_X1 U18580 ( .B1(n15421), .B2(n15408), .A(n15407), .ZN(n15409) );
  AOI21_X1 U18581 ( .B1(n16307), .B2(n15410), .A(n15409), .ZN(n15411) );
  OAI211_X1 U18582 ( .C1(n15427), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        n15414) );
  AOI21_X1 U18583 ( .B1(n15415), .B2(n16295), .A(n15414), .ZN(n15416) );
  OAI21_X1 U18584 ( .B1(n15417), .B2(n16299), .A(n15416), .ZN(P2_U3020) );
  INV_X1 U18585 ( .A(n15418), .ZN(n15429) );
  NOR2_X1 U18586 ( .A1(n16318), .A2(n15419), .ZN(n15423) );
  OAI21_X1 U18587 ( .B1(n15421), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15420), .ZN(n15422) );
  AOI211_X1 U18588 ( .C1(n15424), .C2(n16294), .A(n15423), .B(n15422), .ZN(
        n15425) );
  OAI21_X1 U18589 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15428) );
  AOI21_X1 U18590 ( .B1(n15429), .B2(n16326), .A(n15428), .ZN(n15430) );
  OAI21_X1 U18591 ( .B1(n15431), .B2(n16330), .A(n15430), .ZN(P2_U3021) );
  NAND2_X1 U18592 ( .A1(n15432), .A2(n16295), .ZN(n15442) );
  NOR2_X1 U18593 ( .A1(n15434), .A2(n15433), .ZN(n15437) );
  NAND2_X1 U18594 ( .A1(n16307), .A2(n15435), .ZN(n15436) );
  OAI211_X1 U18595 ( .C1(n15438), .C2(n16319), .A(n15437), .B(n15436), .ZN(
        n15439) );
  AOI21_X1 U18596 ( .B1(n15440), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15439), .ZN(n15441) );
  OAI211_X1 U18597 ( .C1(n15443), .C2(n16299), .A(n15442), .B(n15441), .ZN(
        P2_U3022) );
  OAI211_X1 U18598 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15458), .B(n15444), .ZN(
        n15445) );
  OAI211_X1 U18599 ( .C1(n16318), .C2(n15447), .A(n15446), .B(n15445), .ZN(
        n15450) );
  INV_X1 U18600 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15448) );
  NOR2_X1 U18601 ( .A1(n15462), .A2(n15448), .ZN(n15449) );
  AOI211_X1 U18602 ( .C1(n15451), .C2(n16294), .A(n15450), .B(n15449), .ZN(
        n15454) );
  OR2_X1 U18603 ( .A1(n15452), .A2(n16299), .ZN(n15453) );
  OAI211_X1 U18604 ( .C1(n15455), .C2(n16330), .A(n15454), .B(n15453), .ZN(
        P2_U3023) );
  NAND3_X1 U18605 ( .A1(n15457), .A2(n16295), .A3(n15456), .ZN(n15467) );
  NAND2_X1 U18606 ( .A1(n15458), .A2(n15461), .ZN(n15459) );
  OAI211_X1 U18607 ( .C1(n16318), .C2(n16183), .A(n15460), .B(n15459), .ZN(
        n15464) );
  NOR2_X1 U18608 ( .A1(n15462), .A2(n15461), .ZN(n15463) );
  AOI211_X1 U18609 ( .C1(n15465), .C2(n16294), .A(n15464), .B(n15463), .ZN(
        n15466) );
  OAI211_X1 U18610 ( .C1(n15468), .C2(n16299), .A(n15467), .B(n15466), .ZN(
        P2_U3024) );
  NAND2_X1 U18611 ( .A1(n15479), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15474) );
  NOR2_X1 U18612 ( .A1(n16318), .A2(n18926), .ZN(n15469) );
  AOI211_X1 U18613 ( .C1(n15472), .C2(n15471), .A(n15470), .B(n15469), .ZN(
        n15473) );
  OAI211_X1 U18614 ( .C1(n18919), .C2(n16319), .A(n15474), .B(n15473), .ZN(
        n15475) );
  AOI21_X1 U18615 ( .B1(n15476), .B2(n16295), .A(n15475), .ZN(n15477) );
  OAI21_X1 U18616 ( .B1(n15478), .B2(n16299), .A(n15477), .ZN(P2_U3027) );
  NAND2_X1 U18617 ( .A1(n15479), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15485) );
  INV_X1 U18618 ( .A(n18939), .ZN(n15483) );
  NOR2_X1 U18619 ( .A1(n15480), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15481) );
  AOI211_X1 U18620 ( .C1(n16307), .C2(n15483), .A(n15482), .B(n15481), .ZN(
        n15484) );
  OAI211_X1 U18621 ( .C1(n18934), .C2(n16319), .A(n15485), .B(n15484), .ZN(
        n15486) );
  AOI21_X1 U18622 ( .B1(n15487), .B2(n16295), .A(n15486), .ZN(n15488) );
  OAI21_X1 U18623 ( .B1(n15489), .B2(n16299), .A(n15488), .ZN(P2_U3028) );
  AND2_X1 U18624 ( .A1(n16330), .A2(n15490), .ZN(n15491) );
  OR2_X1 U18625 ( .A1(n15492), .A2(n15491), .ZN(n15498) );
  AND2_X1 U18626 ( .A1(n16322), .A2(n9785), .ZN(n15494) );
  OR2_X1 U18627 ( .A1(n15562), .A2(n15494), .ZN(n16271) );
  NOR2_X1 U18628 ( .A1(n15495), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15496) );
  NOR2_X1 U18629 ( .A1(n16271), .A2(n15496), .ZN(n15497) );
  NAND2_X1 U18630 ( .A1(n15498), .A2(n15497), .ZN(n15519) );
  AOI21_X1 U18631 ( .B1(n15502), .B2(n16322), .A(n15519), .ZN(n15508) );
  NAND2_X1 U18632 ( .A1(n15499), .A2(n16326), .ZN(n15506) );
  OAI22_X1 U18633 ( .A1(n16318), .A2(n18954), .B1(n10856), .B2(n19757), .ZN(
        n15504) );
  INV_X1 U18634 ( .A(n16268), .ZN(n15500) );
  AOI22_X1 U18635 ( .A1(n15501), .A2(n16295), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15500), .ZN(n15517) );
  NOR3_X1 U18636 ( .A1(n15517), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15502), .ZN(n15503) );
  AOI211_X1 U18637 ( .C1(n18945), .C2(n16294), .A(n15504), .B(n15503), .ZN(
        n15505) );
  OAI211_X1 U18638 ( .C1(n15508), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        P2_U3029) );
  NOR2_X1 U18639 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  NOR2_X1 U18640 ( .A1(n15512), .A2(n15511), .ZN(n19074) );
  OAI22_X1 U18641 ( .A1(n16319), .A2(n15514), .B1(n18941), .B2(n15513), .ZN(
        n15515) );
  AOI21_X1 U18642 ( .B1(n16307), .B2(n19074), .A(n15515), .ZN(n15516) );
  OAI21_X1 U18643 ( .B1(n15517), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15516), .ZN(n15518) );
  AOI21_X1 U18644 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15519), .A(
        n15518), .ZN(n15520) );
  OAI21_X1 U18645 ( .B1(n15521), .B2(n16299), .A(n15520), .ZN(P2_U3030) );
  AND2_X1 U18646 ( .A1(n15522), .A2(n15579), .ZN(n16281) );
  OAI211_X1 U18647 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n16281), .B(n15523), .ZN(
        n15534) );
  AND2_X1 U18648 ( .A1(n16322), .A2(n15524), .ZN(n15525) );
  OR2_X1 U18649 ( .A1(n15562), .A2(n15525), .ZN(n16276) );
  INV_X1 U18650 ( .A(n15526), .ZN(n15527) );
  AOI21_X1 U18651 ( .B1(n16294), .B2(n15528), .A(n15527), .ZN(n15531) );
  NAND2_X1 U18652 ( .A1(n16295), .A2(n15529), .ZN(n15530) );
  OAI211_X1 U18653 ( .C1(n16318), .C2(n19086), .A(n15531), .B(n15530), .ZN(
        n15532) );
  AOI21_X1 U18654 ( .B1(n16276), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15532), .ZN(n15533) );
  OAI211_X1 U18655 ( .C1(n15535), .C2(n16299), .A(n15534), .B(n15533), .ZN(
        P2_U3033) );
  INV_X1 U18656 ( .A(n15536), .ZN(n15537) );
  AOI21_X1 U18657 ( .B1(n15555), .B2(n15539), .A(n15537), .ZN(n16206) );
  NAND2_X1 U18658 ( .A1(n16206), .A2(n16295), .ZN(n15553) );
  NOR2_X1 U18659 ( .A1(n10792), .A2(n18941), .ZN(n15538) );
  AOI221_X1 U18660 ( .B1(n16281), .B2(n15539), .C1(n16276), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15538), .ZN(n15552) );
  XNOR2_X1 U18661 ( .A(n15540), .B(n15541), .ZN(n19089) );
  INV_X1 U18662 ( .A(n19089), .ZN(n15542) );
  AOI22_X1 U18663 ( .A1(n16307), .A2(n15542), .B1(n16294), .B2(n18982), .ZN(
        n15551) );
  NAND2_X1 U18664 ( .A1(n15557), .A2(n15559), .ZN(n15545) );
  INV_X1 U18665 ( .A(n15543), .ZN(n15544) );
  NAND2_X1 U18666 ( .A1(n15545), .A2(n15544), .ZN(n15549) );
  OR2_X1 U18667 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  XNOR2_X1 U18668 ( .A(n15549), .B(n15548), .ZN(n16207) );
  NAND2_X1 U18669 ( .A1(n16207), .A2(n16326), .ZN(n15550) );
  NAND4_X1 U18670 ( .A1(n15553), .A2(n15552), .A3(n15551), .A4(n15550), .ZN(
        P2_U3034) );
  INV_X1 U18671 ( .A(n15554), .ZN(n16215) );
  OAI21_X1 U18672 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16215), .A(
        n15555), .ZN(n16211) );
  NAND2_X1 U18673 ( .A1(n16219), .A2(n16217), .ZN(n15556) );
  OR2_X1 U18674 ( .A1(n15557), .A2(n15556), .ZN(n15561) );
  AND2_X1 U18675 ( .A1(n15559), .A2(n15558), .ZN(n15560) );
  XNOR2_X1 U18676 ( .A(n15561), .B(n15560), .ZN(n16210) );
  AOI21_X1 U18677 ( .B1(n15563), .B2(n15579), .A(n15562), .ZN(n16288) );
  INV_X1 U18678 ( .A(n16288), .ZN(n15580) );
  NOR2_X1 U18679 ( .A1(n10779), .A2(n18941), .ZN(n15566) );
  NAND2_X1 U18680 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15579), .ZN(
        n16290) );
  AOI221_X1 U18681 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n16289), .C2(n15564), .A(
        n16290), .ZN(n15565) );
  AOI211_X1 U18682 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15580), .A(
        n15566), .B(n15565), .ZN(n15571) );
  OAI21_X1 U18683 ( .B1(n15568), .B2(n15567), .A(n15540), .ZN(n19091) );
  INV_X1 U18684 ( .A(n19091), .ZN(n15569) );
  AOI22_X1 U18685 ( .A1(n16307), .A2(n15569), .B1(n16294), .B2(n18991), .ZN(
        n15570) );
  OAI211_X1 U18686 ( .C1(n16210), .C2(n16299), .A(n15571), .B(n15570), .ZN(
        n15572) );
  INV_X1 U18687 ( .A(n15572), .ZN(n15573) );
  OAI21_X1 U18688 ( .B1(n16211), .B2(n16330), .A(n15573), .ZN(P2_U3035) );
  INV_X1 U18689 ( .A(n15574), .ZN(n16216) );
  OAI21_X1 U18690 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15575), .A(
        n16216), .ZN(n16230) );
  NAND2_X1 U18691 ( .A1(n9685), .A2(n16217), .ZN(n15576) );
  XNOR2_X1 U18692 ( .A(n15577), .B(n15576), .ZN(n16229) );
  NOR2_X1 U18693 ( .A1(n10787), .A2(n18941), .ZN(n15578) );
  AOI221_X1 U18694 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15580), .C1(
        n15579), .C2(n15580), .A(n15578), .ZN(n15585) );
  OAI21_X1 U18695 ( .B1(n15582), .B2(n15581), .A(n13614), .ZN(n19097) );
  OAI22_X1 U18696 ( .A1(n19097), .A2(n16318), .B1(n16319), .B2(n19002), .ZN(
        n15583) );
  INV_X1 U18697 ( .A(n15583), .ZN(n15584) );
  OAI211_X1 U18698 ( .C1(n16229), .C2(n16299), .A(n15585), .B(n15584), .ZN(
        n15586) );
  INV_X1 U18699 ( .A(n15586), .ZN(n15587) );
  OAI21_X1 U18700 ( .B1(n16230), .B2(n16330), .A(n15587), .ZN(P2_U3037) );
  NOR2_X1 U18701 ( .A1(n16302), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15596) );
  OR2_X1 U18702 ( .A1(n15589), .A2(n15588), .ZN(n15590) );
  NAND2_X1 U18703 ( .A1(n15590), .A2(n13410), .ZN(n19102) );
  INV_X1 U18704 ( .A(n16316), .ZN(n15608) );
  NOR2_X1 U18705 ( .A1(n10771), .A2(n10856), .ZN(n15591) );
  AOI21_X1 U18706 ( .B1(n15608), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15591), .ZN(n15594) );
  INV_X1 U18707 ( .A(n19013), .ZN(n15592) );
  NAND2_X1 U18708 ( .A1(n15592), .A2(n16294), .ZN(n15593) );
  OAI211_X1 U18709 ( .C1(n19102), .C2(n16318), .A(n15594), .B(n15593), .ZN(
        n15595) );
  AOI211_X1 U18710 ( .C1(n15597), .C2(n16326), .A(n15596), .B(n15595), .ZN(
        n15598) );
  OAI21_X1 U18711 ( .B1(n15599), .B2(n16330), .A(n15598), .ZN(P2_U3039) );
  INV_X1 U18712 ( .A(n15600), .ZN(n15616) );
  INV_X1 U18713 ( .A(n15601), .ZN(n15614) );
  INV_X1 U18714 ( .A(n15602), .ZN(n15604) );
  NOR3_X1 U18715 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15604), .A3(
        n15603), .ZN(n15613) );
  XNOR2_X1 U18716 ( .A(n15605), .B(n15606), .ZN(n19104) );
  NOR2_X1 U18717 ( .A1(n10767), .A2(n10856), .ZN(n15607) );
  AOI21_X1 U18718 ( .B1(n15608), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15607), .ZN(n15611) );
  NAND2_X1 U18719 ( .A1(n15609), .A2(n16294), .ZN(n15610) );
  OAI211_X1 U18720 ( .C1(n19104), .C2(n16318), .A(n15611), .B(n15610), .ZN(
        n15612) );
  AOI211_X1 U18721 ( .C1(n15614), .C2(n16326), .A(n15613), .B(n15612), .ZN(
        n15615) );
  OAI21_X1 U18722 ( .B1(n15616), .B2(n16330), .A(n15615), .ZN(P2_U3040) );
  XNOR2_X1 U18723 ( .A(n15618), .B(n15617), .ZN(n16251) );
  NAND2_X1 U18724 ( .A1(n15622), .A2(n15621), .ZN(n15623) );
  OAI21_X1 U18725 ( .B1(n10881), .B2(n15624), .A(n15623), .ZN(n15625) );
  OAI21_X1 U18726 ( .B1(n15626), .B2(n10881), .A(n15625), .ZN(n16252) );
  INV_X1 U18727 ( .A(n16252), .ZN(n15638) );
  OAI21_X1 U18728 ( .B1(n9687), .B2(n15628), .A(n15627), .ZN(n19113) );
  NOR2_X1 U18729 ( .A1(n10761), .A2(n10856), .ZN(n15633) );
  AOI221_X1 U18730 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n15631), .C2(n15630), .A(
        n15629), .ZN(n15632) );
  AOI211_X1 U18731 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15634), .A(
        n15633), .B(n15632), .ZN(n15636) );
  NAND2_X1 U18732 ( .A1(n19040), .A2(n16294), .ZN(n15635) );
  OAI211_X1 U18733 ( .C1(n19113), .C2(n16318), .A(n15636), .B(n15635), .ZN(
        n15637) );
  AOI21_X1 U18734 ( .B1(n15638), .B2(n16295), .A(n15637), .ZN(n15639) );
  OAI21_X1 U18735 ( .B1(n16299), .B2(n16251), .A(n15639), .ZN(P2_U3041) );
  OAI22_X1 U18736 ( .A1(n16319), .A2(n15641), .B1(n15640), .B2(n16318), .ZN(
        n15644) );
  OAI22_X1 U18737 ( .A1(n16320), .A2(n15642), .B1(n10037), .B2(n18941), .ZN(
        n15643) );
  NOR2_X1 U18738 ( .A1(n15644), .A2(n15643), .ZN(n15650) );
  AOI22_X1 U18739 ( .A1(n16295), .A2(n15646), .B1(n16326), .B2(n15645), .ZN(
        n15649) );
  OAI211_X1 U18740 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n16322), .B(n15647), .ZN(n15648) );
  NAND3_X1 U18741 ( .A1(n15650), .A2(n15649), .A3(n15648), .ZN(P2_U3045) );
  OR2_X1 U18742 ( .A1(n19058), .A2(n15651), .ZN(n15656) );
  INV_X1 U18743 ( .A(n10743), .ZN(n15652) );
  NAND2_X1 U18744 ( .A1(n15653), .A2(n15652), .ZN(n15661) );
  INV_X1 U18745 ( .A(n15661), .ZN(n15654) );
  INV_X1 U18746 ( .A(n15676), .ZN(n15670) );
  MUX2_X1 U18747 ( .A(n15654), .B(n15670), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15655) );
  NAND2_X1 U18748 ( .A1(n15656), .A2(n15655), .ZN(n16347) );
  AOI21_X1 U18749 ( .B1(n16347), .B2(n19240), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n15657) );
  OAI22_X1 U18750 ( .A1(n15660), .A2(n15657), .B1(n13219), .B2(n15692), .ZN(
        n15658) );
  MUX2_X1 U18751 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15658), .S(
        n15685), .Z(P2_U3601) );
  INV_X1 U18752 ( .A(n15660), .ZN(n15667) );
  INV_X1 U18753 ( .A(n19799), .ZN(n15684) );
  OAI21_X1 U18754 ( .B1(n10145), .B2(n15662), .A(n15661), .ZN(n15663) );
  OAI21_X1 U18755 ( .B1(n15670), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15663), .ZN(n15664) );
  AOI21_X1 U18756 ( .B1(n15665), .B2(n15683), .A(n15664), .ZN(n16351) );
  OAI222_X1 U18757 ( .A1(n19817), .A2(n15692), .B1(n15667), .B2(n15666), .C1(
        n15684), .C2(n16351), .ZN(n15668) );
  MUX2_X1 U18758 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15668), .S(
        n15685), .Z(P2_U3600) );
  INV_X1 U18759 ( .A(n15669), .ZN(n15675) );
  OAI22_X1 U18760 ( .A1(n15671), .A2(n15674), .B1(n15670), .B2(n15675), .ZN(
        n15680) );
  NAND2_X1 U18761 ( .A1(n15673), .A2(n9638), .ZN(n15678) );
  AOI21_X1 U18762 ( .B1(n15676), .B2(n15675), .A(n15674), .ZN(n15677) );
  NAND2_X1 U18763 ( .A1(n15678), .A2(n15677), .ZN(n15679) );
  MUX2_X1 U18764 ( .A(n15680), .B(n15679), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15681) );
  AOI211_X1 U18765 ( .C1(n12379), .C2(n15683), .A(n15682), .B(n15681), .ZN(
        n16331) );
  OAI22_X1 U18766 ( .A1(n19801), .A2(n15692), .B1(n16331), .B2(n15684), .ZN(
        n15686) );
  MUX2_X1 U18767 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15686), .S(
        n15685), .Z(P2_U3596) );
  NOR3_X1 U18768 ( .A1(n19710), .A2(n19266), .A3(n19795), .ZN(n15687) );
  NOR2_X1 U18769 ( .A1(n19795), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19798) );
  NOR2_X1 U18770 ( .A1(n15687), .A2(n19798), .ZN(n15705) );
  INV_X1 U18771 ( .A(n15705), .ZN(n15695) );
  INV_X1 U18772 ( .A(n15688), .ZN(n15689) );
  AND2_X1 U18773 ( .A1(n15689), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19706) );
  NOR2_X1 U18774 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19272) );
  INV_X1 U18775 ( .A(n19272), .ZN(n19301) );
  NOR2_X1 U18776 ( .A1(n19441), .A2(n19301), .ZN(n19231) );
  NOR2_X1 U18777 ( .A1(n19706), .A2(n19231), .ZN(n15704) );
  AOI211_X1 U18778 ( .C1(n10282), .C2(n19240), .A(n19800), .B(n19231), .ZN(
        n15694) );
  NAND2_X1 U18779 ( .A1(n15690), .A2(n15903), .ZN(n15691) );
  INV_X1 U18780 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15709) );
  AOI22_X1 U18781 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19233), .ZN(n19656) );
  INV_X1 U18782 ( .A(n19656), .ZN(n19608) );
  AOI22_X1 U18783 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19233), .ZN(n19611) );
  INV_X1 U18784 ( .A(n19266), .ZN(n15701) );
  NAND2_X1 U18785 ( .A1(n15699), .A2(n19229), .ZN(n19255) );
  INV_X1 U18786 ( .A(n19231), .ZN(n15700) );
  OAI22_X1 U18787 ( .A1(n19611), .A2(n15701), .B1(n19255), .B2(n15700), .ZN(
        n15702) );
  AOI21_X1 U18788 ( .B1(n19710), .B2(n19608), .A(n15702), .ZN(n15708) );
  OAI21_X1 U18789 ( .B1(n10282), .B2(n19231), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15703) );
  NAND2_X1 U18790 ( .A1(n19235), .A2(n15706), .ZN(n15707) );
  OAI211_X1 U18791 ( .C1(n19239), .C2(n15709), .A(n15708), .B(n15707), .ZN(
        P2_U3051) );
  NAND2_X1 U18792 ( .A1(n19801), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19796) );
  NAND2_X1 U18793 ( .A1(n15721), .A2(n19807), .ZN(n19391) );
  OAI21_X1 U18794 ( .B1(n19796), .B2(n19794), .A(n19391), .ZN(n15713) );
  NAND2_X1 U18795 ( .A1(n9653), .A2(n19240), .ZN(n15711) );
  AND2_X1 U18796 ( .A1(n19795), .A2(n15714), .ZN(n15710) );
  AOI21_X1 U18797 ( .B1(n15711), .B2(n15710), .A(n19563), .ZN(n15712) );
  NAND2_X1 U18798 ( .A1(n15713), .A2(n15712), .ZN(n19438) );
  INV_X1 U18799 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U18800 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19233), .ZN(n19651) );
  INV_X1 U18801 ( .A(n19651), .ZN(n19574) );
  AOI22_X1 U18802 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19233), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19234), .ZN(n19577) );
  AOI22_X1 U18803 ( .A1(n19462), .A2(n19574), .B1(n19437), .B2(n19648), .ZN(
        n15719) );
  INV_X1 U18804 ( .A(n15714), .ZN(n19446) );
  OAI21_X1 U18805 ( .B1(n9653), .B2(n19446), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15715) );
  OAI21_X1 U18806 ( .B1(n19391), .B2(n19795), .A(n15715), .ZN(n19436) );
  NOR2_X2 U18807 ( .A1(n15717), .A2(n19220), .ZN(n19647) );
  AOI22_X1 U18808 ( .A1(n19436), .A2(n15716), .B1(n19446), .B2(n19647), .ZN(
        n15718) );
  OAI211_X1 U18809 ( .C1(n19435), .C2(n15720), .A(n15719), .B(n15718), .ZN(
        P2_U3106) );
  NAND2_X1 U18810 ( .A1(n15727), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19597) );
  NAND2_X1 U18811 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15721), .ZN(
        n19628) );
  OAI21_X1 U18812 ( .B1(n19597), .B2(n19794), .A(n19628), .ZN(n15724) );
  OAI21_X1 U18813 ( .B1(n15725), .B2(n19852), .A(n19240), .ZN(n15722) );
  INV_X1 U18814 ( .A(n19706), .ZN(n15734) );
  AOI21_X1 U18815 ( .B1(n15722), .B2(n15734), .A(n19563), .ZN(n15723) );
  NAND2_X1 U18816 ( .A1(n15724), .A2(n15723), .ZN(n19711) );
  INV_X1 U18817 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15732) );
  OAI21_X1 U18818 ( .B1(n15725), .B2(n19706), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15726) );
  OAI21_X1 U18819 ( .B1(n19628), .B2(n19795), .A(n15726), .ZN(n19708) );
  INV_X1 U18820 ( .A(n19647), .ZN(n15729) );
  AOI22_X1 U18821 ( .A1(n19700), .A2(n19648), .B1(n19710), .B2(n19574), .ZN(
        n15728) );
  OAI21_X1 U18822 ( .B1(n15729), .B2(n15734), .A(n15728), .ZN(n15730) );
  AOI21_X1 U18823 ( .B1(n19708), .B2(n15716), .A(n15730), .ZN(n15731) );
  OAI21_X1 U18824 ( .B1(n19704), .B2(n15732), .A(n15731), .ZN(P2_U3170) );
  INV_X1 U18825 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15737) );
  AOI22_X1 U18826 ( .A1(n19710), .A2(n19653), .B1(n19700), .B2(n19608), .ZN(
        n15733) );
  OAI21_X1 U18827 ( .B1(n19255), .B2(n15734), .A(n15733), .ZN(n15735) );
  AOI21_X1 U18828 ( .B1(n19708), .B2(n15706), .A(n15735), .ZN(n15736) );
  OAI21_X1 U18829 ( .B1(n19704), .B2(n15737), .A(n15736), .ZN(P2_U3171) );
  INV_X1 U18830 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16952) );
  INV_X1 U18831 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16951) );
  INV_X1 U18832 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16953) );
  INV_X1 U18833 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17019) );
  INV_X1 U18834 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17064) );
  INV_X1 U18835 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20777) );
  NAND3_X1 U18836 ( .A1(n17232), .A2(n15739), .A3(n15738), .ZN(n15742) );
  INV_X1 U18837 ( .A(n18688), .ZN(n15740) );
  NAND2_X1 U18838 ( .A1(n15741), .A2(n15740), .ZN(n15828) );
  INV_X1 U18839 ( .A(n17263), .ZN(n17260) );
  INV_X1 U18840 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16731) );
  INV_X1 U18841 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20880) );
  NAND2_X1 U18842 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17252) );
  NOR2_X1 U18843 ( .A1(n20880), .A2(n17252), .ZN(n17249) );
  NAND2_X1 U18844 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17249), .ZN(n17244) );
  NAND3_X1 U18845 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17109) );
  NAND3_X1 U18846 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n17107) );
  NAND4_X1 U18847 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n15743) );
  NOR4_X1 U18848 ( .A1(n17244), .A2(n17109), .A3(n17107), .A4(n15743), .ZN(
        n15744) );
  NAND4_X1 U18849 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(n15744), .ZN(n17089) );
  NOR2_X1 U18850 ( .A1(n16731), .A2(n17089), .ZN(n17090) );
  NAND3_X1 U18851 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17260), .A3(n17090), 
        .ZN(n20776) );
  NAND2_X1 U18852 ( .A1(n17232), .A2(n20775), .ZN(n17063) );
  NOR2_X1 U18853 ( .A1(n17064), .A2(n17063), .ZN(n17047) );
  NAND2_X1 U18854 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17047), .ZN(n17018) );
  NOR3_X1 U18855 ( .A1(n16953), .A2(n17019), .A3(n17018), .ZN(n17017) );
  NAND2_X1 U18856 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17017), .ZN(n17007) );
  NOR3_X1 U18857 ( .A1(n16952), .A2(n16951), .A3(n17007), .ZN(n17003) );
  NAND2_X1 U18858 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17003), .ZN(n16996) );
  INV_X1 U18859 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U18860 ( .A1(n18274), .A2(n17263), .ZN(n17257) );
  NAND2_X1 U18861 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16950) );
  NOR2_X2 U18862 ( .A1(n17232), .A2(n17263), .ZN(n20780) );
  NOR2_X1 U18863 ( .A1(n20780), .A2(n17003), .ZN(n17000) );
  AOI21_X1 U18864 ( .B1(n17257), .B2(n16950), .A(n17000), .ZN(n16989) );
  AOI22_X1 U18865 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U18866 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U18867 ( .A1(n12686), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15746) );
  AOI22_X1 U18868 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15745) );
  NAND4_X1 U18869 ( .A1(n15748), .A2(n15747), .A3(n15746), .A4(n15745), .ZN(
        n15754) );
  AOI22_X1 U18870 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15752) );
  AOI22_X1 U18871 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U18872 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18873 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15749) );
  NAND4_X1 U18874 ( .A1(n15752), .A2(n15751), .A3(n15750), .A4(n15749), .ZN(
        n15753) );
  NOR2_X1 U18875 ( .A1(n15754), .A2(n15753), .ZN(n15818) );
  AOI22_X1 U18876 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15758) );
  AOI22_X1 U18877 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15757) );
  AOI22_X1 U18878 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15756) );
  AOI22_X1 U18879 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15755) );
  NAND4_X1 U18880 ( .A1(n15758), .A2(n15757), .A3(n15756), .A4(n15755), .ZN(
        n15764) );
  AOI22_X1 U18881 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U18882 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15761) );
  AOI22_X1 U18883 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U18884 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15759) );
  NAND4_X1 U18885 ( .A1(n15762), .A2(n15761), .A3(n15760), .A4(n15759), .ZN(
        n15763) );
  NOR2_X1 U18886 ( .A1(n15764), .A2(n15763), .ZN(n16999) );
  AOI22_X1 U18887 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17342), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17170), .ZN(n15768) );
  AOI22_X1 U18888 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17340), .ZN(n15767) );
  AOI22_X1 U18889 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17214), .ZN(n15766) );
  AOI22_X1 U18890 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17201), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15765) );
  NAND4_X1 U18891 ( .A1(n15768), .A2(n15767), .A3(n15766), .A4(n15765), .ZN(
        n15774) );
  AOI22_X1 U18892 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17331), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U18893 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17329), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17330), .ZN(n15771) );
  AOI22_X1 U18894 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17328), .ZN(n15770) );
  AOI22_X1 U18895 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17219), .ZN(n15769) );
  NAND4_X1 U18896 ( .A1(n15772), .A2(n15771), .A3(n15770), .A4(n15769), .ZN(
        n15773) );
  NOR2_X1 U18897 ( .A1(n15774), .A2(n15773), .ZN(n17009) );
  AOI22_X1 U18898 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U18899 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15783) );
  INV_X1 U18900 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U18901 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15775) );
  OAI21_X1 U18902 ( .B1(n17188), .B2(n17216), .A(n15775), .ZN(n15781) );
  AOI22_X1 U18903 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15779) );
  AOI22_X1 U18904 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18905 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15777) );
  AOI22_X1 U18906 ( .A1(n15786), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15776) );
  NAND4_X1 U18907 ( .A1(n15779), .A2(n15778), .A3(n15777), .A4(n15776), .ZN(
        n15780) );
  AOI211_X1 U18908 ( .C1(n16971), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15781), .B(n15780), .ZN(n15782) );
  NAND3_X1 U18909 ( .A1(n15784), .A2(n15783), .A3(n15782), .ZN(n17014) );
  AOI22_X1 U18910 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15795) );
  AOI22_X1 U18911 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15794) );
  AOI22_X1 U18912 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15785) );
  OAI21_X1 U18913 ( .B1(n12718), .B2(n20794), .A(n15785), .ZN(n15792) );
  AOI22_X1 U18914 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U18915 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15789) );
  AOI22_X1 U18916 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U18917 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17201), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15787) );
  NAND4_X1 U18918 ( .A1(n15790), .A2(n15789), .A3(n15788), .A4(n15787), .ZN(
        n15791) );
  AOI211_X1 U18919 ( .C1(n17329), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n15792), .B(n15791), .ZN(n15793) );
  NAND3_X1 U18920 ( .A1(n15795), .A2(n15794), .A3(n15793), .ZN(n17015) );
  NAND2_X1 U18921 ( .A1(n17014), .A2(n17015), .ZN(n17013) );
  NOR2_X1 U18922 ( .A1(n17009), .A2(n17013), .ZN(n17008) );
  AOI22_X1 U18923 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17332), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15806) );
  AOI22_X1 U18924 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15805) );
  AOI22_X1 U18925 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15796) );
  OAI21_X1 U18926 ( .B1(n15797), .B2(n20851), .A(n15796), .ZN(n15803) );
  AOI22_X1 U18927 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15801) );
  AOI22_X1 U18928 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U18929 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15799) );
  AOI22_X1 U18930 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12684), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15798) );
  NAND4_X1 U18931 ( .A1(n15801), .A2(n15800), .A3(n15799), .A4(n15798), .ZN(
        n15802) );
  AOI211_X1 U18932 ( .C1(n17329), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15803), .B(n15802), .ZN(n15804) );
  NAND3_X1 U18933 ( .A1(n15806), .A2(n15805), .A3(n15804), .ZN(n17005) );
  NAND2_X1 U18934 ( .A1(n17008), .A2(n17005), .ZN(n17004) );
  NOR2_X1 U18935 ( .A1(n16999), .A2(n17004), .ZN(n16998) );
  AOI22_X1 U18936 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15817) );
  AOI22_X1 U18937 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U18938 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15807) );
  OAI21_X1 U18939 ( .B1(n15808), .B2(n20867), .A(n15807), .ZN(n15814) );
  AOI22_X1 U18940 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18941 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15811) );
  AOI22_X1 U18942 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U18943 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15809) );
  NAND4_X1 U18944 ( .A1(n15812), .A2(n15811), .A3(n15810), .A4(n15809), .ZN(
        n15813) );
  AOI211_X1 U18945 ( .C1(n17058), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15814), .B(n15813), .ZN(n15815) );
  NAND3_X1 U18946 ( .A1(n15817), .A2(n15816), .A3(n15815), .ZN(n16995) );
  NAND2_X1 U18947 ( .A1(n16998), .A2(n16995), .ZN(n16994) );
  NOR2_X1 U18948 ( .A1(n15818), .A2(n16994), .ZN(n16988) );
  AOI21_X1 U18949 ( .B1(n15818), .B2(n16994), .A(n16988), .ZN(n17281) );
  NAND2_X1 U18950 ( .A1(n17281), .A2(n20780), .ZN(n15819) );
  OAI221_X1 U18951 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16996), .C1(n20898), 
        .C2(n16989), .A(n15819), .ZN(P3_U2675) );
  NAND2_X1 U18952 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18416) );
  AOI221_X1 U18953 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18416), .C1(n15821), 
        .C2(n18416), .A(n15820), .ZN(n18235) );
  NOR2_X1 U18954 ( .A1(n15822), .A2(n20892), .ZN(n15823) );
  OAI21_X1 U18955 ( .B1(n15823), .B2(n18243), .A(n18236), .ZN(n18233) );
  AOI22_X1 U18956 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18235), .B1(
        n18233), .B2(n18240), .ZN(P3_U2865) );
  NOR2_X1 U18957 ( .A1(n15824), .A2(n18750), .ZN(n15832) );
  INV_X1 U18958 ( .A(n15825), .ZN(n18666) );
  NAND2_X1 U18959 ( .A1(n15826), .A2(n18666), .ZN(n16559) );
  OAI21_X1 U18960 ( .B1(n18877), .B2(n17494), .A(n16559), .ZN(n15827) );
  NAND3_X1 U18961 ( .A1(n18682), .A2(n18878), .A3(n15827), .ZN(n15908) );
  NAND3_X1 U18962 ( .A1(n15829), .A2(n15908), .A3(n15828), .ZN(n15830) );
  AOI21_X1 U18963 ( .B1(n15832), .B2(n15831), .A(n15830), .ZN(n18692) );
  INV_X1 U18964 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18231) );
  OR2_X1 U18965 ( .A1(n18231), .A2(n18829), .ZN(n15833) );
  NAND2_X1 U18966 ( .A1(n16561), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18237) );
  OAI211_X1 U18967 ( .C1(n18725), .C2(n18692), .A(n15833), .B(n18237), .ZN(
        n18855) );
  INV_X1 U18968 ( .A(n18852), .ZN(n15837) );
  OAI21_X1 U18969 ( .B1(n18849), .B2(n15834), .A(n18716), .ZN(n15835) );
  INV_X1 U18970 ( .A(n15835), .ZN(n15836) );
  NOR2_X1 U18971 ( .A1(n15836), .A2(n16559), .ZN(n18691) );
  NAND3_X1 U18972 ( .A1(n18855), .A2(n15837), .A3(n18691), .ZN(n15838) );
  OAI21_X1 U18973 ( .B1(n18855), .B2(n18716), .A(n15838), .ZN(P3_U3284) );
  NAND2_X1 U18974 ( .A1(n15840), .A2(n15839), .ZN(n15841) );
  XNOR2_X1 U18975 ( .A(n15841), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16409) );
  AOI21_X1 U18976 ( .B1(n18073), .B2(n16415), .A(n15842), .ZN(n16421) );
  OAI22_X1 U18977 ( .A1(n16394), .A2(n18139), .B1(n16405), .B2(n18187), .ZN(
        n15843) );
  NOR2_X1 U18978 ( .A1(n18204), .A2(n15843), .ZN(n15894) );
  NAND2_X1 U18979 ( .A1(n18210), .A2(n16425), .ZN(n15844) );
  OAI211_X1 U18980 ( .C1(n16421), .C2(n18182), .A(n15894), .B(n15844), .ZN(
        n15845) );
  AOI22_X1 U18981 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15845), .B1(
        n18209), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15849) );
  OR2_X1 U18982 ( .A1(n17909), .A2(n18187), .ZN(n15846) );
  OAI211_X1 U18983 ( .C1(n18139), .C2(n17908), .A(n15847), .B(n15846), .ZN(
        n15897) );
  NAND3_X1 U18984 ( .A1(n16393), .A2(n16396), .A3(n15897), .ZN(n15848) );
  OAI211_X1 U18985 ( .C1(n16409), .C2(n18127), .A(n15849), .B(n15848), .ZN(
        P3_U2833) );
  INV_X1 U18986 ( .A(n15850), .ZN(n15852) );
  NOR3_X1 U18987 ( .A1(n15852), .A2(n15851), .A3(n20493), .ZN(n15857) );
  INV_X1 U18988 ( .A(n15853), .ZN(n15855) );
  NAND2_X1 U18989 ( .A1(n15855), .A2(n15854), .ZN(n15856) );
  AOI222_X1 U18990 ( .A1(n15857), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .B1(n15857), .B2(n15856), .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C2(n15856), .ZN(n15858) );
  AOI222_X1 U18991 ( .A1(n15859), .A2(n20320), .B1(n15859), .B2(n15858), .C1(
        n20320), .C2(n15858), .ZN(n15863) );
  INV_X1 U18992 ( .A(n15863), .ZN(n15861) );
  OAI21_X1 U18993 ( .B1(n15861), .B2(n20125), .A(n15860), .ZN(n15862) );
  OAI21_X1 U18994 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15863), .A(
        n15862), .ZN(n15873) );
  INV_X1 U18995 ( .A(n15864), .ZN(n15872) );
  INV_X1 U18996 ( .A(n15865), .ZN(n15869) );
  OAI21_X1 U18997 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15866), .ZN(n15867) );
  NAND4_X1 U18998 ( .A1(n15870), .A2(n15869), .A3(n15868), .A4(n15867), .ZN(
        n15871) );
  AOI211_X1 U18999 ( .C1(n15873), .C2(n20029), .A(n15872), .B(n15871), .ZN(
        n15888) );
  INV_X1 U19000 ( .A(n15888), .ZN(n15879) );
  OAI21_X1 U19001 ( .B1(n20741), .B2(n15875), .A(n15874), .ZN(n15876) );
  OAI21_X1 U19002 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(n16146) );
  AOI221_X1 U19003 ( .B1(n20635), .B2(n20634), .C1(n15879), .C2(n20634), .A(
        n16146), .ZN(n16151) );
  NOR2_X1 U19004 ( .A1(n16149), .A2(n15880), .ZN(n15881) );
  NOR2_X1 U19005 ( .A1(n16151), .A2(n15881), .ZN(n15885) );
  AOI21_X1 U19006 ( .B1(n15899), .B2(n20638), .A(n15882), .ZN(n15883) );
  NAND2_X1 U19007 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15883), .ZN(n15884) );
  OAI22_X1 U19008 ( .A1(n15885), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n16151), 
        .B2(n15884), .ZN(n15886) );
  OAI211_X1 U19009 ( .C1(n15888), .C2(n19870), .A(n15887), .B(n15886), .ZN(
        P1_U3161) );
  NOR2_X1 U19010 ( .A1(n15890), .A2(n15889), .ZN(n15891) );
  XNOR2_X1 U19011 ( .A(n15891), .B(n15893), .ZN(n16391) );
  NOR2_X1 U19012 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15892), .ZN(
        n16387) );
  AOI21_X1 U19013 ( .B1(n15895), .B2(n15894), .A(n15893), .ZN(n15896) );
  AOI21_X1 U19014 ( .B1(n16387), .B2(n15897), .A(n15896), .ZN(n15898) );
  NAND2_X1 U19015 ( .A1(n18209), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16382) );
  OAI211_X1 U19016 ( .C1(n16391), .C2(n18127), .A(n15898), .B(n16382), .ZN(
        P3_U2832) );
  INV_X1 U19017 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20653) );
  INV_X1 U19018 ( .A(HOLD), .ZN(n19734) );
  NOR2_X1 U19019 ( .A1(n20653), .A2(n19734), .ZN(n20642) );
  AOI22_X1 U19020 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15901) );
  NAND2_X1 U19021 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15899), .ZN(n20640) );
  OAI211_X1 U19022 ( .C1(n20642), .C2(n15901), .A(n15900), .B(n20640), .ZN(
        P1_U3195) );
  AND2_X1 U19023 ( .A1(n15902), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19024 ( .A(n15903), .ZN(n19854) );
  NOR3_X1 U19025 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19716), .A3(n19861), 
        .ZN(n16365) );
  NOR4_X1 U19026 ( .A1(n15904), .A2(n19854), .A3(n16379), .A4(n16365), .ZN(
        P2_U3178) );
  INV_X1 U19027 ( .A(n15905), .ZN(n19840) );
  INV_X1 U19028 ( .A(n19834), .ZN(n19831) );
  NOR2_X1 U19029 ( .A1(n16358), .A2(n19831), .ZN(P2_U3047) );
  NAND3_X1 U19030 ( .A1(n17433), .A2(n18877), .A3(n15906), .ZN(n15907) );
  NAND2_X1 U19031 ( .A1(n17232), .A2(n17266), .ZN(n17401) );
  INV_X1 U19032 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17491) );
  NAND2_X1 U19033 ( .A1(n18694), .A2(n20913), .ZN(n17425) );
  INV_X1 U19034 ( .A(n17425), .ZN(n17429) );
  AOI22_X1 U19035 ( .A1(n17429), .A2(BUF2_REG_0__SCAN_IN), .B1(n17397), .B2(
        n15910), .ZN(n15911) );
  OAI221_X1 U19036 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17401), .C1(n17491), 
        .C2(n17266), .A(n15911), .ZN(P3_U2735) );
  AOI22_X1 U19037 ( .A1(n19955), .A2(P1_EBX_REG_26__SCAN_IN), .B1(n15912), 
        .B2(n19909), .ZN(n15921) );
  AOI22_X1 U19038 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19953), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n15913), .ZN(n15920) );
  INV_X1 U19039 ( .A(n15914), .ZN(n15917) );
  INV_X1 U19040 ( .A(n15915), .ZN(n15916) );
  AOI22_X1 U19041 ( .A1(n15917), .A2(n19902), .B1(n15916), .B2(n19936), .ZN(
        n15919) );
  INV_X1 U19042 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20698) );
  NAND3_X1 U19043 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15925), .A3(n20698), 
        .ZN(n15918) );
  NAND4_X1 U19044 ( .A1(n15921), .A2(n15920), .A3(n15919), .A4(n15918), .ZN(
        P1_U2814) );
  AOI22_X1 U19045 ( .A1(n19955), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19953), .ZN(n15931) );
  INV_X1 U19046 ( .A(n15922), .ZN(n15924) );
  AOI22_X1 U19047 ( .A1(n15924), .A2(n19909), .B1(n15923), .B2(n19936), .ZN(
        n15930) );
  INV_X1 U19048 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20696) );
  AOI22_X1 U19049 ( .A1(n15926), .A2(n19902), .B1(n15925), .B2(n20696), .ZN(
        n15929) );
  OAI21_X1 U19050 ( .B1(n15927), .B2(n15937), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15928) );
  NAND4_X1 U19051 ( .A1(n15931), .A2(n15930), .A3(n15929), .A4(n15928), .ZN(
        P1_U2815) );
  INV_X1 U19052 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15933) );
  OAI22_X1 U19053 ( .A1(n15933), .A2(n19919), .B1(n19965), .B2(n15932), .ZN(
        n15934) );
  AOI21_X1 U19054 ( .B1(n19955), .B2(P1_EBX_REG_23__SCAN_IN), .A(n15934), .ZN(
        n15941) );
  INV_X1 U19055 ( .A(n15935), .ZN(n16024) );
  INV_X1 U19056 ( .A(n15936), .ZN(n16022) );
  AOI22_X1 U19057 ( .A1(n16024), .A2(n19902), .B1(n16022), .B2(n19936), .ZN(
        n15940) );
  OAI21_X1 U19058 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n15938), .A(n15937), 
        .ZN(n15939) );
  NAND3_X1 U19059 ( .A1(n15941), .A2(n15940), .A3(n15939), .ZN(P1_U2817) );
  AOI22_X1 U19060 ( .A1(n19955), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19953), .ZN(n15952) );
  INV_X1 U19061 ( .A(n15942), .ZN(n15943) );
  AOI22_X1 U19062 ( .A1(n15943), .A2(n19909), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15957), .ZN(n15951) );
  INV_X1 U19063 ( .A(n15944), .ZN(n15947) );
  INV_X1 U19064 ( .A(n15945), .ZN(n15946) );
  AOI22_X1 U19065 ( .A1(n15947), .A2(n19902), .B1(n15946), .B2(n19936), .ZN(
        n15950) );
  INV_X1 U19066 ( .A(n15948), .ZN(n15949) );
  NAND4_X1 U19067 ( .A1(n15952), .A2(n15951), .A3(n15950), .A4(n15949), .ZN(
        P1_U2819) );
  AOI22_X1 U19068 ( .A1(n19955), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19909), 
        .B2(n15953), .ZN(n15958) );
  OAI21_X1 U19069 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15960), .ZN(n15966) );
  AND2_X1 U19070 ( .A1(n19932), .A2(n15961), .ZN(n15978) );
  AOI22_X1 U19071 ( .A1(n15978), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n19955), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n15962) );
  OAI21_X1 U19072 ( .B1(n16035), .B2(n19965), .A(n15962), .ZN(n15963) );
  AOI211_X1 U19073 ( .C1(n19953), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19952), .B(n15963), .ZN(n15965) );
  AOI22_X1 U19074 ( .A1(n16032), .A2(n19902), .B1(n16074), .B2(n19936), .ZN(
        n15964) );
  OAI211_X1 U19075 ( .C1(n15975), .C2(n15966), .A(n15965), .B(n15964), .ZN(
        P1_U2821) );
  AOI22_X1 U19076 ( .A1(n15978), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n19955), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15967) );
  OAI211_X1 U19077 ( .C1(n19919), .C2(n15968), .A(n15967), .B(n19933), .ZN(
        n15972) );
  OAI22_X1 U19078 ( .A1(n15970), .A2(n19924), .B1(n19948), .B2(n15969), .ZN(
        n15971) );
  AOI211_X1 U19079 ( .C1(n15973), .C2(n19909), .A(n15972), .B(n15971), .ZN(
        n15974) );
  OAI21_X1 U19080 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15975), .A(n15974), 
        .ZN(P1_U2822) );
  AOI22_X1 U19081 ( .A1(n19955), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19953), .ZN(n15983) );
  AOI21_X1 U19082 ( .B1(n19909), .B2(n16036), .A(n19952), .ZN(n15982) );
  INV_X1 U19083 ( .A(n15976), .ZN(n15977) );
  AOI22_X1 U19084 ( .A1(n16037), .A2(n19902), .B1(n15977), .B2(n19936), .ZN(
        n15981) );
  OAI221_X1 U19085 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15979), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(P1_REIP_REG_16__SCAN_IN), .A(n15978), 
        .ZN(n15980) );
  NAND4_X1 U19086 ( .A1(n15983), .A2(n15982), .A3(n15981), .A4(n15980), .ZN(
        P1_U2823) );
  AOI22_X1 U19087 ( .A1(n16042), .A2(n19902), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15984), .ZN(n15994) );
  OAI22_X1 U19088 ( .A1(n15987), .A2(n19948), .B1(n15986), .B2(n15985), .ZN(
        n15988) );
  INV_X1 U19089 ( .A(n15988), .ZN(n15989) );
  OAI211_X1 U19090 ( .C1(n19919), .C2(n15990), .A(n15989), .B(n19933), .ZN(
        n15991) );
  AOI211_X1 U19091 ( .C1(n19909), .C2(n16041), .A(n15992), .B(n15991), .ZN(
        n15993) );
  NAND2_X1 U19092 ( .A1(n15994), .A2(n15993), .ZN(P1_U2825) );
  NAND2_X1 U19093 ( .A1(n19932), .A2(n15995), .ZN(n16005) );
  AOI22_X1 U19094 ( .A1(n16084), .A2(n19936), .B1(n19955), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U19095 ( .C1(n19919), .C2(n14740), .A(n15996), .B(n19933), .ZN(
        n16000) );
  OAI22_X1 U19096 ( .A1(n15998), .A2(n19924), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15997), .ZN(n15999) );
  AOI211_X1 U19097 ( .C1(n16001), .C2(n19909), .A(n16000), .B(n15999), .ZN(
        n16002) );
  OAI21_X1 U19098 ( .B1(n20675), .B2(n16005), .A(n16002), .ZN(P1_U2827) );
  AOI22_X1 U19099 ( .A1(n19955), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19953), .ZN(n16011) );
  AOI21_X1 U19100 ( .B1(n16003), .B2(n19936), .A(n19952), .ZN(n16010) );
  INV_X1 U19101 ( .A(n16004), .ZN(n16046) );
  AOI22_X1 U19102 ( .A1(n16047), .A2(n19909), .B1(n19902), .B2(n16046), .ZN(
        n16009) );
  INV_X1 U19103 ( .A(n16005), .ZN(n16006) );
  OAI21_X1 U19104 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n16007), .A(n16006), 
        .ZN(n16008) );
  NAND4_X1 U19105 ( .A1(n16011), .A2(n16010), .A3(n16009), .A4(n16008), .ZN(
        P1_U2828) );
  INV_X1 U19106 ( .A(n16012), .ZN(n16090) );
  AOI22_X1 U19107 ( .A1(n19936), .A2(n16090), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n16013), .ZN(n16014) );
  NAND2_X1 U19108 ( .A1(n19933), .A2(n16014), .ZN(n16016) );
  OAI22_X1 U19109 ( .A1(n11657), .A2(n19919), .B1(n19965), .B2(n16060), .ZN(
        n16015) );
  AOI211_X1 U19110 ( .C1(n19955), .C2(P1_EBX_REG_11__SCAN_IN), .A(n16016), .B(
        n16015), .ZN(n16017) );
  INV_X1 U19111 ( .A(n16017), .ZN(n16018) );
  AOI21_X1 U19112 ( .B1(n16057), .B2(n19902), .A(n16018), .ZN(n16019) );
  OAI21_X1 U19113 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16020), .A(n16019), 
        .ZN(P1_U2829) );
  AOI22_X1 U19114 ( .A1(n16024), .A2(n16023), .B1(n16022), .B2(n16021), .ZN(
        n16025) );
  OAI21_X1 U19115 ( .B1(n14535), .B2(n20759), .A(n16025), .ZN(P1_U2849) );
  AOI22_X1 U19116 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16034) );
  INV_X1 U19117 ( .A(n16026), .ZN(n16029) );
  NAND3_X1 U19118 ( .A1(n16031), .A2(n16030), .A3(n16027), .ZN(n16028) );
  OAI211_X1 U19119 ( .C1(n16031), .C2(n16030), .A(n16029), .B(n16028), .ZN(
        n16075) );
  AOI22_X1 U19120 ( .A1(n16075), .A2(n19981), .B1(n19980), .B2(n16032), .ZN(
        n16033) );
  OAI211_X1 U19121 ( .C1(n19985), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        P1_U2980) );
  AOI22_X1 U19122 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19952), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U19123 ( .A1(n16037), .A2(n19980), .B1(n16036), .B2(n16048), .ZN(
        n16038) );
  OAI211_X1 U19124 ( .C1(n19877), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P1_U2982) );
  AOI22_X1 U19125 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16044) );
  AOI22_X1 U19126 ( .A1(n16042), .A2(n19980), .B1(n16041), .B2(n16048), .ZN(
        n16043) );
  OAI211_X1 U19127 ( .C1(n16045), .C2(n19877), .A(n16044), .B(n16043), .ZN(
        P1_U2984) );
  AOI22_X1 U19128 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U19129 ( .A1(n16048), .A2(n16047), .B1(n19980), .B2(n16046), .ZN(
        n16049) );
  OAI211_X1 U19130 ( .C1(n16051), .C2(n19877), .A(n16050), .B(n16049), .ZN(
        P1_U2987) );
  AOI22_X1 U19131 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19952), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16059) );
  NOR3_X1 U19132 ( .A1(n16053), .A2(n16052), .A3(n14747), .ZN(n16055) );
  NOR2_X1 U19133 ( .A1(n16055), .A2(n16054), .ZN(n16056) );
  XNOR2_X1 U19134 ( .A(n16056), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16092) );
  AOI22_X1 U19135 ( .A1(n19981), .A2(n16092), .B1(n19980), .B2(n16057), .ZN(
        n16058) );
  OAI211_X1 U19136 ( .C1(n19985), .C2(n16060), .A(n16059), .B(n16058), .ZN(
        P1_U2988) );
  AOI22_X1 U19137 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16067) );
  INV_X1 U19138 ( .A(n16061), .ZN(n16063) );
  NAND2_X1 U19139 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  XNOR2_X1 U19140 ( .A(n16065), .B(n16064), .ZN(n16129) );
  AOI22_X1 U19141 ( .A1(n16129), .A2(n19981), .B1(n19980), .B2(n19903), .ZN(
        n16066) );
  OAI211_X1 U19142 ( .C1(n19985), .C2(n19907), .A(n16067), .B(n16066), .ZN(
        P1_U2992) );
  AOI22_X1 U19143 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16072) );
  OAI21_X1 U19144 ( .B1(n13918), .B2(n16069), .A(n16068), .ZN(n16070) );
  INV_X1 U19145 ( .A(n16070), .ZN(n16135) );
  AOI22_X1 U19146 ( .A1(n16135), .A2(n19981), .B1(n19980), .B2(n19942), .ZN(
        n16071) );
  OAI211_X1 U19147 ( .C1(n19985), .C2(n19947), .A(n16072), .B(n16071), .ZN(
        P1_U2994) );
  AOI22_X1 U19148 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16073), .B1(
        n19973), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16077) );
  AOI22_X1 U19149 ( .A1(n16075), .A2(n20013), .B1(n20021), .B2(n16074), .ZN(
        n16076) );
  OAI211_X1 U19150 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16078), .A(
        n16077), .B(n16076), .ZN(P1_U3012) );
  NOR2_X1 U19151 ( .A1(n19933), .A2(n20675), .ZN(n16080) );
  AOI211_X1 U19152 ( .C1(n16082), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16087) );
  INV_X1 U19153 ( .A(n16083), .ZN(n16085) );
  AOI22_X1 U19154 ( .A1(n16085), .A2(n20013), .B1(n20021), .B2(n16084), .ZN(
        n16086) );
  OAI211_X1 U19155 ( .C1(n16089), .C2(n16088), .A(n16087), .B(n16086), .ZN(
        P1_U3018) );
  INV_X1 U19156 ( .A(n20003), .ZN(n16096) );
  AOI22_X1 U19157 ( .A1(n16090), .A2(n20021), .B1(n19973), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16094) );
  AOI22_X1 U19158 ( .A1(n16092), .A2(n20013), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16091), .ZN(n16093) );
  OAI211_X1 U19159 ( .C1(n16096), .C2(n16095), .A(n16094), .B(n16093), .ZN(
        P1_U3020) );
  AOI221_X1 U19160 ( .B1(n16102), .B2(n16118), .C1(n16098), .C2(n16118), .A(
        n16097), .ZN(n16116) );
  OAI22_X1 U19161 ( .A1(n16099), .A2(n19993), .B1(n20671), .B2(n19933), .ZN(
        n16100) );
  AOI21_X1 U19162 ( .B1(n16101), .B2(n20013), .A(n16100), .ZN(n16104) );
  NOR2_X1 U19163 ( .A1(n16102), .A2(n16123), .ZN(n16111) );
  OAI221_X1 U19164 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14747), .C2(n16115), .A(
        n16111), .ZN(n16103) );
  OAI211_X1 U19165 ( .C1(n16116), .C2(n14747), .A(n16104), .B(n16103), .ZN(
        P1_U3021) );
  NAND2_X1 U19166 ( .A1(n16106), .A2(n16105), .ZN(n16107) );
  NAND2_X1 U19167 ( .A1(n16108), .A2(n16107), .ZN(n19966) );
  INV_X1 U19168 ( .A(n19966), .ZN(n19895) );
  INV_X1 U19169 ( .A(n16109), .ZN(n16110) );
  AOI21_X1 U19170 ( .B1(n19895), .B2(n20021), .A(n16110), .ZN(n16114) );
  AOI22_X1 U19171 ( .A1(n16112), .A2(n20013), .B1(n16111), .B2(n16115), .ZN(
        n16113) );
  OAI211_X1 U19172 ( .C1(n16116), .C2(n16115), .A(n16114), .B(n16113), .ZN(
        P1_U3022) );
  AOI21_X1 U19173 ( .B1(n13932), .B2(n16118), .A(n16117), .ZN(n16133) );
  INV_X1 U19174 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16126) );
  INV_X1 U19175 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20665) );
  OAI222_X1 U19176 ( .A1(n16121), .A2(n19993), .B1(n19933), .B2(n20665), .C1(
        n16120), .C2(n16119), .ZN(n16122) );
  INV_X1 U19177 ( .A(n16122), .ZN(n16125) );
  INV_X1 U19178 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16132) );
  NOR2_X1 U19179 ( .A1(n13932), .A2(n16123), .ZN(n16128) );
  OAI221_X1 U19180 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16126), .C2(n16132), .A(
        n16128), .ZN(n16124) );
  OAI211_X1 U19181 ( .C1(n16133), .C2(n16126), .A(n16125), .B(n16124), .ZN(
        P1_U3023) );
  INV_X1 U19182 ( .A(n16127), .ZN(n19906) );
  AOI22_X1 U19183 ( .A1(n19906), .A2(n20021), .B1(n19973), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U19184 ( .A1(n16129), .A2(n20013), .B1(n16128), .B2(n16132), .ZN(
        n16130) );
  OAI211_X1 U19185 ( .C1(n16133), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        P1_U3024) );
  AOI22_X1 U19186 ( .A1(n19937), .A2(n20021), .B1(n19973), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16137) );
  AOI22_X1 U19187 ( .A1(n16135), .A2(n20013), .B1(n20003), .B2(n16134), .ZN(
        n16136) );
  OAI211_X1 U19188 ( .C1(n16139), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        P1_U3026) );
  NAND2_X1 U19189 ( .A1(n20724), .A2(n16140), .ZN(n16142) );
  OAI22_X1 U19190 ( .A1(n16143), .A2(n16142), .B1(n16141), .B2(n20727), .ZN(
        P1_U3468) );
  NAND4_X1 U19191 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20638), .A4(n20741), .ZN(n16144) );
  NAND2_X1 U19192 ( .A1(n16145), .A2(n16144), .ZN(n20636) );
  OAI21_X1 U19193 ( .B1(n16147), .B2(n20636), .A(n16146), .ZN(n16148) );
  OAI221_X1 U19194 ( .B1(n16149), .B2(n20451), .C1(n16149), .C2(n20741), .A(
        n16148), .ZN(n16150) );
  AOI221_X1 U19195 ( .B1(n16151), .B2(n20634), .C1(n20635), .C2(n20634), .A(
        n16150), .ZN(P1_U3162) );
  NOR2_X1 U19196 ( .A1(n16151), .A2(n20635), .ZN(n16153) );
  OAI22_X1 U19197 ( .A1(n20451), .A2(n16153), .B1(n16152), .B2(n20635), .ZN(
        P1_U3466) );
  AOI21_X1 U19198 ( .B1(n16155), .B2(n16154), .A(n14259), .ZN(n16162) );
  INV_X1 U19199 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U19200 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19049), .ZN(n16156) );
  OAI21_X1 U19201 ( .B1(n19030), .B2(n19779), .A(n16156), .ZN(n16157) );
  AOI21_X1 U19202 ( .B1(n16158), .B2(n19041), .A(n16157), .ZN(n16159) );
  OAI21_X1 U19203 ( .B1(n16160), .B2(n19052), .A(n16159), .ZN(n16161) );
  AOI21_X1 U19204 ( .B1(n19042), .B2(n16162), .A(n16161), .ZN(n16163) );
  OAI21_X1 U19205 ( .B1(n16164), .B2(n19046), .A(n16163), .ZN(P2_U2826) );
  AOI21_X1 U19206 ( .B1(n16167), .B2(n16166), .A(n16165), .ZN(n16179) );
  NAND2_X1 U19207 ( .A1(n19036), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16168) );
  OAI21_X1 U19208 ( .B1(n19030), .B2(n19775), .A(n16168), .ZN(n16175) );
  INV_X1 U19209 ( .A(n16169), .ZN(n16173) );
  INV_X1 U19210 ( .A(n16170), .ZN(n16171) );
  AOI211_X1 U19211 ( .C1(n16173), .C2(n16172), .A(n19052), .B(n16171), .ZN(
        n16174) );
  AOI211_X1 U19212 ( .C1(P2_EBX_REG_27__SCAN_IN), .C2(n19049), .A(n16175), .B(
        n16174), .ZN(n16176) );
  OAI21_X1 U19213 ( .B1(n16177), .B2(n19057), .A(n16176), .ZN(n16178) );
  AOI21_X1 U19214 ( .B1(n19042), .B2(n16179), .A(n16178), .ZN(n16180) );
  OAI21_X1 U19215 ( .B1(n16181), .B2(n19046), .A(n16180), .ZN(P2_U2828) );
  AOI22_X1 U19216 ( .A1(n19071), .A2(n16182), .B1(n19129), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16188) );
  AOI22_X1 U19217 ( .A1(n19073), .A2(BUF1_REG_22__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16187) );
  INV_X1 U19218 ( .A(n16183), .ZN(n16184) );
  AOI22_X1 U19219 ( .A1(n16185), .A2(n19108), .B1(n19130), .B2(n16184), .ZN(
        n16186) );
  NAND3_X1 U19220 ( .A1(n16188), .A2(n16187), .A3(n16186), .ZN(P2_U2897) );
  AOI22_X1 U19221 ( .A1(n19071), .A2(n16189), .B1(n19129), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16196) );
  AOI22_X1 U19222 ( .A1(n19073), .A2(BUF1_REG_20__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16195) );
  NOR2_X1 U19223 ( .A1(n16191), .A2(n16190), .ZN(n16192) );
  AOI21_X1 U19224 ( .B1(n16193), .B2(n19108), .A(n16192), .ZN(n16194) );
  NAND3_X1 U19225 ( .A1(n16196), .A2(n16195), .A3(n16194), .ZN(P2_U2899) );
  AOI22_X1 U19226 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19176), .ZN(n16204) );
  INV_X1 U19227 ( .A(n14193), .ZN(n16197) );
  AOI21_X1 U19228 ( .B1(n9709), .B2(n16198), .A(n16197), .ZN(n16279) );
  NAND2_X1 U19229 ( .A1(n16200), .A2(n16199), .ZN(n16202) );
  XOR2_X1 U19230 ( .A(n16202), .B(n16201), .Z(n16278) );
  AOI222_X1 U19231 ( .A1(n16279), .A2(n9578), .B1(n19180), .B2(n16278), .C1(
        n19198), .C2(n16277), .ZN(n16203) );
  OAI211_X1 U19232 ( .C1(n19191), .C2(n16205), .A(n16204), .B(n16203), .ZN(
        P2_U3000) );
  AOI22_X1 U19233 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19176), .ZN(n16209) );
  AOI222_X1 U19234 ( .A1(n16207), .A2(n19180), .B1(n19198), .B2(n18982), .C1(
        n9578), .C2(n16206), .ZN(n16208) );
  OAI211_X1 U19235 ( .C1(n19191), .C2(n18980), .A(n16209), .B(n16208), .ZN(
        P2_U3002) );
  AOI22_X1 U19236 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19176), .B1(n16258), 
        .B2(n18987), .ZN(n16214) );
  OAI22_X1 U19237 ( .A1(n16211), .A2(n19192), .B1(n16210), .B2(n19194), .ZN(
        n16212) );
  AOI21_X1 U19238 ( .B1(n19198), .B2(n18991), .A(n16212), .ZN(n16213) );
  OAI211_X1 U19239 ( .C1(n19202), .C2(n10778), .A(n16214), .B(n16213), .ZN(
        P2_U3003) );
  AOI22_X1 U19240 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19176), .ZN(n16227) );
  AOI21_X1 U19241 ( .B1(n16289), .B2(n16216), .A(n16215), .ZN(n16296) );
  NAND2_X1 U19242 ( .A1(n16218), .A2(n16217), .ZN(n16223) );
  INV_X1 U19243 ( .A(n16219), .ZN(n16220) );
  NOR2_X1 U19244 ( .A1(n16221), .A2(n16220), .ZN(n16222) );
  XNOR2_X1 U19245 ( .A(n16223), .B(n16222), .ZN(n16300) );
  OAI22_X1 U19246 ( .A1(n16300), .A2(n19194), .B1(n19185), .B2(n16224), .ZN(
        n16225) );
  AOI21_X1 U19247 ( .B1(n16296), .B2(n9578), .A(n16225), .ZN(n16226) );
  OAI211_X1 U19248 ( .C1(n19191), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        P2_U3004) );
  AOI22_X1 U19249 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19176), .B1(n16258), 
        .B2(n18998), .ZN(n16234) );
  INV_X1 U19250 ( .A(n19002), .ZN(n16232) );
  OAI22_X1 U19251 ( .A1(n16230), .A2(n19192), .B1(n19194), .B2(n16229), .ZN(
        n16231) );
  AOI21_X1 U19252 ( .B1(n19198), .B2(n16232), .A(n16231), .ZN(n16233) );
  OAI211_X1 U19253 ( .C1(n19202), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        P2_U3005) );
  AOI22_X1 U19254 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19176), .ZN(n16249) );
  AOI21_X1 U19255 ( .B1(n15348), .B2(n16237), .A(n16236), .ZN(n16242) );
  INV_X1 U19256 ( .A(n16238), .ZN(n16239) );
  NOR2_X1 U19257 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  XNOR2_X1 U19258 ( .A(n16242), .B(n16241), .ZN(n16312) );
  INV_X1 U19259 ( .A(n16309), .ZN(n16247) );
  AND2_X1 U19260 ( .A1(n16244), .A2(n16243), .ZN(n16245) );
  XOR2_X1 U19261 ( .A(n16246), .B(n16245), .Z(n16308) );
  AOI222_X1 U19262 ( .A1(n16312), .A2(n19180), .B1(n19198), .B2(n16247), .C1(
        n9578), .C2(n16308), .ZN(n16248) );
  OAI211_X1 U19263 ( .C1(n19191), .C2(n16250), .A(n16249), .B(n16248), .ZN(
        P2_U3006) );
  AOI22_X1 U19264 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19176), .B1(n16258), 
        .B2(n19039), .ZN(n16255) );
  OAI22_X1 U19265 ( .A1(n19192), .A2(n16252), .B1(n16251), .B2(n19194), .ZN(
        n16253) );
  AOI21_X1 U19266 ( .B1(n19198), .B2(n19040), .A(n16253), .ZN(n16254) );
  OAI211_X1 U19267 ( .C1(n19202), .C2(n16256), .A(n16255), .B(n16254), .ZN(
        P2_U3009) );
  AOI22_X1 U19268 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19176), .B1(n16258), 
        .B2(n16257), .ZN(n16265) );
  NAND3_X1 U19269 ( .A1(n16259), .A2(n9578), .A3(n13811), .ZN(n16260) );
  OAI21_X1 U19270 ( .B1(n19185), .B2(n16261), .A(n16260), .ZN(n16262) );
  AOI21_X1 U19271 ( .B1(n16263), .B2(n19180), .A(n16262), .ZN(n16264) );
  OAI211_X1 U19272 ( .C1(n10080), .C2(n19202), .A(n16265), .B(n16264), .ZN(
        P2_U3011) );
  NOR2_X1 U19273 ( .A1(n15326), .A2(n18941), .ZN(n16270) );
  INV_X1 U19274 ( .A(n15509), .ZN(n16266) );
  OAI21_X1 U19275 ( .B1(n16267), .B2(n9643), .A(n16266), .ZN(n19080) );
  OAI22_X1 U19276 ( .A1(n16318), .A2(n19080), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16268), .ZN(n16269) );
  AOI211_X1 U19277 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16271), .A(
        n16270), .B(n16269), .ZN(n16274) );
  AOI22_X1 U19278 ( .A1(n16272), .A2(n16295), .B1(n16294), .B2(n18972), .ZN(
        n16273) );
  OAI211_X1 U19279 ( .C1(n16275), .C2(n16299), .A(n16274), .B(n16273), .ZN(
        P2_U3031) );
  AOI22_X1 U19280 ( .A1(n16276), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16307), .B2(n19081), .ZN(n16286) );
  AOI222_X1 U19281 ( .A1(n16279), .A2(n16295), .B1(n16326), .B2(n16278), .C1(
        n16294), .C2(n16277), .ZN(n16285) );
  NAND2_X1 U19282 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19176), .ZN(n16284) );
  OAI211_X1 U19283 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16282), .A(
        n16281), .B(n16280), .ZN(n16283) );
  NAND4_X1 U19284 ( .A1(n16286), .A2(n16285), .A3(n16284), .A4(n16283), .ZN(
        P2_U3032) );
  NAND2_X1 U19285 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19176), .ZN(n16287) );
  OAI221_X1 U19286 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16290), 
        .C1(n16289), .C2(n16288), .A(n16287), .ZN(n16291) );
  AOI21_X1 U19287 ( .B1(n16292), .B2(n16307), .A(n16291), .ZN(n16298) );
  AOI22_X1 U19288 ( .A1(n16296), .A2(n16295), .B1(n16294), .B2(n16293), .ZN(
        n16297) );
  OAI211_X1 U19289 ( .C1(n16300), .C2(n16299), .A(n16298), .B(n16297), .ZN(
        P2_U3036) );
  INV_X1 U19290 ( .A(n16301), .ZN(n16303) );
  AOI211_X1 U19291 ( .C1(n16315), .C2(n16304), .A(n16303), .B(n16302), .ZN(
        n16306) );
  NOR2_X1 U19292 ( .A1(n10856), .A2(n13413), .ZN(n16305) );
  AOI211_X1 U19293 ( .C1(n16307), .C2(n19098), .A(n16306), .B(n16305), .ZN(
        n16314) );
  INV_X1 U19294 ( .A(n16308), .ZN(n16310) );
  OAI22_X1 U19295 ( .A1(n16310), .A2(n16330), .B1(n16319), .B2(n16309), .ZN(
        n16311) );
  AOI21_X1 U19296 ( .B1(n16326), .B2(n16312), .A(n16311), .ZN(n16313) );
  OAI211_X1 U19297 ( .C1(n16316), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        P2_U3038) );
  OAI22_X1 U19298 ( .A1(n16319), .A2(n19058), .B1(n16318), .B2(n16317), .ZN(
        n16324) );
  INV_X1 U19299 ( .A(n16320), .ZN(n16321) );
  MUX2_X1 U19300 ( .A(n16322), .B(n16321), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n16323) );
  AOI211_X1 U19301 ( .C1(n16326), .C2(n16325), .A(n16324), .B(n16323), .ZN(
        n16328) );
  OAI211_X1 U19302 ( .C1(n16330), .C2(n16329), .A(n16328), .B(n16327), .ZN(
        P2_U3046) );
  MUX2_X1 U19303 ( .A(n16331), .B(n9999), .S(n16357), .Z(n16364) );
  INV_X1 U19304 ( .A(n16357), .ZN(n16332) );
  MUX2_X1 U19305 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16333), .S(
        n16332), .Z(n16359) );
  INV_X1 U19306 ( .A(n16359), .ZN(n16363) );
  OAI21_X1 U19307 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16335), .ZN(n16338) );
  INV_X1 U19308 ( .A(n16336), .ZN(n16337) );
  OAI211_X1 U19309 ( .C1(n9627), .C2(n16339), .A(n16338), .B(n16337), .ZN(
        n16346) );
  AOI22_X1 U19310 ( .A1(n16345), .A2(n16342), .B1(n9707), .B2(n16341), .ZN(
        n16343) );
  OAI21_X1 U19311 ( .B1(n16345), .B2(n16344), .A(n16343), .ZN(n19841) );
  AOI211_X1 U19312 ( .C1(n16357), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16346), .B(n19841), .ZN(n16362) );
  INV_X1 U19313 ( .A(n16364), .ZN(n16355) );
  INV_X1 U19314 ( .A(n16347), .ZN(n16348) );
  NAND2_X1 U19315 ( .A1(n16348), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16349) );
  NAND2_X1 U19316 ( .A1(n16349), .A2(n19824), .ZN(n16352) );
  INV_X1 U19317 ( .A(n16349), .ZN(n16350) );
  AOI22_X1 U19318 ( .A1(n16352), .A2(n16351), .B1(n16350), .B2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16354) );
  NAND2_X1 U19319 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16363), .ZN(
        n16353) );
  OAI211_X1 U19320 ( .C1(n16355), .C2(n19807), .A(n16354), .B(n16353), .ZN(
        n16356) );
  OAI22_X1 U19321 ( .A1(n16357), .A2(n16356), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16364), .ZN(n16360) );
  OAI221_X1 U19322 ( .B1(n16360), .B2(n16359), .C1(n16360), .C2(n19272), .A(
        n16358), .ZN(n16361) );
  OAI211_X1 U19323 ( .C1(n16364), .C2(n16363), .A(n16362), .B(n16361), .ZN(
        n16374) );
  AOI211_X1 U19324 ( .C1(n19721), .C2(n16374), .A(n16366), .B(n16365), .ZN(
        n16377) );
  NAND3_X1 U19325 ( .A1(n16368), .A2(n10566), .A3(n16367), .ZN(n16370) );
  NOR2_X1 U19326 ( .A1(n16369), .A2(n19852), .ZN(n19857) );
  AND2_X1 U19327 ( .A1(n16370), .A2(n19857), .ZN(n16372) );
  AOI22_X1 U19328 ( .A1(n19853), .A2(n16372), .B1(n19854), .B2(n16371), .ZN(
        n16375) );
  INV_X1 U19329 ( .A(n16372), .ZN(n16373) );
  AOI221_X1 U19330 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16374), .C1(
        P2_STATE2_REG_0__SCAN_IN), .C2(P2_STATE2_REG_1__SCAN_IN), .A(n16373), 
        .ZN(n19718) );
  INV_X1 U19331 ( .A(n19718), .ZN(n19719) );
  NAND2_X1 U19332 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19719), .ZN(n16380) );
  OAI21_X1 U19333 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16375), .A(n16380), 
        .ZN(n16376) );
  OAI211_X1 U19334 ( .C1(n19840), .C2(n16378), .A(n16377), .B(n16376), .ZN(
        P2_U3176) );
  AOI21_X1 U19335 ( .B1(n16380), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16379), 
        .ZN(n16381) );
  INV_X1 U19336 ( .A(n16381), .ZN(P2_U3593) );
  XOR2_X1 U19337 ( .A(n16397), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16594) );
  INV_X1 U19338 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16384) );
  OAI221_X1 U19339 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16385), .C1(
        n16384), .C2(n16383), .A(n16382), .ZN(n16386) );
  AOI21_X1 U19340 ( .B1(n17754), .B2(n16594), .A(n16386), .ZN(n16390) );
  OAI22_X1 U19341 ( .A1(n9602), .A2(n17905), .B1(n16394), .B2(n17745), .ZN(
        n16388) );
  NOR2_X1 U19342 ( .A1(n16413), .A2(n17704), .ZN(n17600) );
  INV_X1 U19343 ( .A(n17600), .ZN(n17616) );
  NOR2_X1 U19344 ( .A1(n16414), .A2(n17616), .ZN(n17567) );
  AOI22_X1 U19345 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16388), .B1(
        n16387), .B2(n17567), .ZN(n16389) );
  OAI211_X1 U19346 ( .C1(n16391), .C2(n17778), .A(n16390), .B(n16389), .ZN(
        P3_U2800) );
  OAI21_X1 U19347 ( .B1(n18278), .B2(n16392), .A(n16610), .ZN(n16402) );
  INV_X1 U19348 ( .A(n16393), .ZN(n16404) );
  NOR2_X1 U19349 ( .A1(n16404), .A2(n17908), .ZN(n16420) );
  INV_X1 U19350 ( .A(n16420), .ZN(n16395) );
  AOI211_X1 U19351 ( .C1(n16396), .C2(n16395), .A(n16394), .B(n17745), .ZN(
        n16401) );
  INV_X1 U19352 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18811) );
  AOI21_X1 U19353 ( .B1(n16572), .B2(n16610), .A(n16397), .ZN(n16604) );
  OAI21_X1 U19354 ( .B1(n17754), .B2(n16398), .A(n16604), .ZN(n16399) );
  OAI21_X1 U19355 ( .B1(n18811), .B2(n18175), .A(n16399), .ZN(n16400) );
  AOI211_X1 U19356 ( .C1(n16403), .C2(n16402), .A(n16401), .B(n16400), .ZN(
        n16408) );
  NOR2_X1 U19357 ( .A1(n17909), .A2(n16404), .ZN(n16422) );
  NOR2_X1 U19358 ( .A1(n9602), .A2(n17905), .ZN(n16406) );
  OAI21_X1 U19359 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16422), .A(
        n16406), .ZN(n16407) );
  OAI211_X1 U19360 ( .C1(n16409), .C2(n17778), .A(n16408), .B(n16407), .ZN(
        P3_U2801) );
  INV_X1 U19361 ( .A(n18201), .ZN(n18687) );
  AOI22_X1 U19362 ( .A1(n18687), .A2(n16411), .B1(n16410), .B2(n18097), .ZN(
        n18012) );
  INV_X1 U19363 ( .A(n18194), .ZN(n18009) );
  AOI22_X1 U19364 ( .A1(n18689), .A2(n17926), .B1(n18017), .B2(n18009), .ZN(
        n17929) );
  OAI21_X1 U19365 ( .B1(n18012), .B2(n16412), .A(n17929), .ZN(n17954) );
  NAND2_X1 U19366 ( .A1(n18218), .A2(n17954), .ZN(n17980) );
  NOR2_X1 U19367 ( .A1(n16413), .A2(n17980), .ZN(n17948) );
  NOR3_X1 U19368 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16415), .A3(
        n16414), .ZN(n17554) );
  AOI22_X1 U19369 ( .A1(n18209), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17948), 
        .B2(n17554), .ZN(n16430) );
  AOI21_X1 U19370 ( .B1(n17811), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16416), .ZN(n17557) );
  OAI21_X1 U19371 ( .B1(n17563), .B2(n12810), .A(n16426), .ZN(n17556) );
  NAND2_X1 U19372 ( .A1(n17557), .A2(n17556), .ZN(n17555) );
  NAND2_X1 U19373 ( .A1(n17811), .A2(n17563), .ZN(n16417) );
  NAND2_X1 U19374 ( .A1(n17555), .A2(n16417), .ZN(n16418) );
  AOI221_X1 U19375 ( .B1(n17402), .B2(n16420), .C1(n16419), .C2(n16418), .A(
        n18684), .ZN(n16424) );
  OAI211_X1 U19376 ( .C1(n16422), .C2(n18201), .A(n16421), .B(n18221), .ZN(
        n16423) );
  OAI211_X1 U19377 ( .C1(n16424), .C2(n16423), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18175), .ZN(n16429) );
  NAND4_X1 U19378 ( .A1(n17811), .A2(n17563), .A3(n18227), .A4(n16425), .ZN(
        n16428) );
  OR3_X1 U19379 ( .A1(n18127), .A2(n16426), .A3(n17557), .ZN(n16427) );
  NAND4_X1 U19380 ( .A1(n16430), .A2(n16429), .A3(n16428), .A4(n16427), .ZN(
        P3_U2834) );
  NOR3_X1 U19381 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16432) );
  NOR4_X1 U19382 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16431) );
  NAND4_X1 U19383 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16432), .A3(n16431), .A4(
        U215), .ZN(U213) );
  INV_X1 U19384 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16529) );
  NOR2_X1 U19385 ( .A1(n16486), .A2(n16433), .ZN(n16484) );
  INV_X1 U19386 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16530) );
  OAI222_X1 U19387 ( .A1(U212), .A2(n16529), .B1(n16491), .B2(n16434), .C1(
        U214), .C2(n16530), .ZN(U216) );
  INV_X1 U19388 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U19389 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16489), .ZN(n16435) );
  OAI21_X1 U19390 ( .B1(n16436), .B2(n16491), .A(n16435), .ZN(U217) );
  INV_X1 U19391 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16489), .ZN(n16437) );
  OAI21_X1 U19393 ( .B1(n16438), .B2(n16491), .A(n16437), .ZN(U218) );
  INV_X1 U19394 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U19395 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16489), .ZN(n16439) );
  OAI21_X1 U19396 ( .B1(n16440), .B2(n16491), .A(n16439), .ZN(U219) );
  INV_X1 U19397 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16489), .ZN(n16441) );
  OAI21_X1 U19399 ( .B1(n16442), .B2(n16491), .A(n16441), .ZN(U220) );
  INV_X1 U19400 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19401 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16489), .ZN(n16443) );
  OAI21_X1 U19402 ( .B1(n16444), .B2(n16491), .A(n16443), .ZN(U221) );
  INV_X1 U19403 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16446) );
  AOI22_X1 U19404 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16489), .ZN(n16445) );
  OAI21_X1 U19405 ( .B1(n16446), .B2(n16491), .A(n16445), .ZN(U222) );
  INV_X1 U19406 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U19407 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16489), .ZN(n16447) );
  OAI21_X1 U19408 ( .B1(n16448), .B2(n16491), .A(n16447), .ZN(U223) );
  AOI22_X1 U19409 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16489), .ZN(n16449) );
  OAI21_X1 U19410 ( .B1(n16450), .B2(n16491), .A(n16449), .ZN(U224) );
  INV_X1 U19411 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U19412 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16489), .ZN(n16451) );
  OAI21_X1 U19413 ( .B1(n16452), .B2(n16491), .A(n16451), .ZN(U225) );
  INV_X1 U19414 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U19415 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16489), .ZN(n16453) );
  OAI21_X1 U19416 ( .B1(n16454), .B2(n16491), .A(n16453), .ZN(U226) );
  INV_X1 U19417 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19418 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16489), .ZN(n16455) );
  OAI21_X1 U19419 ( .B1(n16456), .B2(n16491), .A(n16455), .ZN(U227) );
  INV_X1 U19420 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16458) );
  AOI22_X1 U19421 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16489), .ZN(n16457) );
  OAI21_X1 U19422 ( .B1(n16458), .B2(n16491), .A(n16457), .ZN(U228) );
  INV_X1 U19423 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16460) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16489), .ZN(n16459) );
  OAI21_X1 U19425 ( .B1(n16460), .B2(n16491), .A(n16459), .ZN(U229) );
  INV_X1 U19426 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19427 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16489), .ZN(n16461) );
  OAI21_X1 U19428 ( .B1(n16462), .B2(n16491), .A(n16461), .ZN(U230) );
  INV_X1 U19429 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16464) );
  AOI22_X1 U19430 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16489), .ZN(n16463) );
  OAI21_X1 U19431 ( .B1(n16464), .B2(n16491), .A(n16463), .ZN(U231) );
  AOI22_X1 U19432 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16484), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16489), .ZN(n16465) );
  OAI21_X1 U19433 ( .B1(n13658), .B2(U214), .A(n16465), .ZN(U232) );
  INV_X1 U19434 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16509) );
  AOI22_X1 U19435 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16486), .ZN(n16466) );
  OAI21_X1 U19436 ( .B1(n16509), .B2(U212), .A(n16466), .ZN(U233) );
  AOI22_X1 U19437 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16489), .ZN(n16467) );
  OAI21_X1 U19438 ( .B1(n16468), .B2(n16491), .A(n16467), .ZN(U234) );
  AOI22_X1 U19439 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16489), .ZN(n16469) );
  OAI21_X1 U19440 ( .B1(n16470), .B2(n16491), .A(n16469), .ZN(U235) );
  INV_X1 U19441 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16505) );
  AOI22_X1 U19442 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16486), .ZN(n16471) );
  OAI21_X1 U19443 ( .B1(n16505), .B2(U212), .A(n16471), .ZN(U236) );
  AOI22_X1 U19444 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16489), .ZN(n16472) );
  OAI21_X1 U19445 ( .B1(n16473), .B2(n16491), .A(n16472), .ZN(U237) );
  AOI22_X1 U19446 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16489), .ZN(n16474) );
  OAI21_X1 U19447 ( .B1(n16475), .B2(n16491), .A(n16474), .ZN(U238) );
  INV_X1 U19448 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16501) );
  OAI222_X1 U19449 ( .A1(U212), .A2(n16501), .B1(n16491), .B2(n16476), .C1(
        U214), .C2(n13765), .ZN(U239) );
  INV_X1 U19450 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19451 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16486), .ZN(n16477) );
  OAI21_X1 U19452 ( .B1(n16500), .B2(U212), .A(n16477), .ZN(U240) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16489), .ZN(n16478) );
  OAI21_X1 U19454 ( .B1(n16479), .B2(n16491), .A(n16478), .ZN(U241) );
  INV_X1 U19455 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16498) );
  AOI22_X1 U19456 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16486), .ZN(n16480) );
  OAI21_X1 U19457 ( .B1(n16498), .B2(U212), .A(n16480), .ZN(U242) );
  AOI22_X1 U19458 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16489), .ZN(n16481) );
  OAI21_X1 U19459 ( .B1(n16482), .B2(n16491), .A(n16481), .ZN(U243) );
  INV_X1 U19460 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16496) );
  AOI22_X1 U19461 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16486), .ZN(n16483) );
  OAI21_X1 U19462 ( .B1(n16496), .B2(U212), .A(n16483), .ZN(U244) );
  INV_X1 U19463 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16495) );
  AOI22_X1 U19464 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16484), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16486), .ZN(n16485) );
  OAI21_X1 U19465 ( .B1(n16495), .B2(U212), .A(n16485), .ZN(U245) );
  AOI22_X1 U19466 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16489), .ZN(n16487) );
  OAI21_X1 U19467 ( .B1(n16488), .B2(n16491), .A(n16487), .ZN(U246) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16486), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16489), .ZN(n16490) );
  OAI21_X1 U19469 ( .B1(n16492), .B2(n16491), .A(n16490), .ZN(U247) );
  INV_X1 U19470 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16493) );
  AOI22_X1 U19471 ( .A1(n16527), .A2(n16493), .B1(n18241), .B2(U215), .ZN(U251) );
  OAI22_X1 U19472 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16527), .ZN(n16494) );
  INV_X1 U19473 ( .A(n16494), .ZN(U252) );
  INV_X1 U19474 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18252) );
  AOI22_X1 U19475 ( .A1(n16527), .A2(n16495), .B1(n18252), .B2(U215), .ZN(U253) );
  INV_X1 U19476 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U19477 ( .A1(n16527), .A2(n16496), .B1(n18257), .B2(U215), .ZN(U254) );
  INV_X1 U19478 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U19479 ( .A1(n16521), .A2(n16497), .B1(n18261), .B2(U215), .ZN(U255) );
  INV_X1 U19480 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18266) );
  AOI22_X1 U19481 ( .A1(n16521), .A2(n16498), .B1(n18266), .B2(U215), .ZN(U256) );
  INV_X1 U19482 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16499) );
  INV_X1 U19483 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U19484 ( .A1(n16521), .A2(n16499), .B1(n18271), .B2(U215), .ZN(U257) );
  INV_X1 U19485 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U19486 ( .A1(n16527), .A2(n16500), .B1(n18276), .B2(U215), .ZN(U258) );
  INV_X1 U19487 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U19488 ( .A1(n16521), .A2(n16501), .B1(n17524), .B2(U215), .ZN(U259) );
  INV_X1 U19489 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16502) );
  INV_X1 U19490 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U19491 ( .A1(n16527), .A2(n16502), .B1(n17526), .B2(U215), .ZN(U260) );
  INV_X1 U19492 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16503) );
  INV_X1 U19493 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U19494 ( .A1(n16527), .A2(n16503), .B1(n17528), .B2(U215), .ZN(U261) );
  INV_X1 U19495 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19496 ( .A1(n16521), .A2(n16505), .B1(n16504), .B2(U215), .ZN(U262) );
  INV_X1 U19497 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16506) );
  INV_X1 U19498 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U19499 ( .A1(n16527), .A2(n16506), .B1(n17532), .B2(U215), .ZN(U263) );
  INV_X1 U19500 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16507) );
  INV_X1 U19501 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U19502 ( .A1(n16521), .A2(n16507), .B1(n17537), .B2(U215), .ZN(U264) );
  INV_X1 U19503 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16508) );
  AOI22_X1 U19504 ( .A1(n16521), .A2(n16509), .B1(n16508), .B2(U215), .ZN(U265) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16527), .ZN(n16510) );
  INV_X1 U19506 ( .A(n16510), .ZN(U266) );
  OAI22_X1 U19507 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16527), .ZN(n16511) );
  INV_X1 U19508 ( .A(n16511), .ZN(U267) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16527), .ZN(n16512) );
  INV_X1 U19510 ( .A(n16512), .ZN(U268) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16527), .ZN(n16513) );
  INV_X1 U19512 ( .A(n16513), .ZN(U269) );
  INV_X1 U19513 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16514) );
  INV_X1 U19514 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U19515 ( .A1(n16527), .A2(n16514), .B1(n18256), .B2(U215), .ZN(U270) );
  INV_X1 U19516 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16515) );
  INV_X1 U19517 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U19518 ( .A1(n16527), .A2(n16515), .B1(n20883), .B2(U215), .ZN(U271) );
  INV_X1 U19519 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16516) );
  INV_X1 U19520 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18265) );
  AOI22_X1 U19521 ( .A1(n16527), .A2(n16516), .B1(n18265), .B2(U215), .ZN(U272) );
  OAI22_X1 U19522 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16527), .ZN(n16517) );
  INV_X1 U19523 ( .A(n16517), .ZN(U273) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16527), .ZN(n16518) );
  INV_X1 U19525 ( .A(n16518), .ZN(U274) );
  OAI22_X1 U19526 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16521), .ZN(n16519) );
  INV_X1 U19527 ( .A(n16519), .ZN(U275) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16521), .ZN(n16520) );
  INV_X1 U19529 ( .A(n16520), .ZN(U276) );
  OAI22_X1 U19530 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16521), .ZN(n16522) );
  INV_X1 U19531 ( .A(n16522), .ZN(U277) );
  OAI22_X1 U19532 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16527), .ZN(n16523) );
  INV_X1 U19533 ( .A(n16523), .ZN(U278) );
  OAI22_X1 U19534 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16527), .ZN(n16524) );
  INV_X1 U19535 ( .A(n16524), .ZN(U279) );
  OAI22_X1 U19536 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16527), .ZN(n16525) );
  INV_X1 U19537 ( .A(n16525), .ZN(U280) );
  INV_X1 U19538 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16526) );
  INV_X1 U19539 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U19540 ( .A1(n16527), .A2(n16526), .B1(n18270), .B2(U215), .ZN(U281) );
  INV_X1 U19541 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U19542 ( .A1(n16527), .A2(n16529), .B1(n18277), .B2(U215), .ZN(U282) );
  INV_X1 U19543 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16528) );
  AOI222_X1 U19544 ( .A1(n16530), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16529), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16528), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16531) );
  INV_X1 U19545 ( .A(n16533), .ZN(n16532) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18775) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19548 ( .A1(n16532), .A2(n18775), .B1(n19752), .B2(n16533), .ZN(
        U347) );
  INV_X1 U19549 ( .A(n16533), .ZN(n16534) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18773) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19552 ( .A1(n16534), .A2(n18773), .B1(n19751), .B2(n16533), .ZN(
        U348) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18771) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19555 ( .A1(n16532), .A2(n18771), .B1(n19750), .B2(n16533), .ZN(
        U349) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18769) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19558 ( .A1(n16532), .A2(n18769), .B1(n19749), .B2(n16533), .ZN(
        U350) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18767) );
  INV_X1 U19560 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19561 ( .A1(n16532), .A2(n18767), .B1(n19748), .B2(n16533), .ZN(
        U351) );
  INV_X1 U19562 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18764) );
  INV_X1 U19563 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19564 ( .A1(n16532), .A2(n18764), .B1(n19747), .B2(n16533), .ZN(
        U352) );
  INV_X1 U19565 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18763) );
  INV_X1 U19566 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19567 ( .A1(n16534), .A2(n18763), .B1(n19746), .B2(n16533), .ZN(
        U353) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18761) );
  AOI22_X1 U19569 ( .A1(n16532), .A2(n18761), .B1(n19745), .B2(n16533), .ZN(
        U354) );
  INV_X1 U19570 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18814) );
  INV_X1 U19571 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19572 ( .A1(n16532), .A2(n18814), .B1(n19782), .B2(n16533), .ZN(
        U355) );
  INV_X1 U19573 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18812) );
  INV_X1 U19574 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19575 ( .A1(n16532), .A2(n18812), .B1(n19780), .B2(n16533), .ZN(
        U356) );
  INV_X1 U19576 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18808) );
  INV_X1 U19577 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19578 ( .A1(n16532), .A2(n18808), .B1(n19777), .B2(n16533), .ZN(
        U357) );
  INV_X1 U19579 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18807) );
  INV_X1 U19580 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20886) );
  AOI22_X1 U19581 ( .A1(n16532), .A2(n18807), .B1(n20886), .B2(n16533), .ZN(
        U358) );
  INV_X1 U19582 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18805) );
  INV_X1 U19583 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19584 ( .A1(n16532), .A2(n18805), .B1(n19774), .B2(n16533), .ZN(
        U359) );
  INV_X1 U19585 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20877) );
  INV_X1 U19586 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U19587 ( .A1(n16532), .A2(n20877), .B1(n19772), .B2(n16533), .ZN(
        U360) );
  INV_X1 U19588 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18801) );
  INV_X1 U19589 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19590 ( .A1(n16532), .A2(n18801), .B1(n19770), .B2(n16533), .ZN(
        U361) );
  INV_X1 U19591 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18798) );
  INV_X1 U19592 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19593 ( .A1(n16532), .A2(n18798), .B1(n19769), .B2(n16533), .ZN(
        U362) );
  INV_X1 U19594 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18797) );
  INV_X1 U19595 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19596 ( .A1(n16532), .A2(n18797), .B1(n19767), .B2(n16533), .ZN(
        U363) );
  INV_X1 U19597 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20846) );
  INV_X1 U19598 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19599 ( .A1(n16532), .A2(n20846), .B1(n19766), .B2(n16533), .ZN(
        U364) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18759) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19602 ( .A1(n16532), .A2(n18759), .B1(n19744), .B2(n16533), .ZN(
        U365) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18794) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19605 ( .A1(n16532), .A2(n18794), .B1(n19764), .B2(n16533), .ZN(
        U366) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18792) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19608 ( .A1(n16532), .A2(n18792), .B1(n19762), .B2(n16533), .ZN(
        U367) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18790) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U19611 ( .A1(n16532), .A2(n18790), .B1(n19760), .B2(n16533), .ZN(
        U368) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18788) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U19614 ( .A1(n16532), .A2(n18788), .B1(n19758), .B2(n16533), .ZN(
        U369) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18787) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19756) );
  AOI22_X1 U19617 ( .A1(n16532), .A2(n18787), .B1(n19756), .B2(n16533), .ZN(
        U370) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18785) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19620 ( .A1(n16534), .A2(n18785), .B1(n19755), .B2(n16533), .ZN(
        U371) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18782) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U19623 ( .A1(n16534), .A2(n18782), .B1(n20868), .B2(n16533), .ZN(
        U372) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18781) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19626 ( .A1(n16534), .A2(n18781), .B1(n19754), .B2(n16533), .ZN(
        U373) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18779) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19629 ( .A1(n16534), .A2(n18779), .B1(n19753), .B2(n16533), .ZN(
        U374) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18777) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U19632 ( .A1(n16534), .A2(n18777), .B1(n20785), .B2(n16533), .ZN(
        U375) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18757) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U19635 ( .A1(n16534), .A2(n18757), .B1(n19743), .B2(n16533), .ZN(
        U376) );
  INV_X1 U19636 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16536) );
  INV_X1 U19637 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18756) );
  NAND2_X1 U19638 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18756), .ZN(n18746) );
  INV_X1 U19639 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n16535) );
  NAND2_X1 U19640 ( .A1(n18741), .A2(n16535), .ZN(n18742) );
  OAI21_X1 U19641 ( .B1(n18746), .B2(n16535), .A(n18742), .ZN(n18827) );
  INV_X1 U19642 ( .A(n18827), .ZN(n18824) );
  OAI21_X1 U19643 ( .B1(n18741), .B2(n16536), .A(n18824), .ZN(P3_U2633) );
  INV_X1 U19644 ( .A(n18887), .ZN(n16539) );
  NAND2_X1 U19645 ( .A1(n18682), .A2(n16537), .ZN(n16542) );
  OAI21_X1 U19646 ( .B1(n18725), .B2(n16542), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16538) );
  OAI21_X1 U19647 ( .B1(n16539), .B2(n16561), .A(n16538), .ZN(P3_U2634) );
  AOI22_X1 U19648 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18885), .B1(n16541), .B2(
        n18741), .ZN(n16540) );
  OAI21_X1 U19649 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18885), .A(n16540), 
        .ZN(P3_U2635) );
  OAI21_X1 U19650 ( .B1(n16541), .B2(BS16), .A(n18827), .ZN(n18825) );
  OAI21_X1 U19651 ( .B1(n18827), .B2(n18876), .A(n18825), .ZN(P3_U2636) );
  NOR2_X1 U19652 ( .A1(n16543), .A2(n16542), .ZN(n18693) );
  NOR2_X1 U19653 ( .A1(n18693), .A2(n18725), .ZN(n18868) );
  OAI21_X1 U19654 ( .B1(n18868), .B2(n18231), .A(n16544), .ZN(P3_U2637) );
  NOR4_X1 U19655 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16548) );
  NOR4_X1 U19656 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16547) );
  NOR4_X1 U19657 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16546) );
  NOR4_X1 U19658 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16545) );
  NAND4_X1 U19659 ( .A1(n16548), .A2(n16547), .A3(n16546), .A4(n16545), .ZN(
        n16554) );
  NOR4_X1 U19660 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16552) );
  AOI211_X1 U19661 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16551) );
  NOR4_X1 U19662 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16550) );
  NOR4_X1 U19663 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16549) );
  NAND4_X1 U19664 ( .A1(n16552), .A2(n16551), .A3(n16550), .A4(n16549), .ZN(
        n16553) );
  NOR2_X1 U19665 ( .A1(n16554), .A2(n16553), .ZN(n18862) );
  INV_X1 U19666 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16556) );
  NOR3_X1 U19667 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n16557) );
  OAI21_X1 U19668 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16557), .A(n18862), .ZN(
        n16555) );
  OAI21_X1 U19669 ( .B1(n18862), .B2(n16556), .A(n16555), .ZN(P3_U2638) );
  INV_X1 U19670 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18858) );
  INV_X1 U19671 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18826) );
  AOI21_X1 U19672 ( .B1(n18858), .B2(n18826), .A(n16557), .ZN(n16558) );
  INV_X1 U19673 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18818) );
  INV_X1 U19674 ( .A(n18862), .ZN(n18865) );
  AOI22_X1 U19675 ( .A1(n18862), .A2(n16558), .B1(n18818), .B2(n18865), .ZN(
        P3_U2639) );
  NAND2_X1 U19676 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16562), .ZN(n18729) );
  NOR2_X1 U19677 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18729), .ZN(n18722) );
  NAND4_X1 U19678 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n16562), .A3(n16561), 
        .A4(n18876), .ZN(n18734) );
  NAND2_X1 U19679 ( .A1(n18175), .A2(n18734), .ZN(n16563) );
  NOR2_X2 U19680 ( .A1(n16933), .A2(n18830), .ZN(n16897) );
  OAI211_X1 U19681 ( .C1(n16564), .C2(n18248), .A(n18878), .B(n18876), .ZN(
        n18720) );
  INV_X1 U19682 ( .A(n18720), .ZN(n16565) );
  AOI211_X4 U19683 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18248), .A(n16565), .B(
        n16567), .ZN(n16921) );
  AOI22_X1 U19684 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16897), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16921), .ZN(n16590) );
  NAND2_X1 U19685 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18248), .ZN(n16566) );
  AOI211_X4 U19686 ( .C1(n18876), .C2(n18878), .A(n16567), .B(n16566), .ZN(
        n16890) );
  NOR2_X1 U19687 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16944), .ZN(n16586) );
  NOR2_X1 U19688 ( .A1(n16931), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n16917) );
  INV_X1 U19689 ( .A(n16917), .ZN(n16899) );
  NOR2_X1 U19690 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16899), .ZN(n16898) );
  INV_X1 U19691 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17105) );
  NAND2_X1 U19692 ( .A1(n16898), .A2(n17105), .ZN(n16889) );
  NOR2_X1 U19693 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16889), .ZN(n16871) );
  INV_X1 U19694 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U19695 ( .A1(n16871), .A2(n17233), .ZN(n16862) );
  INV_X1 U19696 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16844) );
  NAND2_X1 U19697 ( .A1(n16847), .A2(n16844), .ZN(n16843) );
  INV_X1 U19698 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17108) );
  NAND2_X1 U19699 ( .A1(n16821), .A2(n17108), .ZN(n16813) );
  INV_X1 U19700 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17127) );
  NAND2_X1 U19701 ( .A1(n16795), .A2(n17127), .ZN(n16792) );
  INV_X1 U19702 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17140) );
  NAND2_X1 U19703 ( .A1(n16772), .A2(n17140), .ZN(n16764) );
  INV_X1 U19704 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17111) );
  NAND2_X1 U19705 ( .A1(n16753), .A2(n17111), .ZN(n16746) );
  INV_X1 U19706 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17076) );
  NAND2_X1 U19707 ( .A1(n16726), .A2(n17076), .ZN(n16721) );
  NAND2_X1 U19708 ( .A1(n16704), .A2(n17064), .ZN(n16696) );
  NAND2_X1 U19709 ( .A1(n16682), .A2(n17019), .ZN(n16675) );
  NOR2_X1 U19710 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16675), .ZN(n16662) );
  INV_X1 U19711 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16954) );
  NAND2_X1 U19712 ( .A1(n16662), .A2(n16954), .ZN(n16655) );
  NOR2_X1 U19713 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16655), .ZN(n16641) );
  NAND2_X1 U19714 ( .A1(n16641), .A2(n16952), .ZN(n16635) );
  NOR2_X1 U19715 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16635), .ZN(n16621) );
  NAND2_X1 U19716 ( .A1(n16621), .A2(n20898), .ZN(n16615) );
  NOR2_X1 U19717 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16615), .ZN(n16600) );
  NAND2_X1 U19718 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16611) );
  NOR2_X1 U19719 ( .A1(n18811), .A2(n16611), .ZN(n16569) );
  NOR2_X1 U19720 ( .A1(n16926), .A2(n16933), .ZN(n16949) );
  INV_X1 U19721 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18800) );
  INV_X1 U19722 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18795) );
  INV_X1 U19723 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18796) );
  INV_X1 U19724 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20801) );
  INV_X1 U19725 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18783) );
  INV_X1 U19726 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18778) );
  INV_X1 U19727 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18774) );
  INV_X1 U19728 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18770) );
  INV_X1 U19729 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18762) );
  NAND3_X1 U19730 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16907) );
  NOR2_X1 U19731 ( .A1(n18762), .A2(n16907), .ZN(n16872) );
  NAND2_X1 U19732 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16872), .ZN(n16860) );
  NAND2_X1 U19733 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16838) );
  NOR3_X1 U19734 ( .A1(n18770), .A2(n16860), .A3(n16838), .ZN(n16827) );
  NAND2_X1 U19735 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16827), .ZN(n16812) );
  NOR2_X1 U19736 ( .A1(n18774), .A2(n16812), .ZN(n16796) );
  NAND2_X1 U19737 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16796), .ZN(n16773) );
  NOR2_X1 U19738 ( .A1(n18778), .A2(n16773), .ZN(n16776) );
  NAND2_X1 U19739 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16776), .ZN(n16738) );
  NOR2_X1 U19740 ( .A1(n18783), .A2(n16738), .ZN(n16737) );
  NAND3_X1 U19741 ( .A1(n16737), .A2(P3_REIP_REG_16__SCAN_IN), .A3(
        P3_REIP_REG_15__SCAN_IN), .ZN(n16730) );
  NOR2_X1 U19742 ( .A1(n20801), .A2(n16730), .ZN(n16728) );
  NAND4_X1 U19743 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16728), .ZN(n16676) );
  NOR3_X1 U19744 ( .A1(n18795), .A2(n18796), .A3(n16676), .ZN(n16661) );
  NAND2_X1 U19745 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16661), .ZN(n16650) );
  NOR2_X1 U19746 ( .A1(n18800), .A2(n16650), .ZN(n16631) );
  AND3_X1 U19747 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16631), .ZN(n16568) );
  OAI21_X1 U19748 ( .B1(n16937), .B2(n16568), .A(n16946), .ZN(n16634) );
  INV_X1 U19749 ( .A(n16634), .ZN(n16630) );
  OAI21_X1 U19750 ( .B1(n16569), .B2(n16949), .A(n16630), .ZN(n16607) );
  INV_X1 U19751 ( .A(n16607), .ZN(n16571) );
  NAND2_X1 U19752 ( .A1(n16926), .A2(n16568), .ZN(n16622) );
  INV_X1 U19753 ( .A(n16569), .ZN(n16570) );
  NOR2_X1 U19754 ( .A1(n16622), .A2(n16570), .ZN(n16587) );
  INV_X1 U19755 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18815) );
  NAND2_X1 U19756 ( .A1(n16587), .A2(n18815), .ZN(n16595) );
  AOI21_X1 U19757 ( .B1(n16571), .B2(n16595), .A(n18813), .ZN(n16585) );
  INV_X1 U19758 ( .A(n16604), .ZN(n16602) );
  OAI21_X1 U19759 ( .B1(n16573), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16572), .ZN(n17551) );
  AOI21_X1 U19760 ( .B1(n16574), .B2(n17546), .A(n16573), .ZN(n17562) );
  INV_X1 U19761 ( .A(n17562), .ZN(n16627) );
  OAI21_X1 U19762 ( .B1(n17548), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16574), .ZN(n17574) );
  INV_X1 U19763 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16651) );
  NOR2_X1 U19764 ( .A1(n16578), .A2(n16651), .ZN(n16576) );
  INV_X1 U19765 ( .A(n17548), .ZN(n16575) );
  OAI21_X1 U19766 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16576), .A(
        n16575), .ZN(n17586) );
  INV_X1 U19767 ( .A(n16578), .ZN(n16577) );
  AOI22_X1 U19768 ( .A1(n16577), .A2(n16651), .B1(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16578), .ZN(n17594) );
  NAND2_X1 U19769 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17620) );
  NAND2_X1 U19770 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17619), .ZN(
        n16582) );
  NOR2_X1 U19771 ( .A1(n17620), .A2(n16582), .ZN(n17581) );
  OAI21_X1 U19772 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17581), .A(
        n16578), .ZN(n17611) );
  INV_X1 U19773 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16687) );
  NOR2_X1 U19774 ( .A1(n16687), .A2(n16582), .ZN(n16580) );
  INV_X1 U19775 ( .A(n17581), .ZN(n16579) );
  OAI21_X1 U19776 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16580), .A(
        n16579), .ZN(n17622) );
  INV_X1 U19777 ( .A(n16582), .ZN(n16581) );
  AOI22_X1 U19778 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16582), .B1(
        n16581), .B2(n16687), .ZN(n17632) );
  NOR2_X1 U19779 ( .A1(n17894), .A2(n17643), .ZN(n17617) );
  OAI21_X1 U19780 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17617), .A(
        n16582), .ZN(n17644) );
  NAND2_X1 U19781 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17653) );
  INV_X1 U19782 ( .A(n17720), .ZN(n17737) );
  NAND2_X1 U19783 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17737), .ZN(
        n17739) );
  NOR2_X1 U19784 ( .A1(n17695), .A2(n17739), .ZN(n17693) );
  NAND3_X1 U19785 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17693), .ZN(n16739) );
  NOR2_X1 U19786 ( .A1(n17680), .A2(n16739), .ZN(n17652) );
  NAND2_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17693), .ZN(
        n16750) );
  NOR2_X1 U19788 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16750), .ZN(
        n16741) );
  NAND2_X1 U19789 ( .A1(n17652), .A2(n16741), .ZN(n16714) );
  OAI21_X1 U19790 ( .B1(n17653), .B2(n16714), .A(n16903), .ZN(n16695) );
  NAND2_X1 U19791 ( .A1(n17644), .A2(n16695), .ZN(n16694) );
  NAND2_X1 U19792 ( .A1(n16903), .A2(n16694), .ZN(n16684) );
  NAND2_X1 U19793 ( .A1(n17632), .A2(n16684), .ZN(n16683) );
  NAND2_X1 U19794 ( .A1(n16903), .A2(n16683), .ZN(n16674) );
  NAND2_X1 U19795 ( .A1(n17622), .A2(n16674), .ZN(n16673) );
  NAND2_X1 U19796 ( .A1(n16903), .A2(n16673), .ZN(n16666) );
  NAND2_X1 U19797 ( .A1(n17611), .A2(n16666), .ZN(n16665) );
  NAND2_X1 U19798 ( .A1(n16903), .A2(n16665), .ZN(n16657) );
  NAND2_X1 U19799 ( .A1(n17594), .A2(n16657), .ZN(n16656) );
  NAND2_X1 U19800 ( .A1(n16903), .A2(n16656), .ZN(n16646) );
  NAND2_X1 U19801 ( .A1(n17586), .A2(n16646), .ZN(n16645) );
  NAND2_X1 U19802 ( .A1(n16903), .A2(n16645), .ZN(n16637) );
  NAND2_X1 U19803 ( .A1(n17574), .A2(n16637), .ZN(n16636) );
  NAND2_X1 U19804 ( .A1(n16903), .A2(n16636), .ZN(n16626) );
  NAND2_X1 U19805 ( .A1(n16627), .A2(n16626), .ZN(n16625) );
  NAND2_X1 U19806 ( .A1(n16903), .A2(n16625), .ZN(n16617) );
  NAND2_X1 U19807 ( .A1(n17551), .A2(n16617), .ZN(n16616) );
  NAND2_X1 U19808 ( .A1(n16903), .A2(n16616), .ZN(n16601) );
  OAI21_X1 U19809 ( .B1(n16602), .B2(n16583), .A(n16601), .ZN(n16593) );
  INV_X1 U19810 ( .A(n18734), .ZN(n16904) );
  NAND2_X1 U19811 ( .A1(n16903), .A2(n16904), .ZN(n16935) );
  NOR3_X1 U19812 ( .A1(n16594), .A2(n16593), .A3(n16935), .ZN(n16584) );
  AOI211_X1 U19813 ( .C1(n16586), .C2(n16600), .A(n16585), .B(n16584), .ZN(
        n16589) );
  NAND3_X1 U19814 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16587), .A3(n18813), 
        .ZN(n16588) );
  NAND3_X1 U19815 ( .A1(n16590), .A2(n16589), .A3(n16588), .ZN(P3_U2640) );
  AOI22_X1 U19816 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16897), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16607), .ZN(n16598) );
  XNOR2_X1 U19817 ( .A(P3_EBX_REG_30__SCAN_IN), .B(n16600), .ZN(n16591) );
  AOI22_X1 U19818 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16921), .B1(n16890), 
        .B2(n16591), .ZN(n16597) );
  AOI21_X1 U19819 ( .B1(n16594), .B2(n16593), .A(n18734), .ZN(n16592) );
  OAI21_X1 U19820 ( .B1(n16594), .B2(n16593), .A(n16592), .ZN(n16596) );
  NAND4_X1 U19821 ( .A1(n16598), .A2(n16597), .A3(n16596), .A4(n16595), .ZN(
        P3_U2641) );
  NOR3_X1 U19822 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16622), .A3(n16611), 
        .ZN(n16599) );
  AOI21_X1 U19823 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16921), .A(n16599), .ZN(
        n16609) );
  AOI211_X1 U19824 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16615), .A(n16600), .B(
        n16944), .ZN(n16606) );
  INV_X1 U19825 ( .A(n16601), .ZN(n16603) );
  AOI221_X1 U19826 ( .B1(n16604), .B2(n16603), .C1(n16602), .C2(n16601), .A(
        n18734), .ZN(n16605) );
  AOI211_X1 U19827 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16607), .A(n16606), 
        .B(n16605), .ZN(n16608) );
  OAI211_X1 U19828 ( .C1(n16610), .C2(n16934), .A(n16609), .B(n16608), .ZN(
        P3_U2642) );
  INV_X1 U19829 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18809) );
  INV_X1 U19830 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18806) );
  INV_X1 U19831 ( .A(n16611), .ZN(n16612) );
  AOI211_X1 U19832 ( .C1(n18809), .C2(n18806), .A(n16612), .B(n16622), .ZN(
        n16614) );
  INV_X1 U19833 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17545) );
  OAI22_X1 U19834 ( .A1(n17545), .A2(n16934), .B1(n16943), .B2(n20898), .ZN(
        n16613) );
  AOI211_X1 U19835 ( .C1(n16634), .C2(P3_REIP_REG_28__SCAN_IN), .A(n16614), 
        .B(n16613), .ZN(n16620) );
  OAI211_X1 U19836 ( .C1(n16621), .C2(n20898), .A(n16890), .B(n16615), .ZN(
        n16619) );
  OAI211_X1 U19837 ( .C1(n17551), .C2(n16617), .A(n16904), .B(n16616), .ZN(
        n16618) );
  NAND3_X1 U19838 ( .A1(n16620), .A2(n16619), .A3(n16618), .ZN(P3_U2643) );
  AOI211_X1 U19839 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16635), .A(n16621), .B(
        n16944), .ZN(n16624) );
  OAI22_X1 U19840 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16622), .B1(n17546), 
        .B2(n16934), .ZN(n16623) );
  AOI211_X1 U19841 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16921), .A(n16624), .B(
        n16623), .ZN(n16629) );
  OAI211_X1 U19842 ( .C1(n16627), .C2(n16626), .A(n16904), .B(n16625), .ZN(
        n16628) );
  OAI211_X1 U19843 ( .C1(n16630), .C2(n18806), .A(n16629), .B(n16628), .ZN(
        P3_U2644) );
  INV_X1 U19844 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18802) );
  NAND2_X1 U19845 ( .A1(n16926), .A2(n16631), .ZN(n16642) );
  NOR3_X1 U19846 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18802), .A3(n16642), 
        .ZN(n16633) );
  OAI22_X1 U19847 ( .A1(n17573), .A2(n16934), .B1(n16943), .B2(n16952), .ZN(
        n16632) );
  AOI211_X1 U19848 ( .C1(n16634), .C2(P3_REIP_REG_26__SCAN_IN), .A(n16633), 
        .B(n16632), .ZN(n16640) );
  OAI211_X1 U19849 ( .C1(n16641), .C2(n16952), .A(n16890), .B(n16635), .ZN(
        n16639) );
  OAI211_X1 U19850 ( .C1(n17574), .C2(n16637), .A(n16904), .B(n16636), .ZN(
        n16638) );
  NAND3_X1 U19851 ( .A1(n16640), .A2(n16639), .A3(n16638), .ZN(P3_U2645) );
  AOI21_X1 U19852 ( .B1(n16650), .B2(n16926), .A(n16933), .ZN(n16670) );
  INV_X1 U19853 ( .A(n16670), .ZN(n16654) );
  AOI21_X1 U19854 ( .B1(n16926), .B2(n18800), .A(n16654), .ZN(n16649) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16655), .A(n16641), .B(
        n16944), .ZN(n16644) );
  OAI22_X1 U19856 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16642), .B1(n16951), 
        .B2(n16943), .ZN(n16643) );
  AOI211_X1 U19857 ( .C1(n16897), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16644), .B(n16643), .ZN(n16648) );
  OAI211_X1 U19858 ( .C1(n17586), .C2(n16646), .A(n16904), .B(n16645), .ZN(
        n16647) );
  OAI211_X1 U19859 ( .C1(n16649), .C2(n18802), .A(n16648), .B(n16647), .ZN(
        P3_U2646) );
  NOR3_X1 U19860 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16937), .A3(n16650), 
        .ZN(n16653) );
  OAI22_X1 U19861 ( .A1(n16651), .A2(n16934), .B1(n16943), .B2(n16954), .ZN(
        n16652) );
  AOI211_X1 U19862 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16654), .A(n16653), 
        .B(n16652), .ZN(n16660) );
  OAI211_X1 U19863 ( .C1(n16662), .C2(n16954), .A(n16890), .B(n16655), .ZN(
        n16659) );
  OAI211_X1 U19864 ( .C1(n17594), .C2(n16657), .A(n16904), .B(n16656), .ZN(
        n16658) );
  NAND3_X1 U19865 ( .A1(n16660), .A2(n16659), .A3(n16658), .ZN(P3_U2647) );
  AOI21_X1 U19866 ( .B1(n16926), .B2(n16661), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n16669) );
  AOI211_X1 U19867 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16675), .A(n16662), .B(
        n16944), .ZN(n16664) );
  NOR2_X1 U19868 ( .A1(n17609), .A2(n16934), .ZN(n16663) );
  AOI211_X1 U19869 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16921), .A(n16664), .B(
        n16663), .ZN(n16668) );
  OAI211_X1 U19870 ( .C1(n17611), .C2(n16666), .A(n16904), .B(n16665), .ZN(
        n16667) );
  OAI211_X1 U19871 ( .C1(n16670), .C2(n16669), .A(n16668), .B(n16667), .ZN(
        P3_U2648) );
  OR3_X1 U19872 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16937), .A3(n16676), .ZN(
        n16686) );
  AOI21_X1 U19873 ( .B1(n16676), .B2(n16926), .A(n16933), .ZN(n16691) );
  AOI22_X1 U19874 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16897), .B1(
        n16921), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16671) );
  OAI221_X1 U19875 ( .B1(n16686), .B2(n18796), .C1(n16691), .C2(n18796), .A(
        n16671), .ZN(n16672) );
  INV_X1 U19876 ( .A(n16672), .ZN(n16681) );
  OAI211_X1 U19877 ( .C1(n17622), .C2(n16674), .A(n16904), .B(n16673), .ZN(
        n16680) );
  OAI211_X1 U19878 ( .C1(n16682), .C2(n17019), .A(n16890), .B(n16675), .ZN(
        n16679) );
  NOR2_X1 U19879 ( .A1(n16937), .A2(n16676), .ZN(n16677) );
  NAND3_X1 U19880 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16677), .A3(n18796), 
        .ZN(n16678) );
  NAND4_X1 U19881 ( .A1(n16681), .A2(n16680), .A3(n16679), .A4(n16678), .ZN(
        P3_U2649) );
  AOI211_X1 U19882 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16696), .A(n16682), .B(
        n16944), .ZN(n16689) );
  OAI211_X1 U19883 ( .C1(n17632), .C2(n16684), .A(n16904), .B(n16683), .ZN(
        n16685) );
  OAI211_X1 U19884 ( .C1(n16934), .C2(n16687), .A(n16686), .B(n16685), .ZN(
        n16688) );
  AOI211_X1 U19885 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16921), .A(n16689), .B(
        n16688), .ZN(n16690) );
  OAI21_X1 U19886 ( .B1(n16691), .B2(n18795), .A(n16690), .ZN(P3_U2650) );
  INV_X1 U19887 ( .A(n16691), .ZN(n16693) );
  OAI22_X1 U19888 ( .A1(n20809), .A2(n16934), .B1(n16943), .B2(n17064), .ZN(
        n16692) );
  AOI21_X1 U19889 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16693), .A(n16692), 
        .ZN(n16700) );
  OAI211_X1 U19890 ( .C1(n17644), .C2(n16695), .A(n16904), .B(n16694), .ZN(
        n16699) );
  OAI211_X1 U19891 ( .C1(n16704), .C2(n17064), .A(n16890), .B(n16696), .ZN(
        n16698) );
  INV_X1 U19892 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18791) );
  INV_X1 U19893 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18789) );
  NAND2_X1 U19894 ( .A1(n16926), .A2(n16728), .ZN(n16709) );
  OR4_X1 U19895 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18791), .A3(n18789), .A4(
        n16709), .ZN(n16697) );
  NAND4_X1 U19896 ( .A1(n16700), .A2(n16699), .A3(n16698), .A4(n16697), .ZN(
        P3_U2651) );
  INV_X1 U19897 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16724) );
  INV_X1 U19898 ( .A(n17652), .ZN(n16713) );
  NOR2_X1 U19899 ( .A1(n16724), .A2(n16713), .ZN(n16702) );
  INV_X1 U19900 ( .A(n17617), .ZN(n16701) );
  OAI21_X1 U19901 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16702), .A(
        n16701), .ZN(n17654) );
  OAI21_X1 U19902 ( .B1(n16724), .B2(n16714), .A(n16903), .ZN(n16703) );
  XNOR2_X1 U19903 ( .A(n17654), .B(n16703), .ZN(n16712) );
  AOI211_X1 U19904 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16721), .A(n16704), .B(
        n16944), .ZN(n16708) );
  NOR3_X1 U19905 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18789), .A3(n16709), 
        .ZN(n16707) );
  INV_X1 U19906 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16705) );
  OAI22_X1 U19907 ( .A1(n16705), .A2(n16934), .B1(n16943), .B2(n20777), .ZN(
        n16706) );
  NOR4_X1 U19908 ( .A1(n18209), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        n16711) );
  NOR2_X1 U19909 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16709), .ZN(n16717) );
  OAI21_X1 U19910 ( .B1(n16728), .B2(n16937), .A(n16946), .ZN(n16733) );
  OAI21_X1 U19911 ( .B1(n16717), .B2(n16733), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16710) );
  OAI211_X1 U19912 ( .C1(n16712), .C2(n18734), .A(n16711), .B(n16710), .ZN(
        P3_U2652) );
  AOI22_X1 U19913 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16713), .B1(
        n17652), .B2(n16724), .ZN(n17666) );
  NAND2_X1 U19914 ( .A1(n16903), .A2(n16714), .ZN(n16716) );
  OAI21_X1 U19915 ( .B1(n17666), .B2(n16716), .A(n16904), .ZN(n16715) );
  AOI21_X1 U19916 ( .B1(n17666), .B2(n16716), .A(n16715), .ZN(n16720) );
  INV_X1 U19917 ( .A(n16717), .ZN(n16718) );
  OAI211_X1 U19918 ( .C1(n16943), .C2(n17076), .A(n18175), .B(n16718), .ZN(
        n16719) );
  AOI211_X1 U19919 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n16733), .A(n16720), 
        .B(n16719), .ZN(n16723) );
  OAI211_X1 U19920 ( .C1(n16726), .C2(n17076), .A(n16890), .B(n16721), .ZN(
        n16722) );
  OAI211_X1 U19921 ( .C1(n16934), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        P3_U2653) );
  AOI21_X1 U19922 ( .B1(n17680), .B2(n16739), .A(n17652), .ZN(n17684) );
  AOI21_X1 U19923 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16741), .A(
        n16874), .ZN(n16725) );
  XNOR2_X1 U19924 ( .A(n17684), .B(n16725), .ZN(n16736) );
  AOI211_X1 U19925 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16746), .A(n16726), .B(
        n16944), .ZN(n16727) );
  AOI21_X1 U19926 ( .B1(n16897), .B2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16727), .ZN(n16735) );
  OR2_X1 U19927 ( .A1(n16937), .A2(n16728), .ZN(n16729) );
  OAI22_X1 U19928 ( .A1(n16943), .A2(n16731), .B1(n16730), .B2(n16729), .ZN(
        n16732) );
  AOI211_X1 U19929 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n16733), .A(n18209), 
        .B(n16732), .ZN(n16734) );
  OAI211_X1 U19930 ( .C1(n18734), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P3_U2654) );
  AOI22_X1 U19931 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16897), .B1(
        n16921), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16749) );
  OAI21_X1 U19932 ( .B1(n16737), .B2(n16937), .A(n16946), .ZN(n16770) );
  INV_X1 U19933 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18786) );
  INV_X1 U19934 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18784) );
  NOR2_X1 U19935 ( .A1(n16937), .A2(n16738), .ZN(n16769) );
  NAND2_X1 U19936 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16769), .ZN(n16761) );
  AOI221_X1 U19937 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n18786), .C2(n18784), .A(n16761), .ZN(n16745) );
  INV_X1 U19938 ( .A(n16750), .ZN(n16740) );
  OAI21_X1 U19939 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16740), .A(
        n16739), .ZN(n17699) );
  INV_X1 U19940 ( .A(n17699), .ZN(n16743) );
  NOR2_X1 U19941 ( .A1(n16741), .A2(n16874), .ZN(n16754) );
  INV_X1 U19942 ( .A(n16754), .ZN(n16742) );
  AOI221_X1 U19943 ( .B1(n16743), .B2(n16754), .C1(n17699), .C2(n16742), .A(
        n18734), .ZN(n16744) );
  AOI211_X1 U19944 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16770), .A(n16745), 
        .B(n16744), .ZN(n16748) );
  OAI211_X1 U19945 ( .C1(n16753), .C2(n17111), .A(n16890), .B(n16746), .ZN(
        n16747) );
  NAND4_X1 U19946 ( .A1(n16749), .A2(n16748), .A3(n18175), .A4(n16747), .ZN(
        P3_U2655) );
  AOI21_X1 U19947 ( .B1(n16903), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18734), .ZN(n16940) );
  INV_X1 U19948 ( .A(n17693), .ZN(n16751) );
  OAI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17693), .A(
        n16750), .ZN(n17709) );
  AOI21_X1 U19950 ( .B1(n16903), .B2(n16751), .A(n17709), .ZN(n16752) );
  AOI22_X1 U19951 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16897), .B1(
        n16940), .B2(n16752), .ZN(n16760) );
  AOI211_X1 U19952 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16764), .A(n16753), .B(
        n16944), .ZN(n16758) );
  INV_X1 U19953 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16756) );
  NAND3_X1 U19954 ( .A1(n16904), .A2(n16754), .A3(n17709), .ZN(n16755) );
  OAI211_X1 U19955 ( .C1(n16943), .C2(n16756), .A(n18175), .B(n16755), .ZN(
        n16757) );
  AOI211_X1 U19956 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n16770), .A(n16758), 
        .B(n16757), .ZN(n16759) );
  OAI211_X1 U19957 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n16761), .A(n16760), 
        .B(n16759), .ZN(P3_U2656) );
  INV_X1 U19958 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16767) );
  INV_X1 U19959 ( .A(n17739), .ZN(n16799) );
  NAND2_X1 U19960 ( .A1(n17736), .A2(n16799), .ZN(n16774) );
  AOI21_X1 U19961 ( .B1(n16767), .B2(n16774), .A(n17693), .ZN(n17729) );
  INV_X1 U19962 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16800) );
  NOR2_X1 U19963 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17894), .ZN(
        n16924) );
  NAND2_X1 U19964 ( .A1(n17775), .A2(n16924), .ZN(n16801) );
  OAI21_X1 U19965 ( .B1(n16800), .B2(n16801), .A(n16903), .ZN(n16786) );
  OAI21_X1 U19966 ( .B1(n17736), .B2(n16874), .A(n16786), .ZN(n16782) );
  INV_X1 U19967 ( .A(n17729), .ZN(n16763) );
  INV_X1 U19968 ( .A(n16782), .ZN(n16762) );
  OAI221_X1 U19969 ( .B1(n17729), .B2(n16782), .C1(n16763), .C2(n16762), .A(
        n16904), .ZN(n16766) );
  OAI211_X1 U19970 ( .C1(n16772), .C2(n17140), .A(n16890), .B(n16764), .ZN(
        n16765) );
  OAI211_X1 U19971 ( .C1(n16934), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        n16768) );
  AOI221_X1 U19972 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16770), .C1(n16769), 
        .C2(n16770), .A(n16768), .ZN(n16771) );
  OAI211_X1 U19973 ( .C1(n16943), .C2(n17140), .A(n16771), .B(n18175), .ZN(
        P3_U2657) );
  AOI211_X1 U19974 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16792), .A(n16772), .B(
        n16944), .ZN(n16781) );
  INV_X1 U19975 ( .A(n16773), .ZN(n16788) );
  OAI21_X1 U19976 ( .B1(n16788), .B2(n16937), .A(n16946), .ZN(n16797) );
  NOR2_X1 U19977 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16937), .ZN(n16787) );
  OAI21_X1 U19978 ( .B1(n16797), .B2(n16787), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16779) );
  NOR2_X1 U19979 ( .A1(n17750), .A2(n17739), .ZN(n16785) );
  OAI21_X1 U19980 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16785), .A(
        n16774), .ZN(n17740) );
  INV_X1 U19981 ( .A(n17740), .ZN(n16775) );
  OAI211_X1 U19982 ( .C1(n17742), .C2(n16874), .A(n16775), .B(n16940), .ZN(
        n16778) );
  INV_X1 U19983 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18780) );
  NAND3_X1 U19984 ( .A1(n16926), .A2(n16776), .A3(n18780), .ZN(n16777) );
  NAND4_X1 U19985 ( .A1(n18175), .A2(n16779), .A3(n16778), .A4(n16777), .ZN(
        n16780) );
  AOI211_X1 U19986 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16921), .A(n16781), .B(
        n16780), .ZN(n16784) );
  NAND3_X1 U19987 ( .A1(n16904), .A2(n17740), .A3(n16782), .ZN(n16783) );
  OAI211_X1 U19988 ( .C1(n16934), .C2(n17742), .A(n16784), .B(n16783), .ZN(
        P3_U2658) );
  AOI21_X1 U19989 ( .B1(n17750), .B2(n17739), .A(n16785), .ZN(n17753) );
  XOR2_X1 U19990 ( .A(n17753), .B(n16786), .Z(n16790) );
  AOI22_X1 U19991 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16897), .B1(
        n16788), .B2(n16787), .ZN(n16789) );
  OAI211_X1 U19992 ( .C1(n18734), .C2(n16790), .A(n16789), .B(n18175), .ZN(
        n16791) );
  AOI21_X1 U19993 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16797), .A(n16791), 
        .ZN(n16794) );
  OAI211_X1 U19994 ( .C1(n16795), .C2(n17127), .A(n16890), .B(n16792), .ZN(
        n16793) );
  OAI211_X1 U19995 ( .C1(n17127), .C2(n16943), .A(n16794), .B(n16793), .ZN(
        P3_U2659) );
  INV_X1 U19996 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16809) );
  AOI211_X1 U19997 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16813), .A(n16795), .B(
        n16944), .ZN(n16807) );
  AOI21_X1 U19998 ( .B1(n16926), .B2(n16796), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16805) );
  INV_X1 U19999 ( .A(n16797), .ZN(n16804) );
  NOR2_X1 U20000 ( .A1(n17894), .A2(n17845), .ZN(n16875) );
  INV_X1 U20001 ( .A(n16875), .ZN(n16884) );
  NOR2_X1 U20002 ( .A1(n17844), .A2(n16884), .ZN(n16873) );
  NAND2_X1 U20003 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16873), .ZN(
        n16859) );
  OR2_X1 U20004 ( .A1(n16798), .A2(n16859), .ZN(n16810) );
  AOI21_X1 U20005 ( .B1(n16800), .B2(n16810), .A(n16799), .ZN(n17767) );
  NAND2_X1 U20006 ( .A1(n16903), .A2(n16801), .ZN(n16802) );
  XOR2_X1 U20007 ( .A(n17767), .B(n16802), .Z(n16803) );
  OAI22_X1 U20008 ( .A1(n16805), .A2(n16804), .B1(n18734), .B2(n16803), .ZN(
        n16806) );
  AOI211_X1 U20009 ( .C1(n16897), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16807), .B(n16806), .ZN(n16808) );
  OAI211_X1 U20010 ( .C1(n16943), .C2(n16809), .A(n16808), .B(n18175), .ZN(
        P3_U2660) );
  INV_X1 U20011 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17787) );
  NOR2_X1 U20012 ( .A1(n17820), .A2(n16859), .ZN(n16848) );
  NAND2_X1 U20013 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16848), .ZN(
        n16835) );
  NOR2_X1 U20014 ( .A1(n17787), .A2(n16835), .ZN(n16822) );
  OAI21_X1 U20015 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16822), .A(
        n16810), .ZN(n17784) );
  NOR2_X1 U20016 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16859), .ZN(
        n16858) );
  NAND2_X1 U20017 ( .A1(n17802), .A2(n16858), .ZN(n16823) );
  INV_X1 U20018 ( .A(n16823), .ZN(n16811) );
  AOI21_X1 U20019 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16811), .A(
        n16874), .ZN(n16825) );
  XOR2_X1 U20020 ( .A(n17784), .B(n16825), .Z(n16820) );
  NOR3_X1 U20021 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16937), .A3(n16812), 
        .ZN(n16817) );
  INV_X1 U20022 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16815) );
  OAI211_X1 U20023 ( .C1(n16821), .C2(n17108), .A(n16890), .B(n16813), .ZN(
        n16814) );
  OAI211_X1 U20024 ( .C1(n16815), .C2(n16934), .A(n18175), .B(n16814), .ZN(
        n16816) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16921), .A(n16817), .B(
        n16816), .ZN(n16819) );
  NOR2_X1 U20026 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16937), .ZN(n16826) );
  OAI21_X1 U20027 ( .B1(n16827), .B2(n16937), .A(n16946), .ZN(n16842) );
  OAI21_X1 U20028 ( .B1(n16826), .B2(n16842), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16818) );
  OAI211_X1 U20029 ( .C1(n16820), .C2(n18734), .A(n16819), .B(n16818), .ZN(
        P3_U2661) );
  INV_X1 U20030 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16834) );
  AOI211_X1 U20031 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16843), .A(n16821), .B(
        n16944), .ZN(n16832) );
  INV_X1 U20032 ( .A(n16842), .ZN(n16830) );
  INV_X1 U20033 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18772) );
  AOI21_X1 U20034 ( .B1(n17787), .B2(n16835), .A(n16822), .ZN(n17791) );
  NOR2_X1 U20035 ( .A1(n16903), .A2(n18734), .ZN(n16886) );
  AOI21_X1 U20036 ( .B1(n17791), .B2(n16823), .A(n18734), .ZN(n16824) );
  OAI22_X1 U20037 ( .A1(n17791), .A2(n16825), .B1(n16886), .B2(n16824), .ZN(
        n16829) );
  NAND2_X1 U20038 ( .A1(n16827), .A2(n16826), .ZN(n16828) );
  OAI211_X1 U20039 ( .C1(n16830), .C2(n18772), .A(n16829), .B(n16828), .ZN(
        n16831) );
  AOI211_X1 U20040 ( .C1(n16897), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16832), .B(n16831), .ZN(n16833) );
  OAI211_X1 U20041 ( .C1(n16943), .C2(n16834), .A(n16833), .B(n18175), .ZN(
        P3_U2662) );
  OAI21_X1 U20042 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16848), .A(
        n16835), .ZN(n17807) );
  OR2_X1 U20043 ( .A1(n17804), .A2(n17820), .ZN(n17803) );
  INV_X1 U20044 ( .A(n16924), .ZN(n16836) );
  OAI21_X1 U20045 ( .B1(n17803), .B2(n16836), .A(n16903), .ZN(n16850) );
  OAI21_X1 U20046 ( .B1(n17807), .B2(n16850), .A(n16904), .ZN(n16837) );
  AOI21_X1 U20047 ( .B1(n17807), .B2(n16850), .A(n16837), .ZN(n16841) );
  OR4_X1 U20048 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16937), .A3(n16860), .A4(
        n16838), .ZN(n16839) );
  OAI211_X1 U20049 ( .C1(n16943), .C2(n16844), .A(n18175), .B(n16839), .ZN(
        n16840) );
  AOI211_X1 U20050 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16842), .A(n16841), .B(
        n16840), .ZN(n16846) );
  OAI211_X1 U20051 ( .C1(n16847), .C2(n16844), .A(n16890), .B(n16843), .ZN(
        n16845) );
  OAI211_X1 U20052 ( .C1(n16934), .C2(n17806), .A(n16846), .B(n16845), .ZN(
        P3_U2663) );
  INV_X1 U20053 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18766) );
  AOI221_X1 U20054 ( .B1(n16860), .B2(n16926), .C1(n18766), .C2(n16926), .A(
        n16933), .ZN(n16857) );
  INV_X1 U20055 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18768) );
  AOI22_X1 U20056 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16897), .B1(
        n16921), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16856) );
  AOI211_X1 U20057 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16862), .A(n16847), .B(
        n16944), .ZN(n16854) );
  NOR2_X1 U20058 ( .A1(n16858), .A2(n16874), .ZN(n16851) );
  AOI21_X1 U20059 ( .B1(n17820), .B2(n16859), .A(n16848), .ZN(n17827) );
  INV_X1 U20060 ( .A(n17827), .ZN(n16849) );
  AOI221_X1 U20061 ( .B1(n16851), .B2(n17827), .C1(n16850), .C2(n16849), .A(
        n18734), .ZN(n16853) );
  NOR4_X1 U20062 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16860), .A3(n16937), .A4(
        n18766), .ZN(n16852) );
  NOR4_X1 U20063 ( .A1(n18209), .A2(n16854), .A3(n16853), .A4(n16852), .ZN(
        n16855) );
  OAI211_X1 U20064 ( .C1(n16857), .C2(n18768), .A(n16856), .B(n16855), .ZN(
        P3_U2664) );
  AOI21_X1 U20065 ( .B1(n16926), .B2(n16860), .A(n16933), .ZN(n16878) );
  NOR2_X1 U20066 ( .A1(n16858), .A2(n16935), .ZN(n16867) );
  OAI21_X1 U20067 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16873), .A(
        n16859), .ZN(n17837) );
  INV_X1 U20068 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17836) );
  OAI21_X1 U20069 ( .B1(n17836), .B2(n16934), .A(n18175), .ZN(n16866) );
  NOR2_X1 U20070 ( .A1(n16937), .A2(n16860), .ZN(n16861) );
  NAND2_X1 U20071 ( .A1(n16861), .A2(n18766), .ZN(n16864) );
  OAI211_X1 U20072 ( .C1(n16871), .C2(n17233), .A(n16890), .B(n16862), .ZN(
        n16863) );
  OAI211_X1 U20073 ( .C1(n17233), .C2(n16943), .A(n16864), .B(n16863), .ZN(
        n16865) );
  AOI211_X1 U20074 ( .C1(n16867), .C2(n17837), .A(n16866), .B(n16865), .ZN(
        n16870) );
  INV_X1 U20075 ( .A(n17837), .ZN(n16868) );
  OAI211_X1 U20076 ( .C1(n16873), .C2(n16886), .A(n16868), .B(n16940), .ZN(
        n16869) );
  OAI211_X1 U20077 ( .C1(n16878), .C2(n18766), .A(n16870), .B(n16869), .ZN(
        P3_U2665) );
  INV_X1 U20078 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16882) );
  AOI211_X1 U20079 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16889), .A(n16871), .B(
        n16944), .ZN(n16880) );
  AOI21_X1 U20080 ( .B1(n16926), .B2(n16872), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16877) );
  AOI21_X1 U20081 ( .B1(n17844), .B2(n16884), .A(n16873), .ZN(n17852) );
  INV_X1 U20082 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16936) );
  AOI21_X1 U20083 ( .B1(n16936), .B2(n16875), .A(n16874), .ZN(n16885) );
  XNOR2_X1 U20084 ( .A(n17852), .B(n16885), .ZN(n16876) );
  OAI22_X1 U20085 ( .A1(n16878), .A2(n16877), .B1(n18734), .B2(n16876), .ZN(
        n16879) );
  AOI211_X1 U20086 ( .C1(n16897), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16880), .B(n16879), .ZN(n16881) );
  OAI211_X1 U20087 ( .C1(n16943), .C2(n16882), .A(n16881), .B(n18175), .ZN(
        P3_U2666) );
  NOR2_X1 U20088 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16883), .ZN(
        n17857) );
  NOR2_X1 U20089 ( .A1(n17894), .A2(n16883), .ZN(n16900) );
  OAI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16900), .A(
        n16884), .ZN(n17863) );
  AOI22_X1 U20091 ( .A1(n16924), .A2(n17857), .B1(n16885), .B2(n17863), .ZN(
        n16896) );
  NAND2_X1 U20092 ( .A1(n17433), .A2(n18890), .ZN(n16916) );
  INV_X1 U20093 ( .A(n16886), .ZN(n16918) );
  OAI22_X1 U20094 ( .A1(n16943), .A2(n17105), .B1(n17863), .B2(n16918), .ZN(
        n16887) );
  INV_X1 U20095 ( .A(n16887), .ZN(n16888) );
  OAI221_X1 U20096 ( .B1(n16916), .B2(n18663), .C1(n16916), .C2(n18716), .A(
        n16888), .ZN(n16894) );
  OR2_X1 U20097 ( .A1(n16937), .A2(n16907), .ZN(n16892) );
  AOI21_X1 U20098 ( .B1(n16926), .B2(n16907), .A(n16933), .ZN(n16914) );
  OAI211_X1 U20099 ( .C1(n16898), .C2(n17105), .A(n16890), .B(n16889), .ZN(
        n16891) );
  OAI221_X1 U20100 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16892), .C1(n18762), 
        .C2(n16914), .A(n16891), .ZN(n16893) );
  AOI211_X1 U20101 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16897), .A(
        n16894), .B(n16893), .ZN(n16895) );
  OAI211_X1 U20102 ( .C1(n16896), .C2(n18734), .A(n16895), .B(n18175), .ZN(
        P3_U2667) );
  INV_X1 U20103 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18760) );
  AOI22_X1 U20104 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16897), .B1(
        n16921), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16913) );
  AOI211_X1 U20105 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16899), .A(n16898), .B(
        n16944), .ZN(n16911) );
  INV_X1 U20106 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17887) );
  NOR2_X1 U20107 ( .A1(n17894), .A2(n17887), .ZN(n16902) );
  INV_X1 U20108 ( .A(n16900), .ZN(n16901) );
  OAI21_X1 U20109 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16902), .A(
        n16901), .ZN(n17873) );
  NAND2_X1 U20110 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16924), .ZN(
        n16922) );
  NAND2_X1 U20111 ( .A1(n16922), .A2(n16903), .ZN(n16906) );
  OAI21_X1 U20112 ( .B1(n17873), .B2(n16906), .A(n16904), .ZN(n16905) );
  AOI21_X1 U20113 ( .B1(n17873), .B2(n16906), .A(n16905), .ZN(n16910) );
  NOR2_X1 U20114 ( .A1(n9714), .A2(n18849), .ZN(n18667) );
  NAND2_X1 U20115 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18667), .ZN(
        n16915) );
  AOI21_X1 U20116 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16915), .A(
        n17155), .ZN(n18833) );
  NAND2_X1 U20117 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16925) );
  NAND2_X1 U20118 ( .A1(n16926), .A2(n16907), .ZN(n16908) );
  OAI22_X1 U20119 ( .A1(n18833), .A2(n16916), .B1(n16925), .B2(n16908), .ZN(
        n16909) );
  NOR3_X1 U20120 ( .A1(n16911), .A2(n16910), .A3(n16909), .ZN(n16912) );
  OAI211_X1 U20121 ( .C1(n16914), .C2(n18760), .A(n16913), .B(n16912), .ZN(
        P3_U2668) );
  NAND2_X1 U20122 ( .A1(n9714), .A2(n18675), .ZN(n18659) );
  NAND2_X1 U20123 ( .A1(n18659), .A2(n16915), .ZN(n18681) );
  INV_X1 U20124 ( .A(n18681), .ZN(n18839) );
  INV_X1 U20125 ( .A(n16916), .ZN(n18892) );
  AOI22_X1 U20126 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16933), .B1(n18839), 
        .B2(n18892), .ZN(n16930) );
  AOI211_X1 U20127 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16931), .A(n16917), .B(
        n16944), .ZN(n16920) );
  AOI22_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17887), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17894), .ZN(n17884) );
  OAI22_X1 U20129 ( .A1(n17887), .A2(n16934), .B1(n17884), .B2(n16918), .ZN(
        n16919) );
  AOI211_X1 U20130 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16921), .A(n16920), .B(
        n16919), .ZN(n16929) );
  INV_X1 U20131 ( .A(n16935), .ZN(n16923) );
  OAI211_X1 U20132 ( .C1(n16924), .C2(n17884), .A(n16923), .B(n16922), .ZN(
        n16928) );
  OAI211_X1 U20133 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16926), .B(n16925), .ZN(n16927) );
  NAND4_X1 U20134 ( .A1(n16930), .A2(n16929), .A3(n16928), .A4(n16927), .ZN(
        P3_U2669) );
  NAND2_X1 U20135 ( .A1(n16931), .A2(n17252), .ZN(n17262) );
  AND2_X1 U20136 ( .A1(n18675), .A2(n16932), .ZN(n18846) );
  AOI22_X1 U20137 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16933), .B1(n18846), 
        .B2(n18892), .ZN(n16942) );
  OAI21_X1 U20138 ( .B1(n16936), .B2(n16935), .A(n16934), .ZN(n16939) );
  INV_X1 U20139 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17261) );
  OAI22_X1 U20140 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16937), .B1(n16943), 
        .B2(n17261), .ZN(n16938) );
  AOI221_X1 U20141 ( .B1(n16940), .B2(n17894), .C1(n16939), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16938), .ZN(n16941) );
  OAI211_X1 U20142 ( .C1(n16944), .C2(n17262), .A(n16942), .B(n16941), .ZN(
        P3_U2670) );
  INV_X1 U20143 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U20144 ( .A1(n16944), .A2(n16943), .ZN(n16945) );
  AOI22_X1 U20145 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16945), .B1(n18892), .B2(
        n12933), .ZN(n16948) );
  NAND3_X1 U20146 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18852), .A3(
        n16946), .ZN(n16947) );
  OAI211_X1 U20147 ( .C1(n16949), .C2(n18864), .A(n16948), .B(n16947), .ZN(
        P3_U2671) );
  INV_X1 U20148 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16959) );
  NOR3_X1 U20149 ( .A1(n16952), .A2(n16951), .A3(n16950), .ZN(n16991) );
  NAND2_X1 U20150 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20775), .ZN(n17045) );
  NOR4_X1 U20151 ( .A1(n16954), .A2(n16953), .A3(n17019), .A4(n17045), .ZN(
        n16955) );
  NAND4_X1 U20152 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16991), .A4(n16955), .ZN(n16958) );
  NOR2_X1 U20153 ( .A1(n16959), .A2(n16958), .ZN(n16985) );
  NAND2_X1 U20154 ( .A1(n17258), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16957) );
  NAND2_X1 U20155 ( .A1(n16985), .A2(n17232), .ZN(n16956) );
  OAI22_X1 U20156 ( .A1(n16985), .A2(n16957), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16956), .ZN(P3_U2672) );
  NAND2_X1 U20157 ( .A1(n16959), .A2(n16958), .ZN(n16960) );
  NAND2_X1 U20158 ( .A1(n16960), .A2(n17258), .ZN(n16984) );
  AOI22_X1 U20159 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20160 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12684), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20161 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20162 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16961) );
  NAND4_X1 U20163 ( .A1(n16964), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        n16970) );
  AOI22_X1 U20164 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20165 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20166 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20167 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16965) );
  NAND4_X1 U20168 ( .A1(n16968), .A2(n16967), .A3(n16966), .A4(n16965), .ZN(
        n16969) );
  NOR2_X1 U20169 ( .A1(n16970), .A2(n16969), .ZN(n16983) );
  AOI22_X1 U20170 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20171 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20172 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16972) );
  OAI21_X1 U20173 ( .B1(n17188), .B2(n17238), .A(n16972), .ZN(n16979) );
  AOI22_X1 U20174 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20175 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20176 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16973), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20177 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16974) );
  NAND4_X1 U20178 ( .A1(n16977), .A2(n16976), .A3(n16975), .A4(n16974), .ZN(
        n16978) );
  AOI211_X1 U20179 ( .C1(n17330), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n16979), .B(n16978), .ZN(n16980) );
  NAND3_X1 U20180 ( .A1(n16982), .A2(n16981), .A3(n16980), .ZN(n16987) );
  NAND2_X1 U20181 ( .A1(n16988), .A2(n16987), .ZN(n16986) );
  XNOR2_X1 U20182 ( .A(n16983), .B(n16986), .ZN(n17273) );
  OAI22_X1 U20183 ( .A1(n16985), .A2(n16984), .B1(n17273), .B2(n17258), .ZN(
        P3_U2673) );
  OAI21_X1 U20184 ( .B1(n16988), .B2(n16987), .A(n16986), .ZN(n17280) );
  INV_X1 U20185 ( .A(n16989), .ZN(n16992) );
  NOR2_X1 U20186 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17007), .ZN(n16990) );
  AOI22_X1 U20187 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16992), .B1(n16991), 
        .B2(n16990), .ZN(n16993) );
  OAI21_X1 U20188 ( .B1(n17280), .B2(n17258), .A(n16993), .ZN(P3_U2674) );
  OAI21_X1 U20189 ( .B1(n16998), .B2(n16995), .A(n16994), .ZN(n17290) );
  OAI211_X1 U20190 ( .C1(n17003), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17258), .B(
        n16996), .ZN(n16997) );
  OAI21_X1 U20191 ( .B1(n17258), .B2(n17290), .A(n16997), .ZN(P3_U2676) );
  INV_X1 U20192 ( .A(n17007), .ZN(n17012) );
  NAND2_X1 U20193 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17012), .ZN(n17002) );
  AOI21_X1 U20194 ( .B1(n16999), .B2(n17004), .A(n16998), .ZN(n17291) );
  AOI22_X1 U20195 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17000), .B1(n17291), 
        .B2(n20780), .ZN(n17001) );
  OAI21_X1 U20196 ( .B1(n17003), .B2(n17002), .A(n17001), .ZN(P3_U2677) );
  OAI21_X1 U20197 ( .B1(n17008), .B2(n17005), .A(n17004), .ZN(n17300) );
  NAND3_X1 U20198 ( .A1(n17007), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n17258), 
        .ZN(n17006) );
  OAI221_X1 U20199 ( .B1(n17007), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17258), 
        .C2(n17300), .A(n17006), .ZN(P3_U2678) );
  AOI21_X1 U20200 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17258), .A(n17017), .ZN(
        n17011) );
  AOI21_X1 U20201 ( .B1(n17009), .B2(n17013), .A(n17008), .ZN(n17301) );
  INV_X1 U20202 ( .A(n17301), .ZN(n17010) );
  OAI22_X1 U20203 ( .A1(n17012), .A2(n17011), .B1(n17010), .B2(n17258), .ZN(
        P3_U2679) );
  NOR2_X1 U20204 ( .A1(n17019), .A2(n17018), .ZN(n17034) );
  AOI21_X1 U20205 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17258), .A(n17034), .ZN(
        n17016) );
  OAI21_X1 U20206 ( .B1(n17015), .B2(n17014), .A(n17013), .ZN(n17310) );
  OAI22_X1 U20207 ( .A1(n17017), .A2(n17016), .B1(n17310), .B2(n17258), .ZN(
        P3_U2680) );
  OAI21_X1 U20208 ( .B1(n17019), .B2(n20780), .A(n17018), .ZN(n17020) );
  INV_X1 U20209 ( .A(n17020), .ZN(n17033) );
  AOI22_X1 U20210 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20211 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20212 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17021) );
  OAI21_X1 U20213 ( .B1(n17022), .B2(n17238), .A(n17021), .ZN(n17028) );
  AOI22_X1 U20214 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20215 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20216 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20217 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17023) );
  NAND4_X1 U20218 ( .A1(n17026), .A2(n17025), .A3(n17024), .A4(n17023), .ZN(
        n17027) );
  AOI211_X1 U20219 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17028), .B(n17027), .ZN(n17029) );
  NAND3_X1 U20220 ( .A1(n17031), .A2(n17030), .A3(n17029), .ZN(n17311) );
  INV_X1 U20221 ( .A(n17311), .ZN(n17032) );
  OAI22_X1 U20222 ( .A1(n17034), .A2(n17033), .B1(n17032), .B2(n17258), .ZN(
        P3_U2681) );
  AOI22_X1 U20223 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20224 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20225 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20226 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17035) );
  NAND4_X1 U20227 ( .A1(n17038), .A2(n17037), .A3(n17036), .A4(n17035), .ZN(
        n17044) );
  AOI22_X1 U20228 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20229 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20230 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20231 ( .A1(n17340), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20232 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17043) );
  NOR2_X1 U20233 ( .A1(n17044), .A2(n17043), .ZN(n17319) );
  NAND2_X1 U20234 ( .A1(n17258), .A2(n17045), .ZN(n17065) );
  INV_X1 U20235 ( .A(n17065), .ZN(n17048) );
  INV_X1 U20236 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20237 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17048), .B1(n17047), 
        .B2(n17046), .ZN(n17049) );
  OAI21_X1 U20238 ( .B1(n17319), .B2(n17258), .A(n17049), .ZN(P3_U2682) );
  AOI22_X1 U20239 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20240 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20241 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17050) );
  OAI21_X1 U20242 ( .B1(n17051), .B2(n20867), .A(n17050), .ZN(n17057) );
  AOI22_X1 U20243 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20244 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20245 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20246 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17052) );
  NAND4_X1 U20247 ( .A1(n17055), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17056) );
  AOI211_X1 U20248 ( .C1(n17058), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17057), .B(n17056), .ZN(n17059) );
  NAND3_X1 U20249 ( .A1(n17061), .A2(n17060), .A3(n17059), .ZN(n17322) );
  NAND2_X1 U20250 ( .A1(n20780), .A2(n17322), .ZN(n17062) );
  OAI221_X1 U20251 ( .B1(n17065), .B2(n17064), .C1(n17065), .C2(n17063), .A(
        n17062), .ZN(P3_U2683) );
  NAND2_X1 U20252 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20776), .ZN(n17078) );
  AOI22_X1 U20253 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20254 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20255 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20256 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17066) );
  NAND4_X1 U20257 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17075) );
  AOI22_X1 U20258 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20259 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20260 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20261 ( .A1(n17058), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20262 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20263 ( .A1(n17075), .A2(n17074), .ZN(n17358) );
  NAND3_X1 U20264 ( .A1(n17090), .A2(n17257), .A3(n17076), .ZN(n17077) );
  OAI221_X1 U20265 ( .B1(n20780), .B2(n17078), .C1(n17258), .C2(n17358), .A(
        n17077), .ZN(P3_U2685) );
  AOI22_X1 U20266 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17341), .B1(
        n15786), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20267 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20268 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17170), .ZN(n17080) );
  AOI22_X1 U20269 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20270 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17088) );
  AOI22_X1 U20271 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17214), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17331), .ZN(n17086) );
  AOI22_X1 U20272 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17328), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17340), .ZN(n17085) );
  AOI22_X1 U20273 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n12904), .ZN(n17084) );
  AOI22_X1 U20274 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17339), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17342), .ZN(n17083) );
  NAND4_X1 U20275 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20276 ( .A1(n17088), .A2(n17087), .ZN(n17363) );
  AOI21_X1 U20277 ( .B1(n17232), .B2(n17089), .A(n17263), .ZN(n17092) );
  NAND2_X1 U20278 ( .A1(n17090), .A2(n17257), .ZN(n17091) );
  OAI21_X1 U20279 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17092), .A(n17091), .ZN(
        n17093) );
  AOI21_X1 U20280 ( .B1(n17363), .B2(n20780), .A(n17093), .ZN(P3_U2686) );
  AOI22_X1 U20281 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20282 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17094), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20283 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20284 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17095) );
  NAND4_X1 U20285 ( .A1(n17098), .A2(n17097), .A3(n17096), .A4(n17095), .ZN(
        n17104) );
  AOI22_X1 U20286 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20287 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12686), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20288 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20289 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12904), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U20290 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17103) );
  NOR2_X1 U20291 ( .A1(n17104), .A2(n17103), .ZN(n17369) );
  NOR3_X1 U20292 ( .A1(n17105), .A2(n17263), .A3(n17244), .ZN(n17248) );
  INV_X1 U20293 ( .A(n17248), .ZN(n17106) );
  NOR2_X1 U20294 ( .A1(n17107), .A2(n17106), .ZN(n17236) );
  NAND2_X1 U20295 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17231), .ZN(n17212) );
  NOR2_X1 U20296 ( .A1(n17108), .A2(n17212), .ZN(n17200) );
  NAND2_X1 U20297 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17200), .ZN(n17181) );
  NOR2_X1 U20298 ( .A1(n17109), .A2(n17181), .ZN(n17124) );
  NAND2_X1 U20299 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17124), .ZN(n17123) );
  OAI21_X1 U20300 ( .B1(n20780), .B2(n17111), .A(n17123), .ZN(n17110) );
  OAI221_X1 U20301 ( .B1(n17232), .B2(n17123), .C1(n17123), .C2(n17111), .A(
        n17110), .ZN(n17112) );
  OAI21_X1 U20302 ( .B1(n17369), .B2(n17258), .A(n17112), .ZN(P3_U2687) );
  AOI22_X1 U20303 ( .A1(n12677), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20304 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20305 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20306 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17113) );
  NAND4_X1 U20307 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n17122) );
  AOI22_X1 U20308 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20309 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12904), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20310 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20311 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17117) );
  NAND4_X1 U20312 ( .A1(n17120), .A2(n17119), .A3(n17118), .A4(n17117), .ZN(
        n17121) );
  NOR2_X1 U20313 ( .A1(n17122), .A2(n17121), .ZN(n17373) );
  OAI211_X1 U20314 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17124), .A(n17123), .B(
        n17258), .ZN(n17125) );
  OAI21_X1 U20315 ( .B1(n17373), .B2(n17258), .A(n17125), .ZN(P3_U2688) );
  INV_X1 U20316 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17126) );
  NOR2_X1 U20317 ( .A1(n17127), .A2(n17181), .ZN(n17141) );
  NOR2_X1 U20318 ( .A1(n20780), .A2(n17141), .ZN(n17167) );
  AOI21_X1 U20319 ( .B1(n17257), .B2(n17126), .A(n17167), .ZN(n17154) );
  NOR4_X1 U20320 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18274), .A3(n17127), .A4(
        n17181), .ZN(n17138) );
  AOI22_X1 U20321 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20322 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20323 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17128) );
  OAI21_X1 U20324 ( .B1(n12760), .B2(n17238), .A(n17128), .ZN(n17134) );
  AOI22_X1 U20325 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20326 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20327 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20328 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20329 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  AOI211_X1 U20330 ( .C1(n17218), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17134), .B(n17133), .ZN(n17135) );
  NAND3_X1 U20331 ( .A1(n17137), .A2(n17136), .A3(n17135), .ZN(n17374) );
  AOI22_X1 U20332 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17138), .B1(n20780), 
        .B2(n17374), .ZN(n17139) );
  OAI21_X1 U20333 ( .B1(n17154), .B2(n17140), .A(n17139), .ZN(P3_U2689) );
  NOR2_X1 U20334 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17141), .ZN(n17153) );
  AOI22_X1 U20335 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20336 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12686), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20337 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20338 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17142) );
  NAND4_X1 U20339 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17152) );
  AOI22_X1 U20340 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20341 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20342 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17146), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20343 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17147) );
  NAND4_X1 U20344 ( .A1(n17150), .A2(n17149), .A3(n17148), .A4(n17147), .ZN(
        n17151) );
  NOR2_X1 U20345 ( .A1(n17152), .A2(n17151), .ZN(n17379) );
  OAI22_X1 U20346 ( .A1(n17154), .A2(n17153), .B1(n17379), .B2(n17258), .ZN(
        P3_U2690) );
  AOI22_X1 U20347 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20348 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20349 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17157) );
  AOI22_X1 U20350 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17156) );
  NAND4_X1 U20351 ( .A1(n17159), .A2(n17158), .A3(n17157), .A4(n17156), .ZN(
        n17166) );
  AOI22_X1 U20352 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20353 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20354 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20355 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17161) );
  NAND4_X1 U20356 ( .A1(n17164), .A2(n17163), .A3(n17162), .A4(n17161), .ZN(
        n17165) );
  NOR2_X1 U20357 ( .A1(n17166), .A2(n17165), .ZN(n17383) );
  INV_X1 U20358 ( .A(n17181), .ZN(n17168) );
  OAI21_X1 U20359 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17168), .A(n17167), .ZN(
        n17169) );
  OAI21_X1 U20360 ( .B1(n17383), .B2(n17258), .A(n17169), .ZN(P3_U2691) );
  AOI22_X1 U20361 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20362 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20363 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20364 ( .B1(n12760), .B2(n17251), .A(n17171), .ZN(n17177) );
  AOI22_X1 U20365 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20366 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20367 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20368 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17172) );
  NAND4_X1 U20369 ( .A1(n17175), .A2(n17174), .A3(n17173), .A4(n17172), .ZN(
        n17176) );
  AOI211_X1 U20370 ( .C1(n17334), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17177), .B(n17176), .ZN(n17178) );
  NAND3_X1 U20371 ( .A1(n17180), .A2(n17179), .A3(n17178), .ZN(n17386) );
  INV_X1 U20372 ( .A(n17386), .ZN(n17183) );
  OAI21_X1 U20373 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17200), .A(n17181), .ZN(
        n17182) );
  AOI22_X1 U20374 ( .A1(n20780), .A2(n17183), .B1(n17182), .B2(n17258), .ZN(
        P3_U2692) );
  INV_X1 U20375 ( .A(n17212), .ZN(n17184) );
  OAI21_X1 U20376 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17184), .A(n17258), .ZN(
        n17199) );
  AOI22_X1 U20377 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20378 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20379 ( .A1(n17186), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17187) );
  OAI21_X1 U20380 ( .B1(n17188), .B2(n20851), .A(n17187), .ZN(n17194) );
  AOI22_X1 U20381 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20382 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20383 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17329), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20384 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17189) );
  NAND4_X1 U20385 ( .A1(n17192), .A2(n17191), .A3(n17190), .A4(n17189), .ZN(
        n17193) );
  AOI211_X1 U20386 ( .C1(n17330), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17194), .B(n17193), .ZN(n17195) );
  NAND3_X1 U20387 ( .A1(n17197), .A2(n17196), .A3(n17195), .ZN(n17389) );
  INV_X1 U20388 ( .A(n17389), .ZN(n17198) );
  OAI22_X1 U20389 ( .A1(n17200), .A2(n17199), .B1(n17198), .B2(n17258), .ZN(
        P3_U2693) );
  AOI22_X1 U20390 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17331), .ZN(n17205) );
  AOI22_X1 U20391 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17339), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17340), .ZN(n17204) );
  AOI22_X1 U20392 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20393 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17341), .ZN(n17202) );
  NAND4_X1 U20394 ( .A1(n17205), .A2(n17204), .A3(n17203), .A4(n17202), .ZN(
        n17211) );
  AOI22_X1 U20395 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17332), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20396 ( .A1(n17328), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9599), .ZN(n17208) );
  AOI22_X1 U20397 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17342), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20398 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17329), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17170), .ZN(n17206) );
  NAND4_X1 U20399 ( .A1(n17209), .A2(n17208), .A3(n17207), .A4(n17206), .ZN(
        n17210) );
  NOR2_X1 U20400 ( .A1(n17211), .A2(n17210), .ZN(n17393) );
  OAI21_X1 U20401 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17231), .A(n17212), .ZN(
        n17213) );
  AOI22_X1 U20402 ( .A1(n20780), .A2(n17393), .B1(n17213), .B2(n17258), .ZN(
        P3_U2694) );
  OAI21_X1 U20403 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17236), .A(n17258), .ZN(
        n17230) );
  AOI22_X1 U20404 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20405 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17170), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20406 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17215) );
  OAI21_X1 U20407 ( .B1(n12760), .B2(n17216), .A(n17215), .ZN(n17225) );
  AOI22_X1 U20408 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20409 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17217), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20410 ( .A1(n17330), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20411 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17220) );
  NAND4_X1 U20412 ( .A1(n17223), .A2(n17222), .A3(n17221), .A4(n17220), .ZN(
        n17224) );
  AOI211_X1 U20413 ( .C1(n16971), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17225), .B(n17224), .ZN(n17226) );
  NAND3_X1 U20414 ( .A1(n17228), .A2(n17227), .A3(n17226), .ZN(n17396) );
  INV_X1 U20415 ( .A(n17396), .ZN(n17229) );
  OAI22_X1 U20416 ( .A1(n17231), .A2(n17230), .B1(n17229), .B2(n17258), .ZN(
        P3_U2695) );
  NAND3_X1 U20417 ( .A1(n17232), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n17248), .ZN(
        n17241) );
  NOR2_X1 U20418 ( .A1(n17233), .A2(n17241), .ZN(n17240) );
  AOI21_X1 U20419 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17258), .A(n17240), .ZN(
        n17235) );
  INV_X1 U20420 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17234) );
  OAI22_X1 U20421 ( .A1(n17236), .A2(n17235), .B1(n17234), .B2(n17258), .ZN(
        P3_U2696) );
  INV_X1 U20422 ( .A(n17241), .ZN(n17237) );
  AOI21_X1 U20423 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17258), .A(n17237), .ZN(
        n17239) );
  OAI22_X1 U20424 ( .A1(n17240), .A2(n17239), .B1(n17238), .B2(n17258), .ZN(
        P3_U2697) );
  INV_X1 U20425 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17243) );
  OAI21_X1 U20426 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17248), .A(n17241), .ZN(
        n17242) );
  AOI22_X1 U20427 ( .A1(n20780), .A2(n17243), .B1(n17242), .B2(n17258), .ZN(
        P3_U2698) );
  NOR2_X1 U20428 ( .A1(n17263), .A2(n17244), .ZN(n17245) );
  OAI21_X1 U20429 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17245), .A(n17258), .ZN(
        n17247) );
  INV_X1 U20430 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17246) );
  OAI22_X1 U20431 ( .A1(n17248), .A2(n17247), .B1(n17246), .B2(n17258), .ZN(
        P3_U2699) );
  NAND2_X1 U20432 ( .A1(n17249), .A2(n17257), .ZN(n17253) );
  NAND3_X1 U20433 ( .A1(n17253), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17258), .ZN(
        n17250) );
  OAI221_X1 U20434 ( .B1(n17253), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17258), 
        .C2(n17251), .A(n17250), .ZN(P3_U2700) );
  OAI21_X1 U20435 ( .B1(n17263), .B2(n17252), .A(n20880), .ZN(n17255) );
  AND2_X1 U20436 ( .A1(n17258), .A2(n17253), .ZN(n17254) );
  AOI22_X1 U20437 ( .A1(n17255), .A2(n17254), .B1(
        P3_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n20780), .ZN(n17256) );
  INV_X1 U20438 ( .A(n17256), .ZN(P3_U2701) );
  INV_X1 U20439 ( .A(n17257), .ZN(n17265) );
  INV_X1 U20440 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17259) );
  OAI222_X1 U20441 ( .A1(n17262), .A2(n17265), .B1(n17261), .B2(n17260), .C1(
        n17259), .C2(n17258), .ZN(P3_U2702) );
  AOI22_X1 U20442 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20780), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17263), .ZN(n17264) );
  OAI21_X1 U20443 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17265), .A(n17264), .ZN(
        P3_U2703) );
  INV_X1 U20444 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17438) );
  INV_X1 U20445 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17442) );
  INV_X1 U20446 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17448) );
  INV_X1 U20447 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17544) );
  INV_X1 U20448 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17516) );
  INV_X1 U20449 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17480) );
  INV_X1 U20450 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17482) );
  INV_X1 U20451 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17484) );
  INV_X1 U20452 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17486) );
  NOR4_X1 U20453 ( .A1(n17480), .A2(n17482), .A3(n17484), .A4(n17486), .ZN(
        n17267) );
  NAND4_X1 U20454 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17268)
         );
  NAND4_X1 U20455 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17269), .ZN(n17375) );
  AND4_X1 U20456 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n17312)
         );
  NAND2_X1 U20457 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17312), .ZN(n17313) );
  INV_X1 U20458 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17513) );
  OR2_X1 U20459 ( .A1(n17277), .A2(n17513), .ZN(n17271) );
  NAND2_X1 U20460 ( .A1(n18269), .A2(n20913), .ZN(n17349) );
  OAI21_X1 U20461 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17271), .A(n17270), .ZN(
        P3_U2704) );
  NAND2_X1 U20462 ( .A1(n17272), .A2(n20913), .ZN(n17318) );
  OAI22_X1 U20463 ( .A1(n17273), .A2(n17431), .B1(n18270), .B2(n17349), .ZN(
        n17274) );
  AOI21_X1 U20464 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17365), .A(n17274), .ZN(
        n17275) );
  OAI221_X1 U20465 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17277), .C1(n17513), 
        .C2(n17276), .A(n17275), .ZN(P3_U2705) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17364), .ZN(n17279) );
  OAI211_X1 U20467 ( .C1(n17282), .C2(P3_EAX_REG_29__SCAN_IN), .A(n9582), .B(
        n17277), .ZN(n17278) );
  OAI211_X1 U20468 ( .C1(n17280), .C2(n17431), .A(n17279), .B(n17278), .ZN(
        P3_U2706) );
  AOI22_X1 U20469 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17364), .B1(n17397), .B2(
        n17281), .ZN(n17285) );
  AOI211_X1 U20470 ( .C1(n17438), .C2(n17286), .A(n17282), .B(n20913), .ZN(
        n17283) );
  INV_X1 U20471 ( .A(n17283), .ZN(n17284) );
  OAI211_X1 U20472 ( .C1(n17318), .C2(n17532), .A(n17285), .B(n17284), .ZN(
        P3_U2707) );
  AOI22_X1 U20473 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17364), .ZN(n17289) );
  OAI211_X1 U20474 ( .C1(n17287), .C2(P3_EAX_REG_27__SCAN_IN), .A(n9582), .B(
        n17286), .ZN(n17288) );
  OAI211_X1 U20475 ( .C1(n17290), .C2(n17431), .A(n17289), .B(n17288), .ZN(
        P3_U2708) );
  AOI22_X1 U20476 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17364), .B1(n17397), .B2(
        n17291), .ZN(n17294) );
  OAI211_X1 U20477 ( .C1(n17296), .C2(P3_EAX_REG_26__SCAN_IN), .A(n9582), .B(
        n17292), .ZN(n17293) );
  OAI211_X1 U20478 ( .C1(n17318), .C2(n17528), .A(n17294), .B(n17293), .ZN(
        P3_U2709) );
  AOI22_X1 U20479 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17364), .ZN(n17299) );
  AOI211_X1 U20480 ( .C1(n17442), .C2(n17302), .A(n17296), .B(n20913), .ZN(
        n17297) );
  INV_X1 U20481 ( .A(n17297), .ZN(n17298) );
  OAI211_X1 U20482 ( .C1(n17300), .C2(n17431), .A(n17299), .B(n17298), .ZN(
        P3_U2710) );
  AOI22_X1 U20483 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17364), .B1(n17397), .B2(
        n17301), .ZN(n17305) );
  OAI211_X1 U20484 ( .C1(n17303), .C2(P3_EAX_REG_24__SCAN_IN), .A(n9582), .B(
        n17302), .ZN(n17304) );
  OAI211_X1 U20485 ( .C1(n17318), .C2(n17524), .A(n17305), .B(n17304), .ZN(
        P3_U2711) );
  AOI22_X1 U20486 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17364), .ZN(n17309) );
  OAI211_X1 U20487 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17307), .A(n9582), .B(
        n17306), .ZN(n17308) );
  OAI211_X1 U20488 ( .C1(n17310), .C2(n17431), .A(n17309), .B(n17308), .ZN(
        P3_U2712) );
  AOI22_X1 U20489 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17364), .B1(n17397), .B2(
        n17311), .ZN(n17317) );
  NOR2_X1 U20490 ( .A1(n18274), .A2(n17366), .ZN(n17360) );
  NAND2_X1 U20491 ( .A1(n17312), .A2(n17360), .ZN(n17324) );
  NAND2_X1 U20492 ( .A1(n9582), .A2(n17324), .ZN(n17327) );
  OAI21_X1 U20493 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17401), .A(n17327), .ZN(
        n17315) );
  NOR2_X1 U20494 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17313), .ZN(n17314) );
  AOI22_X1 U20495 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17315), .B1(n17360), 
        .B2(n17314), .ZN(n17316) );
  OAI211_X1 U20496 ( .C1(n18271), .C2(n17318), .A(n17317), .B(n17316), .ZN(
        P3_U2713) );
  INV_X1 U20497 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17450) );
  OAI22_X1 U20498 ( .A1(n17319), .A2(n17431), .B1(n18265), .B2(n17349), .ZN(
        n17320) );
  AOI21_X1 U20499 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17365), .A(n17320), .ZN(
        n17321) );
  OAI221_X1 U20500 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17324), .C1(n17450), 
        .C2(n17327), .A(n17321), .ZN(P3_U2714) );
  INV_X1 U20501 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17364), .B1(n17397), .B2(
        n17322), .ZN(n17326) );
  NAND2_X1 U20503 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17323) );
  NAND2_X1 U20504 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17360), .ZN(n17359) );
  NOR2_X1 U20505 ( .A1(n17323), .A2(n17359), .ZN(n17351) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17365), .B1(n17351), .B2(
        n17324), .ZN(n17325) );
  OAI211_X1 U20507 ( .C1(n17452), .C2(n17327), .A(n17326), .B(n17325), .ZN(
        P3_U2715) );
  AOI22_X1 U20508 ( .A1(n17329), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17328), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20509 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17330), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20510 ( .A1(n17332), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20511 ( .A1(n17334), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17333), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17335) );
  NAND4_X1 U20512 ( .A1(n17338), .A2(n17337), .A3(n17336), .A4(n17335), .ZN(
        n17348) );
  AOI22_X1 U20513 ( .A1(n17218), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20514 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U20515 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U20516 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17343) );
  NAND4_X1 U20517 ( .A1(n17346), .A2(n17345), .A3(n17344), .A4(n17343), .ZN(
        n17347) );
  NOR2_X1 U20518 ( .A1(n17348), .A2(n17347), .ZN(n20774) );
  INV_X1 U20519 ( .A(n17359), .ZN(n17355) );
  AOI22_X1 U20520 ( .A1(n17355), .A2(P3_EAX_REG_18__SCAN_IN), .B1(
        P3_EAX_REG_19__SCAN_IN), .B2(n9582), .ZN(n17350) );
  OAI22_X1 U20521 ( .A1(n17351), .A2(n17350), .B1(n18256), .B2(n17349), .ZN(
        n17352) );
  AOI21_X1 U20522 ( .B1(BUF2_REG_3__SCAN_IN), .B2(n17365), .A(n17352), .ZN(
        n17353) );
  OAI21_X1 U20523 ( .B1(n20774), .B2(n17431), .A(n17353), .ZN(P3_U2716) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17364), .ZN(n17357) );
  NAND2_X1 U20525 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17355), .ZN(n17354) );
  OAI211_X1 U20526 ( .C1(n17355), .C2(P3_EAX_REG_18__SCAN_IN), .A(n9582), .B(
        n17354), .ZN(n17356) );
  OAI211_X1 U20527 ( .C1(n17358), .C2(n17431), .A(n17357), .B(n17356), .ZN(
        P3_U2717) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17364), .ZN(n17362) );
  OAI211_X1 U20529 ( .C1(n17360), .C2(P3_EAX_REG_17__SCAN_IN), .A(n9582), .B(
        n17359), .ZN(n17361) );
  OAI211_X1 U20530 ( .C1(n17363), .C2(n17431), .A(n17362), .B(n17361), .ZN(
        P3_U2718) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17365), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17364), .ZN(n17368) );
  OAI211_X1 U20532 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17370), .A(n9582), .B(
        n17366), .ZN(n17367) );
  OAI211_X1 U20533 ( .C1(n17369), .C2(n17431), .A(n17368), .B(n17367), .ZN(
        P3_U2719) );
  AOI21_X1 U20534 ( .B1(n17544), .B2(n17375), .A(n17370), .ZN(n17371) );
  AOI22_X1 U20535 ( .A1(n17429), .A2(BUF2_REG_15__SCAN_IN), .B1(n17371), .B2(
        n9582), .ZN(n17372) );
  OAI21_X1 U20536 ( .B1(n17373), .B2(n17431), .A(n17372), .ZN(P3_U2720) );
  INV_X1 U20537 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17530) );
  NOR2_X1 U20538 ( .A1(n18274), .A2(n17398), .ZN(n17404) );
  NAND3_X1 U20539 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17404), .ZN(n17391) );
  INV_X1 U20540 ( .A(n17391), .ZN(n17395) );
  NAND2_X1 U20541 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17395), .ZN(n17388) );
  NOR2_X1 U20542 ( .A1(n17530), .A2(n17388), .ZN(n17382) );
  AND2_X1 U20543 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17382), .ZN(n17385) );
  NAND2_X1 U20544 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17385), .ZN(n17378) );
  AOI22_X1 U20545 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17429), .B1(n17397), .B2(
        n17374), .ZN(n17377) );
  NAND3_X1 U20546 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n9582), .A3(n17375), .ZN(
        n17376) );
  OAI211_X1 U20547 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17378), .A(n17377), .B(
        n17376), .ZN(P3_U2721) );
  INV_X1 U20548 ( .A(n17378), .ZN(n17381) );
  AOI21_X1 U20549 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n9582), .A(n17385), .ZN(
        n17380) );
  OAI222_X1 U20550 ( .A1(n17425), .A2(n17537), .B1(n17381), .B2(n17380), .C1(
        n17431), .C2(n17379), .ZN(P3_U2722) );
  AOI21_X1 U20551 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n9582), .A(n17382), .ZN(
        n17384) );
  OAI222_X1 U20552 ( .A1(n17425), .A2(n17532), .B1(n17385), .B2(n17384), .C1(
        n17431), .C2(n17383), .ZN(P3_U2723) );
  NAND2_X1 U20553 ( .A1(n9582), .A2(n17388), .ZN(n17392) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17429), .B1(n17397), .B2(
        n17386), .ZN(n17387) );
  OAI221_X1 U20555 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17388), .C1(n17530), 
        .C2(n17392), .A(n17387), .ZN(P3_U2724) );
  INV_X1 U20556 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20557 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17429), .B1(n17397), .B2(
        n17389), .ZN(n17390) );
  OAI221_X1 U20558 ( .B1(n17392), .B2(n17470), .C1(n17392), .C2(n17391), .A(
        n17390), .ZN(P3_U2725) );
  AOI22_X1 U20559 ( .A1(n17404), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n9582), .ZN(n17394) );
  OAI222_X1 U20560 ( .A1(n17425), .A2(n17526), .B1(n17395), .B2(n17394), .C1(
        n17431), .C2(n17393), .ZN(P3_U2726) );
  INV_X1 U20561 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20562 ( .A1(n17397), .A2(n17396), .B1(n17404), .B2(n17474), .ZN(
        n17400) );
  NAND3_X1 U20563 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n9582), .A3(n17398), .ZN(
        n17399) );
  OAI211_X1 U20564 ( .C1(n17425), .C2(n17524), .A(n17400), .B(n17399), .ZN(
        P3_U2727) );
  INV_X1 U20565 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17478) );
  NOR3_X1 U20566 ( .A1(n17516), .A2(n17491), .A3(n17401), .ZN(n17420) );
  AND2_X1 U20567 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17420), .ZN(n17424) );
  NAND2_X1 U20568 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17424), .ZN(n17412) );
  NOR2_X1 U20569 ( .A1(n17482), .A2(n17412), .ZN(n17415) );
  NAND2_X1 U20570 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17415), .ZN(n17405) );
  NOR2_X1 U20571 ( .A1(n17478), .A2(n17405), .ZN(n17408) );
  AOI21_X1 U20572 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n9582), .A(n17408), .ZN(
        n17403) );
  OAI222_X1 U20573 ( .A1(n17425), .A2(n18276), .B1(n17404), .B2(n17403), .C1(
        n17431), .C2(n17402), .ZN(P3_U2728) );
  INV_X1 U20574 ( .A(n17405), .ZN(n17411) );
  AOI21_X1 U20575 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n9582), .A(n17411), .ZN(
        n17407) );
  OAI222_X1 U20576 ( .A1(n18271), .A2(n17425), .B1(n17408), .B2(n17407), .C1(
        n17431), .C2(n17406), .ZN(P3_U2729) );
  AOI21_X1 U20577 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n9582), .A(n17415), .ZN(
        n17410) );
  OAI222_X1 U20578 ( .A1(n18266), .A2(n17425), .B1(n17411), .B2(n17410), .C1(
        n17431), .C2(n17409), .ZN(P3_U2730) );
  INV_X1 U20579 ( .A(n17412), .ZN(n17419) );
  AOI21_X1 U20580 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n9582), .A(n17419), .ZN(
        n17414) );
  OAI222_X1 U20581 ( .A1(n18261), .A2(n17425), .B1(n17415), .B2(n17414), .C1(
        n17431), .C2(n17413), .ZN(P3_U2731) );
  AOI21_X1 U20582 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n9582), .A(n17424), .ZN(
        n17418) );
  OAI222_X1 U20583 ( .A1(n18257), .A2(n17425), .B1(n17419), .B2(n17418), .C1(
        n17431), .C2(n17417), .ZN(P3_U2732) );
  AOI21_X1 U20584 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n9582), .A(n17420), .ZN(
        n17423) );
  INV_X1 U20585 ( .A(n17421), .ZN(n17422) );
  OAI222_X1 U20586 ( .A1(n18252), .A2(n17425), .B1(n17424), .B2(n17423), .C1(
        n17431), .C2(n17422), .ZN(P3_U2733) );
  AOI21_X1 U20587 ( .B1(n17516), .B2(n17427), .A(n17426), .ZN(n17428) );
  AOI22_X1 U20588 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17429), .B1(n17428), .B2(
        n9582), .ZN(n17430) );
  OAI21_X1 U20589 ( .B1(n17432), .B2(n17431), .A(n17430), .ZN(P3_U2734) );
  NOR2_X1 U20590 ( .A1(n17490), .A2(n17433), .ZN(n17453) );
  AOI22_X1 U20591 ( .A1(n9600), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20592 ( .B1(n17513), .B2(n17460), .A(n17434), .ZN(P3_U2737) );
  INV_X1 U20593 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20594 ( .A1(n9600), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(
        P3_DATAO_REG_29__SCAN_IN), .B2(n17488), .ZN(n17435) );
  OAI21_X1 U20595 ( .B1(n17436), .B2(n17460), .A(n17435), .ZN(P3_U2738) );
  AOI22_X1 U20596 ( .A1(n9600), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20597 ( .B1(n17438), .B2(n17460), .A(n17437), .ZN(P3_U2739) );
  INV_X1 U20598 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20599 ( .A1(n9600), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20600 ( .B1(n17509), .B2(n17460), .A(n17439), .ZN(P3_U2740) );
  AOI22_X1 U20601 ( .A1(n9600), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20602 ( .B1(n9713), .B2(n17460), .A(n17440), .ZN(P3_U2741) );
  AOI22_X1 U20603 ( .A1(n9600), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20604 ( .B1(n17442), .B2(n17460), .A(n17441), .ZN(P3_U2742) );
  INV_X1 U20605 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20606 ( .A1(n9600), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20607 ( .B1(n17444), .B2(n17460), .A(n17443), .ZN(P3_U2743) );
  INV_X1 U20608 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U20609 ( .A1(n9600), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20610 ( .B1(n17446), .B2(n17460), .A(n17445), .ZN(P3_U2744) );
  AOI22_X1 U20611 ( .A1(n9600), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20612 ( .B1(n17448), .B2(n17460), .A(n17447), .ZN(P3_U2745) );
  AOI22_X1 U20613 ( .A1(n9600), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20614 ( .B1(n17450), .B2(n17460), .A(n17449), .ZN(P3_U2746) );
  AOI22_X1 U20615 ( .A1(n9600), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20616 ( .B1(n17452), .B2(n17460), .A(n17451), .ZN(P3_U2747) );
  INV_X1 U20617 ( .A(P3_UWORD_REG_3__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U20618 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17453), .B1(n17488), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U20619 ( .B1(n17457), .B2(n20882), .A(n17454), .ZN(P3_U2748) );
  INV_X1 U20620 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20621 ( .A1(n9600), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20622 ( .B1(n17456), .B2(n17460), .A(n17455), .ZN(P3_U2749) );
  INV_X1 U20623 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20624 ( .A1(n9600), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20625 ( .B1(n17497), .B2(n17460), .A(n17458), .ZN(P3_U2750) );
  INV_X1 U20626 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U20627 ( .A1(n9600), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20628 ( .B1(n17461), .B2(n17460), .A(n17459), .ZN(P3_U2751) );
  AOI22_X1 U20629 ( .A1(n9600), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20630 ( .B1(n17544), .B2(n17490), .A(n17462), .ZN(P3_U2752) );
  INV_X1 U20631 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U20632 ( .A1(n9600), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20633 ( .B1(n17539), .B2(n17490), .A(n17463), .ZN(P3_U2753) );
  INV_X1 U20634 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U20635 ( .A1(n9600), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20636 ( .B1(n17465), .B2(n17490), .A(n17464), .ZN(P3_U2754) );
  INV_X1 U20637 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U20638 ( .A1(n9600), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20639 ( .B1(n17467), .B2(n17490), .A(n17466), .ZN(P3_U2755) );
  AOI22_X1 U20640 ( .A1(n9600), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20641 ( .B1(n17530), .B2(n17490), .A(n17468), .ZN(P3_U2756) );
  AOI22_X1 U20642 ( .A1(n9600), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20643 ( .B1(n17470), .B2(n17490), .A(n17469), .ZN(P3_U2757) );
  INV_X1 U20644 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20645 ( .A1(n9600), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20646 ( .B1(n17472), .B2(n17490), .A(n17471), .ZN(P3_U2758) );
  AOI22_X1 U20647 ( .A1(n9600), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17473) );
  OAI21_X1 U20648 ( .B1(n17474), .B2(n17490), .A(n17473), .ZN(P3_U2759) );
  INV_X1 U20649 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20650 ( .A1(n9600), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17475) );
  OAI21_X1 U20651 ( .B1(n17476), .B2(n17490), .A(n17475), .ZN(P3_U2760) );
  AOI22_X1 U20652 ( .A1(n9600), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17477) );
  OAI21_X1 U20653 ( .B1(n17478), .B2(n17490), .A(n17477), .ZN(P3_U2761) );
  AOI22_X1 U20654 ( .A1(n9600), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17479) );
  OAI21_X1 U20655 ( .B1(n17480), .B2(n17490), .A(n17479), .ZN(P3_U2762) );
  AOI22_X1 U20656 ( .A1(n9600), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20657 ( .B1(n17482), .B2(n17490), .A(n17481), .ZN(P3_U2763) );
  AOI22_X1 U20658 ( .A1(n9600), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20659 ( .B1(n17484), .B2(n17490), .A(n17483), .ZN(P3_U2764) );
  AOI22_X1 U20660 ( .A1(n9600), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17485) );
  OAI21_X1 U20661 ( .B1(n17486), .B2(n17490), .A(n17485), .ZN(P3_U2765) );
  AOI22_X1 U20662 ( .A1(n9600), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20663 ( .B1(n17516), .B2(n17490), .A(n17487), .ZN(P3_U2766) );
  AOI22_X1 U20664 ( .A1(n9600), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17488), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17489) );
  OAI21_X1 U20665 ( .B1(n17491), .B2(n17490), .A(n17489), .ZN(P3_U2767) );
  OAI211_X1 U20666 ( .C1(n18878), .C2(n18877), .A(n18718), .B(n17492), .ZN(
        n17540) );
  AOI22_X1 U20667 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17533), .ZN(n17495) );
  OAI21_X1 U20668 ( .B1(n18241), .B2(n17536), .A(n17495), .ZN(P3_U2768) );
  AOI22_X1 U20669 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17541), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17533), .ZN(n17496) );
  OAI21_X1 U20670 ( .B1(n17497), .B2(n17543), .A(n17496), .ZN(P3_U2769) );
  AOI22_X1 U20671 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17533), .ZN(n17498) );
  OAI21_X1 U20672 ( .B1(n18252), .B2(n17536), .A(n17498), .ZN(P3_U2770) );
  AOI22_X1 U20673 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17533), .ZN(n17499) );
  OAI21_X1 U20674 ( .B1(n18257), .B2(n17536), .A(n17499), .ZN(P3_U2771) );
  AOI22_X1 U20675 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17533), .ZN(n17500) );
  OAI21_X1 U20676 ( .B1(n18261), .B2(n17536), .A(n17500), .ZN(P3_U2772) );
  AOI22_X1 U20677 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17533), .ZN(n17501) );
  OAI21_X1 U20678 ( .B1(n18266), .B2(n17536), .A(n17501), .ZN(P3_U2773) );
  AOI22_X1 U20679 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17533), .ZN(n17502) );
  OAI21_X1 U20680 ( .B1(n18271), .B2(n17536), .A(n17502), .ZN(P3_U2774) );
  AOI22_X1 U20681 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17503), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17533), .ZN(n17504) );
  OAI21_X1 U20682 ( .B1(n18276), .B2(n17536), .A(n17504), .ZN(P3_U2775) );
  AOI22_X1 U20683 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17533), .ZN(n17505) );
  OAI21_X1 U20684 ( .B1(n17524), .B2(n17536), .A(n17505), .ZN(P3_U2776) );
  AOI22_X1 U20685 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17533), .ZN(n17506) );
  OAI21_X1 U20686 ( .B1(n17526), .B2(n17536), .A(n17506), .ZN(P3_U2777) );
  AOI22_X1 U20687 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17533), .ZN(n17507) );
  OAI21_X1 U20688 ( .B1(n17528), .B2(n17536), .A(n17507), .ZN(P3_U2778) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17541), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17533), .ZN(n17508) );
  OAI21_X1 U20690 ( .B1(n17509), .B2(n17543), .A(n17508), .ZN(P3_U2779) );
  AOI22_X1 U20691 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17533), .ZN(n17510) );
  OAI21_X1 U20692 ( .B1(n17532), .B2(n17536), .A(n17510), .ZN(P3_U2780) );
  AOI22_X1 U20693 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17534), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17533), .ZN(n17511) );
  OAI21_X1 U20694 ( .B1(n17537), .B2(n17536), .A(n17511), .ZN(P3_U2781) );
  AOI22_X1 U20695 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17541), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17533), .ZN(n17512) );
  OAI21_X1 U20696 ( .B1(n17513), .B2(n17543), .A(n17512), .ZN(P3_U2782) );
  AOI22_X1 U20697 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17533), .ZN(n17514) );
  OAI21_X1 U20698 ( .B1(n18241), .B2(n17536), .A(n17514), .ZN(P3_U2783) );
  AOI22_X1 U20699 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17541), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17533), .ZN(n17515) );
  OAI21_X1 U20700 ( .B1(n17516), .B2(n17543), .A(n17515), .ZN(P3_U2784) );
  AOI22_X1 U20701 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17533), .ZN(n17517) );
  OAI21_X1 U20702 ( .B1(n18252), .B2(n17536), .A(n17517), .ZN(P3_U2785) );
  AOI22_X1 U20703 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17540), .ZN(n17518) );
  OAI21_X1 U20704 ( .B1(n18257), .B2(n17536), .A(n17518), .ZN(P3_U2786) );
  AOI22_X1 U20705 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17540), .ZN(n17519) );
  OAI21_X1 U20706 ( .B1(n18261), .B2(n17536), .A(n17519), .ZN(P3_U2787) );
  AOI22_X1 U20707 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17540), .ZN(n17520) );
  OAI21_X1 U20708 ( .B1(n18266), .B2(n17536), .A(n17520), .ZN(P3_U2788) );
  AOI22_X1 U20709 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17540), .ZN(n17521) );
  OAI21_X1 U20710 ( .B1(n18271), .B2(n17536), .A(n17521), .ZN(P3_U2789) );
  AOI22_X1 U20711 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17540), .ZN(n17522) );
  OAI21_X1 U20712 ( .B1(n18276), .B2(n17536), .A(n17522), .ZN(P3_U2790) );
  AOI22_X1 U20713 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17540), .ZN(n17523) );
  OAI21_X1 U20714 ( .B1(n17524), .B2(n17536), .A(n17523), .ZN(P3_U2791) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17540), .ZN(n17525) );
  OAI21_X1 U20716 ( .B1(n17526), .B2(n17536), .A(n17525), .ZN(P3_U2792) );
  AOI22_X1 U20717 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17533), .ZN(n17527) );
  OAI21_X1 U20718 ( .B1(n17528), .B2(n17536), .A(n17527), .ZN(P3_U2793) );
  AOI22_X1 U20719 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17541), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17540), .ZN(n17529) );
  OAI21_X1 U20720 ( .B1(n17530), .B2(n17543), .A(n17529), .ZN(P3_U2794) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17533), .ZN(n17531) );
  OAI21_X1 U20722 ( .B1(n17532), .B2(n17536), .A(n17531), .ZN(P3_U2795) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17534), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17533), .ZN(n17535) );
  OAI21_X1 U20724 ( .B1(n17537), .B2(n17536), .A(n17535), .ZN(P3_U2796) );
  AOI22_X1 U20725 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17541), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17540), .ZN(n17538) );
  OAI21_X1 U20726 ( .B1(n17539), .B2(n17543), .A(n17538), .ZN(P3_U2797) );
  AOI22_X1 U20727 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17541), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17540), .ZN(n17542) );
  OAI21_X1 U20728 ( .B1(n17544), .B2(n17543), .A(n17542), .ZN(P3_U2798) );
  NAND2_X1 U20729 ( .A1(n17547), .A2(n17694), .ZN(n17566) );
  AOI221_X1 U20730 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n17546), .C2(n17545), .A(
        n17566), .ZN(n17553) );
  OAI22_X1 U20731 ( .A1(n17548), .A2(n18739), .B1(n17547), .B2(n17858), .ZN(
        n17549) );
  NOR2_X1 U20732 ( .A1(n17888), .A2(n17549), .ZN(n17571) );
  OAI21_X1 U20733 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17678), .A(
        n17571), .ZN(n17561) );
  AOI22_X1 U20734 ( .A1(n18209), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17561), .ZN(n17550) );
  OAI21_X1 U20735 ( .B1(n17741), .B2(n17551), .A(n17550), .ZN(n17552) );
  AOI211_X1 U20736 ( .C1(n17600), .C2(n17554), .A(n17553), .B(n17552), .ZN(
        n17560) );
  NAND2_X1 U20737 ( .A1(n17905), .A2(n17745), .ZN(n17624) );
  INV_X1 U20738 ( .A(n17745), .ZN(n17813) );
  AOI22_X1 U20739 ( .A1(n17893), .A2(n17909), .B1(n17813), .B2(n17908), .ZN(
        n17578) );
  NAND2_X1 U20740 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17578), .ZN(
        n17568) );
  NAND3_X1 U20741 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17624), .A3(
        n17568), .ZN(n17559) );
  OAI211_X1 U20742 ( .C1(n17557), .C2(n17556), .A(n17812), .B(n17555), .ZN(
        n17558) );
  NAND3_X1 U20743 ( .A1(n17560), .A2(n17559), .A3(n17558), .ZN(P3_U2802) );
  AOI22_X1 U20744 ( .A1(n17754), .A2(n17562), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17561), .ZN(n17569) );
  NOR2_X1 U20745 ( .A1(n17564), .A2(n17563), .ZN(n17565) );
  INV_X1 U20746 ( .A(n17704), .ZN(n17685) );
  NAND2_X1 U20747 ( .A1(n17955), .A2(n17907), .ZN(n17928) );
  NOR2_X1 U20748 ( .A1(n17930), .A2(n17928), .ZN(n17920) );
  NAND2_X1 U20749 ( .A1(n17685), .A2(n17920), .ZN(n17579) );
  OAI21_X1 U20750 ( .B1(n9670), .B2(n20800), .A(n17570), .ZN(n17921) );
  AOI221_X1 U20751 ( .B1(n18278), .B2(n17573), .C1(n17572), .C2(n17573), .A(
        n17571), .ZN(n17576) );
  NAND2_X1 U20752 ( .A1(n18209), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17922) );
  OAI221_X1 U20753 ( .B1(n17574), .B2(n17741), .C1(n17574), .C2(n17678), .A(
        n17922), .ZN(n17575) );
  AOI211_X1 U20754 ( .C1(n17812), .C2(n17921), .A(n17576), .B(n17575), .ZN(
        n17577) );
  OAI221_X1 U20755 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17579), 
        .C1(n20800), .C2(n17578), .A(n17577), .ZN(P3_U2804) );
  XNOR2_X1 U20756 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17580), .ZN(
        n17939) );
  OAI22_X1 U20757 ( .A1(n17583), .A2(n18278), .B1(n17581), .B2(n18739), .ZN(
        n17582) );
  NOR2_X1 U20758 ( .A1(n17888), .A2(n17582), .ZN(n17608) );
  OAI21_X1 U20759 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17678), .A(
        n17608), .ZN(n17597) );
  NOR2_X1 U20760 ( .A1(n18175), .A2(n18802), .ZN(n17934) );
  NAND2_X1 U20761 ( .A1(n17583), .A2(n17694), .ZN(n17595) );
  OAI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17584), .ZN(n17585) );
  OAI22_X1 U20763 ( .A1(n17741), .A2(n17586), .B1(n17595), .B2(n17585), .ZN(
        n17587) );
  AOI211_X1 U20764 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17597), .A(
        n17934), .B(n17587), .ZN(n17593) );
  XNOR2_X1 U20765 ( .A(n17588), .B(n17930), .ZN(n17936) );
  OAI21_X1 U20766 ( .B1(n17811), .B2(n17590), .A(n17589), .ZN(n17591) );
  XNOR2_X1 U20767 ( .A(n17591), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17935) );
  AOI22_X1 U20768 ( .A1(n17893), .A2(n17936), .B1(n17812), .B2(n17935), .ZN(
        n17592) );
  OAI211_X1 U20769 ( .C1(n17745), .C2(n17939), .A(n17593), .B(n17592), .ZN(
        P3_U2805) );
  AOI22_X1 U20770 ( .A1(n17893), .A2(n17941), .B1(n17813), .B2(n17940), .ZN(
        n17615) );
  NOR2_X1 U20771 ( .A1(n18175), .A2(n18800), .ZN(n17950) );
  OAI22_X1 U20772 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17595), .B1(
        n17741), .B2(n17594), .ZN(n17596) );
  AOI211_X1 U20773 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17597), .A(
        n17950), .B(n17596), .ZN(n17602) );
  OAI21_X1 U20774 ( .B1(n17599), .B2(n17603), .A(n17598), .ZN(n17949) );
  NOR2_X1 U20775 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17958), .ZN(
        n17947) );
  AOI22_X1 U20776 ( .A1(n17812), .A2(n17949), .B1(n17600), .B2(n17947), .ZN(
        n17601) );
  OAI211_X1 U20777 ( .C1(n17615), .C2(n17603), .A(n17602), .B(n17601), .ZN(
        P3_U2806) );
  OAI22_X1 U20778 ( .A1(n17811), .A2(n17973), .B1(n17604), .B2(n17627), .ZN(
        n17606) );
  NOR2_X1 U20779 ( .A1(n17606), .A2(n17605), .ZN(n17607) );
  XNOR2_X1 U20780 ( .A(n17607), .B(n17958), .ZN(n17960) );
  AOI221_X1 U20781 ( .B1(n17610), .B2(n17609), .C1(n18278), .C2(n17609), .A(
        n17608), .ZN(n17613) );
  NAND2_X1 U20782 ( .A1(n18209), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17962) );
  OAI221_X1 U20783 ( .B1(n17611), .B2(n17741), .C1(n17611), .C2(n17678), .A(
        n17962), .ZN(n17612) );
  AOI211_X1 U20784 ( .C1(n17960), .C2(n17812), .A(n17613), .B(n17612), .ZN(
        n17614) );
  OAI221_X1 U20785 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17616), 
        .C1(n17958), .C2(n17615), .A(n17614), .ZN(P3_U2807) );
  NAND2_X1 U20786 ( .A1(n17970), .A2(n17973), .ZN(n17979) );
  OAI22_X1 U20787 ( .A1(n17619), .A2(n17858), .B1(n17617), .B2(n18739), .ZN(
        n17618) );
  NOR2_X1 U20788 ( .A1(n17888), .A2(n17618), .ZN(n17642) );
  OAI21_X1 U20789 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17678), .A(
        n17642), .ZN(n17635) );
  NOR2_X1 U20790 ( .A1(n18175), .A2(n18796), .ZN(n17976) );
  NAND2_X1 U20791 ( .A1(n17619), .A2(n17694), .ZN(n17633) );
  OAI21_X1 U20792 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17620), .ZN(n17621) );
  OAI22_X1 U20793 ( .A1(n17741), .A2(n17622), .B1(n17633), .B2(n17621), .ZN(
        n17623) );
  AOI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17635), .A(
        n17976), .B(n17623), .ZN(n17630) );
  INV_X1 U20795 ( .A(n17624), .ZN(n17647) );
  NOR2_X1 U20796 ( .A1(n18045), .A2(n17745), .ZN(n17715) );
  NOR2_X1 U20797 ( .A1(n18044), .A2(n17905), .ZN(n17714) );
  OAI21_X1 U20798 ( .B1(n17970), .B2(n17647), .A(n17702), .ZN(n17639) );
  INV_X1 U20799 ( .A(n17689), .ZN(n17626) );
  INV_X1 U20800 ( .A(n17605), .ZN(n17625) );
  OAI221_X1 U20801 ( .B1(n17627), .B2(n17970), .C1(n17627), .C2(n17626), .A(
        n17625), .ZN(n17628) );
  XNOR2_X1 U20802 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17628), .ZN(
        n17977) );
  AOI22_X1 U20803 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17639), .B1(
        n17812), .B2(n17977), .ZN(n17629) );
  OAI211_X1 U20804 ( .C1(n17704), .C2(n17979), .A(n17630), .B(n17629), .ZN(
        P3_U2808) );
  NAND2_X1 U20805 ( .A1(n17963), .A2(n17986), .ZN(n17992) );
  NOR2_X1 U20806 ( .A1(n17631), .A2(n17671), .ZN(n17981) );
  NAND2_X1 U20807 ( .A1(n17685), .A2(n17981), .ZN(n17664) );
  NOR2_X1 U20808 ( .A1(n18175), .A2(n18795), .ZN(n17989) );
  OAI22_X1 U20809 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17633), .B1(
        n17741), .B2(n17632), .ZN(n17634) );
  AOI211_X1 U20810 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17635), .A(
        n17989), .B(n17634), .ZN(n17641) );
  NAND3_X1 U20811 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17811), .A3(
        n17636), .ZN(n17658) );
  INV_X1 U20812 ( .A(n17672), .ZN(n17659) );
  OAI22_X1 U20813 ( .A1(n17985), .A2(n17658), .B1(n17659), .B2(n17637), .ZN(
        n17638) );
  XOR2_X1 U20814 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17638), .Z(
        n17990) );
  AOI22_X1 U20815 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17639), .B1(
        n17812), .B2(n17990), .ZN(n17640) );
  OAI211_X1 U20816 ( .C1(n17992), .C2(n17664), .A(n17641), .B(n17640), .ZN(
        P3_U2809) );
  NAND2_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17968), .ZN(
        n18001) );
  AOI221_X1 U20818 ( .B1(n17643), .B2(n20809), .C1(n18278), .C2(n20809), .A(
        n17642), .ZN(n17646) );
  AOI21_X1 U20819 ( .B1(n17741), .B2(n17678), .A(n17644), .ZN(n17645) );
  AOI211_X1 U20820 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18209), .A(n17646), 
        .B(n17645), .ZN(n17650) );
  INV_X1 U20821 ( .A(n17981), .ZN(n17965) );
  NOR2_X1 U20822 ( .A1(n18006), .A2(n17965), .ZN(n17993) );
  OAI21_X1 U20823 ( .B1(n17647), .B2(n17993), .A(n17702), .ZN(n17661) );
  AOI221_X1 U20824 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17658), 
        .C1(n18006), .C2(n17670), .A(n17605), .ZN(n17648) );
  XNOR2_X1 U20825 ( .A(n17648), .B(n17968), .ZN(n17997) );
  AOI22_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17661), .B1(
        n17812), .B2(n17997), .ZN(n17649) );
  OAI211_X1 U20827 ( .C1(n17664), .C2(n18001), .A(n17650), .B(n17649), .ZN(
        P3_U2810) );
  INV_X1 U20828 ( .A(n17665), .ZN(n17651) );
  OAI21_X1 U20829 ( .B1(n17888), .B2(n17651), .A(n17896), .ZN(n17679) );
  OAI21_X1 U20830 ( .B1(n17652), .B2(n18739), .A(n17679), .ZN(n17669) );
  NOR2_X1 U20831 ( .A1(n18175), .A2(n18791), .ZN(n18002) );
  INV_X1 U20832 ( .A(n17653), .ZN(n17656) );
  OAI211_X1 U20833 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17665), .B(n17694), .ZN(n17655) );
  OAI22_X1 U20834 ( .A1(n17656), .A2(n17655), .B1(n17741), .B2(n17654), .ZN(
        n17657) );
  AOI211_X1 U20835 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17669), .A(
        n18002), .B(n17657), .ZN(n17663) );
  OAI21_X1 U20836 ( .B1(n17659), .B2(n17670), .A(n17658), .ZN(n17660) );
  XNOR2_X1 U20837 ( .A(n17660), .B(n18006), .ZN(n18003) );
  AOI22_X1 U20838 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17661), .B1(
        n17812), .B2(n18003), .ZN(n17662) );
  OAI211_X1 U20839 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17664), .A(
        n17663), .B(n17662), .ZN(P3_U2811) );
  NAND2_X1 U20840 ( .A1(n18022), .A2(n17671), .ZN(n18026) );
  NOR2_X1 U20841 ( .A1(n18175), .A2(n18789), .ZN(n18014) );
  NAND2_X1 U20842 ( .A1(n17665), .A2(n17694), .ZN(n17667) );
  OAI22_X1 U20843 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17667), .B1(
        n17741), .B2(n17666), .ZN(n17668) );
  AOI211_X1 U20844 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17669), .A(
        n18014), .B(n17668), .ZN(n17675) );
  OAI21_X1 U20845 ( .B1(n18022), .B2(n17704), .A(n17702), .ZN(n17686) );
  OAI21_X1 U20846 ( .B1(n17671), .B2(n12810), .A(n17670), .ZN(n17673) );
  XNOR2_X1 U20847 ( .A(n17673), .B(n17672), .ZN(n18015) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17686), .B1(
        n17812), .B2(n18015), .ZN(n17674) );
  OAI211_X1 U20849 ( .C1(n17704), .C2(n18026), .A(n17675), .B(n17674), .ZN(
        P3_U2812) );
  AOI21_X1 U20850 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17677), .A(
        n17676), .ZN(n18032) );
  NOR2_X1 U20851 ( .A1(n18175), .A2(n20801), .ZN(n17683) );
  AOI221_X1 U20852 ( .B1(n17681), .B2(n17680), .C1(n18278), .C2(n17680), .A(
        n17679), .ZN(n17682) );
  AOI211_X1 U20853 ( .C1(n17684), .C2(n17895), .A(n17683), .B(n17682), .ZN(
        n17688) );
  NOR2_X1 U20854 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17703), .ZN(
        n18027) );
  AOI22_X1 U20855 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17686), .B1(
        n17685), .B2(n18027), .ZN(n17687) );
  OAI211_X1 U20856 ( .C1(n18032), .C2(n17778), .A(n17688), .B(n17687), .ZN(
        P3_U2813) );
  NOR2_X1 U20857 ( .A1(n12810), .A2(n18096), .ZN(n17793) );
  AOI22_X1 U20858 ( .A1(n17793), .A2(n18013), .B1(n17689), .B2(n12810), .ZN(
        n17690) );
  XNOR2_X1 U20859 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17690), .ZN(
        n18037) );
  INV_X1 U20860 ( .A(n17691), .ZN(n17692) );
  AOI21_X1 U20861 ( .B1(n17805), .B2(n17692), .A(n17888), .ZN(n17722) );
  OAI21_X1 U20862 ( .B1(n17693), .B2(n18739), .A(n17722), .ZN(n17711) );
  AOI22_X1 U20863 ( .A1(n18209), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17711), .ZN(n17698) );
  NAND2_X1 U20864 ( .A1(n17737), .A2(n17694), .ZN(n17751) );
  NOR2_X1 U20865 ( .A1(n17695), .A2(n17751), .ZN(n17713) );
  NAND2_X1 U20866 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17696) );
  OAI211_X1 U20867 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17713), .B(n17696), .ZN(n17697) );
  OAI211_X1 U20868 ( .C1(n17741), .C2(n17699), .A(n17698), .B(n17697), .ZN(
        n17700) );
  AOI21_X1 U20869 ( .B1(n17812), .B2(n18037), .A(n17700), .ZN(n17701) );
  OAI221_X1 U20870 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17704), 
        .C1(n17703), .C2(n17702), .A(n17701), .ZN(P3_U2814) );
  OAI21_X1 U20871 ( .B1(n17706), .B2(n17732), .A(n17705), .ZN(n17707) );
  OAI221_X1 U20872 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18060), 
        .C1(n12793), .C2(n17811), .A(n17707), .ZN(n17708) );
  XOR2_X1 U20873 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17708), .Z(
        n18053) );
  INV_X1 U20874 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17712) );
  NAND2_X1 U20875 ( .A1(n18209), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18056) );
  OAI21_X1 U20876 ( .B1(n17741), .B2(n17709), .A(n18056), .ZN(n17710) );
  AOI221_X1 U20877 ( .B1(n17713), .B2(n17712), .C1(n17711), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17710), .ZN(n17717) );
  NOR2_X1 U20878 ( .A1(n18086), .A2(n18096), .ZN(n18075) );
  AND2_X1 U20879 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18075), .ZN(
        n17726) );
  NAND2_X1 U20880 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17726), .ZN(
        n17725) );
  NAND2_X1 U20881 ( .A1(n18058), .A2(n17725), .ZN(n18046) );
  NAND2_X1 U20882 ( .A1(n17718), .A2(n18058), .ZN(n18048) );
  AOI22_X1 U20883 ( .A1(n17715), .A2(n18046), .B1(n17714), .B2(n18048), .ZN(
        n17716) );
  OAI211_X1 U20884 ( .C1(n17778), .C2(n18053), .A(n17717), .B(n17716), .ZN(
        P3_U2815) );
  OAI21_X1 U20885 ( .B1(n17719), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17718), .ZN(n18071) );
  NOR2_X1 U20886 ( .A1(n17720), .A2(n18278), .ZN(n17765) );
  AOI21_X1 U20887 ( .B1(n17736), .B2(n17765), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17721) );
  OAI22_X1 U20888 ( .A1(n17722), .A2(n17721), .B1(n18175), .B2(n18783), .ZN(
        n17728) );
  INV_X1 U20889 ( .A(n17793), .ZN(n17773) );
  NAND3_X1 U20890 ( .A1(n17758), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18042) );
  OAI21_X1 U20891 ( .B1(n17773), .B2(n18042), .A(n17723), .ZN(n17724) );
  XNOR2_X1 U20892 ( .A(n17724), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18067) );
  OAI21_X1 U20893 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17726), .A(
        n17725), .ZN(n18066) );
  OAI22_X1 U20894 ( .A1(n18067), .A2(n17778), .B1(n17745), .B2(n18066), .ZN(
        n17727) );
  AOI211_X1 U20895 ( .C1(n17729), .C2(n17895), .A(n17728), .B(n17727), .ZN(
        n17730) );
  OAI21_X1 U20896 ( .B1(n17905), .B2(n18071), .A(n17730), .ZN(P3_U2816) );
  OAI22_X1 U20897 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17811), .B1(
        n17732), .B2(n18086), .ZN(n17733) );
  OAI21_X1 U20898 ( .B1(n17811), .B2(n17731), .A(n17733), .ZN(n17735) );
  XNOR2_X1 U20899 ( .A(n17735), .B(n17734), .ZN(n18083) );
  AOI211_X1 U20900 ( .C1(n17750), .C2(n17742), .A(n17736), .B(n17751), .ZN(
        n17744) );
  OAI21_X1 U20901 ( .B1(n17737), .B2(n17858), .A(n18739), .ZN(n17738) );
  AOI21_X1 U20902 ( .B1(n17739), .B2(n17738), .A(n17888), .ZN(n17749) );
  OAI22_X1 U20903 ( .A1(n17749), .A2(n17742), .B1(n17741), .B2(n17740), .ZN(
        n17743) );
  AOI211_X1 U20904 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18209), .A(n17744), 
        .B(n17743), .ZN(n17748) );
  OAI22_X1 U20905 ( .A1(n17746), .A2(n17905), .B1(n18075), .B2(n17745), .ZN(
        n17757) );
  NOR2_X1 U20906 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18086), .ZN(
        n18072) );
  AOI22_X1 U20907 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17757), .B1(
        n18072), .B2(n17795), .ZN(n17747) );
  OAI211_X1 U20908 ( .C1(n17778), .C2(n18083), .A(n17748), .B(n17747), .ZN(
        P3_U2817) );
  NAND2_X1 U20909 ( .A1(n18209), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18093) );
  OAI221_X1 U20910 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17751), .C1(
        n17750), .C2(n17749), .A(n18093), .ZN(n17752) );
  AOI21_X1 U20911 ( .B1(n17754), .B2(n17753), .A(n17752), .ZN(n17761) );
  INV_X1 U20912 ( .A(n17758), .ZN(n18084) );
  OAI21_X1 U20913 ( .B1(n18084), .B2(n17773), .A(n17755), .ZN(n17756) );
  XNOR2_X1 U20914 ( .A(n17756), .B(n12793), .ZN(n18092) );
  AOI22_X1 U20915 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17757), .B1(
        n17812), .B2(n18092), .ZN(n17760) );
  NAND3_X1 U20916 ( .A1(n17758), .A2(n12793), .A3(n17795), .ZN(n17759) );
  NAND3_X1 U20917 ( .A1(n17761), .A2(n17760), .A3(n17759), .ZN(P3_U2818) );
  INV_X1 U20918 ( .A(n18107), .ZN(n17768) );
  AOI21_X1 U20919 ( .B1(n17793), .B2(n17768), .A(n17762), .ZN(n17763) );
  XNOR2_X1 U20920 ( .A(n17763), .B(n18108), .ZN(n18114) );
  AOI22_X1 U20921 ( .A1(n18607), .A2(n17775), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17896), .ZN(n17764) );
  NAND2_X1 U20922 ( .A1(n18209), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18112) );
  OAI21_X1 U20923 ( .B1(n17765), .B2(n17764), .A(n18112), .ZN(n17766) );
  AOI21_X1 U20924 ( .B1(n17767), .B2(n17895), .A(n17766), .ZN(n17770) );
  INV_X1 U20925 ( .A(n17795), .ZN(n17771) );
  AOI22_X1 U20926 ( .A1(n17893), .A2(n18098), .B1(n17813), .B2(n18096), .ZN(
        n17799) );
  OAI21_X1 U20927 ( .B1(n17768), .B2(n17771), .A(n17799), .ZN(n17781) );
  NOR2_X1 U20928 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18107), .ZN(
        n18111) );
  AOI22_X1 U20929 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17781), .B1(
        n18111), .B2(n17795), .ZN(n17769) );
  OAI211_X1 U20930 ( .C1(n18114), .C2(n17778), .A(n17770), .B(n17769), .ZN(
        P3_U2819) );
  INV_X1 U20931 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18118) );
  OAI21_X1 U20932 ( .B1(n17771), .B2(n18122), .A(n18118), .ZN(n17780) );
  OAI21_X1 U20933 ( .B1(n18122), .B2(n17773), .A(n17772), .ZN(n17774) );
  XNOR2_X1 U20934 ( .A(n17774), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18121) );
  AND2_X1 U20935 ( .A1(n17775), .A2(n18607), .ZN(n17777) );
  NAND4_X1 U20936 ( .A1(n17819), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17802), .A4(n18607), .ZN(n17788) );
  NOR2_X1 U20937 ( .A1(n17787), .A2(n17788), .ZN(n17785) );
  AOI21_X1 U20938 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17896), .A(
        n17785), .ZN(n17776) );
  OAI22_X1 U20939 ( .A1(n18121), .A2(n17778), .B1(n17777), .B2(n17776), .ZN(
        n17779) );
  AOI21_X1 U20940 ( .B1(n17781), .B2(n17780), .A(n17779), .ZN(n17783) );
  NAND2_X1 U20941 ( .A1(n18209), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17782) );
  OAI211_X1 U20942 ( .C1(n17885), .C2(n17784), .A(n17783), .B(n17782), .ZN(
        P3_U2820) );
  INV_X1 U20943 ( .A(n17896), .ZN(n17786) );
  AOI211_X1 U20944 ( .C1(n17788), .C2(n17787), .A(n17786), .B(n17785), .ZN(
        n17790) );
  NOR2_X1 U20945 ( .A1(n18175), .A2(n18772), .ZN(n17789) );
  AOI211_X1 U20946 ( .C1(n17791), .C2(n17895), .A(n17790), .B(n17789), .ZN(
        n17798) );
  NOR2_X1 U20947 ( .A1(n17793), .A2(n17792), .ZN(n17794) );
  XNOR2_X1 U20948 ( .A(n17794), .B(n18122), .ZN(n18128) );
  INV_X1 U20949 ( .A(n18128), .ZN(n17796) );
  AOI22_X1 U20950 ( .A1(n17812), .A2(n17796), .B1(n18122), .B2(n17795), .ZN(
        n17797) );
  OAI211_X1 U20951 ( .C1(n17799), .C2(n18122), .A(n17798), .B(n17797), .ZN(
        P3_U2821) );
  OAI21_X1 U20952 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17801), .A(
        n17800), .ZN(n18146) );
  AOI211_X1 U20953 ( .C1(n17806), .C2(n17803), .A(n17802), .B(n18278), .ZN(
        n17809) );
  AOI21_X1 U20954 ( .B1(n17805), .B2(n17804), .A(n17888), .ZN(n17818) );
  OAI22_X1 U20955 ( .A1(n17885), .A2(n17807), .B1(n17806), .B2(n17818), .ZN(
        n17808) );
  AOI211_X1 U20956 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18209), .A(n17809), .B(
        n17808), .ZN(n17815) );
  OAI21_X1 U20957 ( .B1(n17811), .B2(n18143), .A(n17810), .ZN(n18140) );
  AOI22_X1 U20958 ( .A1(n17813), .A2(n18143), .B1(n17812), .B2(n18140), .ZN(
        n17814) );
  OAI211_X1 U20959 ( .C1(n17905), .C2(n18146), .A(n17815), .B(n17814), .ZN(
        P3_U2822) );
  OAI21_X1 U20960 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17817), .A(
        n17816), .ZN(n18149) );
  INV_X1 U20961 ( .A(n17818), .ZN(n17822) );
  NAND2_X1 U20962 ( .A1(n17819), .A2(n18607), .ZN(n17835) );
  NOR2_X1 U20963 ( .A1(n17836), .A2(n17835), .ZN(n17821) );
  NOR2_X1 U20964 ( .A1(n18175), .A2(n18768), .ZN(n18148) );
  AOI221_X1 U20965 ( .B1(n17822), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17821), .C2(n17820), .A(n18148), .ZN(n17829) );
  AOI21_X1 U20966 ( .B1(n17825), .B2(n17824), .A(n17823), .ZN(n17826) );
  XNOR2_X1 U20967 ( .A(n17826), .B(n18130), .ZN(n18151) );
  AOI22_X1 U20968 ( .A1(n17893), .A2(n18151), .B1(n17827), .B2(n17895), .ZN(
        n17828) );
  OAI211_X1 U20969 ( .C1(n17904), .C2(n18149), .A(n17829), .B(n17828), .ZN(
        P3_U2823) );
  OAI21_X1 U20970 ( .B1(n17831), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17830), .ZN(n18162) );
  OAI21_X1 U20971 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n18157) );
  OAI22_X1 U20972 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17835), .B1(
        n17904), .B2(n18157), .ZN(n17839) );
  NAND2_X1 U20973 ( .A1(n17896), .A2(n17835), .ZN(n17849) );
  OAI22_X1 U20974 ( .A1(n17885), .A2(n17837), .B1(n17836), .B2(n17849), .ZN(
        n17838) );
  AOI211_X1 U20975 ( .C1(n18209), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17839), .B(
        n17838), .ZN(n17840) );
  OAI21_X1 U20976 ( .B1(n17905), .B2(n18162), .A(n17840), .ZN(P3_U2824) );
  OAI21_X1 U20977 ( .B1(n17843), .B2(n17842), .A(n17841), .ZN(n18169) );
  OAI21_X1 U20978 ( .B1(n17845), .B2(n17888), .A(n17844), .ZN(n17846) );
  INV_X1 U20979 ( .A(n17846), .ZN(n17850) );
  OAI21_X1 U20980 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17848), .A(
        n17847), .ZN(n18163) );
  OAI22_X1 U20981 ( .A1(n17850), .A2(n17849), .B1(n17904), .B2(n18163), .ZN(
        n17851) );
  AOI21_X1 U20982 ( .B1(n17852), .B2(n17895), .A(n17851), .ZN(n17853) );
  NAND2_X1 U20983 ( .A1(n18209), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18167) );
  OAI211_X1 U20984 ( .C1(n17905), .C2(n18169), .A(n17853), .B(n18167), .ZN(
        P3_U2825) );
  OAI21_X1 U20985 ( .B1(n17856), .B2(n17855), .A(n17854), .ZN(n18174) );
  AOI22_X1 U20986 ( .A1(n18209), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18607), 
        .B2(n17857), .ZN(n17866) );
  OAI21_X1 U20987 ( .B1(n17859), .B2(n17858), .A(n17901), .ZN(n17876) );
  OAI21_X1 U20988 ( .B1(n17862), .B2(n17861), .A(n17860), .ZN(n18181) );
  OAI22_X1 U20989 ( .A1(n17885), .A2(n17863), .B1(n17904), .B2(n18181), .ZN(
        n17864) );
  AOI21_X1 U20990 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17876), .A(
        n17864), .ZN(n17865) );
  OAI211_X1 U20991 ( .C1(n17905), .C2(n18174), .A(n17866), .B(n17865), .ZN(
        P3_U2826) );
  OAI21_X1 U20992 ( .B1(n17869), .B2(n17868), .A(n17867), .ZN(n18186) );
  NOR2_X1 U20993 ( .A1(n17888), .A2(n17887), .ZN(n17875) );
  OAI21_X1 U20994 ( .B1(n17872), .B2(n17871), .A(n17870), .ZN(n18185) );
  OAI22_X1 U20995 ( .A1(n17885), .A2(n17873), .B1(n17904), .B2(n18185), .ZN(
        n17874) );
  AOI221_X1 U20996 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17876), .C1(
        n17875), .C2(n17876), .A(n17874), .ZN(n17877) );
  NAND2_X1 U20997 ( .A1(n18209), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18190) );
  OAI211_X1 U20998 ( .C1(n17905), .C2(n18186), .A(n17877), .B(n18190), .ZN(
        P3_U2827) );
  OAI21_X1 U20999 ( .B1(n17880), .B2(n17879), .A(n17878), .ZN(n18202) );
  OAI21_X1 U21000 ( .B1(n17883), .B2(n17882), .A(n17881), .ZN(n18207) );
  OAI22_X1 U21001 ( .A1(n17885), .A2(n17884), .B1(n17904), .B2(n18207), .ZN(
        n17886) );
  AOI221_X1 U21002 ( .B1(n17888), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18607), .C2(n17887), .A(n17886), .ZN(n17889) );
  NAND2_X1 U21003 ( .A1(n18209), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18205) );
  OAI211_X1 U21004 ( .C1(n17905), .C2(n18202), .A(n17889), .B(n18205), .ZN(
        P3_U2828) );
  OAI21_X1 U21005 ( .B1(n17891), .B2(n17899), .A(n17890), .ZN(n18214) );
  NAND2_X1 U21006 ( .A1(n18222), .A2(n17900), .ZN(n17892) );
  XNOR2_X1 U21007 ( .A(n17892), .B(n17891), .ZN(n18216) );
  AOI22_X1 U21008 ( .A1(n17893), .A2(n18216), .B1(n18209), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U21009 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17896), .B1(
        n17895), .B2(n17894), .ZN(n17897) );
  OAI211_X1 U21010 ( .C1(n17904), .C2(n18214), .A(n17898), .B(n17897), .ZN(
        P3_U2829) );
  AOI21_X1 U21011 ( .B1(n17900), .B2(n18222), .A(n17899), .ZN(n18226) );
  INV_X1 U21012 ( .A(n18226), .ZN(n18224) );
  OAI21_X1 U21013 ( .B1(n18731), .B2(n18880), .A(n17901), .ZN(n17902) );
  AOI22_X1 U21014 ( .A1(n18209), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17902), .ZN(n17903) );
  OAI221_X1 U21015 ( .B1(n18226), .B2(n17905), .C1(n18224), .C2(n17904), .A(
        n17903), .ZN(P3_U2830) );
  NOR2_X1 U21016 ( .A1(n18699), .A2(n18668), .ZN(n18193) );
  INV_X1 U21017 ( .A(n18193), .ZN(n18019) );
  INV_X1 U21018 ( .A(n18668), .ZN(n18695) );
  NOR2_X1 U21019 ( .A1(n18695), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18197) );
  AOI21_X1 U21020 ( .B1(n17906), .B2(n18019), .A(n18197), .ZN(n17943) );
  OAI21_X1 U21021 ( .B1(n17907), .B2(n18193), .A(n17943), .ZN(n17927) );
  AOI22_X1 U21022 ( .A1(n18687), .A2(n17909), .B1(n18097), .B2(n17908), .ZN(
        n17911) );
  OAI211_X1 U21023 ( .C1(n17912), .C2(n18193), .A(n17911), .B(n17910), .ZN(
        n17913) );
  NOR2_X1 U21024 ( .A1(n17927), .A2(n17913), .ZN(n17925) );
  AOI22_X1 U21025 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18218), .B1(
        n17914), .B2(n17948), .ZN(n17915) );
  AOI21_X1 U21026 ( .B1(n17925), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17915), .ZN(n17916) );
  AOI21_X1 U21027 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18204), .A(
        n17916), .ZN(n17918) );
  NAND2_X1 U21028 ( .A1(n18209), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17917) );
  OAI211_X1 U21029 ( .C1(n17919), .C2(n18127), .A(n17918), .B(n17917), .ZN(
        P3_U2835) );
  INV_X1 U21030 ( .A(n17980), .ZN(n17982) );
  AOI22_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18218), .B1(
        n17982), .B2(n17920), .ZN(n17924) );
  AOI22_X1 U21032 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18204), .B1(
        n18141), .B2(n17921), .ZN(n17923) );
  OAI211_X1 U21033 ( .C1(n17925), .C2(n17924), .A(n17923), .B(n17922), .ZN(
        P3_U2836) );
  INV_X1 U21034 ( .A(n17926), .ZN(n17966) );
  AOI221_X1 U21035 ( .B1(n17966), .B2(n18689), .C1(n17928), .C2(n18689), .A(
        n17927), .ZN(n17932) );
  OR2_X1 U21036 ( .A1(n17929), .A2(n17928), .ZN(n17931) );
  AOI221_X1 U21037 ( .B1(n17932), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17931), .C2(n17930), .A(n18182), .ZN(n17933) );
  AOI211_X1 U21038 ( .C1(n18204), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17934), .B(n17933), .ZN(n17938) );
  AOI22_X1 U21039 ( .A1(n18225), .A2(n17936), .B1(n18141), .B2(n17935), .ZN(
        n17937) );
  OAI211_X1 U21040 ( .C1(n18139), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        P3_U2837) );
  AOI22_X1 U21041 ( .A1(n18687), .A2(n17941), .B1(n18097), .B2(n17940), .ZN(
        n17942) );
  NAND3_X1 U21042 ( .A1(n17943), .A2(n17942), .A3(n18221), .ZN(n17946) );
  OAI21_X1 U21043 ( .B1(n17944), .B2(n18670), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17945) );
  OAI21_X1 U21044 ( .B1(n17946), .B2(n17945), .A(n18175), .ZN(n17956) );
  OAI21_X1 U21045 ( .B1(n17972), .B2(n17946), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17953) );
  AOI22_X1 U21046 ( .A1(n18141), .A2(n17949), .B1(n17948), .B2(n17947), .ZN(
        n17952) );
  INV_X1 U21047 ( .A(n17950), .ZN(n17951) );
  OAI211_X1 U21048 ( .C1(n17956), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2838) );
  NAND3_X1 U21049 ( .A1(n17955), .A2(n18221), .A3(n17954), .ZN(n17957) );
  AOI21_X1 U21050 ( .B1(n17958), .B2(n17957), .A(n17956), .ZN(n17959) );
  AOI21_X1 U21051 ( .B1(n17960), .B2(n18141), .A(n17959), .ZN(n17961) );
  NAND2_X1 U21052 ( .A1(n17962), .A2(n17961), .ZN(P3_U2839) );
  NAND2_X1 U21053 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17963), .ZN(
        n17971) );
  INV_X1 U21054 ( .A(n18097), .ZN(n18074) );
  OAI22_X1 U21055 ( .A1(n18044), .A2(n18201), .B1(n18045), .B2(n18074), .ZN(
        n17983) );
  NOR2_X1 U21056 ( .A1(n18687), .A2(n18097), .ZN(n18095) );
  AOI21_X1 U21057 ( .B1(n18017), .B2(n17993), .A(n18100), .ZN(n17964) );
  AOI221_X1 U21058 ( .B1(n17966), .B2(n18689), .C1(n17965), .C2(n18689), .A(
        n17964), .ZN(n17967) );
  OAI221_X1 U21059 ( .B1(n18695), .B2(n18033), .C1(n18695), .C2(n17981), .A(
        n17967), .ZN(n17995) );
  AOI21_X1 U21060 ( .B1(n18699), .B2(n17968), .A(n17995), .ZN(n17969) );
  OAI21_X1 U21061 ( .B1(n17970), .B2(n18095), .A(n17969), .ZN(n17984) );
  AOI211_X1 U21062 ( .C1(n17972), .C2(n17971), .A(n17983), .B(n17984), .ZN(
        n17974) );
  AOI221_X1 U21063 ( .B1(n17974), .B2(n18221), .C1(n18182), .C2(n18221), .A(
        n17973), .ZN(n17975) );
  AOI211_X1 U21064 ( .C1(n17977), .C2(n18141), .A(n17976), .B(n17975), .ZN(
        n17978) );
  OAI21_X1 U21065 ( .B1(n17980), .B2(n17979), .A(n17978), .ZN(P3_U2840) );
  NAND2_X1 U21066 ( .A1(n17982), .A2(n17981), .ZN(n18007) );
  NAND2_X1 U21067 ( .A1(n18695), .A2(n18670), .ZN(n18208) );
  AOI21_X1 U21068 ( .B1(n17985), .B2(n18208), .A(n17984), .ZN(n17987) );
  AOI211_X1 U21069 ( .C1(n18036), .C2(n17987), .A(n18209), .B(n17986), .ZN(
        n17988) );
  AOI211_X1 U21070 ( .C1(n18141), .C2(n17990), .A(n17989), .B(n17988), .ZN(
        n17991) );
  OAI21_X1 U21071 ( .B1(n17992), .B2(n18007), .A(n17991), .ZN(P3_U2841) );
  NAND3_X1 U21072 ( .A1(n18006), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18208), 
        .ZN(n17996) );
  OAI21_X1 U21073 ( .B1(n17993), .B2(n18095), .A(n18036), .ZN(n17994) );
  OAI21_X1 U21074 ( .B1(n17995), .B2(n17994), .A(n18175), .ZN(n18005) );
  NAND2_X1 U21075 ( .A1(n17996), .A2(n18005), .ZN(n17998) );
  AOI22_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17998), .B1(
        n18141), .B2(n17997), .ZN(n18000) );
  NAND2_X1 U21077 ( .A1(n18209), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17999) );
  OAI211_X1 U21078 ( .C1(n18001), .C2(n18007), .A(n18000), .B(n17999), .ZN(
        P3_U2842) );
  AOI21_X1 U21079 ( .B1(n18141), .B2(n18003), .A(n18002), .ZN(n18004) );
  OAI221_X1 U21080 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18007), 
        .C1(n18006), .C2(n18005), .A(n18004), .ZN(P3_U2843) );
  INV_X1 U21081 ( .A(n18198), .ZN(n18170) );
  INV_X1 U21082 ( .A(n18008), .ZN(n18171) );
  AOI22_X1 U21083 ( .A1(n18689), .A2(n18170), .B1(n18171), .B2(n18009), .ZN(
        n18184) );
  NOR2_X1 U21084 ( .A1(n18184), .A2(n18010), .ZN(n18147) );
  NAND2_X1 U21085 ( .A1(n18011), .A2(n18147), .ZN(n18043) );
  AND2_X1 U21086 ( .A1(n18012), .A2(n18043), .ZN(n18085) );
  NAND2_X1 U21087 ( .A1(n18013), .A2(n18123), .ZN(n18041) );
  AOI21_X1 U21088 ( .B1(n18015), .B2(n18141), .A(n18014), .ZN(n18025) );
  NOR2_X1 U21089 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18193), .ZN(
        n18023) );
  INV_X1 U21090 ( .A(n18197), .ZN(n18016) );
  NAND3_X1 U21091 ( .A1(n18017), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18016), .ZN(n18018) );
  AOI22_X1 U21092 ( .A1(n18689), .A2(n18020), .B1(n18019), .B2(n18018), .ZN(
        n18021) );
  OAI211_X1 U21093 ( .C1(n18022), .C2(n18095), .A(n18036), .B(n18021), .ZN(
        n18029) );
  OAI211_X1 U21094 ( .C1(n18023), .C2(n18029), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n18175), .ZN(n18024) );
  OAI211_X1 U21095 ( .C1(n18041), .C2(n18026), .A(n18025), .B(n18024), .ZN(
        P3_U2844) );
  INV_X1 U21096 ( .A(n18041), .ZN(n18028) );
  AOI22_X1 U21097 ( .A1(n18209), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18028), 
        .B2(n18027), .ZN(n18031) );
  NAND3_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18175), .A3(
        n18029), .ZN(n18030) );
  OAI211_X1 U21099 ( .C1(n18032), .C2(n18127), .A(n18031), .B(n18030), .ZN(
        P3_U2845) );
  AOI21_X1 U21100 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18695), .A(
        n18033), .ZN(n18035) );
  NAND2_X1 U21101 ( .A1(n18689), .A2(n18034), .ZN(n18103) );
  OAI21_X1 U21102 ( .B1(n18100), .B2(n18099), .A(n18103), .ZN(n18077) );
  AOI211_X1 U21103 ( .C1(n18073), .C2(n18059), .A(n18035), .B(n18077), .ZN(
        n18052) );
  AOI221_X1 U21104 ( .B1(n18135), .B2(n18036), .C1(n18052), .C2(n18036), .A(
        n18209), .ZN(n18038) );
  AOI22_X1 U21105 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18038), .B1(
        n18141), .B2(n18037), .ZN(n18040) );
  NAND2_X1 U21106 ( .A1(n18209), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18039) );
  OAI211_X1 U21107 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18041), .A(
        n18040), .B(n18039), .ZN(P3_U2846) );
  NOR2_X1 U21108 ( .A1(n18043), .A2(n18042), .ZN(n18064) );
  AOI21_X1 U21109 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18064), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18051) );
  NOR2_X1 U21110 ( .A1(n18044), .A2(n18201), .ZN(n18049) );
  NOR2_X1 U21111 ( .A1(n18045), .A2(n18074), .ZN(n18047) );
  AOI22_X1 U21112 ( .A1(n18049), .A2(n18048), .B1(n18047), .B2(n18046), .ZN(
        n18050) );
  OAI21_X1 U21113 ( .B1(n18052), .B2(n18051), .A(n18050), .ZN(n18055) );
  INV_X1 U21114 ( .A(n18053), .ZN(n18054) );
  AOI22_X1 U21115 ( .A1(n18218), .A2(n18055), .B1(n18141), .B2(n18054), .ZN(
        n18057) );
  OAI211_X1 U21116 ( .C1(n18221), .C2(n18058), .A(n18057), .B(n18056), .ZN(
        P3_U2847) );
  INV_X1 U21117 ( .A(n18208), .ZN(n18062) );
  OAI21_X1 U21118 ( .B1(n18060), .B2(n18073), .A(n18059), .ZN(n18061) );
  OAI21_X1 U21119 ( .B1(n18086), .B2(n18101), .A(n18668), .ZN(n18079) );
  OAI211_X1 U21120 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18062), .A(
        n18061), .B(n18079), .ZN(n18063) );
  OAI22_X1 U21121 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18064), .B1(
        n18063), .B2(n18077), .ZN(n18065) );
  OAI22_X1 U21122 ( .A1(n18175), .A2(n18783), .B1(n18182), .B2(n18065), .ZN(
        n18069) );
  OAI22_X1 U21123 ( .A1(n18067), .A2(n18127), .B1(n18139), .B2(n18066), .ZN(
        n18068) );
  AOI211_X1 U21124 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18204), .A(
        n18069), .B(n18068), .ZN(n18070) );
  OAI21_X1 U21125 ( .B1(n18187), .B2(n18071), .A(n18070), .ZN(P3_U2848) );
  AOI22_X1 U21126 ( .A1(n18209), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18123), 
        .B2(n18072), .ZN(n18082) );
  INV_X1 U21127 ( .A(n18073), .ZN(n18116) );
  AOI21_X1 U21128 ( .B1(n18699), .B2(n18108), .A(n12793), .ZN(n18088) );
  AOI22_X1 U21129 ( .A1(n18689), .A2(n18084), .B1(n18699), .B2(n18107), .ZN(
        n18109) );
  OAI21_X1 U21130 ( .B1(n18075), .B2(n18074), .A(n18109), .ZN(n18076) );
  AOI211_X1 U21131 ( .C1(n18687), .C2(n18078), .A(n18077), .B(n18076), .ZN(
        n18087) );
  OAI211_X1 U21132 ( .C1(n18116), .C2(n18088), .A(n18087), .B(n18079), .ZN(
        n18080) );
  OAI211_X1 U21133 ( .C1(n18182), .C2(n18080), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18175), .ZN(n18081) );
  OAI211_X1 U21134 ( .C1(n18127), .C2(n18083), .A(n18082), .B(n18081), .ZN(
        P3_U2849) );
  AOI221_X1 U21135 ( .B1(n18085), .B2(n12793), .C1(n18084), .C2(n12793), .A(
        n18182), .ZN(n18091) );
  NOR2_X1 U21136 ( .A1(n18086), .A2(n18101), .ZN(n18089) );
  OAI211_X1 U21137 ( .C1(n18089), .C2(n18695), .A(n18088), .B(n18087), .ZN(
        n18090) );
  AOI22_X1 U21138 ( .A1(n18141), .A2(n18092), .B1(n18091), .B2(n18090), .ZN(
        n18094) );
  OAI211_X1 U21139 ( .C1(n18221), .C2(n12793), .A(n18094), .B(n18093), .ZN(
        P3_U2850) );
  INV_X1 U21140 ( .A(n18095), .ZN(n18106) );
  AOI22_X1 U21141 ( .A1(n18687), .A2(n18098), .B1(n18097), .B2(n18096), .ZN(
        n18105) );
  NOR2_X1 U21142 ( .A1(n18100), .A2(n18099), .ZN(n18102) );
  OAI21_X1 U21143 ( .B1(n18102), .B2(n18668), .A(n18101), .ZN(n18104) );
  NAND4_X1 U21144 ( .A1(n18218), .A2(n18105), .A3(n18104), .A4(n18103), .ZN(
        n18124) );
  AOI221_X1 U21145 ( .B1(n18668), .B2(n18107), .C1(n18106), .C2(n18107), .A(
        n18124), .ZN(n18115) );
  AOI211_X1 U21146 ( .C1(n18109), .C2(n18115), .A(n18209), .B(n18108), .ZN(
        n18110) );
  AOI21_X1 U21147 ( .B1(n18123), .B2(n18111), .A(n18110), .ZN(n18113) );
  OAI211_X1 U21148 ( .C1(n18114), .C2(n18127), .A(n18113), .B(n18112), .ZN(
        P3_U2851) );
  AOI221_X1 U21149 ( .B1(n18116), .B2(n18115), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18115), .A(n18209), .ZN(
        n18117) );
  AOI22_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18117), .B1(
        n18209), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18120) );
  NAND3_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18123), .A3(
        n18118), .ZN(n18119) );
  OAI211_X1 U21152 ( .C1(n18121), .C2(n18127), .A(n18120), .B(n18119), .ZN(
        P3_U2852) );
  AOI22_X1 U21153 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18209), .B1(n18123), 
        .B2(n18122), .ZN(n18126) );
  NAND3_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18175), .A3(
        n18124), .ZN(n18125) );
  OAI211_X1 U21155 ( .C1(n18128), .C2(n18127), .A(n18126), .B(n18125), .ZN(
        P3_U2853) );
  NOR3_X1 U21156 ( .A1(n18184), .A2(n18182), .A3(n12774), .ZN(n18179) );
  NAND3_X1 U21157 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18179), .ZN(n18158) );
  NOR3_X1 U21158 ( .A1(n18130), .A2(n18129), .A3(n18158), .ZN(n18138) );
  OAI22_X1 U21159 ( .A1(n18132), .A2(n18670), .B1(n18131), .B2(n18193), .ZN(
        n18133) );
  NOR2_X1 U21160 ( .A1(n18197), .A2(n18133), .ZN(n18156) );
  OAI211_X1 U21161 ( .C1(n18135), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18156), .ZN(n18134) );
  NAND2_X1 U21162 ( .A1(n18218), .A2(n18134), .ZN(n18154) );
  OAI21_X1 U21163 ( .B1(n18135), .B2(n18154), .A(n18221), .ZN(n18137) );
  NOR2_X1 U21164 ( .A1(n18175), .A2(n18770), .ZN(n18136) );
  AOI221_X1 U21165 ( .B1(n18138), .B2(n9811), .C1(n18137), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18136), .ZN(n18145) );
  INV_X1 U21166 ( .A(n18139), .ZN(n18142) );
  AOI22_X1 U21167 ( .A1(n18143), .A2(n18142), .B1(n18141), .B2(n18140), .ZN(
        n18144) );
  OAI211_X1 U21168 ( .C1(n18187), .C2(n18146), .A(n18145), .B(n18144), .ZN(
        P3_U2854) );
  AOI21_X1 U21169 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18147), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18155) );
  AOI21_X1 U21170 ( .B1(n18204), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18148), .ZN(n18153) );
  INV_X1 U21171 ( .A(n18149), .ZN(n18150) );
  AOI22_X1 U21172 ( .A1(n18225), .A2(n18151), .B1(n18227), .B2(n18150), .ZN(
        n18152) );
  OAI211_X1 U21173 ( .C1(n18155), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        P3_U2855) );
  OAI21_X1 U21174 ( .B1(n18156), .B2(n18182), .A(n18221), .ZN(n18166) );
  NOR2_X1 U21175 ( .A1(n18175), .A2(n18766), .ZN(n18160) );
  INV_X1 U21176 ( .A(n18227), .ZN(n18213) );
  OAI22_X1 U21177 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18158), .B1(
        n18157), .B2(n18213), .ZN(n18159) );
  AOI211_X1 U21178 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18166), .A(
        n18160), .B(n18159), .ZN(n18161) );
  OAI21_X1 U21179 ( .B1(n18187), .B2(n18162), .A(n18161), .ZN(P3_U2856) );
  NAND2_X1 U21180 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18179), .ZN(
        n18164) );
  OAI22_X1 U21181 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18164), .B1(
        n18163), .B2(n18213), .ZN(n18165) );
  AOI21_X1 U21182 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18166), .A(
        n18165), .ZN(n18168) );
  OAI211_X1 U21183 ( .C1(n18187), .C2(n18169), .A(n18168), .B(n18167), .ZN(
        P3_U2857) );
  OAI22_X1 U21184 ( .A1(n18171), .A2(n18193), .B1(n18670), .B2(n18170), .ZN(
        n18172) );
  NOR3_X1 U21185 ( .A1(n18197), .A2(n12774), .A3(n18172), .ZN(n18183) );
  OAI21_X1 U21186 ( .B1(n18183), .B2(n18173), .A(n18221), .ZN(n18177) );
  OAI22_X1 U21187 ( .A1(n18175), .A2(n18762), .B1(n18187), .B2(n18174), .ZN(
        n18176) );
  AOI221_X1 U21188 ( .B1(n18179), .B2(n18178), .C1(n18177), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18176), .ZN(n18180) );
  OAI21_X1 U21189 ( .B1(n18213), .B2(n18181), .A(n18180), .ZN(P3_U2858) );
  AOI211_X1 U21190 ( .C1(n18184), .C2(n12774), .A(n18183), .B(n18182), .ZN(
        n18189) );
  OAI22_X1 U21191 ( .A1(n18187), .A2(n18186), .B1(n18213), .B2(n18185), .ZN(
        n18188) );
  NOR2_X1 U21192 ( .A1(n18189), .A2(n18188), .ZN(n18191) );
  OAI211_X1 U21193 ( .C1(n18221), .C2(n12774), .A(n18191), .B(n18190), .ZN(
        P3_U2859) );
  NAND2_X1 U21194 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18192) );
  OAI22_X1 U21195 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18193), .B1(
        n18670), .B2(n18192), .ZN(n18196) );
  INV_X1 U21196 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18836) );
  NOR3_X1 U21197 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18836), .A3(
        n18194), .ZN(n18195) );
  AOI221_X1 U21198 ( .B1(n18197), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18196), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18195), .ZN(
        n18200) );
  NAND2_X1 U21199 ( .A1(n18689), .A2(n18198), .ZN(n18199) );
  OAI211_X1 U21200 ( .C1(n18202), .C2(n18201), .A(n18200), .B(n18199), .ZN(
        n18203) );
  AOI22_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18204), .B1(
        n18218), .B2(n18203), .ZN(n18206) );
  OAI211_X1 U21202 ( .C1(n18207), .C2(n18213), .A(n18206), .B(n18205), .ZN(
        P3_U2860) );
  NAND3_X1 U21203 ( .A1(n18218), .A2(n18222), .A3(n18208), .ZN(n18219) );
  NAND2_X1 U21204 ( .A1(n18209), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18212) );
  OAI211_X1 U21205 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18699), .A(
        n18210), .B(n18836), .ZN(n18211) );
  OAI211_X1 U21206 ( .C1(n18214), .C2(n18213), .A(n18212), .B(n18211), .ZN(
        n18215) );
  AOI21_X1 U21207 ( .B1(n18225), .B2(n18216), .A(n18215), .ZN(n18217) );
  OAI221_X1 U21208 ( .B1(n18836), .B2(n18221), .C1(n18836), .C2(n18219), .A(
        n18217), .ZN(P3_U2861) );
  NAND2_X1 U21209 ( .A1(n18218), .A2(n18699), .ZN(n18220) );
  OAI221_X1 U21210 ( .B1(n18222), .B2(n18221), .C1(n18222), .C2(n18220), .A(
        n18219), .ZN(n18223) );
  AOI221_X1 U21211 ( .B1(n18227), .B2(n18226), .C1(n18225), .C2(n18224), .A(
        n18223), .ZN(n18228) );
  OAI21_X1 U21212 ( .B1(n18175), .B2(n18864), .A(n18228), .ZN(P3_U2862) );
  AOI21_X1 U21213 ( .B1(n18231), .B2(n18230), .A(n18229), .ZN(n18721) );
  OAI21_X1 U21214 ( .B1(n18721), .B2(n18284), .A(n18236), .ZN(n18232) );
  OAI221_X1 U21215 ( .B1(n18482), .B2(n18872), .C1(n18482), .C2(n18236), .A(
        n18232), .ZN(P3_U2863) );
  INV_X1 U21216 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18708) );
  NOR2_X1 U21217 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18240), .ZN(
        n18418) );
  NOR2_X1 U21218 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18708), .ZN(
        n18506) );
  NOR2_X1 U21219 ( .A1(n18418), .A2(n18506), .ZN(n18234) );
  OAI22_X1 U21220 ( .A1(n18235), .A2(n18708), .B1(n18234), .B2(n18233), .ZN(
        P3_U2866) );
  NOR2_X1 U21221 ( .A1(n18706), .A2(n18236), .ZN(P3_U2867) );
  NOR2_X1 U21222 ( .A1(n18238), .A2(n18237), .ZN(n18275) );
  NAND2_X1 U21223 ( .A1(n18275), .A2(n18239), .ZN(n18611) );
  NOR2_X1 U21224 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18701) );
  NAND2_X1 U21225 ( .A1(n18240), .A2(n18708), .ZN(n18305) );
  INV_X1 U21226 ( .A(n18305), .ZN(n18328) );
  NAND2_X1 U21227 ( .A1(n18701), .A2(n18328), .ZN(n18283) );
  AND2_X1 U21228 ( .A1(n18607), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18608) );
  NOR2_X1 U21229 ( .A1(n18708), .A2(n18416), .ZN(n18605) );
  NAND2_X1 U21230 ( .A1(n18482), .A2(n18605), .ZN(n18600) );
  INV_X1 U21231 ( .A(n18600), .ZN(n18580) );
  NOR2_X2 U21232 ( .A1(n18285), .A2(n18241), .ZN(n18602) );
  INV_X1 U21233 ( .A(n18729), .ZN(n18574) );
  NOR2_X1 U21234 ( .A1(n20892), .A2(n18482), .ZN(n18700) );
  INV_X1 U21235 ( .A(n18700), .ZN(n18242) );
  NAND2_X1 U21236 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18551) );
  NOR2_X2 U21237 ( .A1(n18242), .A2(n18551), .ZN(n18601) );
  INV_X1 U21238 ( .A(n18283), .ZN(n18343) );
  NOR2_X1 U21239 ( .A1(n18601), .A2(n18343), .ZN(n18306) );
  NOR2_X1 U21240 ( .A1(n18574), .A2(n18306), .ZN(n18279) );
  AOI22_X1 U21241 ( .A1(n18608), .A2(n18580), .B1(n18602), .B2(n18279), .ZN(
        n18247) );
  NAND2_X1 U21242 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20892), .ZN(
        n18370) );
  NOR2_X2 U21243 ( .A1(n18370), .A2(n18551), .ZN(n18650) );
  NOR2_X1 U21244 ( .A1(n18650), .A2(n18580), .ZN(n18575) );
  INV_X1 U21245 ( .A(n18243), .ZN(n18576) );
  OAI22_X1 U21246 ( .A1(n18306), .A2(n18244), .B1(n18575), .B2(n18576), .ZN(
        n18245) );
  NAND2_X1 U21247 ( .A1(n18579), .A2(n18245), .ZN(n18280) );
  AND2_X1 U21248 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18607), .ZN(n18603) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18280), .B1(
        n18603), .B2(n18650), .ZN(n18246) );
  OAI211_X1 U21250 ( .C1(n18611), .C2(n18283), .A(n18247), .B(n18246), .ZN(
        P3_U2868) );
  NAND2_X1 U21251 ( .A1(n18275), .A2(n18248), .ZN(n18617) );
  AND2_X1 U21252 ( .A1(n18607), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18614) );
  AND2_X1 U21253 ( .A1(n18579), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U21254 ( .A1(n18614), .A2(n18580), .B1(n18612), .B2(n18279), .ZN(
        n18250) );
  AND2_X1 U21255 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18607), .ZN(n18613) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18280), .B1(
        n18613), .B2(n18650), .ZN(n18249) );
  OAI211_X1 U21257 ( .C1(n18617), .C2(n18283), .A(n18250), .B(n18249), .ZN(
        P3_U2869) );
  NAND2_X1 U21258 ( .A1(n18275), .A2(n18251), .ZN(n18623) );
  AND2_X1 U21259 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18607), .ZN(n18619) );
  NOR2_X2 U21260 ( .A1(n18285), .A2(n18252), .ZN(n18618) );
  AOI22_X1 U21261 ( .A1(n18619), .A2(n18650), .B1(n18618), .B2(n18279), .ZN(
        n18254) );
  AND2_X1 U21262 ( .A1(n18607), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18280), .B1(
        n18620), .B2(n18580), .ZN(n18253) );
  OAI211_X1 U21264 ( .C1(n18623), .C2(n18283), .A(n18254), .B(n18253), .ZN(
        P3_U2870) );
  NAND2_X1 U21265 ( .A1(n18275), .A2(n18255), .ZN(n18629) );
  NOR2_X2 U21266 ( .A1(n18278), .A2(n18256), .ZN(n18625) );
  NOR2_X2 U21267 ( .A1(n18285), .A2(n18257), .ZN(n18624) );
  AOI22_X1 U21268 ( .A1(n18625), .A2(n18580), .B1(n18624), .B2(n18279), .ZN(
        n18259) );
  AND2_X1 U21269 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18607), .ZN(n18626) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18280), .B1(
        n18626), .B2(n18650), .ZN(n18258) );
  OAI211_X1 U21271 ( .C1(n18629), .C2(n18283), .A(n18259), .B(n18258), .ZN(
        P3_U2871) );
  NAND2_X1 U21272 ( .A1(n18275), .A2(n18260), .ZN(n18635) );
  NOR2_X2 U21273 ( .A1(n18285), .A2(n18261), .ZN(n18631) );
  NOR2_X2 U21274 ( .A1(n18278), .A2(n20883), .ZN(n18630) );
  AOI22_X1 U21275 ( .A1(n18631), .A2(n18279), .B1(n18630), .B2(n18580), .ZN(
        n18263) );
  AND2_X1 U21276 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18607), .ZN(n18632) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18280), .B1(
        n18632), .B2(n18650), .ZN(n18262) );
  OAI211_X1 U21278 ( .C1(n18635), .C2(n18283), .A(n18263), .B(n18262), .ZN(
        P3_U2872) );
  NAND2_X1 U21279 ( .A1(n18275), .A2(n18264), .ZN(n18641) );
  NOR2_X2 U21280 ( .A1(n18278), .A2(n18265), .ZN(n18638) );
  NOR2_X2 U21281 ( .A1(n18285), .A2(n18266), .ZN(n18636) );
  AOI22_X1 U21282 ( .A1(n18638), .A2(n18580), .B1(n18636), .B2(n18279), .ZN(
        n18268) );
  AND2_X1 U21283 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18607), .ZN(n18637) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18280), .B1(
        n18637), .B2(n18650), .ZN(n18267) );
  OAI211_X1 U21285 ( .C1(n18641), .C2(n18283), .A(n18268), .B(n18267), .ZN(
        P3_U2873) );
  NAND2_X1 U21286 ( .A1(n18275), .A2(n18269), .ZN(n18647) );
  NOR2_X2 U21287 ( .A1(n18270), .A2(n18278), .ZN(n18643) );
  NOR2_X2 U21288 ( .A1(n18285), .A2(n18271), .ZN(n18642) );
  AOI22_X1 U21289 ( .A1(n18643), .A2(n18650), .B1(n18642), .B2(n18279), .ZN(
        n18273) );
  AND2_X1 U21290 ( .A1(n18607), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18644) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18280), .B1(
        n18644), .B2(n18580), .ZN(n18272) );
  OAI211_X1 U21292 ( .C1(n18647), .C2(n18283), .A(n18273), .B(n18272), .ZN(
        P3_U2874) );
  NAND2_X1 U21293 ( .A1(n18275), .A2(n18274), .ZN(n18658) );
  NOR2_X2 U21294 ( .A1(n18276), .A2(n18285), .ZN(n18649) );
  NOR2_X2 U21295 ( .A1(n18278), .A2(n18277), .ZN(n18653) );
  AOI22_X1 U21296 ( .A1(n18649), .A2(n18279), .B1(n18653), .B2(n18650), .ZN(
        n18282) );
  AND2_X1 U21297 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18607), .ZN(n18651) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18280), .B1(
        n18651), .B2(n18580), .ZN(n18281) );
  OAI211_X1 U21299 ( .C1(n18658), .C2(n18283), .A(n18282), .B(n18281), .ZN(
        P3_U2875) );
  NOR2_X2 U21300 ( .A1(n18305), .A2(n18370), .ZN(n18365) );
  INV_X1 U21301 ( .A(n18365), .ZN(n18304) );
  NAND2_X1 U21302 ( .A1(n20892), .A2(n18729), .ZN(n18550) );
  NOR2_X1 U21303 ( .A1(n18305), .A2(n18550), .ZN(n18300) );
  AOI22_X1 U21304 ( .A1(n18603), .A2(n18580), .B1(n18602), .B2(n18300), .ZN(
        n18287) );
  NOR2_X1 U21305 ( .A1(n18285), .A2(n18284), .ZN(n18604) );
  INV_X1 U21306 ( .A(n18604), .ZN(n18327) );
  NOR2_X1 U21307 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18327), .ZN(
        n18552) );
  AOI22_X1 U21308 ( .A1(n18607), .A2(n18605), .B1(n18328), .B2(n18552), .ZN(
        n18301) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18301), .B1(
        n18608), .B2(n18601), .ZN(n18286) );
  OAI211_X1 U21310 ( .C1(n18304), .C2(n18611), .A(n18287), .B(n18286), .ZN(
        P3_U2876) );
  AOI22_X1 U21311 ( .A1(n18613), .A2(n18580), .B1(n18612), .B2(n18300), .ZN(
        n18289) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18301), .B1(
        n18614), .B2(n18601), .ZN(n18288) );
  OAI211_X1 U21313 ( .C1(n18304), .C2(n18617), .A(n18289), .B(n18288), .ZN(
        P3_U2877) );
  AOI22_X1 U21314 ( .A1(n18619), .A2(n18580), .B1(n18618), .B2(n18300), .ZN(
        n18291) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18301), .B1(
        n18620), .B2(n18601), .ZN(n18290) );
  OAI211_X1 U21316 ( .C1(n18304), .C2(n18623), .A(n18291), .B(n18290), .ZN(
        P3_U2878) );
  AOI22_X1 U21317 ( .A1(n18626), .A2(n18580), .B1(n18624), .B2(n18300), .ZN(
        n18293) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18301), .B1(
        n18625), .B2(n18601), .ZN(n18292) );
  OAI211_X1 U21319 ( .C1(n18304), .C2(n18629), .A(n18293), .B(n18292), .ZN(
        P3_U2879) );
  AOI22_X1 U21320 ( .A1(n18631), .A2(n18300), .B1(n18630), .B2(n18601), .ZN(
        n18295) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18301), .B1(
        n18632), .B2(n18580), .ZN(n18294) );
  OAI211_X1 U21322 ( .C1(n18304), .C2(n18635), .A(n18295), .B(n18294), .ZN(
        P3_U2880) );
  AOI22_X1 U21323 ( .A1(n18638), .A2(n18601), .B1(n18636), .B2(n18300), .ZN(
        n18297) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18301), .B1(
        n18637), .B2(n18580), .ZN(n18296) );
  OAI211_X1 U21325 ( .C1(n18304), .C2(n18641), .A(n18297), .B(n18296), .ZN(
        P3_U2881) );
  AOI22_X1 U21326 ( .A1(n18642), .A2(n18300), .B1(n18644), .B2(n18601), .ZN(
        n18299) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18301), .B1(
        n18643), .B2(n18580), .ZN(n18298) );
  OAI211_X1 U21328 ( .C1(n18304), .C2(n18647), .A(n18299), .B(n18298), .ZN(
        P3_U2882) );
  AOI22_X1 U21329 ( .A1(n18651), .A2(n18601), .B1(n18649), .B2(n18300), .ZN(
        n18303) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18301), .B1(
        n18653), .B2(n18580), .ZN(n18302) );
  OAI211_X1 U21331 ( .C1(n18304), .C2(n18658), .A(n18303), .B(n18302), .ZN(
        P3_U2883) );
  NOR2_X1 U21332 ( .A1(n20892), .A2(n18305), .ZN(n18373) );
  NAND2_X1 U21333 ( .A1(n18482), .A2(n18373), .ZN(n18326) );
  INV_X1 U21334 ( .A(n18326), .ZN(n18389) );
  NOR2_X1 U21335 ( .A1(n18389), .A2(n18365), .ZN(n18348) );
  NOR2_X1 U21336 ( .A1(n18574), .A2(n18348), .ZN(n18322) );
  AOI22_X1 U21337 ( .A1(n18608), .A2(n18343), .B1(n18602), .B2(n18322), .ZN(
        n18309) );
  OAI21_X1 U21338 ( .B1(n18306), .B2(n18576), .A(n18348), .ZN(n18307) );
  OAI211_X1 U21339 ( .C1(n18389), .C2(n18830), .A(n18579), .B(n18307), .ZN(
        n18323) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18323), .B1(
        n18603), .B2(n18601), .ZN(n18308) );
  OAI211_X1 U21341 ( .C1(n18326), .C2(n18611), .A(n18309), .B(n18308), .ZN(
        P3_U2884) );
  AOI22_X1 U21342 ( .A1(n18614), .A2(n18343), .B1(n18612), .B2(n18322), .ZN(
        n18311) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18323), .B1(
        n18613), .B2(n18601), .ZN(n18310) );
  OAI211_X1 U21344 ( .C1(n18326), .C2(n18617), .A(n18311), .B(n18310), .ZN(
        P3_U2885) );
  AOI22_X1 U21345 ( .A1(n18620), .A2(n18343), .B1(n18618), .B2(n18322), .ZN(
        n18313) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18323), .B1(
        n18619), .B2(n18601), .ZN(n18312) );
  OAI211_X1 U21347 ( .C1(n18326), .C2(n18623), .A(n18313), .B(n18312), .ZN(
        P3_U2886) );
  AOI22_X1 U21348 ( .A1(n18626), .A2(n18601), .B1(n18624), .B2(n18322), .ZN(
        n18315) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18323), .B1(
        n18625), .B2(n18343), .ZN(n18314) );
  OAI211_X1 U21350 ( .C1(n18326), .C2(n18629), .A(n18315), .B(n18314), .ZN(
        P3_U2887) );
  AOI22_X1 U21351 ( .A1(n18632), .A2(n18601), .B1(n18631), .B2(n18322), .ZN(
        n18317) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18323), .B1(
        n18630), .B2(n18343), .ZN(n18316) );
  OAI211_X1 U21353 ( .C1(n18326), .C2(n18635), .A(n18317), .B(n18316), .ZN(
        P3_U2888) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18323), .B1(
        n18636), .B2(n18322), .ZN(n18319) );
  AOI22_X1 U21355 ( .A1(n18638), .A2(n18343), .B1(n18637), .B2(n18601), .ZN(
        n18318) );
  OAI211_X1 U21356 ( .C1(n18326), .C2(n18641), .A(n18319), .B(n18318), .ZN(
        P3_U2889) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18323), .B1(
        n18642), .B2(n18322), .ZN(n18321) );
  AOI22_X1 U21358 ( .A1(n18643), .A2(n18601), .B1(n18644), .B2(n18343), .ZN(
        n18320) );
  OAI211_X1 U21359 ( .C1(n18326), .C2(n18647), .A(n18321), .B(n18320), .ZN(
        P3_U2890) );
  AOI22_X1 U21360 ( .A1(n18649), .A2(n18322), .B1(n18653), .B2(n18601), .ZN(
        n18325) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18323), .B1(
        n18651), .B2(n18343), .ZN(n18324) );
  OAI211_X1 U21362 ( .C1(n18326), .C2(n18658), .A(n18325), .B(n18324), .ZN(
        P3_U2891) );
  NAND2_X1 U21363 ( .A1(n18700), .A2(n18328), .ZN(n18371) );
  AND2_X1 U21364 ( .A1(n18729), .A2(n18373), .ZN(n18344) );
  AOI22_X1 U21365 ( .A1(n18603), .A2(n18343), .B1(n18602), .B2(n18344), .ZN(
        n18330) );
  AOI21_X1 U21366 ( .B1(n20892), .B2(n18576), .A(n18327), .ZN(n18417) );
  NAND2_X1 U21367 ( .A1(n18328), .A2(n18417), .ZN(n18345) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18345), .B1(
        n18608), .B2(n18365), .ZN(n18329) );
  OAI211_X1 U21369 ( .C1(n18371), .C2(n18611), .A(n18330), .B(n18329), .ZN(
        P3_U2892) );
  AOI22_X1 U21370 ( .A1(n18613), .A2(n18343), .B1(n18612), .B2(n18344), .ZN(
        n18332) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18614), .ZN(n18331) );
  OAI211_X1 U21372 ( .C1(n18371), .C2(n18617), .A(n18332), .B(n18331), .ZN(
        P3_U2893) );
  AOI22_X1 U21373 ( .A1(n18365), .A2(n18620), .B1(n18618), .B2(n18344), .ZN(
        n18334) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18345), .B1(
        n18619), .B2(n18343), .ZN(n18333) );
  OAI211_X1 U21375 ( .C1(n18371), .C2(n18623), .A(n18334), .B(n18333), .ZN(
        P3_U2894) );
  AOI22_X1 U21376 ( .A1(n18626), .A2(n18343), .B1(n18624), .B2(n18344), .ZN(
        n18336) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18625), .ZN(n18335) );
  OAI211_X1 U21378 ( .C1(n18371), .C2(n18629), .A(n18336), .B(n18335), .ZN(
        P3_U2895) );
  AOI22_X1 U21379 ( .A1(n18632), .A2(n18343), .B1(n18631), .B2(n18344), .ZN(
        n18338) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18630), .ZN(n18337) );
  OAI211_X1 U21381 ( .C1(n18371), .C2(n18635), .A(n18338), .B(n18337), .ZN(
        P3_U2896) );
  AOI22_X1 U21382 ( .A1(n18637), .A2(n18343), .B1(n18636), .B2(n18344), .ZN(
        n18340) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18638), .ZN(n18339) );
  OAI211_X1 U21384 ( .C1(n18371), .C2(n18641), .A(n18340), .B(n18339), .ZN(
        P3_U2897) );
  AOI22_X1 U21385 ( .A1(n18643), .A2(n18343), .B1(n18642), .B2(n18344), .ZN(
        n18342) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18644), .ZN(n18341) );
  OAI211_X1 U21387 ( .C1(n18371), .C2(n18647), .A(n18342), .B(n18341), .ZN(
        P3_U2898) );
  AOI22_X1 U21388 ( .A1(n18649), .A2(n18344), .B1(n18653), .B2(n18343), .ZN(
        n18347) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18345), .B1(
        n18365), .B2(n18651), .ZN(n18346) );
  OAI211_X1 U21390 ( .C1(n18371), .C2(n18658), .A(n18347), .B(n18346), .ZN(
        P3_U2899) );
  NAND2_X1 U21391 ( .A1(n18701), .A2(n18418), .ZN(n18369) );
  AOI21_X1 U21392 ( .B1(n18369), .B2(n18371), .A(n18574), .ZN(n18364) );
  AOI22_X1 U21393 ( .A1(n18365), .A2(n18603), .B1(n18602), .B2(n18364), .ZN(
        n18351) );
  INV_X1 U21394 ( .A(n18369), .ZN(n18434) );
  AOI221_X1 U21395 ( .B1(n18348), .B2(n18371), .C1(n18576), .C2(n18371), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18349) );
  OAI21_X1 U21396 ( .B1(n18434), .B2(n18349), .A(n18579), .ZN(n18366) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18366), .B1(
        n18608), .B2(n18389), .ZN(n18350) );
  OAI211_X1 U21398 ( .C1(n18369), .C2(n18611), .A(n18351), .B(n18350), .ZN(
        P3_U2900) );
  AOI22_X1 U21399 ( .A1(n18389), .A2(n18614), .B1(n18364), .B2(n18612), .ZN(
        n18353) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18366), .B1(
        n18365), .B2(n18613), .ZN(n18352) );
  OAI211_X1 U21401 ( .C1(n18369), .C2(n18617), .A(n18353), .B(n18352), .ZN(
        P3_U2901) );
  AOI22_X1 U21402 ( .A1(n18389), .A2(n18620), .B1(n18364), .B2(n18618), .ZN(
        n18355) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18366), .B1(
        n18365), .B2(n18619), .ZN(n18354) );
  OAI211_X1 U21404 ( .C1(n18369), .C2(n18623), .A(n18355), .B(n18354), .ZN(
        P3_U2902) );
  AOI22_X1 U21405 ( .A1(n18365), .A2(n18626), .B1(n18364), .B2(n18624), .ZN(
        n18357) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18366), .B1(
        n18389), .B2(n18625), .ZN(n18356) );
  OAI211_X1 U21407 ( .C1(n18369), .C2(n18629), .A(n18357), .B(n18356), .ZN(
        P3_U2903) );
  AOI22_X1 U21408 ( .A1(n18389), .A2(n18630), .B1(n18364), .B2(n18631), .ZN(
        n18359) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18366), .B1(
        n18365), .B2(n18632), .ZN(n18358) );
  OAI211_X1 U21410 ( .C1(n18369), .C2(n18635), .A(n18359), .B(n18358), .ZN(
        P3_U2904) );
  AOI22_X1 U21411 ( .A1(n18365), .A2(n18637), .B1(n18364), .B2(n18636), .ZN(
        n18361) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18366), .B1(
        n18389), .B2(n18638), .ZN(n18360) );
  OAI211_X1 U21413 ( .C1(n18369), .C2(n18641), .A(n18361), .B(n18360), .ZN(
        P3_U2905) );
  AOI22_X1 U21414 ( .A1(n18389), .A2(n18644), .B1(n18364), .B2(n18642), .ZN(
        n18363) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18366), .B1(
        n18365), .B2(n18643), .ZN(n18362) );
  OAI211_X1 U21416 ( .C1(n18369), .C2(n18647), .A(n18363), .B(n18362), .ZN(
        P3_U2906) );
  AOI22_X1 U21417 ( .A1(n18365), .A2(n18653), .B1(n18364), .B2(n18649), .ZN(
        n18368) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18366), .B1(
        n18389), .B2(n18651), .ZN(n18367) );
  OAI211_X1 U21419 ( .C1(n18369), .C2(n18658), .A(n18368), .B(n18367), .ZN(
        P3_U2907) );
  INV_X1 U21420 ( .A(n18370), .ZN(n18461) );
  NAND2_X1 U21421 ( .A1(n18418), .A2(n18461), .ZN(n18393) );
  INV_X1 U21422 ( .A(n18371), .ZN(n18411) );
  INV_X1 U21423 ( .A(n18418), .ZN(n18372) );
  NOR2_X1 U21424 ( .A1(n18372), .A2(n18550), .ZN(n18388) );
  AOI22_X1 U21425 ( .A1(n18608), .A2(n18411), .B1(n18602), .B2(n18388), .ZN(
        n18375) );
  AOI22_X1 U21426 ( .A1(n18607), .A2(n18373), .B1(n18418), .B2(n18552), .ZN(
        n18390) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18390), .B1(
        n18389), .B2(n18603), .ZN(n18374) );
  OAI211_X1 U21428 ( .C1(n18611), .C2(n18393), .A(n18375), .B(n18374), .ZN(
        P3_U2908) );
  AOI22_X1 U21429 ( .A1(n18411), .A2(n18614), .B1(n18612), .B2(n18388), .ZN(
        n18377) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18390), .B1(
        n18389), .B2(n18613), .ZN(n18376) );
  OAI211_X1 U21431 ( .C1(n18617), .C2(n18393), .A(n18377), .B(n18376), .ZN(
        P3_U2909) );
  AOI22_X1 U21432 ( .A1(n18389), .A2(n18619), .B1(n18618), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18390), .B1(
        n18411), .B2(n18620), .ZN(n18378) );
  OAI211_X1 U21434 ( .C1(n18623), .C2(n18393), .A(n18379), .B(n18378), .ZN(
        P3_U2910) );
  AOI22_X1 U21435 ( .A1(n18411), .A2(n18625), .B1(n18624), .B2(n18388), .ZN(
        n18381) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18390), .B1(
        n18389), .B2(n18626), .ZN(n18380) );
  OAI211_X1 U21437 ( .C1(n18629), .C2(n18393), .A(n18381), .B(n18380), .ZN(
        P3_U2911) );
  AOI22_X1 U21438 ( .A1(n18389), .A2(n18632), .B1(n18631), .B2(n18388), .ZN(
        n18383) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18390), .B1(
        n18411), .B2(n18630), .ZN(n18382) );
  OAI211_X1 U21440 ( .C1(n18635), .C2(n18393), .A(n18383), .B(n18382), .ZN(
        P3_U2912) );
  AOI22_X1 U21441 ( .A1(n18389), .A2(n18637), .B1(n18636), .B2(n18388), .ZN(
        n18385) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18390), .B1(
        n18411), .B2(n18638), .ZN(n18384) );
  OAI211_X1 U21443 ( .C1(n18641), .C2(n18393), .A(n18385), .B(n18384), .ZN(
        P3_U2913) );
  AOI22_X1 U21444 ( .A1(n18411), .A2(n18644), .B1(n18642), .B2(n18388), .ZN(
        n18387) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18390), .B1(
        n18389), .B2(n18643), .ZN(n18386) );
  OAI211_X1 U21446 ( .C1(n18647), .C2(n18393), .A(n18387), .B(n18386), .ZN(
        P3_U2914) );
  AOI22_X1 U21447 ( .A1(n18389), .A2(n18653), .B1(n18649), .B2(n18388), .ZN(
        n18392) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18390), .B1(
        n18411), .B2(n18651), .ZN(n18391) );
  OAI211_X1 U21449 ( .C1(n18658), .C2(n18393), .A(n18392), .B(n18391), .ZN(
        P3_U2915) );
  INV_X1 U21450 ( .A(n18477), .ZN(n18415) );
  NOR2_X1 U21451 ( .A1(n18434), .A2(n18411), .ZN(n18394) );
  INV_X1 U21452 ( .A(n18393), .ZN(n18456) );
  NOR2_X1 U21453 ( .A1(n18456), .A2(n18477), .ZN(n18439) );
  OAI21_X1 U21454 ( .B1(n18394), .B2(n18576), .A(n18439), .ZN(n18395) );
  OAI211_X1 U21455 ( .C1(n18477), .C2(n18830), .A(n18579), .B(n18395), .ZN(
        n18412) );
  NOR2_X1 U21456 ( .A1(n18574), .A2(n18439), .ZN(n18410) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18412), .B1(
        n18602), .B2(n18410), .ZN(n18397) );
  AOI22_X1 U21458 ( .A1(n18608), .A2(n18434), .B1(n18411), .B2(n18603), .ZN(
        n18396) );
  OAI211_X1 U21459 ( .C1(n18611), .C2(n18415), .A(n18397), .B(n18396), .ZN(
        P3_U2916) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18412), .B1(
        n18612), .B2(n18410), .ZN(n18399) );
  AOI22_X1 U21461 ( .A1(n18434), .A2(n18614), .B1(n18411), .B2(n18613), .ZN(
        n18398) );
  OAI211_X1 U21462 ( .C1(n18617), .C2(n18415), .A(n18399), .B(n18398), .ZN(
        P3_U2917) );
  AOI22_X1 U21463 ( .A1(n18434), .A2(n18620), .B1(n18618), .B2(n18410), .ZN(
        n18401) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18412), .B1(
        n18411), .B2(n18619), .ZN(n18400) );
  OAI211_X1 U21465 ( .C1(n18623), .C2(n18415), .A(n18401), .B(n18400), .ZN(
        P3_U2918) );
  AOI22_X1 U21466 ( .A1(n18434), .A2(n18625), .B1(n18624), .B2(n18410), .ZN(
        n18403) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18412), .B1(
        n18411), .B2(n18626), .ZN(n18402) );
  OAI211_X1 U21468 ( .C1(n18629), .C2(n18415), .A(n18403), .B(n18402), .ZN(
        P3_U2919) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18412), .B1(
        n18631), .B2(n18410), .ZN(n18405) );
  AOI22_X1 U21470 ( .A1(n18434), .A2(n18630), .B1(n18411), .B2(n18632), .ZN(
        n18404) );
  OAI211_X1 U21471 ( .C1(n18635), .C2(n18415), .A(n18405), .B(n18404), .ZN(
        P3_U2920) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18412), .B1(
        n18636), .B2(n18410), .ZN(n18407) );
  AOI22_X1 U21473 ( .A1(n18434), .A2(n18638), .B1(n18411), .B2(n18637), .ZN(
        n18406) );
  OAI211_X1 U21474 ( .C1(n18641), .C2(n18415), .A(n18407), .B(n18406), .ZN(
        P3_U2921) );
  AOI22_X1 U21475 ( .A1(n18411), .A2(n18643), .B1(n18642), .B2(n18410), .ZN(
        n18409) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18412), .B1(
        n18434), .B2(n18644), .ZN(n18408) );
  OAI211_X1 U21477 ( .C1(n18647), .C2(n18415), .A(n18409), .B(n18408), .ZN(
        P3_U2922) );
  AOI22_X1 U21478 ( .A1(n18434), .A2(n18651), .B1(n18649), .B2(n18410), .ZN(
        n18414) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18412), .B1(
        n18411), .B2(n18653), .ZN(n18413) );
  OAI211_X1 U21480 ( .C1(n18658), .C2(n18415), .A(n18414), .B(n18413), .ZN(
        P3_U2923) );
  NAND2_X1 U21481 ( .A1(n18700), .A2(n18418), .ZN(n18438) );
  NOR2_X1 U21482 ( .A1(n18416), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18462) );
  AND2_X1 U21483 ( .A1(n18729), .A2(n18462), .ZN(n18433) );
  AOI22_X1 U21484 ( .A1(n18608), .A2(n18456), .B1(n18602), .B2(n18433), .ZN(
        n18420) );
  NAND2_X1 U21485 ( .A1(n18418), .A2(n18417), .ZN(n18435) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18603), .ZN(n18419) );
  OAI211_X1 U21487 ( .C1(n18611), .C2(n18438), .A(n18420), .B(n18419), .ZN(
        P3_U2924) );
  AOI22_X1 U21488 ( .A1(n18614), .A2(n18456), .B1(n18612), .B2(n18433), .ZN(
        n18422) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18613), .ZN(n18421) );
  OAI211_X1 U21490 ( .C1(n18617), .C2(n18438), .A(n18422), .B(n18421), .ZN(
        P3_U2925) );
  AOI22_X1 U21491 ( .A1(n18434), .A2(n18619), .B1(n18618), .B2(n18433), .ZN(
        n18424) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18435), .B1(
        n18620), .B2(n18456), .ZN(n18423) );
  OAI211_X1 U21493 ( .C1(n18623), .C2(n18438), .A(n18424), .B(n18423), .ZN(
        P3_U2926) );
  AOI22_X1 U21494 ( .A1(n18625), .A2(n18456), .B1(n18624), .B2(n18433), .ZN(
        n18426) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18626), .ZN(n18425) );
  OAI211_X1 U21496 ( .C1(n18629), .C2(n18438), .A(n18426), .B(n18425), .ZN(
        P3_U2927) );
  AOI22_X1 U21497 ( .A1(n18631), .A2(n18433), .B1(n18630), .B2(n18456), .ZN(
        n18428) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18632), .ZN(n18427) );
  OAI211_X1 U21499 ( .C1(n18635), .C2(n18438), .A(n18428), .B(n18427), .ZN(
        P3_U2928) );
  AOI22_X1 U21500 ( .A1(n18638), .A2(n18456), .B1(n18636), .B2(n18433), .ZN(
        n18430) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18637), .ZN(n18429) );
  OAI211_X1 U21502 ( .C1(n18641), .C2(n18438), .A(n18430), .B(n18429), .ZN(
        P3_U2929) );
  AOI22_X1 U21503 ( .A1(n18434), .A2(n18643), .B1(n18642), .B2(n18433), .ZN(
        n18432) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18435), .B1(
        n18644), .B2(n18456), .ZN(n18431) );
  OAI211_X1 U21505 ( .C1(n18647), .C2(n18438), .A(n18432), .B(n18431), .ZN(
        P3_U2930) );
  AOI22_X1 U21506 ( .A1(n18651), .A2(n18456), .B1(n18649), .B2(n18433), .ZN(
        n18437) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18435), .B1(
        n18434), .B2(n18653), .ZN(n18436) );
  OAI211_X1 U21508 ( .C1(n18658), .C2(n18438), .A(n18437), .B(n18436), .ZN(
        P3_U2931) );
  NAND2_X1 U21509 ( .A1(n18701), .A2(n18506), .ZN(n18460) );
  INV_X1 U21510 ( .A(n18438), .ZN(n18500) );
  INV_X1 U21511 ( .A(n18460), .ZN(n18522) );
  NOR2_X1 U21512 ( .A1(n18500), .A2(n18522), .ZN(n18484) );
  NOR2_X1 U21513 ( .A1(n18574), .A2(n18484), .ZN(n18455) );
  AOI22_X1 U21514 ( .A1(n18603), .A2(n18456), .B1(n18602), .B2(n18455), .ZN(
        n18442) );
  OAI21_X1 U21515 ( .B1(n18439), .B2(n18576), .A(n18484), .ZN(n18440) );
  OAI211_X1 U21516 ( .C1(n18522), .C2(n18830), .A(n18579), .B(n18440), .ZN(
        n18457) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18457), .B1(
        n18608), .B2(n18477), .ZN(n18441) );
  OAI211_X1 U21518 ( .C1(n18611), .C2(n18460), .A(n18442), .B(n18441), .ZN(
        P3_U2932) );
  AOI22_X1 U21519 ( .A1(n18614), .A2(n18477), .B1(n18612), .B2(n18455), .ZN(
        n18444) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18457), .B1(
        n18613), .B2(n18456), .ZN(n18443) );
  OAI211_X1 U21521 ( .C1(n18617), .C2(n18460), .A(n18444), .B(n18443), .ZN(
        P3_U2933) );
  AOI22_X1 U21522 ( .A1(n18619), .A2(n18456), .B1(n18618), .B2(n18455), .ZN(
        n18446) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18457), .B1(
        n18620), .B2(n18477), .ZN(n18445) );
  OAI211_X1 U21524 ( .C1(n18623), .C2(n18460), .A(n18446), .B(n18445), .ZN(
        P3_U2934) );
  AOI22_X1 U21525 ( .A1(n18626), .A2(n18456), .B1(n18624), .B2(n18455), .ZN(
        n18448) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18457), .B1(
        n18625), .B2(n18477), .ZN(n18447) );
  OAI211_X1 U21527 ( .C1(n18629), .C2(n18460), .A(n18448), .B(n18447), .ZN(
        P3_U2935) );
  AOI22_X1 U21528 ( .A1(n18632), .A2(n18456), .B1(n18631), .B2(n18455), .ZN(
        n18450) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18457), .B1(
        n18630), .B2(n18477), .ZN(n18449) );
  OAI211_X1 U21530 ( .C1(n18635), .C2(n18460), .A(n18450), .B(n18449), .ZN(
        P3_U2936) );
  AOI22_X1 U21531 ( .A1(n18638), .A2(n18477), .B1(n18636), .B2(n18455), .ZN(
        n18452) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18457), .B1(
        n18637), .B2(n18456), .ZN(n18451) );
  OAI211_X1 U21533 ( .C1(n18641), .C2(n18460), .A(n18452), .B(n18451), .ZN(
        P3_U2937) );
  AOI22_X1 U21534 ( .A1(n18643), .A2(n18456), .B1(n18642), .B2(n18455), .ZN(
        n18454) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18457), .B1(
        n18644), .B2(n18477), .ZN(n18453) );
  OAI211_X1 U21536 ( .C1(n18647), .C2(n18460), .A(n18454), .B(n18453), .ZN(
        P3_U2938) );
  AOI22_X1 U21537 ( .A1(n18651), .A2(n18477), .B1(n18649), .B2(n18455), .ZN(
        n18459) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18457), .B1(
        n18653), .B2(n18456), .ZN(n18458) );
  OAI211_X1 U21539 ( .C1(n18658), .C2(n18460), .A(n18459), .B(n18458), .ZN(
        P3_U2939) );
  NAND2_X1 U21540 ( .A1(n18461), .A2(n18506), .ZN(n18483) );
  INV_X1 U21541 ( .A(n18506), .ZN(n18481) );
  NOR2_X1 U21542 ( .A1(n18550), .A2(n18481), .ZN(n18507) );
  AOI22_X1 U21543 ( .A1(n18608), .A2(n18500), .B1(n18602), .B2(n18507), .ZN(
        n18464) );
  AOI22_X1 U21544 ( .A1(n18607), .A2(n18462), .B1(n18552), .B2(n18506), .ZN(
        n18478) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18478), .B1(
        n18603), .B2(n18477), .ZN(n18463) );
  OAI211_X1 U21546 ( .C1(n18611), .C2(n18483), .A(n18464), .B(n18463), .ZN(
        P3_U2940) );
  AOI22_X1 U21547 ( .A1(n18614), .A2(n18500), .B1(n18612), .B2(n18507), .ZN(
        n18466) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18478), .B1(
        n18613), .B2(n18477), .ZN(n18465) );
  OAI211_X1 U21549 ( .C1(n18617), .C2(n18483), .A(n18466), .B(n18465), .ZN(
        P3_U2941) );
  AOI22_X1 U21550 ( .A1(n18619), .A2(n18477), .B1(n18618), .B2(n18507), .ZN(
        n18468) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18478), .B1(
        n18620), .B2(n18500), .ZN(n18467) );
  OAI211_X1 U21552 ( .C1(n18623), .C2(n18483), .A(n18468), .B(n18467), .ZN(
        P3_U2942) );
  AOI22_X1 U21553 ( .A1(n18626), .A2(n18477), .B1(n18624), .B2(n18507), .ZN(
        n18470) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18478), .B1(
        n18625), .B2(n18500), .ZN(n18469) );
  OAI211_X1 U21555 ( .C1(n18629), .C2(n18483), .A(n18470), .B(n18469), .ZN(
        P3_U2943) );
  AOI22_X1 U21556 ( .A1(n18632), .A2(n18477), .B1(n18631), .B2(n18507), .ZN(
        n18472) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18478), .B1(
        n18630), .B2(n18500), .ZN(n18471) );
  OAI211_X1 U21558 ( .C1(n18635), .C2(n18483), .A(n18472), .B(n18471), .ZN(
        P3_U2944) );
  AOI22_X1 U21559 ( .A1(n18638), .A2(n18500), .B1(n18636), .B2(n18507), .ZN(
        n18474) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18478), .B1(
        n18637), .B2(n18477), .ZN(n18473) );
  OAI211_X1 U21561 ( .C1(n18641), .C2(n18483), .A(n18474), .B(n18473), .ZN(
        P3_U2945) );
  AOI22_X1 U21562 ( .A1(n18643), .A2(n18477), .B1(n18642), .B2(n18507), .ZN(
        n18476) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18478), .B1(
        n18644), .B2(n18500), .ZN(n18475) );
  OAI211_X1 U21564 ( .C1(n18647), .C2(n18483), .A(n18476), .B(n18475), .ZN(
        P3_U2946) );
  AOI22_X1 U21565 ( .A1(n18649), .A2(n18507), .B1(n18653), .B2(n18477), .ZN(
        n18480) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18478), .B1(
        n18651), .B2(n18500), .ZN(n18479) );
  OAI211_X1 U21567 ( .C1(n18658), .C2(n18483), .A(n18480), .B(n18479), .ZN(
        P3_U2947) );
  NOR2_X1 U21568 ( .A1(n20892), .A2(n18481), .ZN(n18554) );
  NAND2_X1 U21569 ( .A1(n18554), .A2(n18482), .ZN(n18505) );
  INV_X1 U21570 ( .A(n18483), .ZN(n18544) );
  INV_X1 U21571 ( .A(n18505), .ZN(n18569) );
  NOR2_X1 U21572 ( .A1(n18544), .A2(n18569), .ZN(n18528) );
  NOR2_X1 U21573 ( .A1(n18574), .A2(n18528), .ZN(n18501) );
  AOI22_X1 U21574 ( .A1(n18608), .A2(n18522), .B1(n18602), .B2(n18501), .ZN(
        n18487) );
  OAI21_X1 U21575 ( .B1(n18484), .B2(n18576), .A(n18528), .ZN(n18485) );
  OAI211_X1 U21576 ( .C1(n18569), .C2(n18830), .A(n18579), .B(n18485), .ZN(
        n18502) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18502), .B1(
        n18603), .B2(n18500), .ZN(n18486) );
  OAI211_X1 U21578 ( .C1(n18611), .C2(n18505), .A(n18487), .B(n18486), .ZN(
        P3_U2948) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18502), .B1(
        n18612), .B2(n18501), .ZN(n18489) );
  AOI22_X1 U21580 ( .A1(n18613), .A2(n18500), .B1(n18614), .B2(n18522), .ZN(
        n18488) );
  OAI211_X1 U21581 ( .C1(n18617), .C2(n18505), .A(n18489), .B(n18488), .ZN(
        P3_U2949) );
  AOI22_X1 U21582 ( .A1(n18620), .A2(n18522), .B1(n18618), .B2(n18501), .ZN(
        n18491) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18502), .B1(
        n18619), .B2(n18500), .ZN(n18490) );
  OAI211_X1 U21584 ( .C1(n18623), .C2(n18505), .A(n18491), .B(n18490), .ZN(
        P3_U2950) );
  AOI22_X1 U21585 ( .A1(n18626), .A2(n18500), .B1(n18624), .B2(n18501), .ZN(
        n18493) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18502), .B1(
        n18625), .B2(n18522), .ZN(n18492) );
  OAI211_X1 U21587 ( .C1(n18629), .C2(n18505), .A(n18493), .B(n18492), .ZN(
        P3_U2951) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18502), .B1(
        n18631), .B2(n18501), .ZN(n18495) );
  AOI22_X1 U21589 ( .A1(n18632), .A2(n18500), .B1(n18630), .B2(n18522), .ZN(
        n18494) );
  OAI211_X1 U21590 ( .C1(n18635), .C2(n18505), .A(n18495), .B(n18494), .ZN(
        P3_U2952) );
  AOI22_X1 U21591 ( .A1(n18637), .A2(n18500), .B1(n18636), .B2(n18501), .ZN(
        n18497) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18502), .B1(
        n18638), .B2(n18522), .ZN(n18496) );
  OAI211_X1 U21593 ( .C1(n18641), .C2(n18505), .A(n18497), .B(n18496), .ZN(
        P3_U2953) );
  AOI22_X1 U21594 ( .A1(n18642), .A2(n18501), .B1(n18644), .B2(n18522), .ZN(
        n18499) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18502), .B1(
        n18643), .B2(n18500), .ZN(n18498) );
  OAI211_X1 U21596 ( .C1(n18647), .C2(n18505), .A(n18499), .B(n18498), .ZN(
        P3_U2954) );
  AOI22_X1 U21597 ( .A1(n18649), .A2(n18501), .B1(n18653), .B2(n18500), .ZN(
        n18504) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18502), .B1(
        n18651), .B2(n18522), .ZN(n18503) );
  OAI211_X1 U21599 ( .C1(n18658), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2955) );
  NAND2_X1 U21600 ( .A1(n18700), .A2(n18506), .ZN(n18527) );
  AND2_X1 U21601 ( .A1(n18729), .A2(n18554), .ZN(n18523) );
  AOI22_X1 U21602 ( .A1(n18603), .A2(n18522), .B1(n18602), .B2(n18523), .ZN(
        n18509) );
  AOI22_X1 U21603 ( .A1(n18607), .A2(n18507), .B1(n18604), .B2(n18554), .ZN(
        n18524) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18524), .B1(
        n18608), .B2(n18544), .ZN(n18508) );
  OAI211_X1 U21605 ( .C1(n18611), .C2(n18527), .A(n18509), .B(n18508), .ZN(
        P3_U2956) );
  AOI22_X1 U21606 ( .A1(n18614), .A2(n18544), .B1(n18612), .B2(n18523), .ZN(
        n18511) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18524), .B1(
        n18613), .B2(n18522), .ZN(n18510) );
  OAI211_X1 U21608 ( .C1(n18617), .C2(n18527), .A(n18511), .B(n18510), .ZN(
        P3_U2957) );
  AOI22_X1 U21609 ( .A1(n18620), .A2(n18544), .B1(n18618), .B2(n18523), .ZN(
        n18513) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18524), .B1(
        n18619), .B2(n18522), .ZN(n18512) );
  OAI211_X1 U21611 ( .C1(n18623), .C2(n18527), .A(n18513), .B(n18512), .ZN(
        P3_U2958) );
  AOI22_X1 U21612 ( .A1(n18625), .A2(n18544), .B1(n18624), .B2(n18523), .ZN(
        n18515) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18524), .B1(
        n18626), .B2(n18522), .ZN(n18514) );
  OAI211_X1 U21614 ( .C1(n18629), .C2(n18527), .A(n18515), .B(n18514), .ZN(
        P3_U2959) );
  AOI22_X1 U21615 ( .A1(n18632), .A2(n18522), .B1(n18631), .B2(n18523), .ZN(
        n18517) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18524), .B1(
        n18630), .B2(n18544), .ZN(n18516) );
  OAI211_X1 U21617 ( .C1(n18635), .C2(n18527), .A(n18517), .B(n18516), .ZN(
        P3_U2960) );
  AOI22_X1 U21618 ( .A1(n18637), .A2(n18522), .B1(n18636), .B2(n18523), .ZN(
        n18519) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18524), .B1(
        n18638), .B2(n18544), .ZN(n18518) );
  OAI211_X1 U21620 ( .C1(n18641), .C2(n18527), .A(n18519), .B(n18518), .ZN(
        P3_U2961) );
  AOI22_X1 U21621 ( .A1(n18643), .A2(n18522), .B1(n18642), .B2(n18523), .ZN(
        n18521) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18524), .B1(
        n18644), .B2(n18544), .ZN(n18520) );
  OAI211_X1 U21623 ( .C1(n18647), .C2(n18527), .A(n18521), .B(n18520), .ZN(
        P3_U2962) );
  AOI22_X1 U21624 ( .A1(n18649), .A2(n18523), .B1(n18653), .B2(n18522), .ZN(
        n18526) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18524), .B1(
        n18651), .B2(n18544), .ZN(n18525) );
  OAI211_X1 U21626 ( .C1(n18658), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        P3_U2963) );
  INV_X1 U21627 ( .A(n18551), .ZN(n18553) );
  NAND2_X1 U21628 ( .A1(n18701), .A2(n18553), .ZN(n18549) );
  INV_X1 U21629 ( .A(n18527), .ZN(n18595) );
  INV_X1 U21630 ( .A(n18549), .ZN(n18652) );
  NOR2_X1 U21631 ( .A1(n18595), .A2(n18652), .ZN(n18577) );
  NOR2_X1 U21632 ( .A1(n18574), .A2(n18577), .ZN(n18545) );
  AOI22_X1 U21633 ( .A1(n18603), .A2(n18544), .B1(n18602), .B2(n18545), .ZN(
        n18531) );
  OAI21_X1 U21634 ( .B1(n18528), .B2(n18576), .A(n18577), .ZN(n18529) );
  OAI211_X1 U21635 ( .C1(n18652), .C2(n18830), .A(n18579), .B(n18529), .ZN(
        n18546) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18546), .B1(
        n18608), .B2(n18569), .ZN(n18530) );
  OAI211_X1 U21637 ( .C1(n18611), .C2(n18549), .A(n18531), .B(n18530), .ZN(
        P3_U2964) );
  AOI22_X1 U21638 ( .A1(n18614), .A2(n18569), .B1(n18612), .B2(n18545), .ZN(
        n18533) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18546), .B1(
        n18613), .B2(n18544), .ZN(n18532) );
  OAI211_X1 U21640 ( .C1(n18617), .C2(n18549), .A(n18533), .B(n18532), .ZN(
        P3_U2965) );
  AOI22_X1 U21641 ( .A1(n18619), .A2(n18544), .B1(n18618), .B2(n18545), .ZN(
        n18535) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18546), .B1(
        n18620), .B2(n18569), .ZN(n18534) );
  OAI211_X1 U21643 ( .C1(n18623), .C2(n18549), .A(n18535), .B(n18534), .ZN(
        P3_U2966) );
  AOI22_X1 U21644 ( .A1(n18625), .A2(n18569), .B1(n18624), .B2(n18545), .ZN(
        n18537) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18546), .B1(
        n18626), .B2(n18544), .ZN(n18536) );
  OAI211_X1 U21646 ( .C1(n18629), .C2(n18549), .A(n18537), .B(n18536), .ZN(
        P3_U2967) );
  AOI22_X1 U21647 ( .A1(n18632), .A2(n18544), .B1(n18631), .B2(n18545), .ZN(
        n18539) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18546), .B1(
        n18630), .B2(n18569), .ZN(n18538) );
  OAI211_X1 U21649 ( .C1(n18635), .C2(n18549), .A(n18539), .B(n18538), .ZN(
        P3_U2968) );
  AOI22_X1 U21650 ( .A1(n18637), .A2(n18544), .B1(n18636), .B2(n18545), .ZN(
        n18541) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18546), .B1(
        n18638), .B2(n18569), .ZN(n18540) );
  OAI211_X1 U21652 ( .C1(n18641), .C2(n18549), .A(n18541), .B(n18540), .ZN(
        P3_U2969) );
  AOI22_X1 U21653 ( .A1(n18643), .A2(n18544), .B1(n18642), .B2(n18545), .ZN(
        n18543) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18546), .B1(
        n18644), .B2(n18569), .ZN(n18542) );
  OAI211_X1 U21655 ( .C1(n18647), .C2(n18549), .A(n18543), .B(n18542), .ZN(
        P3_U2970) );
  AOI22_X1 U21656 ( .A1(n18649), .A2(n18545), .B1(n18653), .B2(n18544), .ZN(
        n18548) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18546), .B1(
        n18651), .B2(n18569), .ZN(n18547) );
  OAI211_X1 U21658 ( .C1(n18658), .C2(n18549), .A(n18548), .B(n18547), .ZN(
        P3_U2971) );
  INV_X1 U21659 ( .A(n18650), .ZN(n18573) );
  NOR2_X1 U21660 ( .A1(n18551), .A2(n18550), .ZN(n18606) );
  AOI22_X1 U21661 ( .A1(n18603), .A2(n18569), .B1(n18602), .B2(n18606), .ZN(
        n18556) );
  AOI22_X1 U21662 ( .A1(n18607), .A2(n18554), .B1(n18553), .B2(n18552), .ZN(
        n18570) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18570), .B1(
        n18608), .B2(n18595), .ZN(n18555) );
  OAI211_X1 U21664 ( .C1(n18611), .C2(n18573), .A(n18556), .B(n18555), .ZN(
        P3_U2972) );
  AOI22_X1 U21665 ( .A1(n18613), .A2(n18569), .B1(n18612), .B2(n18606), .ZN(
        n18558) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18570), .B1(
        n18614), .B2(n18595), .ZN(n18557) );
  OAI211_X1 U21667 ( .C1(n18617), .C2(n18573), .A(n18558), .B(n18557), .ZN(
        P3_U2973) );
  AOI22_X1 U21668 ( .A1(n18620), .A2(n18595), .B1(n18618), .B2(n18606), .ZN(
        n18560) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18570), .B1(
        n18619), .B2(n18569), .ZN(n18559) );
  OAI211_X1 U21670 ( .C1(n18623), .C2(n18573), .A(n18560), .B(n18559), .ZN(
        P3_U2974) );
  AOI22_X1 U21671 ( .A1(n18625), .A2(n18595), .B1(n18624), .B2(n18606), .ZN(
        n18562) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18570), .B1(
        n18626), .B2(n18569), .ZN(n18561) );
  OAI211_X1 U21673 ( .C1(n18629), .C2(n18573), .A(n18562), .B(n18561), .ZN(
        P3_U2975) );
  AOI22_X1 U21674 ( .A1(n18632), .A2(n18569), .B1(n18631), .B2(n18606), .ZN(
        n18564) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18570), .B1(
        n18630), .B2(n18595), .ZN(n18563) );
  OAI211_X1 U21676 ( .C1(n18635), .C2(n18573), .A(n18564), .B(n18563), .ZN(
        P3_U2976) );
  AOI22_X1 U21677 ( .A1(n18637), .A2(n18569), .B1(n18636), .B2(n18606), .ZN(
        n18566) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18570), .B1(
        n18638), .B2(n18595), .ZN(n18565) );
  OAI211_X1 U21679 ( .C1(n18641), .C2(n18573), .A(n18566), .B(n18565), .ZN(
        P3_U2977) );
  AOI22_X1 U21680 ( .A1(n18642), .A2(n18606), .B1(n18644), .B2(n18595), .ZN(
        n18568) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18570), .B1(
        n18643), .B2(n18569), .ZN(n18567) );
  OAI211_X1 U21682 ( .C1(n18647), .C2(n18573), .A(n18568), .B(n18567), .ZN(
        P3_U2978) );
  AOI22_X1 U21683 ( .A1(n18651), .A2(n18595), .B1(n18649), .B2(n18606), .ZN(
        n18572) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18570), .B1(
        n18653), .B2(n18569), .ZN(n18571) );
  OAI211_X1 U21685 ( .C1(n18658), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2979) );
  NOR2_X1 U21686 ( .A1(n18574), .A2(n18575), .ZN(n18596) );
  AOI22_X1 U21687 ( .A1(n18608), .A2(n18652), .B1(n18602), .B2(n18596), .ZN(
        n18582) );
  OAI21_X1 U21688 ( .B1(n18577), .B2(n18576), .A(n18575), .ZN(n18578) );
  OAI211_X1 U21689 ( .C1(n18580), .C2(n18830), .A(n18579), .B(n18578), .ZN(
        n18597) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18597), .B1(
        n18603), .B2(n18595), .ZN(n18581) );
  OAI211_X1 U21691 ( .C1(n18611), .C2(n18600), .A(n18582), .B(n18581), .ZN(
        P3_U2980) );
  AOI22_X1 U21692 ( .A1(n18613), .A2(n18595), .B1(n18612), .B2(n18596), .ZN(
        n18584) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18597), .B1(
        n18614), .B2(n18652), .ZN(n18583) );
  OAI211_X1 U21694 ( .C1(n18617), .C2(n18600), .A(n18584), .B(n18583), .ZN(
        P3_U2981) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18597), .B1(
        n18618), .B2(n18596), .ZN(n18586) );
  AOI22_X1 U21696 ( .A1(n18619), .A2(n18595), .B1(n18620), .B2(n18652), .ZN(
        n18585) );
  OAI211_X1 U21697 ( .C1(n18623), .C2(n18600), .A(n18586), .B(n18585), .ZN(
        P3_U2982) );
  AOI22_X1 U21698 ( .A1(n18625), .A2(n18652), .B1(n18624), .B2(n18596), .ZN(
        n18588) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18597), .B1(
        n18626), .B2(n18595), .ZN(n18587) );
  OAI211_X1 U21700 ( .C1(n18629), .C2(n18600), .A(n18588), .B(n18587), .ZN(
        P3_U2983) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18597), .B1(
        n18631), .B2(n18596), .ZN(n18590) );
  AOI22_X1 U21702 ( .A1(n18632), .A2(n18595), .B1(n18630), .B2(n18652), .ZN(
        n18589) );
  OAI211_X1 U21703 ( .C1(n18635), .C2(n18600), .A(n18590), .B(n18589), .ZN(
        P3_U2984) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18597), .B1(
        n18636), .B2(n18596), .ZN(n18592) );
  AOI22_X1 U21705 ( .A1(n18638), .A2(n18652), .B1(n18637), .B2(n18595), .ZN(
        n18591) );
  OAI211_X1 U21706 ( .C1(n18641), .C2(n18600), .A(n18592), .B(n18591), .ZN(
        P3_U2985) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18597), .B1(
        n18642), .B2(n18596), .ZN(n18594) );
  AOI22_X1 U21708 ( .A1(n18643), .A2(n18595), .B1(n18644), .B2(n18652), .ZN(
        n18593) );
  OAI211_X1 U21709 ( .C1(n18647), .C2(n18600), .A(n18594), .B(n18593), .ZN(
        P3_U2986) );
  AOI22_X1 U21710 ( .A1(n18649), .A2(n18596), .B1(n18653), .B2(n18595), .ZN(
        n18599) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18597), .B1(
        n18651), .B2(n18652), .ZN(n18598) );
  OAI211_X1 U21712 ( .C1(n18658), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        P3_U2987) );
  INV_X1 U21713 ( .A(n18601), .ZN(n18657) );
  AND2_X1 U21714 ( .A1(n18729), .A2(n18605), .ZN(n18648) );
  AOI22_X1 U21715 ( .A1(n18603), .A2(n18652), .B1(n18602), .B2(n18648), .ZN(
        n18610) );
  AOI22_X1 U21716 ( .A1(n18607), .A2(n18606), .B1(n18605), .B2(n18604), .ZN(
        n18654) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18654), .B1(
        n18608), .B2(n18650), .ZN(n18609) );
  OAI211_X1 U21718 ( .C1(n18611), .C2(n18657), .A(n18610), .B(n18609), .ZN(
        P3_U2988) );
  AOI22_X1 U21719 ( .A1(n18613), .A2(n18652), .B1(n18612), .B2(n18648), .ZN(
        n18616) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18654), .B1(
        n18614), .B2(n18650), .ZN(n18615) );
  OAI211_X1 U21721 ( .C1(n18617), .C2(n18657), .A(n18616), .B(n18615), .ZN(
        P3_U2989) );
  AOI22_X1 U21722 ( .A1(n18619), .A2(n18652), .B1(n18618), .B2(n18648), .ZN(
        n18622) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18654), .B1(
        n18620), .B2(n18650), .ZN(n18621) );
  OAI211_X1 U21724 ( .C1(n18623), .C2(n18657), .A(n18622), .B(n18621), .ZN(
        P3_U2990) );
  AOI22_X1 U21725 ( .A1(n18625), .A2(n18650), .B1(n18624), .B2(n18648), .ZN(
        n18628) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18654), .B1(
        n18626), .B2(n18652), .ZN(n18627) );
  OAI211_X1 U21727 ( .C1(n18629), .C2(n18657), .A(n18628), .B(n18627), .ZN(
        P3_U2991) );
  AOI22_X1 U21728 ( .A1(n18631), .A2(n18648), .B1(n18630), .B2(n18650), .ZN(
        n18634) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18654), .B1(
        n18632), .B2(n18652), .ZN(n18633) );
  OAI211_X1 U21730 ( .C1(n18635), .C2(n18657), .A(n18634), .B(n18633), .ZN(
        P3_U2992) );
  AOI22_X1 U21731 ( .A1(n18637), .A2(n18652), .B1(n18636), .B2(n18648), .ZN(
        n18640) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18654), .B1(
        n18638), .B2(n18650), .ZN(n18639) );
  OAI211_X1 U21733 ( .C1(n18641), .C2(n18657), .A(n18640), .B(n18639), .ZN(
        P3_U2993) );
  AOI22_X1 U21734 ( .A1(n18643), .A2(n18652), .B1(n18642), .B2(n18648), .ZN(
        n18646) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18654), .B1(
        n18644), .B2(n18650), .ZN(n18645) );
  OAI211_X1 U21736 ( .C1(n18647), .C2(n18657), .A(n18646), .B(n18645), .ZN(
        P3_U2994) );
  AOI22_X1 U21737 ( .A1(n18651), .A2(n18650), .B1(n18649), .B2(n18648), .ZN(
        n18656) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18654), .B1(
        n18653), .B2(n18652), .ZN(n18655) );
  OAI211_X1 U21739 ( .C1(n18658), .C2(n18657), .A(n18656), .B(n18655), .ZN(
        P3_U2995) );
  NOR2_X1 U21740 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18715) );
  INV_X1 U21741 ( .A(n18659), .ZN(n18673) );
  OAI21_X1 U21742 ( .B1(n18662), .B2(n18661), .A(n18660), .ZN(n18676) );
  OAI21_X1 U21743 ( .B1(n18674), .B2(n18676), .A(n18663), .ZN(n18664) );
  OAI221_X1 U21744 ( .B1(n18667), .B2(n18666), .C1(n18667), .C2(n18665), .A(
        n18664), .ZN(n18672) );
  INV_X1 U21745 ( .A(n18667), .ZN(n18669) );
  AOI21_X1 U21746 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18668), .A(
        n18699), .ZN(n18696) );
  OAI22_X1 U21747 ( .A1(n18673), .A2(n18670), .B1(n18669), .B2(n18696), .ZN(
        n18671) );
  OAI22_X1 U21748 ( .A1(n18673), .A2(n18672), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18671), .ZN(n18832) );
  INV_X1 U21749 ( .A(n18692), .ZN(n18702) );
  AOI22_X1 U21750 ( .A1(n18692), .A2(n18674), .B1(n18832), .B2(n18702), .ZN(
        n18714) );
  NOR2_X1 U21751 ( .A1(n18849), .A2(n18696), .ZN(n18679) );
  OAI221_X1 U21752 ( .B1(n18676), .B2(n18849), .C1(n18676), .C2(n18699), .A(
        n18675), .ZN(n18677) );
  INV_X1 U21753 ( .A(n18677), .ZN(n18678) );
  MUX2_X1 U21754 ( .A(n18679), .B(n18678), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n18680) );
  AOI21_X1 U21755 ( .B1(n18689), .B2(n18681), .A(n18680), .ZN(n18837) );
  AOI22_X1 U21756 ( .A1(n18692), .A2(n9714), .B1(n18837), .B2(n18702), .ZN(
        n18713) );
  OAI22_X1 U21757 ( .A1(n18685), .A2(n18684), .B1(n18683), .B2(n18682), .ZN(
        n18686) );
  AOI221_X1 U21758 ( .B1(n18689), .B2(n18688), .C1(n18687), .C2(n18688), .A(
        n18686), .ZN(n18870) );
  AOI211_X1 U21759 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18692), .A(
        n18691), .B(n18690), .ZN(n18711) );
  OAI21_X1 U21760 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18693), .ZN(n18710) );
  NAND2_X1 U21761 ( .A1(n18695), .A2(n18694), .ZN(n18698) );
  INV_X1 U21762 ( .A(n18696), .ZN(n18697) );
  AOI22_X1 U21763 ( .A1(n18846), .A2(n18698), .B1(n18697), .B2(n18849), .ZN(
        n18844) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18699), .B1(
        n18698), .B2(n12933), .ZN(n18851) );
  AOI222_X1 U21765 ( .A1(n18844), .A2(n18851), .B1(n18844), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18851), .C2(n18700), .ZN(
        n18703) );
  AOI21_X1 U21766 ( .B1(n18703), .B2(n18702), .A(n18701), .ZN(n18705) );
  INV_X1 U21767 ( .A(n18713), .ZN(n18704) );
  AOI222_X1 U21768 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18705), 
        .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18704), .C1(n18705), 
        .C2(n18704), .ZN(n18707) );
  OAI211_X1 U21769 ( .C1(n18708), .C2(n18714), .A(n18707), .B(n18706), .ZN(
        n18709) );
  NAND4_X1 U21770 ( .A1(n18870), .A2(n18711), .A3(n18710), .A4(n18709), .ZN(
        n18712) );
  AOI221_X1 U21771 ( .B1(n18715), .B2(n18714), .C1(n18713), .C2(n18714), .A(
        n18712), .ZN(n18726) );
  AOI22_X1 U21772 ( .A1(n9600), .A2(n18750), .B1(n18722), .B2(n18716), .ZN(
        n18717) );
  NOR2_X1 U21773 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18717), .ZN(n18724) );
  NOR2_X1 U21774 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18878), .ZN(n18727) );
  NAND2_X1 U21775 ( .A1(n18877), .A2(n18718), .ZN(n18719) );
  OAI211_X1 U21776 ( .C1(n18720), .C2(n18719), .A(n18873), .B(n18726), .ZN(
        n18730) );
  NAND2_X1 U21777 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18730), .ZN(n18828) );
  NOR4_X1 U21778 ( .A1(n18722), .A2(n18727), .A3(n18721), .A4(n18828), .ZN(
        n18723) );
  OAI22_X1 U21779 ( .A1(n18726), .A2(n18725), .B1(n18724), .B2(n18723), .ZN(
        P3_U2996) );
  NAND2_X1 U21780 ( .A1(n18750), .A2(n9600), .ZN(n18733) );
  NAND3_X1 U21781 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18727), .ZN(n18736) );
  INV_X1 U21782 ( .A(n18727), .ZN(n18728) );
  NAND4_X1 U21783 ( .A1(n18731), .A2(n18730), .A3(n18729), .A4(n18728), .ZN(
        n18732) );
  NAND4_X1 U21784 ( .A1(n18734), .A2(n18733), .A3(n18736), .A4(n18732), .ZN(
        P3_U2997) );
  OAI21_X1 U21785 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18735), .ZN(n18738) );
  INV_X1 U21786 ( .A(n18736), .ZN(n18737) );
  AOI21_X1 U21787 ( .B1(n18739), .B2(n18738), .A(n18737), .ZN(P3_U2998) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18824), .ZN(
        P3_U2999) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18824), .ZN(
        P3_U3000) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18824), .ZN(
        P3_U3001) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18824), .ZN(
        P3_U3002) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18824), .ZN(
        P3_U3003) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18824), .ZN(
        P3_U3004) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18824), .ZN(
        P3_U3005) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18824), .ZN(
        P3_U3006) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18824), .ZN(
        P3_U3007) );
  AND2_X1 U21797 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18824), .ZN(
        P3_U3008) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18824), .ZN(
        P3_U3009) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18824), .ZN(
        P3_U3010) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18824), .ZN(
        P3_U3011) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18824), .ZN(
        P3_U3012) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18824), .ZN(
        P3_U3013) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18824), .ZN(
        P3_U3014) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18824), .ZN(
        P3_U3015) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18824), .ZN(
        P3_U3016) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18824), .ZN(
        P3_U3017) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18824), .ZN(
        P3_U3018) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18824), .ZN(
        P3_U3019) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18824), .ZN(
        P3_U3020) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18824), .ZN(P3_U3021) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18824), .ZN(P3_U3022) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18824), .ZN(P3_U3023) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18824), .ZN(P3_U3024) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18824), .ZN(P3_U3025) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18824), .ZN(P3_U3026) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18824), .ZN(P3_U3027) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18824), .ZN(P3_U3028) );
  INV_X1 U21818 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18747) );
  AOI21_X1 U21819 ( .B1(HOLD), .B2(n18740), .A(n18747), .ZN(n18744) );
  AOI21_X1 U21820 ( .B1(n18750), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18741), 
        .ZN(n18755) );
  INV_X1 U21821 ( .A(NA), .ZN(n20646) );
  OAI21_X1 U21822 ( .B1(n20646), .B2(n18742), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18754) );
  INV_X1 U21823 ( .A(n18754), .ZN(n18743) );
  OAI22_X1 U21824 ( .A1(n18822), .A2(n18744), .B1(n18755), .B2(n18743), .ZN(
        P3_U3029) );
  NAND3_X1 U21825 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n18756), .ZN(
        n18745) );
  OAI221_X1 U21826 ( .B1(n18747), .B2(HOLD), .C1(n18747), .C2(n18746), .A(
        n18745), .ZN(n18748) );
  AOI22_X1 U21827 ( .A1(n18750), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18748), .ZN(n18749) );
  NAND2_X1 U21828 ( .A1(n18749), .A2(n18875), .ZN(P3_U3030) );
  NAND2_X1 U21829 ( .A1(n18750), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18751) );
  OAI222_X1 U21830 ( .A1(n18756), .A2(n19734), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18751), .C2(NA), .ZN(n18752)
         );
  OAI211_X1 U21831 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18752), .ZN(n18753) );
  OAI21_X1 U21832 ( .B1(n18755), .B2(n18754), .A(n18753), .ZN(P3_U3031) );
  INV_X1 U21833 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18758) );
  OAI222_X1 U21834 ( .A1(n18858), .A2(n18810), .B1(n18757), .B2(n18822), .C1(
        n18758), .C2(n18803), .ZN(P3_U3032) );
  OAI222_X1 U21835 ( .A1(n18803), .A2(n18760), .B1(n18759), .B2(n18822), .C1(
        n18758), .C2(n18810), .ZN(P3_U3033) );
  OAI222_X1 U21836 ( .A1(n18803), .A2(n18762), .B1(n18761), .B2(n18822), .C1(
        n18760), .C2(n18810), .ZN(P3_U3034) );
  INV_X1 U21837 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18765) );
  OAI222_X1 U21838 ( .A1(n18803), .A2(n18765), .B1(n18763), .B2(n18822), .C1(
        n18762), .C2(n18810), .ZN(P3_U3035) );
  OAI222_X1 U21839 ( .A1(n18765), .A2(n18810), .B1(n18764), .B2(n18822), .C1(
        n18766), .C2(n18803), .ZN(P3_U3036) );
  OAI222_X1 U21840 ( .A1(n18803), .A2(n18768), .B1(n18767), .B2(n18822), .C1(
        n18766), .C2(n18810), .ZN(P3_U3037) );
  OAI222_X1 U21841 ( .A1(n18803), .A2(n18770), .B1(n18769), .B2(n18822), .C1(
        n18768), .C2(n18810), .ZN(P3_U3038) );
  OAI222_X1 U21842 ( .A1(n18803), .A2(n18772), .B1(n18771), .B2(n18822), .C1(
        n18770), .C2(n18810), .ZN(P3_U3039) );
  OAI222_X1 U21843 ( .A1(n18803), .A2(n18774), .B1(n18773), .B2(n18822), .C1(
        n18772), .C2(n18810), .ZN(P3_U3040) );
  INV_X1 U21844 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18776) );
  OAI222_X1 U21845 ( .A1(n18803), .A2(n18776), .B1(n18775), .B2(n18822), .C1(
        n18774), .C2(n18810), .ZN(P3_U3041) );
  OAI222_X1 U21846 ( .A1(n18803), .A2(n18778), .B1(n18777), .B2(n18822), .C1(
        n18776), .C2(n18810), .ZN(P3_U3042) );
  OAI222_X1 U21847 ( .A1(n18803), .A2(n18780), .B1(n18779), .B2(n18822), .C1(
        n18778), .C2(n18810), .ZN(P3_U3043) );
  OAI222_X1 U21848 ( .A1(n18803), .A2(n18783), .B1(n18781), .B2(n18822), .C1(
        n18780), .C2(n18816), .ZN(P3_U3044) );
  OAI222_X1 U21849 ( .A1(n18783), .A2(n18810), .B1(n18782), .B2(n18822), .C1(
        n18784), .C2(n18803), .ZN(P3_U3045) );
  OAI222_X1 U21850 ( .A1(n18803), .A2(n18786), .B1(n18785), .B2(n18822), .C1(
        n18784), .C2(n18816), .ZN(P3_U3046) );
  OAI222_X1 U21851 ( .A1(n18803), .A2(n20801), .B1(n18787), .B2(n18822), .C1(
        n18786), .C2(n18816), .ZN(P3_U3047) );
  OAI222_X1 U21852 ( .A1(n18803), .A2(n18789), .B1(n18788), .B2(n18822), .C1(
        n20801), .C2(n18816), .ZN(P3_U3048) );
  OAI222_X1 U21853 ( .A1(n18803), .A2(n18791), .B1(n18790), .B2(n18822), .C1(
        n18789), .C2(n18816), .ZN(P3_U3049) );
  INV_X1 U21854 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18793) );
  OAI222_X1 U21855 ( .A1(n18803), .A2(n18793), .B1(n18792), .B2(n18822), .C1(
        n18791), .C2(n18816), .ZN(P3_U3050) );
  OAI222_X1 U21856 ( .A1(n18803), .A2(n18795), .B1(n18794), .B2(n18822), .C1(
        n18793), .C2(n18816), .ZN(P3_U3051) );
  OAI222_X1 U21857 ( .A1(n18795), .A2(n18810), .B1(n20846), .B2(n18822), .C1(
        n18796), .C2(n18803), .ZN(P3_U3052) );
  INV_X1 U21858 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18799) );
  OAI222_X1 U21859 ( .A1(n18803), .A2(n18799), .B1(n18797), .B2(n18822), .C1(
        n18796), .C2(n18816), .ZN(P3_U3053) );
  OAI222_X1 U21860 ( .A1(n18799), .A2(n18810), .B1(n18798), .B2(n18822), .C1(
        n18800), .C2(n18803), .ZN(P3_U3054) );
  OAI222_X1 U21861 ( .A1(n18803), .A2(n18802), .B1(n18801), .B2(n18822), .C1(
        n18800), .C2(n18816), .ZN(P3_U3055) );
  INV_X1 U21862 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18804) );
  OAI222_X1 U21863 ( .A1(n18803), .A2(n18804), .B1(n20877), .B2(n18822), .C1(
        n18802), .C2(n18810), .ZN(P3_U3056) );
  OAI222_X1 U21864 ( .A1(n18803), .A2(n18806), .B1(n18805), .B2(n18822), .C1(
        n18804), .C2(n18810), .ZN(P3_U3057) );
  OAI222_X1 U21865 ( .A1(n18803), .A2(n18809), .B1(n18807), .B2(n18822), .C1(
        n18806), .C2(n18810), .ZN(P3_U3058) );
  OAI222_X1 U21866 ( .A1(n18809), .A2(n18810), .B1(n18808), .B2(n18822), .C1(
        n18811), .C2(n18803), .ZN(P3_U3059) );
  OAI222_X1 U21867 ( .A1(n18803), .A2(n18815), .B1(n18812), .B2(n18822), .C1(
        n18811), .C2(n18810), .ZN(P3_U3060) );
  OAI222_X1 U21868 ( .A1(n18816), .A2(n18815), .B1(n18814), .B2(n18822), .C1(
        n18813), .C2(n18803), .ZN(P3_U3061) );
  INV_X1 U21869 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18817) );
  AOI22_X1 U21870 ( .A1(n18822), .A2(n18818), .B1(n18817), .B2(n18885), .ZN(
        P3_U3274) );
  INV_X1 U21871 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18860) );
  INV_X1 U21872 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18819) );
  AOI22_X1 U21873 ( .A1(n18822), .A2(n18860), .B1(n18819), .B2(n18885), .ZN(
        P3_U3275) );
  OAI22_X1 U21874 ( .A1(n18885), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18822), .ZN(n18820) );
  INV_X1 U21875 ( .A(n18820), .ZN(P3_U3276) );
  INV_X1 U21876 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18866) );
  INV_X1 U21877 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18821) );
  AOI22_X1 U21878 ( .A1(n18822), .A2(n18866), .B1(n18821), .B2(n18885), .ZN(
        P3_U3277) );
  INV_X1 U21879 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20885) );
  INV_X1 U21880 ( .A(n18825), .ZN(n18823) );
  AOI21_X1 U21881 ( .B1(n18824), .B2(n20885), .A(n18823), .ZN(P3_U3280) );
  OAI21_X1 U21882 ( .B1(n18827), .B2(n18826), .A(n18825), .ZN(P3_U3281) );
  INV_X1 U21883 ( .A(n18828), .ZN(n18831) );
  OAI21_X1 U21884 ( .B1(n18831), .B2(n18830), .A(n18829), .ZN(P3_U3282) );
  INV_X1 U21885 ( .A(n18847), .ZN(n18850) );
  OAI22_X1 U21886 ( .A1(n18833), .A2(n18850), .B1(n18852), .B2(n18832), .ZN(
        n18834) );
  INV_X1 U21887 ( .A(n18855), .ZN(n18857) );
  MUX2_X1 U21888 ( .A(n18834), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n18857), .Z(P3_U3285) );
  INV_X1 U21889 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18835) );
  AOI22_X1 U21890 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18836), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18835), .ZN(n18841) );
  NAND2_X1 U21891 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18842) );
  OAI22_X1 U21892 ( .A1(n18837), .A2(n18852), .B1(n18841), .B2(n18842), .ZN(
        n18838) );
  AOI21_X1 U21893 ( .B1(n18847), .B2(n18839), .A(n18838), .ZN(n18840) );
  AOI22_X1 U21894 ( .A1(n18857), .A2(n12935), .B1(n18840), .B2(n18855), .ZN(
        P3_U3288) );
  INV_X1 U21895 ( .A(n18841), .ZN(n18843) );
  OAI22_X1 U21896 ( .A1(n18844), .A2(n18852), .B1(n18843), .B2(n18842), .ZN(
        n18845) );
  AOI21_X1 U21897 ( .B1(n18847), .B2(n18846), .A(n18845), .ZN(n18848) );
  AOI22_X1 U21898 ( .A1(n18857), .A2(n18849), .B1(n18848), .B2(n18855), .ZN(
        P3_U3289) );
  OAI222_X1 U21899 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18851), .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(
        n18850), .ZN(n18854) );
  INV_X1 U21900 ( .A(n18854), .ZN(n18856) );
  AOI22_X1 U21901 ( .A1(n18857), .A2(n12933), .B1(n18856), .B2(n18855), .ZN(
        P3_U3290) );
  AOI21_X1 U21902 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18859) );
  AOI22_X1 U21903 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18859), .B2(n18858), .ZN(n18861) );
  AOI22_X1 U21904 ( .A1(n18862), .A2(n18861), .B1(n18860), .B2(n18865), .ZN(
        P3_U3292) );
  NOR2_X1 U21905 ( .A1(n18865), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18863) );
  AOI22_X1 U21906 ( .A1(n18866), .A2(n18865), .B1(n18864), .B2(n18863), .ZN(
        P3_U3293) );
  INV_X1 U21907 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18867) );
  AOI22_X1 U21908 ( .A1(n18822), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18867), 
        .B2(n18885), .ZN(P3_U3294) );
  INV_X1 U21909 ( .A(n18868), .ZN(n18871) );
  NAND2_X1 U21910 ( .A1(n18871), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18869) );
  OAI21_X1 U21911 ( .B1(n18871), .B2(n18870), .A(n18869), .ZN(P3_U3295) );
  NOR2_X1 U21912 ( .A1(n18873), .A2(n18872), .ZN(n18874) );
  AOI211_X1 U21913 ( .C1(n9600), .C2(n18878), .A(n18874), .B(n18890), .ZN(
        n18884) );
  AOI21_X1 U21914 ( .B1(n18877), .B2(n18876), .A(n18875), .ZN(n18879) );
  OAI211_X1 U21915 ( .C1(n18888), .C2(n18879), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18878), .ZN(n18881) );
  AOI21_X1 U21916 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18881), .A(n18880), 
        .ZN(n18883) );
  NAND2_X1 U21917 ( .A1(n18884), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18882) );
  OAI21_X1 U21918 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(P3_U3296) );
  INV_X1 U21919 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18893) );
  INV_X1 U21920 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18886) );
  AOI22_X1 U21921 ( .A1(n18822), .A2(n18893), .B1(n18886), .B2(n18885), .ZN(
        P3_U3297) );
  NOR2_X1 U21922 ( .A1(n18887), .A2(n18890), .ZN(n18894) );
  INV_X1 U21923 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18891) );
  INV_X1 U21924 ( .A(n18888), .ZN(n18889) );
  AOI22_X1 U21925 ( .A1(n18894), .A2(n18891), .B1(n18890), .B2(n18889), .ZN(
        P3_U3298) );
  AOI21_X1 U21926 ( .B1(n18894), .B2(n18893), .A(n18892), .ZN(P3_U3299) );
  INV_X1 U21927 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18895) );
  INV_X1 U21928 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19742) );
  NAND2_X1 U21929 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19742), .ZN(n19735) );
  OR2_X1 U21930 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19731) );
  OAI21_X1 U21931 ( .B1(n20893), .B2(n19735), .A(n19731), .ZN(n19793) );
  INV_X1 U21932 ( .A(n19793), .ZN(n19726) );
  OAI21_X1 U21933 ( .B1(n20893), .B2(n18895), .A(n19726), .ZN(P2_U2815) );
  AOI22_X1 U21934 ( .A1(n19867), .A2(n18896), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19864), .ZN(n18897) );
  OAI21_X1 U21935 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19736), .A(n18897), 
        .ZN(P2_U2817) );
  OAI21_X1 U21936 ( .B1(n19727), .B2(BS16), .A(n19793), .ZN(n19791) );
  OAI21_X1 U21937 ( .B1(n19793), .B2(n19847), .A(n19791), .ZN(P2_U2818) );
  NOR4_X1 U21938 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18907) );
  NOR4_X1 U21939 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18906) );
  NOR4_X1 U21940 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18898) );
  INV_X1 U21941 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20849) );
  INV_X1 U21942 ( .A(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19725) );
  NAND3_X1 U21943 ( .A1(n18898), .A2(n20849), .A3(n19725), .ZN(n18904) );
  NOR4_X1 U21944 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18902) );
  NOR4_X1 U21945 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n18901) );
  NOR4_X1 U21946 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18900) );
  NOR4_X1 U21947 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18899) );
  NAND4_X1 U21948 ( .A1(n18902), .A2(n18901), .A3(n18900), .A4(n18899), .ZN(
        n18903) );
  AOI211_X1 U21949 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18904), .B(n18903), .ZN(n18905) );
  NAND3_X1 U21950 ( .A1(n18907), .A2(n18906), .A3(n18905), .ZN(n18913) );
  NOR2_X1 U21951 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18913), .ZN(n18908) );
  INV_X1 U21952 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U21953 ( .A1(n18908), .A2(n10052), .B1(n18913), .B2(n19789), .ZN(
        P2_U2820) );
  OR3_X1 U21954 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18912) );
  INV_X1 U21955 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U21956 ( .A1(n18908), .A2(n18912), .B1(n18913), .B2(n19787), .ZN(
        P2_U2821) );
  INV_X1 U21957 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19792) );
  NAND2_X1 U21958 ( .A1(n18908), .A2(n19792), .ZN(n18911) );
  INV_X1 U21959 ( .A(n18913), .ZN(n18914) );
  OAI21_X1 U21960 ( .B1(n10037), .B2(n10052), .A(n18914), .ZN(n18909) );
  OAI21_X1 U21961 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18914), .A(n18909), 
        .ZN(n18910) );
  OAI221_X1 U21962 ( .B1(n18911), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18911), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18910), .ZN(P2_U2822) );
  INV_X1 U21963 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20784) );
  OAI221_X1 U21964 ( .B1(n18914), .B2(n20784), .C1(n18913), .C2(n18912), .A(
        n18911), .ZN(P2_U2823) );
  AOI211_X1 U21965 ( .C1(n18917), .C2(n18916), .A(n19724), .B(n18915), .ZN(
        n18924) );
  NOR2_X1 U21966 ( .A1(n18918), .A2(n19052), .ZN(n18923) );
  NOR2_X1 U21967 ( .A1(n18919), .A2(n19057), .ZN(n18922) );
  AOI22_X1 U21968 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19049), .ZN(n18920) );
  OAI211_X1 U21969 ( .C1(n19030), .C2(n19761), .A(n18920), .B(n18941), .ZN(
        n18921) );
  NOR4_X1 U21970 ( .A1(n18924), .A2(n18923), .A3(n18922), .A4(n18921), .ZN(
        n18925) );
  OAI21_X1 U21971 ( .B1(n18926), .B2(n19046), .A(n18925), .ZN(P2_U2836) );
  INV_X1 U21972 ( .A(n18933), .ZN(n18927) );
  NOR3_X1 U21973 ( .A1(n18927), .A2(n19724), .A3(n18936), .ZN(n18932) );
  OAI21_X1 U21974 ( .B1(n19030), .B2(n19759), .A(n18941), .ZN(n18928) );
  AOI21_X1 U21975 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19036), .A(
        n18928), .ZN(n18929) );
  OAI21_X1 U21976 ( .B1(n18930), .B2(n19052), .A(n18929), .ZN(n18931) );
  AOI211_X1 U21977 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19049), .A(n18932), .B(
        n18931), .ZN(n18938) );
  NOR2_X1 U21978 ( .A1(n19724), .A2(n18933), .ZN(n18949) );
  INV_X1 U21979 ( .A(n18934), .ZN(n18935) );
  AOI22_X1 U21980 ( .A1(n18949), .A2(n18936), .B1(n19041), .B2(n18935), .ZN(
        n18937) );
  OAI211_X1 U21981 ( .C1(n18939), .C2(n19046), .A(n18938), .B(n18937), .ZN(
        P2_U2837) );
  NOR2_X1 U21982 ( .A1(n19032), .A2(n10809), .ZN(n18944) );
  AOI22_X1 U21983 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n19048), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19036), .ZN(n18940) );
  OAI211_X1 U21984 ( .C1(n18942), .C2(n18950), .A(n18941), .B(n18940), .ZN(
        n18943) );
  AOI211_X1 U21985 ( .C1(n18945), .C2(n19041), .A(n18944), .B(n18943), .ZN(
        n18946) );
  OAI21_X1 U21986 ( .B1(n18947), .B2(n19052), .A(n18946), .ZN(n18948) );
  INV_X1 U21987 ( .A(n18948), .ZN(n18953) );
  OAI21_X1 U21988 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(n18952) );
  OAI211_X1 U21989 ( .C1(n19046), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        P2_U2838) );
  NOR2_X1 U21990 ( .A1(n12329), .A2(n18955), .ZN(n18957) );
  XOR2_X1 U21991 ( .A(n18957), .B(n18956), .Z(n18964) );
  OAI21_X1 U21992 ( .B1(n15513), .B2(n19030), .A(n18941), .ZN(n18960) );
  OAI22_X1 U21993 ( .A1(n18958), .A2(n19052), .B1(n10804), .B2(n19060), .ZN(
        n18959) );
  AOI211_X1 U21994 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19049), .A(n18960), .B(
        n18959), .ZN(n18963) );
  AOI22_X1 U21995 ( .A1(n18961), .A2(n19041), .B1(n19055), .B2(n19074), .ZN(
        n18962) );
  OAI211_X1 U21996 ( .C1(n19724), .C2(n18964), .A(n18963), .B(n18962), .ZN(
        P2_U2839) );
  OAI21_X1 U21997 ( .B1(n15326), .B2(n19030), .A(n18941), .ZN(n18968) );
  OAI22_X1 U21998 ( .A1(n18966), .A2(n19052), .B1(n19032), .B2(n18965), .ZN(
        n18967) );
  AOI211_X1 U21999 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19036), .A(
        n18968), .B(n18967), .ZN(n18975) );
  NAND2_X1 U22000 ( .A1(n12347), .A2(n18969), .ZN(n18970) );
  XNOR2_X1 U22001 ( .A(n18971), .B(n18970), .ZN(n18973) );
  AOI22_X1 U22002 ( .A1(n18973), .A2(n19042), .B1(n19041), .B2(n18972), .ZN(
        n18974) );
  OAI211_X1 U22003 ( .C1(n19080), .C2(n19046), .A(n18975), .B(n18974), .ZN(
        P2_U2840) );
  AOI22_X1 U22004 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19036), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19049), .ZN(n18976) );
  OAI21_X1 U22005 ( .B1(n18977), .B2(n19052), .A(n18976), .ZN(n18978) );
  AOI211_X1 U22006 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19048), .A(n19176), 
        .B(n18978), .ZN(n18985) );
  NOR2_X1 U22007 ( .A1(n12329), .A2(n18979), .ZN(n18981) );
  XNOR2_X1 U22008 ( .A(n18981), .B(n18980), .ZN(n18983) );
  AOI22_X1 U22009 ( .A1(n18983), .A2(n19042), .B1(n19041), .B2(n18982), .ZN(
        n18984) );
  OAI211_X1 U22010 ( .C1(n19089), .C2(n19046), .A(n18985), .B(n18984), .ZN(
        P2_U2843) );
  NAND2_X1 U22011 ( .A1(n13081), .A2(n18986), .ZN(n18988) );
  XOR2_X1 U22012 ( .A(n18988), .B(n18987), .Z(n18996) );
  AOI22_X1 U22013 ( .A1(n18989), .A2(n12367), .B1(P2_EBX_REG_11__SCAN_IN), 
        .B2(n19049), .ZN(n18990) );
  OAI211_X1 U22014 ( .C1(n10779), .C2(n19030), .A(n18990), .B(n10856), .ZN(
        n18994) );
  INV_X1 U22015 ( .A(n18991), .ZN(n18992) );
  OAI22_X1 U22016 ( .A1(n18992), .A2(n19057), .B1(n19046), .B2(n19091), .ZN(
        n18993) );
  AOI211_X1 U22017 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19036), .A(
        n18994), .B(n18993), .ZN(n18995) );
  OAI21_X1 U22018 ( .B1(n18996), .B2(n19724), .A(n18995), .ZN(P2_U2844) );
  NAND2_X1 U22019 ( .A1(n13081), .A2(n18997), .ZN(n18999) );
  XOR2_X1 U22020 ( .A(n18999), .B(n18998), .Z(n19006) );
  AOI22_X1 U22021 ( .A1(n19000), .A2(n12367), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19049), .ZN(n19001) );
  OAI211_X1 U22022 ( .C1(n10787), .C2(n19030), .A(n19001), .B(n10856), .ZN(
        n19004) );
  OAI22_X1 U22023 ( .A1(n19097), .A2(n19046), .B1(n19057), .B2(n19002), .ZN(
        n19003) );
  AOI211_X1 U22024 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19036), .A(
        n19004), .B(n19003), .ZN(n19005) );
  OAI21_X1 U22025 ( .B1(n19006), .B2(n19724), .A(n19005), .ZN(P2_U2846) );
  NAND2_X1 U22026 ( .A1(n12347), .A2(n19007), .ZN(n19009) );
  XOR2_X1 U22027 ( .A(n19009), .B(n19008), .Z(n19017) );
  INV_X1 U22028 ( .A(n19010), .ZN(n19011) );
  AOI22_X1 U22029 ( .A1(n19011), .A2(n12367), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19049), .ZN(n19012) );
  OAI211_X1 U22030 ( .C1(n10771), .C2(n19030), .A(n19012), .B(n10856), .ZN(
        n19015) );
  OAI22_X1 U22031 ( .A1(n19102), .A2(n19046), .B1(n19057), .B2(n19013), .ZN(
        n19014) );
  AOI211_X1 U22032 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19036), .A(
        n19015), .B(n19014), .ZN(n19016) );
  OAI21_X1 U22033 ( .B1(n19017), .B2(n19724), .A(n19016), .ZN(P2_U2848) );
  INV_X1 U22034 ( .A(n19018), .ZN(n19019) );
  AOI22_X1 U22035 ( .A1(n19019), .A2(n12367), .B1(P2_EBX_REG_6__SCAN_IN), .B2(
        n19049), .ZN(n19020) );
  OAI211_X1 U22036 ( .C1(n10767), .C2(n19030), .A(n10856), .B(n19020), .ZN(
        n19021) );
  INV_X1 U22037 ( .A(n19021), .ZN(n19029) );
  NOR2_X1 U22038 ( .A1(n12329), .A2(n19022), .ZN(n19023) );
  XNOR2_X1 U22039 ( .A(n19024), .B(n19023), .ZN(n19027) );
  OAI22_X1 U22040 ( .A1(n19104), .A2(n19046), .B1(n19057), .B2(n19025), .ZN(
        n19026) );
  AOI21_X1 U22041 ( .B1(n19027), .B2(n19042), .A(n19026), .ZN(n19028) );
  OAI211_X1 U22042 ( .C1(n9739), .C2(n19060), .A(n19029), .B(n19028), .ZN(
        P2_U2849) );
  OAI21_X1 U22043 ( .B1(n10761), .B2(n19030), .A(n18941), .ZN(n19035) );
  OAI22_X1 U22044 ( .A1(n19033), .A2(n19052), .B1(n19032), .B2(n19031), .ZN(
        n19034) );
  AOI211_X1 U22045 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19036), .A(
        n19035), .B(n19034), .ZN(n19045) );
  NAND2_X1 U22046 ( .A1(n12347), .A2(n19037), .ZN(n19038) );
  XNOR2_X1 U22047 ( .A(n19039), .B(n19038), .ZN(n19043) );
  AOI22_X1 U22048 ( .A1(n19043), .A2(n19042), .B1(n19041), .B2(n19040), .ZN(
        n19044) );
  OAI211_X1 U22049 ( .C1(n19046), .C2(n19113), .A(n19045), .B(n19044), .ZN(
        P2_U2850) );
  AOI22_X1 U22050 ( .A1(n19049), .A2(P2_EBX_REG_0__SCAN_IN), .B1(
        P2_REIP_REG_0__SCAN_IN), .B2(n19048), .ZN(n19050) );
  OAI21_X1 U22051 ( .B1(n19052), .B2(n19051), .A(n19050), .ZN(n19053) );
  AOI21_X1 U22052 ( .B1(n19055), .B2(n19054), .A(n19053), .ZN(n19056) );
  OAI21_X1 U22053 ( .B1(n19058), .B2(n19057), .A(n19056), .ZN(n19062) );
  NOR2_X1 U22054 ( .A1(n19060), .A2(n19059), .ZN(n19061) );
  AOI211_X1 U22055 ( .C1(n19064), .C2(n19063), .A(n19062), .B(n19061), .ZN(
        n19065) );
  OAI21_X1 U22056 ( .B1(n19724), .B2(n13791), .A(n19065), .ZN(P2_U2855) );
  INV_X1 U22057 ( .A(n19066), .ZN(n19067) );
  AOI22_X1 U22058 ( .A1(n19067), .A2(n19130), .B1(n19072), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19069) );
  AOI22_X1 U22059 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19129), .B1(n19073), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19068) );
  NAND2_X1 U22060 ( .A1(n19069), .A2(n19068), .ZN(P2_U2888) );
  AOI22_X1 U22061 ( .A1(n19071), .A2(n19070), .B1(n19129), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19078) );
  AOI22_X1 U22062 ( .A1(n19073), .A2(BUF1_REG_16__SCAN_IN), .B1(n19072), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19077) );
  AOI22_X1 U22063 ( .A1(n19075), .A2(n19108), .B1(n19130), .B2(n19074), .ZN(
        n19076) );
  NAND3_X1 U22064 ( .A1(n19078), .A2(n19077), .A3(n19076), .ZN(P2_U2903) );
  OAI222_X1 U22065 ( .A1(n19080), .A2(n19114), .B1(n19141), .B2(n19103), .C1(
        n19079), .C2(n19138), .ZN(P2_U2904) );
  INV_X1 U22066 ( .A(n19081), .ZN(n19084) );
  AOI22_X1 U22067 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19129), .B1(n19082), 
        .B2(n19105), .ZN(n19083) );
  OAI21_X1 U22068 ( .B1(n19114), .B2(n19084), .A(n19083), .ZN(P2_U2905) );
  INV_X1 U22069 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19145) );
  OAI222_X1 U22070 ( .A1(n19086), .A2(n19114), .B1(n19145), .B2(n19103), .C1(
        n19138), .C2(n19085), .ZN(P2_U2906) );
  AOI22_X1 U22071 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19129), .B1(n19087), 
        .B2(n19105), .ZN(n19088) );
  OAI21_X1 U22072 ( .B1(n19114), .B2(n19089), .A(n19088), .ZN(P2_U2907) );
  INV_X1 U22073 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19149) );
  OAI222_X1 U22074 ( .A1(n19091), .A2(n19114), .B1(n19149), .B2(n19103), .C1(
        n19138), .C2(n19090), .ZN(P2_U2908) );
  AOI22_X1 U22075 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19129), .B1(n19092), 
        .B2(n19105), .ZN(n19093) );
  OAI21_X1 U22076 ( .B1(n19114), .B2(n19094), .A(n19093), .ZN(P2_U2909) );
  AOI22_X1 U22077 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19129), .B1(n19095), .B2(
        n19105), .ZN(n19096) );
  OAI21_X1 U22078 ( .B1(n19114), .B2(n19097), .A(n19096), .ZN(P2_U2910) );
  INV_X1 U22079 ( .A(n19098), .ZN(n19101) );
  AOI22_X1 U22080 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19129), .B1(n19099), .B2(
        n19105), .ZN(n19100) );
  OAI21_X1 U22081 ( .B1(n19114), .B2(n19101), .A(n19100), .ZN(P2_U2911) );
  INV_X1 U22082 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19157) );
  OAI222_X1 U22083 ( .A1(n19102), .A2(n19114), .B1(n19157), .B2(n19103), .C1(
        n19138), .C2(n19232), .ZN(P2_U2912) );
  INV_X1 U22084 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19159) );
  OAI222_X1 U22085 ( .A1(n19104), .A2(n19114), .B1(n19159), .B2(n19103), .C1(
        n19138), .C2(n19225), .ZN(P2_U2913) );
  AOI22_X1 U22086 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19129), .B1(n19106), .B2(
        n19105), .ZN(n19112) );
  INV_X1 U22087 ( .A(n19107), .ZN(n19109) );
  NAND3_X1 U22088 ( .A1(n19110), .A2(n19109), .A3(n19108), .ZN(n19111) );
  OAI211_X1 U22089 ( .C1(n19114), .C2(n19113), .A(n19112), .B(n19111), .ZN(
        P2_U2914) );
  AOI22_X1 U22090 ( .A1(n19805), .A2(n19130), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19129), .ZN(n19120) );
  AOI21_X1 U22091 ( .B1(n19117), .B2(n19116), .A(n19115), .ZN(n19118) );
  OR2_X1 U22092 ( .A1(n19118), .A2(n19134), .ZN(n19119) );
  OAI211_X1 U22093 ( .C1(n19121), .C2(n19138), .A(n19120), .B(n19119), .ZN(
        P2_U2916) );
  AOI22_X1 U22094 ( .A1(n19809), .A2(n19130), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19129), .ZN(n19127) );
  AOI21_X1 U22095 ( .B1(n19124), .B2(n19123), .A(n19122), .ZN(n19125) );
  OR2_X1 U22096 ( .A1(n19125), .A2(n19134), .ZN(n19126) );
  OAI211_X1 U22097 ( .C1(n19128), .C2(n19138), .A(n19127), .B(n19126), .ZN(
        P2_U2917) );
  AOI22_X1 U22098 ( .A1(n19130), .A2(n19822), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19129), .ZN(n19137) );
  AOI21_X1 U22099 ( .B1(n19133), .B2(n19132), .A(n19131), .ZN(n19135) );
  OR2_X1 U22100 ( .A1(n19135), .A2(n19134), .ZN(n19136) );
  OAI211_X1 U22101 ( .C1(n19209), .C2(n19138), .A(n19137), .B(n19136), .ZN(
        P2_U2918) );
  AND2_X1 U22102 ( .A1(n19162), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22103 ( .A1(n19860), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22104 ( .B1(n19141), .B2(n19174), .A(n19140), .ZN(P2_U2936) );
  AOI22_X1 U22105 ( .A1(n19860), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22106 ( .B1(n19143), .B2(n19174), .A(n19142), .ZN(P2_U2937) );
  AOI22_X1 U22107 ( .A1(n19860), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22108 ( .B1(n19145), .B2(n19174), .A(n19144), .ZN(P2_U2938) );
  AOI22_X1 U22109 ( .A1(n19165), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U22110 ( .B1(n19147), .B2(n19174), .A(n19146), .ZN(P2_U2939) );
  AOI22_X1 U22111 ( .A1(n19165), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22112 ( .B1(n19149), .B2(n19174), .A(n19148), .ZN(P2_U2940) );
  AOI22_X1 U22113 ( .A1(n19165), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22114 ( .B1(n19151), .B2(n19174), .A(n19150), .ZN(P2_U2941) );
  AOI22_X1 U22115 ( .A1(n19165), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19152) );
  OAI21_X1 U22116 ( .B1(n19153), .B2(n19174), .A(n19152), .ZN(P2_U2942) );
  AOI22_X1 U22117 ( .A1(n19165), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19154) );
  OAI21_X1 U22118 ( .B1(n19155), .B2(n19174), .A(n19154), .ZN(P2_U2943) );
  AOI22_X1 U22119 ( .A1(n19165), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19156) );
  OAI21_X1 U22120 ( .B1(n19157), .B2(n19174), .A(n19156), .ZN(P2_U2944) );
  AOI22_X1 U22121 ( .A1(n19165), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22122 ( .B1(n19159), .B2(n19174), .A(n19158), .ZN(P2_U2945) );
  INV_X1 U22123 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19161) );
  AOI22_X1 U22124 ( .A1(n19165), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19160) );
  OAI21_X1 U22125 ( .B1(n19161), .B2(n19174), .A(n19160), .ZN(P2_U2946) );
  INV_X1 U22126 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22127 ( .A1(n19165), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19162), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U22128 ( .B1(n19164), .B2(n19174), .A(n19163), .ZN(P2_U2947) );
  INV_X1 U22129 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19167) );
  AOI22_X1 U22130 ( .A1(n19165), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19166) );
  OAI21_X1 U22131 ( .B1(n19167), .B2(n19174), .A(n19166), .ZN(P2_U2948) );
  INV_X1 U22132 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19169) );
  AOI22_X1 U22133 ( .A1(n19860), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19168) );
  OAI21_X1 U22134 ( .B1(n19169), .B2(n19174), .A(n19168), .ZN(P2_U2949) );
  INV_X1 U22135 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U22136 ( .A1(n19860), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19170) );
  OAI21_X1 U22137 ( .B1(n19171), .B2(n19174), .A(n19170), .ZN(P2_U2950) );
  INV_X1 U22138 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19175) );
  AOI22_X1 U22139 ( .A1(n19860), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19172), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19173) );
  OAI21_X1 U22140 ( .B1(n19175), .B2(n19174), .A(n19173), .ZN(P2_U2951) );
  AOI22_X1 U22141 ( .A1(n19177), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19176), .ZN(n19188) );
  NAND2_X1 U22142 ( .A1(n19179), .A2(n9578), .ZN(n19183) );
  NAND2_X1 U22143 ( .A1(n19181), .A2(n19180), .ZN(n19182) );
  OAI211_X1 U22144 ( .C1(n19185), .C2(n19184), .A(n19183), .B(n19182), .ZN(
        n19186) );
  INV_X1 U22145 ( .A(n19186), .ZN(n19187) );
  OAI211_X1 U22146 ( .C1(n19191), .C2(n19189), .A(n19188), .B(n19187), .ZN(
        P2_U3010) );
  NOR2_X1 U22147 ( .A1(n19191), .A2(n19190), .ZN(n19197) );
  OAI22_X1 U22148 ( .A1(n19195), .A2(n19194), .B1(n19193), .B2(n19192), .ZN(
        n19196) );
  AOI211_X1 U22149 ( .C1(n19198), .C2(n9595), .A(n19197), .B(n19196), .ZN(
        n19200) );
  OAI211_X1 U22150 ( .C1(n19202), .C2(n19201), .A(n19200), .B(n19199), .ZN(
        P2_U3012) );
  AOI22_X1 U22151 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19233), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19234), .ZN(n19571) );
  INV_X1 U22152 ( .A(n19571), .ZN(n19674) );
  AND2_X1 U22153 ( .A1(n19203), .A2(n19229), .ZN(n19673) );
  AOI22_X1 U22154 ( .A1(n19674), .A2(n19710), .B1(n19231), .B2(n19673), .ZN(
        n19207) );
  AOI22_X1 U22155 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19233), .ZN(n19642) );
  AOI22_X1 U22156 ( .A1(n19205), .A2(n19235), .B1(n19266), .B2(n19675), .ZN(
        n19206) );
  OAI211_X1 U22157 ( .C1(n19239), .C2(n19208), .A(n19207), .B(n19206), .ZN(
        P2_U3048) );
  AOI22_X1 U22158 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19233), .ZN(n19683) );
  NOR2_X2 U22159 ( .A1(n10566), .A2(n19220), .ZN(n19679) );
  AOI22_X1 U22160 ( .A1(n19710), .A2(n19643), .B1(n19231), .B2(n19679), .ZN(
        n19212) );
  AOI22_X1 U22161 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19233), .ZN(n19646) );
  INV_X1 U22162 ( .A(n19646), .ZN(n19680) );
  AOI22_X1 U22163 ( .A1(n19210), .A2(n19235), .B1(n19266), .B2(n19680), .ZN(
        n19211) );
  OAI211_X1 U22164 ( .C1(n19239), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        P2_U3049) );
  INV_X1 U22165 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20852) );
  AOI22_X1 U22166 ( .A1(n19710), .A2(n19648), .B1(n19647), .B2(n19231), .ZN(
        n19215) );
  AOI22_X1 U22167 ( .A1(n15716), .A2(n19235), .B1(n19266), .B2(n19574), .ZN(
        n19214) );
  OAI211_X1 U22168 ( .C1(n19239), .C2(n20852), .A(n19215), .B(n19214), .ZN(
        P2_U3050) );
  AOI22_X1 U22169 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19233), .ZN(n19689) );
  NOR2_X2 U22170 ( .A1(n9967), .A2(n19220), .ZN(n19684) );
  AOI22_X1 U22171 ( .A1(n19658), .A2(n19710), .B1(n19231), .B2(n19684), .ZN(
        n19218) );
  NOR2_X2 U22172 ( .A1(n19216), .A2(n19563), .ZN(n19685) );
  AOI22_X1 U22173 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19233), .ZN(n19661) );
  INV_X1 U22174 ( .A(n19661), .ZN(n19686) );
  AOI22_X1 U22175 ( .A1(n19685), .A2(n19235), .B1(n19266), .B2(n19686), .ZN(
        n19217) );
  OAI211_X1 U22176 ( .C1(n19239), .C2(n19219), .A(n19218), .B(n19217), .ZN(
        P2_U3052) );
  AOI22_X1 U22177 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19233), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19234), .ZN(n19695) );
  INV_X1 U22178 ( .A(n19695), .ZN(n19614) );
  NOR2_X2 U22179 ( .A1(n9585), .A2(n19220), .ZN(n19690) );
  AOI22_X1 U22180 ( .A1(n19614), .A2(n19710), .B1(n19231), .B2(n19690), .ZN(
        n19223) );
  NOR2_X2 U22181 ( .A1(n19221), .A2(n19563), .ZN(n19691) );
  AOI22_X1 U22182 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19233), .ZN(n19617) );
  AOI22_X1 U22183 ( .A1(n19691), .A2(n19235), .B1(n19266), .B2(n19692), .ZN(
        n19222) );
  OAI211_X1 U22184 ( .C1(n19239), .C2(n13580), .A(n19223), .B(n19222), .ZN(
        P2_U3053) );
  AOI22_X1 U22185 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19233), .ZN(n19666) );
  AND2_X1 U22186 ( .A1(n19224), .A2(n19229), .ZN(n19696) );
  AOI22_X1 U22187 ( .A1(n19699), .A2(n19710), .B1(n19231), .B2(n19696), .ZN(
        n19227) );
  NOR2_X2 U22188 ( .A1(n19225), .A2(n19563), .ZN(n19697) );
  AOI22_X1 U22189 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19233), .ZN(n19620) );
  AOI22_X1 U22190 ( .A1(n19697), .A2(n19235), .B1(n19266), .B2(n19698), .ZN(
        n19226) );
  OAI211_X1 U22191 ( .C1(n19239), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        P2_U3054) );
  INV_X1 U22192 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19238) );
  AOI22_X1 U22193 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19233), .ZN(n19715) );
  INV_X1 U22194 ( .A(n19715), .ZN(n19622) );
  AND2_X1 U22195 ( .A1(n19230), .A2(n19229), .ZN(n19705) );
  AOI22_X1 U22196 ( .A1(n19622), .A2(n19710), .B1(n19231), .B2(n19705), .ZN(
        n19237) );
  NOR2_X2 U22197 ( .A1(n19232), .A2(n19563), .ZN(n19707) );
  AOI22_X1 U22198 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19233), .ZN(n19627) );
  AOI22_X1 U22199 ( .A1(n19707), .A2(n19235), .B1(n19266), .B2(n19709), .ZN(
        n19236) );
  OAI211_X1 U22200 ( .C1(n19239), .C2(n19238), .A(n19237), .B(n19236), .ZN(
        P2_U3055) );
  NAND2_X1 U22201 ( .A1(n19272), .A2(n19824), .ZN(n19246) );
  NOR2_X1 U22202 ( .A1(n19833), .A2(n19246), .ZN(n19264) );
  NOR3_X1 U22203 ( .A1(n10281), .A2(n19264), .A3(n19852), .ZN(n19245) );
  INV_X1 U22204 ( .A(n19246), .ZN(n19241) );
  AOI21_X1 U22205 ( .B1(n19241), .B2(n19240), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19242) );
  NOR2_X1 U22206 ( .A1(n19245), .A2(n19242), .ZN(n19265) );
  AOI22_X1 U22207 ( .A1(n19265), .A2(n19205), .B1(n19673), .B2(n19264), .ZN(
        n19250) );
  INV_X1 U22208 ( .A(n19796), .ZN(n19244) );
  INV_X1 U22209 ( .A(n19471), .ZN(n19243) );
  NAND2_X1 U22210 ( .A1(n19244), .A2(n19243), .ZN(n19247) );
  AOI21_X1 U22211 ( .B1(n19247), .B2(n19246), .A(n19245), .ZN(n19248) );
  OAI211_X1 U22212 ( .C1(n19264), .C2(n19240), .A(n19248), .B(n19634), .ZN(
        n19267) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19674), .ZN(n19249) );
  OAI211_X1 U22214 ( .C1(n19642), .C2(n19299), .A(n19250), .B(n19249), .ZN(
        P2_U3056) );
  AOI22_X1 U22215 ( .A1(n19265), .A2(n19210), .B1(n19679), .B2(n19264), .ZN(
        n19252) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19643), .ZN(n19251) );
  OAI211_X1 U22217 ( .C1(n19646), .C2(n19299), .A(n19252), .B(n19251), .ZN(
        P2_U3057) );
  AOI22_X1 U22218 ( .A1(n19265), .A2(n15716), .B1(n19647), .B2(n19264), .ZN(
        n19254) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19648), .ZN(n19253) );
  OAI211_X1 U22220 ( .C1(n19651), .C2(n19299), .A(n19254), .B(n19253), .ZN(
        P2_U3058) );
  AOI22_X1 U22221 ( .A1(n19265), .A2(n15706), .B1(n19652), .B2(n19264), .ZN(
        n19257) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19608), .ZN(n19256) );
  OAI211_X1 U22223 ( .C1(n19611), .C2(n19299), .A(n19257), .B(n19256), .ZN(
        P2_U3059) );
  AOI22_X1 U22224 ( .A1(n19265), .A2(n19685), .B1(n19684), .B2(n19264), .ZN(
        n19259) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19658), .ZN(n19258) );
  OAI211_X1 U22226 ( .C1(n19661), .C2(n19299), .A(n19259), .B(n19258), .ZN(
        P2_U3060) );
  AOI22_X1 U22227 ( .A1(n19265), .A2(n19691), .B1(n19690), .B2(n19264), .ZN(
        n19261) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19614), .ZN(n19260) );
  OAI211_X1 U22229 ( .C1(n19617), .C2(n19299), .A(n19261), .B(n19260), .ZN(
        P2_U3061) );
  AOI22_X1 U22230 ( .A1(n19265), .A2(n19697), .B1(n19696), .B2(n19264), .ZN(
        n19263) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19699), .ZN(n19262) );
  OAI211_X1 U22232 ( .C1(n19620), .C2(n19299), .A(n19263), .B(n19262), .ZN(
        P2_U3062) );
  AOI22_X1 U22233 ( .A1(n19265), .A2(n19707), .B1(n19705), .B2(n19264), .ZN(
        n19269) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19267), .B1(
        n19266), .B2(n19622), .ZN(n19268) );
  OAI211_X1 U22235 ( .C1(n19627), .C2(n19299), .A(n19269), .B(n19268), .ZN(
        P2_U3063) );
  NAND2_X1 U22236 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19272), .ZN(
        n19308) );
  NOR2_X1 U22237 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19308), .ZN(
        n19294) );
  OAI21_X1 U22238 ( .B1(n19270), .B2(n19294), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19273) );
  INV_X1 U22239 ( .A(n19500), .ZN(n19271) );
  NAND2_X1 U22240 ( .A1(n19272), .A2(n19271), .ZN(n19275) );
  NAND2_X1 U22241 ( .A1(n19273), .A2(n19275), .ZN(n19295) );
  AOI22_X1 U22242 ( .A1(n19295), .A2(n19205), .B1(n19673), .B2(n19294), .ZN(
        n19280) );
  AOI21_X1 U22243 ( .B1(n19274), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19278) );
  OAI21_X1 U22244 ( .B1(n19326), .B2(n19287), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19276) );
  NAND3_X1 U22245 ( .A1(n19276), .A2(n19800), .A3(n19275), .ZN(n19277) );
  OAI211_X1 U22246 ( .C1(n19294), .C2(n19278), .A(n19277), .B(n19634), .ZN(
        n19296) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19296), .B1(
        n19326), .B2(n19675), .ZN(n19279) );
  OAI211_X1 U22248 ( .C1(n19571), .C2(n19299), .A(n19280), .B(n19279), .ZN(
        P2_U3064) );
  AOI22_X1 U22249 ( .A1(n19295), .A2(n19210), .B1(n19679), .B2(n19294), .ZN(
        n19282) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19296), .B1(
        n19287), .B2(n19643), .ZN(n19281) );
  OAI211_X1 U22251 ( .C1(n19646), .C2(n19318), .A(n19282), .B(n19281), .ZN(
        P2_U3065) );
  AOI22_X1 U22252 ( .A1(n19295), .A2(n15716), .B1(n19647), .B2(n19294), .ZN(
        n19284) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19296), .B1(
        n19287), .B2(n19648), .ZN(n19283) );
  OAI211_X1 U22254 ( .C1(n19651), .C2(n19318), .A(n19284), .B(n19283), .ZN(
        P2_U3066) );
  AOI22_X1 U22255 ( .A1(n19295), .A2(n15706), .B1(n19652), .B2(n19294), .ZN(
        n19286) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19296), .B1(
        n19326), .B2(n19653), .ZN(n19285) );
  OAI211_X1 U22257 ( .C1(n19656), .C2(n19299), .A(n19286), .B(n19285), .ZN(
        P2_U3067) );
  AOI22_X1 U22258 ( .A1(n19295), .A2(n19685), .B1(n19684), .B2(n19294), .ZN(
        n19289) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19296), .B1(
        n19287), .B2(n19658), .ZN(n19288) );
  OAI211_X1 U22260 ( .C1(n19661), .C2(n19318), .A(n19289), .B(n19288), .ZN(
        P2_U3068) );
  AOI22_X1 U22261 ( .A1(n19295), .A2(n19691), .B1(n19690), .B2(n19294), .ZN(
        n19291) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19296), .B1(
        n19326), .B2(n19692), .ZN(n19290) );
  OAI211_X1 U22263 ( .C1(n19695), .C2(n19299), .A(n19291), .B(n19290), .ZN(
        P2_U3069) );
  AOI22_X1 U22264 ( .A1(n19295), .A2(n19697), .B1(n19696), .B2(n19294), .ZN(
        n19293) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19296), .B1(
        n19326), .B2(n19698), .ZN(n19292) );
  OAI211_X1 U22266 ( .C1(n19666), .C2(n19299), .A(n19293), .B(n19292), .ZN(
        P2_U3070) );
  AOI22_X1 U22267 ( .A1(n19295), .A2(n19707), .B1(n19705), .B2(n19294), .ZN(
        n19298) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19296), .B1(
        n19326), .B2(n19709), .ZN(n19297) );
  OAI211_X1 U22269 ( .C1(n19715), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P2_U3071) );
  NOR2_X1 U22270 ( .A1(n19301), .A2(n19300), .ZN(n19325) );
  AOI22_X1 U22271 ( .A1(n19675), .A2(n19348), .B1(n19325), .B2(n19673), .ZN(
        n19311) );
  OAI21_X1 U22272 ( .B1(n19796), .B2(n19797), .A(n19800), .ZN(n19309) );
  INV_X1 U22273 ( .A(n19308), .ZN(n19305) );
  INV_X1 U22274 ( .A(n19325), .ZN(n19302) );
  OAI211_X1 U22275 ( .C1(n19303), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19795), 
        .B(n19302), .ZN(n19304) );
  OAI211_X1 U22276 ( .C1(n19309), .C2(n19305), .A(n19634), .B(n19304), .ZN(
        n19328) );
  OAI21_X1 U22277 ( .B1(n19306), .B2(n19325), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19307) );
  OAI21_X1 U22278 ( .B1(n19309), .B2(n19308), .A(n19307), .ZN(n19327) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19328), .B1(
        n19205), .B2(n19327), .ZN(n19310) );
  OAI211_X1 U22280 ( .C1(n19571), .C2(n19318), .A(n19311), .B(n19310), .ZN(
        P2_U3072) );
  AOI22_X1 U22281 ( .A1(n19680), .A2(n19348), .B1(n19325), .B2(n19679), .ZN(
        n19313) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19328), .B1(
        n19210), .B2(n19327), .ZN(n19312) );
  OAI211_X1 U22283 ( .C1(n19683), .C2(n19318), .A(n19313), .B(n19312), .ZN(
        P2_U3073) );
  AOI22_X1 U22284 ( .A1(n19648), .A2(n19326), .B1(n19647), .B2(n19325), .ZN(
        n19315) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19328), .B1(
        n15716), .B2(n19327), .ZN(n19314) );
  OAI211_X1 U22286 ( .C1(n19651), .C2(n19360), .A(n19315), .B(n19314), .ZN(
        P2_U3074) );
  AOI22_X1 U22287 ( .A1(n19653), .A2(n19348), .B1(n19652), .B2(n19325), .ZN(
        n19317) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19328), .B1(
        n15706), .B2(n19327), .ZN(n19316) );
  OAI211_X1 U22289 ( .C1(n19656), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P2_U3075) );
  AOI22_X1 U22290 ( .A1(n19658), .A2(n19326), .B1(n19325), .B2(n19684), .ZN(
        n19320) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19328), .B1(
        n19685), .B2(n19327), .ZN(n19319) );
  OAI211_X1 U22292 ( .C1(n19661), .C2(n19360), .A(n19320), .B(n19319), .ZN(
        P2_U3076) );
  AOI22_X1 U22293 ( .A1(n19614), .A2(n19326), .B1(n19325), .B2(n19690), .ZN(
        n19322) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19328), .B1(
        n19691), .B2(n19327), .ZN(n19321) );
  OAI211_X1 U22295 ( .C1(n19617), .C2(n19360), .A(n19322), .B(n19321), .ZN(
        P2_U3077) );
  AOI22_X1 U22296 ( .A1(n19699), .A2(n19326), .B1(n19325), .B2(n19696), .ZN(
        n19324) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19328), .B1(
        n19697), .B2(n19327), .ZN(n19323) );
  OAI211_X1 U22298 ( .C1(n19620), .C2(n19360), .A(n19324), .B(n19323), .ZN(
        P2_U3078) );
  AOI22_X1 U22299 ( .A1(n19622), .A2(n19326), .B1(n19325), .B2(n19705), .ZN(
        n19330) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19328), .B1(
        n19707), .B2(n19327), .ZN(n19329) );
  OAI211_X1 U22301 ( .C1(n19627), .C2(n19360), .A(n19330), .B(n19329), .ZN(
        P2_U3079) );
  INV_X1 U22302 ( .A(n19331), .ZN(n19395) );
  AND2_X1 U22303 ( .A1(n19395), .A2(n19332), .ZN(n19567) );
  NAND2_X1 U22304 ( .A1(n19567), .A2(n19807), .ZN(n19337) );
  NOR2_X1 U22305 ( .A1(n19396), .A2(n19441), .ZN(n19355) );
  OAI21_X1 U22306 ( .B1(n10290), .B2(n19355), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19333) );
  OAI21_X1 U22307 ( .B1(n19337), .B2(n19795), .A(n19333), .ZN(n19356) );
  AOI22_X1 U22308 ( .A1(n19356), .A2(n19205), .B1(n19673), .B2(n19355), .ZN(
        n19341) );
  AOI21_X1 U22309 ( .B1(n19334), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19339) );
  OAI21_X1 U22310 ( .B1(n19348), .B2(n19386), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19336) );
  AOI21_X1 U22311 ( .B1(n19337), .B2(n19336), .A(n19563), .ZN(n19338) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19357), .B1(
        n19386), .B2(n19675), .ZN(n19340) );
  OAI211_X1 U22313 ( .C1(n19571), .C2(n19360), .A(n19341), .B(n19340), .ZN(
        P2_U3080) );
  AOI22_X1 U22314 ( .A1(n19356), .A2(n19210), .B1(n19679), .B2(n19355), .ZN(
        n19343) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19357), .B1(
        n19348), .B2(n19643), .ZN(n19342) );
  OAI211_X1 U22316 ( .C1(n19646), .C2(n19384), .A(n19343), .B(n19342), .ZN(
        P2_U3081) );
  AOI22_X1 U22317 ( .A1(n19356), .A2(n15716), .B1(n19647), .B2(n19355), .ZN(
        n19345) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19357), .B1(
        n19348), .B2(n19648), .ZN(n19344) );
  OAI211_X1 U22319 ( .C1(n19651), .C2(n19384), .A(n19345), .B(n19344), .ZN(
        P2_U3082) );
  AOI22_X1 U22320 ( .A1(n19356), .A2(n15706), .B1(n19652), .B2(n19355), .ZN(
        n19347) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19357), .B1(
        n19386), .B2(n19653), .ZN(n19346) );
  OAI211_X1 U22322 ( .C1(n19656), .C2(n19360), .A(n19347), .B(n19346), .ZN(
        P2_U3083) );
  AOI22_X1 U22323 ( .A1(n19356), .A2(n19685), .B1(n19684), .B2(n19355), .ZN(
        n19350) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19357), .B1(
        n19348), .B2(n19658), .ZN(n19349) );
  OAI211_X1 U22325 ( .C1(n19661), .C2(n19384), .A(n19350), .B(n19349), .ZN(
        P2_U3084) );
  AOI22_X1 U22326 ( .A1(n19356), .A2(n19691), .B1(n19690), .B2(n19355), .ZN(
        n19352) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19357), .B1(
        n19386), .B2(n19692), .ZN(n19351) );
  OAI211_X1 U22328 ( .C1(n19695), .C2(n19360), .A(n19352), .B(n19351), .ZN(
        P2_U3085) );
  AOI22_X1 U22329 ( .A1(n19356), .A2(n19697), .B1(n19696), .B2(n19355), .ZN(
        n19354) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19357), .B1(
        n19386), .B2(n19698), .ZN(n19353) );
  OAI211_X1 U22331 ( .C1(n19666), .C2(n19360), .A(n19354), .B(n19353), .ZN(
        P2_U3086) );
  AOI22_X1 U22332 ( .A1(n19356), .A2(n19707), .B1(n19705), .B2(n19355), .ZN(
        n19359) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19357), .B1(
        n19386), .B2(n19709), .ZN(n19358) );
  OAI211_X1 U22334 ( .C1(n19715), .C2(n19360), .A(n19359), .B(n19358), .ZN(
        P2_U3087) );
  NOR3_X2 U22335 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19833), .A3(
        n19396), .ZN(n19385) );
  AOI22_X1 U22336 ( .A1(n19675), .A2(n19393), .B1(n19673), .B2(n19385), .ZN(
        n19371) );
  OAI21_X1 U22337 ( .B1(n19796), .B2(n19596), .A(n19800), .ZN(n19369) );
  NOR2_X1 U22338 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19396), .ZN(
        n19365) );
  OAI21_X1 U22339 ( .B1(n19366), .B2(n19852), .A(n19240), .ZN(n19363) );
  INV_X1 U22340 ( .A(n19385), .ZN(n19362) );
  AOI21_X1 U22341 ( .B1(n19363), .B2(n19362), .A(n19563), .ZN(n19364) );
  OAI21_X1 U22342 ( .B1(n19369), .B2(n19365), .A(n19364), .ZN(n19388) );
  INV_X1 U22343 ( .A(n19365), .ZN(n19368) );
  OAI21_X1 U22344 ( .B1(n19366), .B2(n19385), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19367) );
  OAI21_X1 U22345 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n19387) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19388), .B1(
        n19205), .B2(n19387), .ZN(n19370) );
  OAI211_X1 U22347 ( .C1(n19571), .C2(n19384), .A(n19371), .B(n19370), .ZN(
        P2_U3088) );
  AOI22_X1 U22348 ( .A1(n19643), .A2(n19386), .B1(n19679), .B2(n19385), .ZN(
        n19373) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19388), .B1(
        n19210), .B2(n19387), .ZN(n19372) );
  OAI211_X1 U22350 ( .C1(n19646), .C2(n19420), .A(n19373), .B(n19372), .ZN(
        P2_U3089) );
  AOI22_X1 U22351 ( .A1(n19574), .A2(n19393), .B1(n19647), .B2(n19385), .ZN(
        n19375) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19388), .B1(
        n15716), .B2(n19387), .ZN(n19374) );
  OAI211_X1 U22353 ( .C1(n19577), .C2(n19384), .A(n19375), .B(n19374), .ZN(
        P2_U3090) );
  AOI22_X1 U22354 ( .A1(n19653), .A2(n19393), .B1(n19652), .B2(n19385), .ZN(
        n19377) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19388), .B1(
        n15706), .B2(n19387), .ZN(n19376) );
  OAI211_X1 U22356 ( .C1(n19656), .C2(n19384), .A(n19377), .B(n19376), .ZN(
        P2_U3091) );
  AOI22_X1 U22357 ( .A1(n19686), .A2(n19393), .B1(n19385), .B2(n19684), .ZN(
        n19379) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19388), .B1(
        n19685), .B2(n19387), .ZN(n19378) );
  OAI211_X1 U22359 ( .C1(n19689), .C2(n19384), .A(n19379), .B(n19378), .ZN(
        P2_U3092) );
  AOI22_X1 U22360 ( .A1(n19692), .A2(n19393), .B1(n19385), .B2(n19690), .ZN(
        n19381) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19388), .B1(
        n19691), .B2(n19387), .ZN(n19380) );
  OAI211_X1 U22362 ( .C1(n19695), .C2(n19384), .A(n19381), .B(n19380), .ZN(
        P2_U3093) );
  AOI22_X1 U22363 ( .A1(n19698), .A2(n19393), .B1(n19385), .B2(n19696), .ZN(
        n19383) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19388), .B1(
        n19697), .B2(n19387), .ZN(n19382) );
  OAI211_X1 U22365 ( .C1(n19666), .C2(n19384), .A(n19383), .B(n19382), .ZN(
        P2_U3094) );
  AOI22_X1 U22366 ( .A1(n19622), .A2(n19386), .B1(n19385), .B2(n19705), .ZN(
        n19390) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19388), .B1(
        n19707), .B2(n19387), .ZN(n19389) );
  OAI211_X1 U22368 ( .C1(n19627), .C2(n19420), .A(n19390), .B(n19389), .ZN(
        P2_U3095) );
  NOR2_X1 U22369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19391), .ZN(
        n19415) );
  OAI21_X1 U22370 ( .B1(n10283), .B2(n19415), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19392) );
  OAI21_X1 U22371 ( .B1(n19396), .B2(n19500), .A(n19392), .ZN(n19416) );
  AOI22_X1 U22372 ( .A1(n19416), .A2(n19205), .B1(n19673), .B2(n19415), .ZN(
        n19402) );
  OAI21_X1 U22373 ( .B1(n19393), .B2(n19437), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19394) );
  OAI21_X1 U22374 ( .B1(n19396), .B2(n19395), .A(n19394), .ZN(n19400) );
  INV_X1 U22375 ( .A(n19415), .ZN(n19397) );
  OAI211_X1 U22376 ( .C1(n19398), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19397), 
        .B(n19795), .ZN(n19399) );
  NAND3_X1 U22377 ( .A1(n19400), .A2(n19634), .A3(n19399), .ZN(n19417) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19675), .ZN(n19401) );
  OAI211_X1 U22379 ( .C1(n19571), .C2(n19420), .A(n19402), .B(n19401), .ZN(
        P2_U3096) );
  AOI22_X1 U22380 ( .A1(n19416), .A2(n19210), .B1(n19679), .B2(n19415), .ZN(
        n19404) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19680), .ZN(n19403) );
  OAI211_X1 U22382 ( .C1(n19683), .C2(n19420), .A(n19404), .B(n19403), .ZN(
        P2_U3097) );
  AOI22_X1 U22383 ( .A1(n19416), .A2(n15716), .B1(n19647), .B2(n19415), .ZN(
        n19406) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19574), .ZN(n19405) );
  OAI211_X1 U22385 ( .C1(n19577), .C2(n19420), .A(n19406), .B(n19405), .ZN(
        P2_U3098) );
  AOI22_X1 U22386 ( .A1(n19416), .A2(n15706), .B1(n19652), .B2(n19415), .ZN(
        n19408) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19653), .ZN(n19407) );
  OAI211_X1 U22388 ( .C1(n19656), .C2(n19420), .A(n19408), .B(n19407), .ZN(
        P2_U3099) );
  AOI22_X1 U22389 ( .A1(n19416), .A2(n19685), .B1(n19684), .B2(n19415), .ZN(
        n19410) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19686), .ZN(n19409) );
  OAI211_X1 U22391 ( .C1(n19689), .C2(n19420), .A(n19410), .B(n19409), .ZN(
        P2_U3100) );
  AOI22_X1 U22392 ( .A1(n19416), .A2(n19691), .B1(n19690), .B2(n19415), .ZN(
        n19412) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19692), .ZN(n19411) );
  OAI211_X1 U22394 ( .C1(n19695), .C2(n19420), .A(n19412), .B(n19411), .ZN(
        P2_U3101) );
  AOI22_X1 U22395 ( .A1(n19416), .A2(n19697), .B1(n19696), .B2(n19415), .ZN(
        n19414) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19698), .ZN(n19413) );
  OAI211_X1 U22397 ( .C1(n19666), .C2(n19420), .A(n19414), .B(n19413), .ZN(
        P2_U3102) );
  AOI22_X1 U22398 ( .A1(n19416), .A2(n19707), .B1(n19705), .B2(n19415), .ZN(
        n19419) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19417), .B1(
        n19437), .B2(n19709), .ZN(n19418) );
  OAI211_X1 U22400 ( .C1(n19715), .C2(n19420), .A(n19419), .B(n19418), .ZN(
        P2_U3103) );
  INV_X1 U22401 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19423) );
  AOI22_X1 U22402 ( .A1(n19436), .A2(n19205), .B1(n19446), .B2(n19673), .ZN(
        n19422) );
  AOI22_X1 U22403 ( .A1(n19462), .A2(n19675), .B1(n19437), .B2(n19674), .ZN(
        n19421) );
  OAI211_X1 U22404 ( .C1(n19435), .C2(n19423), .A(n19422), .B(n19421), .ZN(
        P2_U3104) );
  INV_X1 U22405 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n19426) );
  AOI22_X1 U22406 ( .A1(n19436), .A2(n19210), .B1(n19446), .B2(n19679), .ZN(
        n19425) );
  AOI22_X1 U22407 ( .A1(n19462), .A2(n19680), .B1(n19437), .B2(n19643), .ZN(
        n19424) );
  OAI211_X1 U22408 ( .C1(n19435), .C2(n19426), .A(n19425), .B(n19424), .ZN(
        P2_U3105) );
  AOI22_X1 U22409 ( .A1(n19436), .A2(n15706), .B1(n19446), .B2(n19652), .ZN(
        n19428) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19608), .ZN(n19427) );
  OAI211_X1 U22411 ( .C1(n19611), .C2(n19470), .A(n19428), .B(n19427), .ZN(
        P2_U3107) );
  AOI22_X1 U22412 ( .A1(n19436), .A2(n19685), .B1(n19446), .B2(n19684), .ZN(
        n19430) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19658), .ZN(n19429) );
  OAI211_X1 U22414 ( .C1(n19661), .C2(n19470), .A(n19430), .B(n19429), .ZN(
        P2_U3108) );
  AOI22_X1 U22415 ( .A1(n19436), .A2(n19691), .B1(n19446), .B2(n19690), .ZN(
        n19432) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19614), .ZN(n19431) );
  OAI211_X1 U22417 ( .C1(n19617), .C2(n19470), .A(n19432), .B(n19431), .ZN(
        P2_U3109) );
  AOI22_X1 U22418 ( .A1(n19436), .A2(n19697), .B1(n19446), .B2(n19696), .ZN(
        n19434) );
  AOI22_X1 U22419 ( .A1(n19462), .A2(n19698), .B1(n19437), .B2(n19699), .ZN(
        n19433) );
  OAI211_X1 U22420 ( .C1(n19435), .C2(n20788), .A(n19434), .B(n19433), .ZN(
        P2_U3110) );
  AOI22_X1 U22421 ( .A1(n19436), .A2(n19707), .B1(n19446), .B2(n19705), .ZN(
        n19440) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19438), .B1(
        n19437), .B2(n19622), .ZN(n19439) );
  OAI211_X1 U22423 ( .C1(n19627), .C2(n19470), .A(n19440), .B(n19439), .ZN(
        P2_U3111) );
  NAND2_X1 U22424 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12395), .ZN(
        n19534) );
  NOR2_X1 U22425 ( .A1(n19441), .A2(n19534), .ZN(n19465) );
  AOI22_X1 U22426 ( .A1(n19491), .A2(n19675), .B1(n19673), .B2(n19465), .ZN(
        n19451) );
  NOR3_X1 U22427 ( .A1(n19491), .A2(n19462), .A3(n19795), .ZN(n19442) );
  NOR2_X1 U22428 ( .A1(n19442), .A2(n19798), .ZN(n19449) );
  NOR2_X1 U22429 ( .A1(n19449), .A2(n19446), .ZN(n19443) );
  AOI211_X1 U22430 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19444), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19443), .ZN(n19445) );
  NOR2_X1 U22431 ( .A1(n19446), .A2(n19465), .ZN(n19448) );
  OAI21_X1 U22432 ( .B1(n10181), .B2(n19465), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19447) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19467), .B1(
        n19205), .B2(n19466), .ZN(n19450) );
  OAI211_X1 U22434 ( .C1(n19571), .C2(n19470), .A(n19451), .B(n19450), .ZN(
        P2_U3112) );
  AOI22_X1 U22435 ( .A1(n19643), .A2(n19462), .B1(n19679), .B2(n19465), .ZN(
        n19453) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n19210), .ZN(n19452) );
  OAI211_X1 U22437 ( .C1(n19646), .C2(n19498), .A(n19453), .B(n19452), .ZN(
        P2_U3113) );
  AOI22_X1 U22438 ( .A1(n19648), .A2(n19462), .B1(n19647), .B2(n19465), .ZN(
        n19455) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n15716), .ZN(n19454) );
  OAI211_X1 U22440 ( .C1(n19651), .C2(n19498), .A(n19455), .B(n19454), .ZN(
        P2_U3114) );
  AOI22_X1 U22441 ( .A1(n19491), .A2(n19653), .B1(n19652), .B2(n19465), .ZN(
        n19457) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n15706), .ZN(n19456) );
  OAI211_X1 U22443 ( .C1(n19656), .C2(n19470), .A(n19457), .B(n19456), .ZN(
        P2_U3115) );
  AOI22_X1 U22444 ( .A1(n19686), .A2(n19491), .B1(n19684), .B2(n19465), .ZN(
        n19459) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n19685), .ZN(n19458) );
  OAI211_X1 U22446 ( .C1(n19689), .C2(n19470), .A(n19459), .B(n19458), .ZN(
        P2_U3116) );
  AOI22_X1 U22447 ( .A1(n19692), .A2(n19491), .B1(n19690), .B2(n19465), .ZN(
        n19461) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n19691), .ZN(n19460) );
  OAI211_X1 U22449 ( .C1(n19695), .C2(n19470), .A(n19461), .B(n19460), .ZN(
        P2_U3117) );
  AOI22_X1 U22450 ( .A1(n19699), .A2(n19462), .B1(n19696), .B2(n19465), .ZN(
        n19464) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n19697), .ZN(n19463) );
  OAI211_X1 U22452 ( .C1(n19620), .C2(n19498), .A(n19464), .B(n19463), .ZN(
        P2_U3118) );
  AOI22_X1 U22453 ( .A1(n19709), .A2(n19491), .B1(n19705), .B2(n19465), .ZN(
        n19469) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19467), .B1(
        n19466), .B2(n19707), .ZN(n19468) );
  OAI211_X1 U22455 ( .C1(n19715), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3119) );
  NOR3_X2 U22456 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19833), .A3(
        n19534), .ZN(n19501) );
  AOI22_X1 U22457 ( .A1(n19517), .A2(n19675), .B1(n19673), .B2(n19501), .ZN(
        n19480) );
  OAI21_X1 U22458 ( .B1(n19597), .B2(n19471), .A(n19800), .ZN(n19478) );
  NOR2_X1 U22459 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19534), .ZN(
        n19475) );
  INV_X1 U22460 ( .A(n10289), .ZN(n19473) );
  INV_X1 U22461 ( .A(n19501), .ZN(n19472) );
  OAI211_X1 U22462 ( .C1(n19473), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19795), 
        .B(n19472), .ZN(n19474) );
  OAI211_X1 U22463 ( .C1(n19478), .C2(n19475), .A(n19634), .B(n19474), .ZN(
        n19495) );
  INV_X1 U22464 ( .A(n19475), .ZN(n19477) );
  OAI21_X1 U22465 ( .B1(n10289), .B2(n19501), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19476) );
  OAI21_X1 U22466 ( .B1(n19478), .B2(n19477), .A(n19476), .ZN(n19494) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19495), .B1(
        n19205), .B2(n19494), .ZN(n19479) );
  OAI211_X1 U22468 ( .C1(n19571), .C2(n19498), .A(n19480), .B(n19479), .ZN(
        P2_U3120) );
  AOI22_X1 U22469 ( .A1(n19491), .A2(n19643), .B1(n19679), .B2(n19501), .ZN(
        n19482) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19495), .B1(
        n19210), .B2(n19494), .ZN(n19481) );
  OAI211_X1 U22471 ( .C1(n19646), .C2(n19526), .A(n19482), .B(n19481), .ZN(
        P2_U3121) );
  AOI22_X1 U22472 ( .A1(n19574), .A2(n19517), .B1(n19647), .B2(n19501), .ZN(
        n19484) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19495), .B1(
        n15716), .B2(n19494), .ZN(n19483) );
  OAI211_X1 U22474 ( .C1(n19577), .C2(n19498), .A(n19484), .B(n19483), .ZN(
        P2_U3122) );
  AOI22_X1 U22475 ( .A1(n19608), .A2(n19491), .B1(n19652), .B2(n19501), .ZN(
        n19486) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19495), .B1(
        n15706), .B2(n19494), .ZN(n19485) );
  OAI211_X1 U22477 ( .C1(n19611), .C2(n19526), .A(n19486), .B(n19485), .ZN(
        P2_U3123) );
  AOI22_X1 U22478 ( .A1(n19658), .A2(n19491), .B1(n19684), .B2(n19501), .ZN(
        n19488) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19495), .B1(
        n19685), .B2(n19494), .ZN(n19487) );
  OAI211_X1 U22480 ( .C1(n19661), .C2(n19526), .A(n19488), .B(n19487), .ZN(
        P2_U3124) );
  AOI22_X1 U22481 ( .A1(n19614), .A2(n19491), .B1(n19690), .B2(n19501), .ZN(
        n19490) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19495), .B1(
        n19691), .B2(n19494), .ZN(n19489) );
  OAI211_X1 U22483 ( .C1(n19617), .C2(n19526), .A(n19490), .B(n19489), .ZN(
        P2_U3125) );
  AOI22_X1 U22484 ( .A1(n19699), .A2(n19491), .B1(n19696), .B2(n19501), .ZN(
        n19493) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19495), .B1(
        n19697), .B2(n19494), .ZN(n19492) );
  OAI211_X1 U22486 ( .C1(n19620), .C2(n19526), .A(n19493), .B(n19492), .ZN(
        P2_U3126) );
  AOI22_X1 U22487 ( .A1(n19709), .A2(n19517), .B1(n19705), .B2(n19501), .ZN(
        n19497) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19495), .B1(
        n19707), .B2(n19494), .ZN(n19496) );
  OAI211_X1 U22489 ( .C1(n19715), .C2(n19498), .A(n19497), .B(n19496), .ZN(
        P2_U3127) );
  NOR3_X2 U22490 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19824), .A3(
        n19534), .ZN(n19521) );
  OAI21_X1 U22491 ( .B1(n10288), .B2(n19521), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19499) );
  OAI21_X1 U22492 ( .B1(n19534), .B2(n19500), .A(n19499), .ZN(n19522) );
  AOI22_X1 U22493 ( .A1(n19522), .A2(n19205), .B1(n19673), .B2(n19521), .ZN(
        n19506) );
  AOI221_X1 U22494 ( .B1(n19554), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19517), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19501), .ZN(n19502) );
  AOI211_X1 U22495 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19503), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19502), .ZN(n19504) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19523), .B1(
        n19554), .B2(n19675), .ZN(n19505) );
  OAI211_X1 U22497 ( .C1(n19571), .C2(n19526), .A(n19506), .B(n19505), .ZN(
        P2_U3128) );
  INV_X1 U22498 ( .A(n19554), .ZN(n19520) );
  AOI22_X1 U22499 ( .A1(n19522), .A2(n19210), .B1(n19679), .B2(n19521), .ZN(
        n19508) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19523), .B1(
        n19517), .B2(n19643), .ZN(n19507) );
  OAI211_X1 U22501 ( .C1(n19646), .C2(n19520), .A(n19508), .B(n19507), .ZN(
        P2_U3129) );
  AOI22_X1 U22502 ( .A1(n19522), .A2(n15716), .B1(n19647), .B2(n19521), .ZN(
        n19510) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19523), .B1(
        n19517), .B2(n19648), .ZN(n19509) );
  OAI211_X1 U22504 ( .C1(n19651), .C2(n19520), .A(n19510), .B(n19509), .ZN(
        P2_U3130) );
  AOI22_X1 U22505 ( .A1(n19522), .A2(n15706), .B1(n19652), .B2(n19521), .ZN(
        n19512) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19523), .B1(
        n19554), .B2(n19653), .ZN(n19511) );
  OAI211_X1 U22507 ( .C1(n19656), .C2(n19526), .A(n19512), .B(n19511), .ZN(
        P2_U3131) );
  AOI22_X1 U22508 ( .A1(n19522), .A2(n19685), .B1(n19684), .B2(n19521), .ZN(
        n19514) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19523), .B1(
        n19554), .B2(n19686), .ZN(n19513) );
  OAI211_X1 U22510 ( .C1(n19689), .C2(n19526), .A(n19514), .B(n19513), .ZN(
        P2_U3132) );
  AOI22_X1 U22511 ( .A1(n19522), .A2(n19691), .B1(n19690), .B2(n19521), .ZN(
        n19516) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19523), .B1(
        n19554), .B2(n19692), .ZN(n19515) );
  OAI211_X1 U22513 ( .C1(n19695), .C2(n19526), .A(n19516), .B(n19515), .ZN(
        P2_U3133) );
  AOI22_X1 U22514 ( .A1(n19522), .A2(n19697), .B1(n19696), .B2(n19521), .ZN(
        n19519) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19523), .B1(
        n19517), .B2(n19699), .ZN(n19518) );
  OAI211_X1 U22516 ( .C1(n19620), .C2(n19520), .A(n19519), .B(n19518), .ZN(
        P2_U3134) );
  AOI22_X1 U22517 ( .A1(n19522), .A2(n19707), .B1(n19705), .B2(n19521), .ZN(
        n19525) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19523), .B1(
        n19554), .B2(n19709), .ZN(n19524) );
  OAI211_X1 U22519 ( .C1(n19715), .C2(n19526), .A(n19525), .B(n19524), .ZN(
        P2_U3135) );
  INV_X1 U22520 ( .A(n19527), .ZN(n19530) );
  INV_X1 U22521 ( .A(n19534), .ZN(n19528) );
  NAND2_X1 U22522 ( .A1(n19529), .A2(n19528), .ZN(n19533) );
  NAND3_X1 U22523 ( .A1(n19530), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19533), 
        .ZN(n19535) );
  OR2_X1 U22524 ( .A1(n19824), .A2(n19534), .ZN(n19531) );
  OAI21_X1 U22525 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19531), .A(n19852), 
        .ZN(n19532) );
  AND2_X1 U22526 ( .A1(n19535), .A2(n19532), .ZN(n19553) );
  INV_X1 U22527 ( .A(n19533), .ZN(n19552) );
  AOI22_X1 U22528 ( .A1(n19553), .A2(n19205), .B1(n19552), .B2(n19673), .ZN(
        n19539) );
  NOR3_X1 U22529 ( .A1(n19597), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19797), 
        .ZN(n19537) );
  AOI211_X1 U22530 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19833), .A(n19824), 
        .B(n19534), .ZN(n19536) );
  OAI211_X1 U22531 ( .C1(n19537), .C2(n19536), .A(n19634), .B(n19535), .ZN(
        n19555) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19674), .ZN(n19538) );
  OAI211_X1 U22533 ( .C1(n19642), .C2(n19591), .A(n19539), .B(n19538), .ZN(
        P2_U3136) );
  AOI22_X1 U22534 ( .A1(n19553), .A2(n19210), .B1(n19552), .B2(n19679), .ZN(
        n19541) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19643), .ZN(n19540) );
  OAI211_X1 U22536 ( .C1(n19646), .C2(n19591), .A(n19541), .B(n19540), .ZN(
        P2_U3137) );
  AOI22_X1 U22537 ( .A1(n19553), .A2(n15716), .B1(n19647), .B2(n19552), .ZN(
        n19543) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19648), .ZN(n19542) );
  OAI211_X1 U22539 ( .C1(n19651), .C2(n19591), .A(n19543), .B(n19542), .ZN(
        P2_U3138) );
  AOI22_X1 U22540 ( .A1(n19553), .A2(n15706), .B1(n19652), .B2(n19552), .ZN(
        n19545) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19608), .ZN(n19544) );
  OAI211_X1 U22542 ( .C1(n19611), .C2(n19591), .A(n19545), .B(n19544), .ZN(
        P2_U3139) );
  AOI22_X1 U22543 ( .A1(n19553), .A2(n19685), .B1(n19552), .B2(n19684), .ZN(
        n19547) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19658), .ZN(n19546) );
  OAI211_X1 U22545 ( .C1(n19661), .C2(n19591), .A(n19547), .B(n19546), .ZN(
        P2_U3140) );
  AOI22_X1 U22546 ( .A1(n19553), .A2(n19691), .B1(n19552), .B2(n19690), .ZN(
        n19549) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19614), .ZN(n19548) );
  OAI211_X1 U22548 ( .C1(n19617), .C2(n19591), .A(n19549), .B(n19548), .ZN(
        P2_U3141) );
  AOI22_X1 U22549 ( .A1(n19553), .A2(n19697), .B1(n19552), .B2(n19696), .ZN(
        n19551) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19699), .ZN(n19550) );
  OAI211_X1 U22551 ( .C1(n19620), .C2(n19591), .A(n19551), .B(n19550), .ZN(
        P2_U3142) );
  AOI22_X1 U22552 ( .A1(n19553), .A2(n19707), .B1(n19552), .B2(n19705), .ZN(
        n19557) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19622), .ZN(n19556) );
  OAI211_X1 U22554 ( .C1(n19627), .C2(n19591), .A(n19557), .B(n19556), .ZN(
        P2_U3143) );
  INV_X1 U22555 ( .A(n19558), .ZN(n19561) );
  INV_X1 U22556 ( .A(n19567), .ZN(n19560) );
  NAND3_X1 U22557 ( .A1(n19824), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19595) );
  NOR2_X1 U22558 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19595), .ZN(
        n19586) );
  OAI21_X1 U22559 ( .B1(n10291), .B2(n19586), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19559) );
  OAI21_X1 U22560 ( .B1(n19561), .B2(n19560), .A(n19559), .ZN(n19587) );
  AOI22_X1 U22561 ( .A1(n19587), .A2(n19205), .B1(n19673), .B2(n19586), .ZN(
        n19570) );
  INV_X1 U22562 ( .A(n19623), .ZN(n19605) );
  AOI21_X1 U22563 ( .B1(n19591), .B2(n19605), .A(n19847), .ZN(n19568) );
  OAI21_X1 U22564 ( .B1(n10291), .B2(n19852), .A(n19240), .ZN(n19565) );
  INV_X1 U22565 ( .A(n19586), .ZN(n19564) );
  AOI21_X1 U22566 ( .B1(n19565), .B2(n19564), .A(n19563), .ZN(n19566) );
  OAI211_X1 U22567 ( .C1(n19568), .C2(n19567), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19566), .ZN(n19588) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19675), .ZN(n19569) );
  OAI211_X1 U22569 ( .C1(n19571), .C2(n19591), .A(n19570), .B(n19569), .ZN(
        P2_U3144) );
  AOI22_X1 U22570 ( .A1(n19587), .A2(n19210), .B1(n19679), .B2(n19586), .ZN(
        n19573) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19680), .ZN(n19572) );
  OAI211_X1 U22572 ( .C1(n19683), .C2(n19591), .A(n19573), .B(n19572), .ZN(
        P2_U3145) );
  AOI22_X1 U22573 ( .A1(n19587), .A2(n15716), .B1(n19647), .B2(n19586), .ZN(
        n19576) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19574), .ZN(n19575) );
  OAI211_X1 U22575 ( .C1(n19577), .C2(n19591), .A(n19576), .B(n19575), .ZN(
        P2_U3146) );
  AOI22_X1 U22576 ( .A1(n19587), .A2(n15706), .B1(n19652), .B2(n19586), .ZN(
        n19579) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19653), .ZN(n19578) );
  OAI211_X1 U22578 ( .C1(n19656), .C2(n19591), .A(n19579), .B(n19578), .ZN(
        P2_U3147) );
  AOI22_X1 U22579 ( .A1(n19587), .A2(n19685), .B1(n19684), .B2(n19586), .ZN(
        n19581) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19686), .ZN(n19580) );
  OAI211_X1 U22581 ( .C1(n19689), .C2(n19591), .A(n19581), .B(n19580), .ZN(
        P2_U3148) );
  AOI22_X1 U22582 ( .A1(n19587), .A2(n19691), .B1(n19690), .B2(n19586), .ZN(
        n19583) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19692), .ZN(n19582) );
  OAI211_X1 U22584 ( .C1(n19695), .C2(n19591), .A(n19583), .B(n19582), .ZN(
        P2_U3149) );
  AOI22_X1 U22585 ( .A1(n19587), .A2(n19697), .B1(n19696), .B2(n19586), .ZN(
        n19585) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19698), .ZN(n19584) );
  OAI211_X1 U22587 ( .C1(n19666), .C2(n19591), .A(n19585), .B(n19584), .ZN(
        P2_U3150) );
  AOI22_X1 U22588 ( .A1(n19587), .A2(n19707), .B1(n19705), .B2(n19586), .ZN(
        n19590) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19588), .B1(
        n19623), .B2(n19709), .ZN(n19589) );
  OAI211_X1 U22590 ( .C1(n19715), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3151) );
  NOR2_X1 U22591 ( .A1(n19833), .A2(n19595), .ZN(n19630) );
  OAI21_X1 U22592 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19595), .A(n19852), 
        .ZN(n19594) );
  AND2_X1 U22593 ( .A1(n19598), .A2(n19594), .ZN(n19621) );
  AOI22_X1 U22594 ( .A1(n19621), .A2(n19205), .B1(n19673), .B2(n19630), .ZN(
        n19602) );
  OAI21_X1 U22595 ( .B1(n19597), .B2(n19596), .A(n19595), .ZN(n19599) );
  AND2_X1 U22596 ( .A1(n19599), .A2(n19598), .ZN(n19600) );
  OAI211_X1 U22597 ( .C1(n19630), .C2(n19240), .A(n19600), .B(n19634), .ZN(
        n19624) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19674), .ZN(n19601) );
  OAI211_X1 U22599 ( .C1(n19642), .C2(n19672), .A(n19602), .B(n19601), .ZN(
        P2_U3152) );
  AOI22_X1 U22600 ( .A1(n19621), .A2(n19210), .B1(n19679), .B2(n19630), .ZN(
        n19604) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19624), .B1(
        n19657), .B2(n19680), .ZN(n19603) );
  OAI211_X1 U22602 ( .C1(n19683), .C2(n19605), .A(n19604), .B(n19603), .ZN(
        P2_U3153) );
  AOI22_X1 U22603 ( .A1(n19621), .A2(n15716), .B1(n19647), .B2(n19630), .ZN(
        n19607) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19648), .ZN(n19606) );
  OAI211_X1 U22605 ( .C1(n19651), .C2(n19672), .A(n19607), .B(n19606), .ZN(
        P2_U3154) );
  AOI22_X1 U22606 ( .A1(n19621), .A2(n15706), .B1(n19652), .B2(n19630), .ZN(
        n19610) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19608), .ZN(n19609) );
  OAI211_X1 U22608 ( .C1(n19611), .C2(n19672), .A(n19610), .B(n19609), .ZN(
        P2_U3155) );
  AOI22_X1 U22609 ( .A1(n19621), .A2(n19685), .B1(n19684), .B2(n19630), .ZN(
        n19613) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19658), .ZN(n19612) );
  OAI211_X1 U22611 ( .C1(n19661), .C2(n19672), .A(n19613), .B(n19612), .ZN(
        P2_U3156) );
  AOI22_X1 U22612 ( .A1(n19621), .A2(n19691), .B1(n19690), .B2(n19630), .ZN(
        n19616) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19614), .ZN(n19615) );
  OAI211_X1 U22614 ( .C1(n19617), .C2(n19672), .A(n19616), .B(n19615), .ZN(
        P2_U3157) );
  AOI22_X1 U22615 ( .A1(n19621), .A2(n19697), .B1(n19696), .B2(n19630), .ZN(
        n19619) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19699), .ZN(n19618) );
  OAI211_X1 U22617 ( .C1(n19620), .C2(n19672), .A(n19619), .B(n19618), .ZN(
        P2_U3158) );
  AOI22_X1 U22618 ( .A1(n19621), .A2(n19707), .B1(n19705), .B2(n19630), .ZN(
        n19626) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19624), .B1(
        n19623), .B2(n19622), .ZN(n19625) );
  OAI211_X1 U22620 ( .C1(n19627), .C2(n19672), .A(n19626), .B(n19625), .ZN(
        P2_U3159) );
  NOR2_X1 U22621 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19628), .ZN(
        n19667) );
  AOI22_X1 U22622 ( .A1(n19674), .A2(n19657), .B1(n19673), .B2(n19667), .ZN(
        n19641) );
  NOR3_X1 U22623 ( .A1(n19700), .A2(n19657), .A3(n19795), .ZN(n19629) );
  NOR2_X1 U22624 ( .A1(n19629), .A2(n19798), .ZN(n19639) );
  NOR2_X1 U22625 ( .A1(n19667), .A2(n19630), .ZN(n19638) );
  INV_X1 U22626 ( .A(n19638), .ZN(n19635) );
  INV_X1 U22627 ( .A(n19667), .ZN(n19631) );
  OAI211_X1 U22628 ( .C1(n19632), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19795), 
        .B(n19631), .ZN(n19633) );
  OAI211_X1 U22629 ( .C1(n19639), .C2(n19635), .A(n19634), .B(n19633), .ZN(
        n19669) );
  OAI21_X1 U22630 ( .B1(n19636), .B2(n19667), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19637) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19669), .B1(
        n19205), .B2(n19668), .ZN(n19640) );
  OAI211_X1 U22632 ( .C1(n19642), .C2(n19714), .A(n19641), .B(n19640), .ZN(
        P2_U3160) );
  AOI22_X1 U22633 ( .A1(n19657), .A2(n19643), .B1(n19679), .B2(n19667), .ZN(
        n19645) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19669), .B1(
        n19210), .B2(n19668), .ZN(n19644) );
  OAI211_X1 U22635 ( .C1(n19646), .C2(n19714), .A(n19645), .B(n19644), .ZN(
        P2_U3161) );
  AOI22_X1 U22636 ( .A1(n19657), .A2(n19648), .B1(n19647), .B2(n19667), .ZN(
        n19650) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19669), .B1(
        n15716), .B2(n19668), .ZN(n19649) );
  OAI211_X1 U22638 ( .C1(n19651), .C2(n19714), .A(n19650), .B(n19649), .ZN(
        P2_U3162) );
  AOI22_X1 U22639 ( .A1(n19700), .A2(n19653), .B1(n19652), .B2(n19667), .ZN(
        n19655) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19669), .B1(
        n15706), .B2(n19668), .ZN(n19654) );
  OAI211_X1 U22641 ( .C1(n19656), .C2(n19672), .A(n19655), .B(n19654), .ZN(
        P2_U3163) );
  AOI22_X1 U22642 ( .A1(n19658), .A2(n19657), .B1(n19684), .B2(n19667), .ZN(
        n19660) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19669), .B1(
        n19685), .B2(n19668), .ZN(n19659) );
  OAI211_X1 U22644 ( .C1(n19661), .C2(n19714), .A(n19660), .B(n19659), .ZN(
        P2_U3164) );
  AOI22_X1 U22645 ( .A1(n19692), .A2(n19700), .B1(n19690), .B2(n19667), .ZN(
        n19663) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19669), .B1(
        n19691), .B2(n19668), .ZN(n19662) );
  OAI211_X1 U22647 ( .C1(n19695), .C2(n19672), .A(n19663), .B(n19662), .ZN(
        P2_U3165) );
  AOI22_X1 U22648 ( .A1(n19698), .A2(n19700), .B1(n19696), .B2(n19667), .ZN(
        n19665) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19669), .B1(
        n19697), .B2(n19668), .ZN(n19664) );
  OAI211_X1 U22650 ( .C1(n19666), .C2(n19672), .A(n19665), .B(n19664), .ZN(
        P2_U3166) );
  AOI22_X1 U22651 ( .A1(n19709), .A2(n19700), .B1(n19705), .B2(n19667), .ZN(
        n19671) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19669), .B1(
        n19707), .B2(n19668), .ZN(n19670) );
  OAI211_X1 U22653 ( .C1(n19715), .C2(n19672), .A(n19671), .B(n19670), .ZN(
        P2_U3167) );
  INV_X1 U22654 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19678) );
  AOI22_X1 U22655 ( .A1(n19708), .A2(n19205), .B1(n19706), .B2(n19673), .ZN(
        n19677) );
  AOI22_X1 U22656 ( .A1(n19710), .A2(n19675), .B1(n19700), .B2(n19674), .ZN(
        n19676) );
  OAI211_X1 U22657 ( .C1(n19704), .C2(n19678), .A(n19677), .B(n19676), .ZN(
        P2_U3168) );
  AOI22_X1 U22658 ( .A1(n19708), .A2(n19210), .B1(n19706), .B2(n19679), .ZN(
        n19682) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19680), .ZN(n19681) );
  OAI211_X1 U22660 ( .C1(n19683), .C2(n19714), .A(n19682), .B(n19681), .ZN(
        P2_U3169) );
  AOI22_X1 U22661 ( .A1(n19708), .A2(n19685), .B1(n19706), .B2(n19684), .ZN(
        n19688) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19686), .ZN(n19687) );
  OAI211_X1 U22663 ( .C1(n19689), .C2(n19714), .A(n19688), .B(n19687), .ZN(
        P2_U3172) );
  AOI22_X1 U22664 ( .A1(n19708), .A2(n19691), .B1(n19706), .B2(n19690), .ZN(
        n19694) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19692), .ZN(n19693) );
  OAI211_X1 U22666 ( .C1(n19695), .C2(n19714), .A(n19694), .B(n19693), .ZN(
        P2_U3173) );
  AOI22_X1 U22667 ( .A1(n19708), .A2(n19697), .B1(n19706), .B2(n19696), .ZN(
        n19702) );
  AOI22_X1 U22668 ( .A1(n19700), .A2(n19699), .B1(n19710), .B2(n19698), .ZN(
        n19701) );
  OAI211_X1 U22669 ( .C1(n19704), .C2(n19703), .A(n19702), .B(n19701), .ZN(
        P2_U3174) );
  AOI22_X1 U22670 ( .A1(n19708), .A2(n19707), .B1(n19706), .B2(n19705), .ZN(
        n19713) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19711), .B1(
        n19710), .B2(n19709), .ZN(n19712) );
  OAI211_X1 U22672 ( .C1(n19715), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3175) );
  NOR2_X1 U22673 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19716), .ZN(n19717) );
  OAI211_X1 U22674 ( .C1(n19718), .C2(n19717), .A(n19853), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19723) );
  NOR4_X1 U22675 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n19853), .A4(n19716), .ZN(n19720) );
  OAI21_X1 U22676 ( .B1(n19721), .B2(n19720), .A(n19719), .ZN(n19722) );
  NAND3_X1 U22677 ( .A1(n19724), .A2(n19723), .A3(n19722), .ZN(P2_U3177) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19726), .ZN(
        P2_U3179) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19726), .ZN(
        P2_U3180) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19726), .ZN(
        P2_U3181) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19726), .ZN(
        P2_U3182) );
  NOR2_X1 U22682 ( .A1(n19725), .A2(n19793), .ZN(P2_U3183) );
  AND2_X1 U22683 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19726), .ZN(
        P2_U3184) );
  AND2_X1 U22684 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19726), .ZN(
        P2_U3185) );
  AND2_X1 U22685 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19726), .ZN(
        P2_U3186) );
  AND2_X1 U22686 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19726), .ZN(
        P2_U3187) );
  AND2_X1 U22687 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19726), .ZN(
        P2_U3188) );
  NOR2_X1 U22688 ( .A1(n20849), .A2(n19793), .ZN(P2_U3189) );
  AND2_X1 U22689 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19726), .ZN(
        P2_U3190) );
  AND2_X1 U22690 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19726), .ZN(
        P2_U3191) );
  AND2_X1 U22691 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19726), .ZN(
        P2_U3192) );
  AND2_X1 U22692 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19726), .ZN(
        P2_U3193) );
  AND2_X1 U22693 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19726), .ZN(
        P2_U3194) );
  AND2_X1 U22694 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19726), .ZN(
        P2_U3195) );
  AND2_X1 U22695 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19726), .ZN(
        P2_U3196) );
  AND2_X1 U22696 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19726), .ZN(
        P2_U3197) );
  AND2_X1 U22697 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19726), .ZN(
        P2_U3198) );
  AND2_X1 U22698 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19726), .ZN(
        P2_U3199) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19726), .ZN(
        P2_U3200) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19726), .ZN(P2_U3201) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19726), .ZN(P2_U3202) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19726), .ZN(P2_U3203) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19726), .ZN(P2_U3204) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19726), .ZN(P2_U3205) );
  AND2_X1 U22705 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19726), .ZN(P2_U3206) );
  AND2_X1 U22706 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19726), .ZN(P2_U3207) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19726), .ZN(P2_U3208) );
  OAI21_X1 U22708 ( .B1(n20646), .B2(n19731), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19741) );
  NAND2_X1 U22709 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19853), .ZN(n19739) );
  NAND3_X1 U22710 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19739), .ZN(n19729) );
  AOI211_X1 U22711 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n19734), .A(
        n19867), .B(n19727), .ZN(n19728) );
  AOI21_X1 U22712 ( .B1(n19741), .B2(n19729), .A(n19728), .ZN(n19730) );
  INV_X1 U22713 ( .A(n19730), .ZN(P2_U3209) );
  AND2_X1 U22714 ( .A1(n19848), .A2(n19739), .ZN(n19733) );
  NOR2_X1 U22715 ( .A1(HOLD), .A2(n20893), .ZN(n19740) );
  OAI211_X1 U22716 ( .C1(n19740), .C2(n19742), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19731), .ZN(n19732) );
  OAI211_X1 U22717 ( .C1(n19735), .C2(n19734), .A(n19733), .B(n19732), .ZN(
        P2_U3210) );
  OAI22_X1 U22718 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19736), .B1(NA), 
        .B2(n19739), .ZN(n19737) );
  OAI211_X1 U22719 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19737), .ZN(n19738) );
  OAI221_X1 U22720 ( .B1(n19741), .B2(n19740), .C1(n19741), .C2(n19739), .A(
        n19738), .ZN(P2_U3211) );
  OAI222_X1 U22721 ( .A1(n19784), .A2(n13281), .B1(n19743), .B2(n19867), .C1(
        n10037), .C2(n19778), .ZN(P2_U3212) );
  OAI222_X1 U22722 ( .A1(n19784), .A2(n10081), .B1(n19744), .B2(n19867), .C1(
        n13281), .C2(n19778), .ZN(P2_U3213) );
  OAI222_X1 U22723 ( .A1(n19784), .A2(n10755), .B1(n19745), .B2(n19867), .C1(
        n10081), .C2(n19778), .ZN(P2_U3214) );
  OAI222_X1 U22724 ( .A1(n19784), .A2(n10761), .B1(n19746), .B2(n19867), .C1(
        n10755), .C2(n19778), .ZN(P2_U3215) );
  OAI222_X1 U22725 ( .A1(n19784), .A2(n10767), .B1(n19747), .B2(n19867), .C1(
        n10761), .C2(n19778), .ZN(P2_U3216) );
  OAI222_X1 U22726 ( .A1(n19784), .A2(n10771), .B1(n19748), .B2(n19867), .C1(
        n10767), .C2(n19778), .ZN(P2_U3217) );
  OAI222_X1 U22727 ( .A1(n19784), .A2(n13413), .B1(n19749), .B2(n19867), .C1(
        n10771), .C2(n19778), .ZN(P2_U3218) );
  OAI222_X1 U22728 ( .A1(n19784), .A2(n10787), .B1(n19750), .B2(n19867), .C1(
        n13413), .C2(n19778), .ZN(P2_U3219) );
  OAI222_X1 U22729 ( .A1(n19784), .A2(n13620), .B1(n19751), .B2(n19867), .C1(
        n10787), .C2(n19781), .ZN(P2_U3220) );
  OAI222_X1 U22730 ( .A1(n19784), .A2(n10779), .B1(n19752), .B2(n19867), .C1(
        n13620), .C2(n19781), .ZN(P2_U3221) );
  OAI222_X1 U22731 ( .A1(n19784), .A2(n10792), .B1(n20785), .B2(n19867), .C1(
        n10779), .C2(n19781), .ZN(P2_U3222) );
  OAI222_X1 U22732 ( .A1(n19784), .A2(n15336), .B1(n19753), .B2(n19867), .C1(
        n10792), .C2(n19781), .ZN(P2_U3223) );
  OAI222_X1 U22733 ( .A1(n19784), .A2(n13960), .B1(n19754), .B2(n19867), .C1(
        n15336), .C2(n19781), .ZN(P2_U3224) );
  OAI222_X1 U22734 ( .A1(n19784), .A2(n15326), .B1(n20868), .B2(n19867), .C1(
        n13960), .C2(n19781), .ZN(P2_U3225) );
  OAI222_X1 U22735 ( .A1(n19784), .A2(n15513), .B1(n19755), .B2(n19867), .C1(
        n15326), .C2(n19781), .ZN(P2_U3226) );
  OAI222_X1 U22736 ( .A1(n19784), .A2(n19757), .B1(n19756), .B2(n19867), .C1(
        n15513), .C2(n19781), .ZN(P2_U3227) );
  OAI222_X1 U22737 ( .A1(n19784), .A2(n19759), .B1(n19758), .B2(n19867), .C1(
        n19757), .C2(n19781), .ZN(P2_U3228) );
  OAI222_X1 U22738 ( .A1(n19784), .A2(n19761), .B1(n19760), .B2(n19867), .C1(
        n19759), .C2(n19781), .ZN(P2_U3229) );
  OAI222_X1 U22739 ( .A1(n19784), .A2(n19763), .B1(n19762), .B2(n19867), .C1(
        n19761), .C2(n19778), .ZN(P2_U3230) );
  OAI222_X1 U22740 ( .A1(n19784), .A2(n19765), .B1(n19764), .B2(n19867), .C1(
        n19763), .C2(n19778), .ZN(P2_U3231) );
  OAI222_X1 U22741 ( .A1(n19784), .A2(n15042), .B1(n19766), .B2(n19867), .C1(
        n19765), .C2(n19778), .ZN(P2_U3232) );
  OAI222_X1 U22742 ( .A1(n19784), .A2(n19768), .B1(n19767), .B2(n19867), .C1(
        n15042), .C2(n19778), .ZN(P2_U3233) );
  OAI222_X1 U22743 ( .A1(n19784), .A2(n15253), .B1(n19769), .B2(n19867), .C1(
        n19768), .C2(n19778), .ZN(P2_U3234) );
  OAI222_X1 U22744 ( .A1(n19784), .A2(n19771), .B1(n19770), .B2(n19867), .C1(
        n15253), .C2(n19778), .ZN(P2_U3235) );
  OAI222_X1 U22745 ( .A1(n19784), .A2(n19773), .B1(n19772), .B2(n19867), .C1(
        n19771), .C2(n19778), .ZN(P2_U3236) );
  OAI222_X1 U22746 ( .A1(n19784), .A2(n19775), .B1(n19774), .B2(n19867), .C1(
        n19773), .C2(n19778), .ZN(P2_U3237) );
  OAI222_X1 U22747 ( .A1(n19781), .A2(n19775), .B1(n20886), .B2(n19867), .C1(
        n19776), .C2(n19784), .ZN(P2_U3238) );
  OAI222_X1 U22748 ( .A1(n19784), .A2(n19779), .B1(n19777), .B2(n19867), .C1(
        n19776), .C2(n19778), .ZN(P2_U3239) );
  OAI222_X1 U22749 ( .A1(n19784), .A2(n10857), .B1(n19780), .B2(n19867), .C1(
        n19779), .C2(n19778), .ZN(P2_U3240) );
  INV_X1 U22750 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19783) );
  OAI222_X1 U22751 ( .A1(n19784), .A2(n19783), .B1(n19782), .B2(n19867), .C1(
        n10857), .C2(n19781), .ZN(P2_U3241) );
  INV_X1 U22752 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U22753 ( .A1(n19867), .A2(n20784), .B1(n19785), .B2(n19864), .ZN(
        P2_U3585) );
  MUX2_X1 U22754 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19867), .Z(P2_U3586) );
  INV_X1 U22755 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U22756 ( .A1(n19867), .A2(n19787), .B1(n19786), .B2(n19864), .ZN(
        P2_U3587) );
  INV_X1 U22757 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U22758 ( .A1(n19867), .A2(n19789), .B1(n19788), .B2(n19864), .ZN(
        P2_U3588) );
  OAI21_X1 U22759 ( .B1(n19793), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19791), 
        .ZN(n19790) );
  INV_X1 U22760 ( .A(n19790), .ZN(P2_U3591) );
  OAI21_X1 U22761 ( .B1(n19793), .B2(n19792), .A(n19791), .ZN(P2_U3592) );
  NOR3_X1 U22762 ( .A1(n19796), .A2(n19795), .A3(n19794), .ZN(n19804) );
  NAND2_X1 U22763 ( .A1(n19800), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19819) );
  NOR2_X1 U22764 ( .A1(n19797), .A2(n19819), .ZN(n19812) );
  INV_X1 U22765 ( .A(n19812), .ZN(n19802) );
  AOI211_X1 U22766 ( .C1(n19817), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        n19808) );
  AOI21_X1 U22767 ( .B1(n19802), .B2(n19808), .A(n19801), .ZN(n19803) );
  AOI211_X1 U22768 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19805), .A(n19804), 
        .B(n19803), .ZN(n19806) );
  AOI22_X1 U22769 ( .A1(n19834), .A2(n19807), .B1(n19806), .B2(n19831), .ZN(
        P2_U3602) );
  INV_X1 U22770 ( .A(n19808), .ZN(n19811) );
  AOI22_X1 U22771 ( .A1(n19811), .A2(n19810), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19809), .ZN(n19814) );
  NOR2_X1 U22772 ( .A1(n19834), .A2(n19812), .ZN(n19813) );
  AOI22_X1 U22773 ( .A1(n12395), .A2(n19834), .B1(n19814), .B2(n19813), .ZN(
        P2_U3603) );
  INV_X1 U22774 ( .A(n19815), .ZN(n19826) );
  OR3_X1 U22775 ( .A1(n19817), .A2(n19826), .A3(n19816), .ZN(n19818) );
  OAI21_X1 U22776 ( .B1(n19820), .B2(n19819), .A(n19818), .ZN(n19821) );
  AOI21_X1 U22777 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19822), .A(n19821), 
        .ZN(n19823) );
  AOI22_X1 U22778 ( .A1(n19834), .A2(n19824), .B1(n19823), .B2(n19831), .ZN(
        P2_U3604) );
  NAND2_X1 U22779 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19833), .ZN(n19825) );
  OAI21_X1 U22780 ( .B1(n19827), .B2(n19826), .A(n19825), .ZN(n19828) );
  AOI21_X1 U22781 ( .B1(n19830), .B2(n19829), .A(n19828), .ZN(n19832) );
  AOI22_X1 U22782 ( .A1(n19834), .A2(n19833), .B1(n19832), .B2(n19831), .ZN(
        P2_U3605) );
  INV_X1 U22783 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19835) );
  AOI22_X1 U22784 ( .A1(n19867), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19835), 
        .B2(n19864), .ZN(P2_U3608) );
  INV_X1 U22785 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19845) );
  INV_X1 U22786 ( .A(n19836), .ZN(n19844) );
  AOI22_X1 U22787 ( .A1(n19840), .A2(n19839), .B1(n19838), .B2(n19837), .ZN(
        n19843) );
  NOR2_X1 U22788 ( .A1(n19844), .A2(n19841), .ZN(n19842) );
  AOI22_X1 U22789 ( .A1(n19845), .A2(n19844), .B1(n19843), .B2(n19842), .ZN(
        P2_U3609) );
  OAI21_X1 U22790 ( .B1(n19848), .B2(n19847), .A(n19846), .ZN(n19851) );
  NAND3_X1 U22791 ( .A1(n19848), .A2(n9627), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19850) );
  MUX2_X1 U22792 ( .A(n19851), .B(n19850), .S(n19849), .Z(n19856) );
  OAI22_X1 U22793 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19854), .B1(n19853), 
        .B2(n19852), .ZN(n19855) );
  NAND2_X1 U22794 ( .A1(n19856), .A2(n19855), .ZN(n19863) );
  NOR2_X1 U22795 ( .A1(n19857), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19859) );
  AOI211_X1 U22796 ( .C1(n19861), .C2(n19860), .A(n19859), .B(n19858), .ZN(
        n19862) );
  MUX2_X1 U22797 ( .A(n19863), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19862), 
        .Z(P2_U3610) );
  INV_X1 U22798 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19865) );
  AOI22_X1 U22799 ( .A1(n19867), .A2(n19866), .B1(n19865), .B2(n19864), .ZN(
        P2_U3611) );
  AOI21_X1 U22800 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20653), .A(n20650), 
        .ZN(n19875) );
  INV_X1 U22801 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19869) );
  INV_X2 U22802 ( .A(n20737), .ZN(n20750) );
  AOI21_X1 U22803 ( .B1(n19875), .B2(n19869), .A(n20750), .ZN(P1_U2802) );
  NAND2_X1 U22804 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20745), .ZN(n19873) );
  OAI21_X1 U22805 ( .B1(n19871), .B2(n19870), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19872) );
  OAI21_X1 U22806 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n19873), .A(n19872), 
        .ZN(P1_U2803) );
  NOR2_X1 U22807 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19876) );
  OAI21_X1 U22808 ( .B1(n19876), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20737), .ZN(
        n19874) );
  OAI21_X1 U22809 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20737), .A(n19874), 
        .ZN(P1_U2804) );
  NOR2_X1 U22810 ( .A1(n20750), .A2(n19875), .ZN(n20721) );
  OAI21_X1 U22811 ( .B1(BS16), .B2(n19876), .A(n20721), .ZN(n20719) );
  OAI21_X1 U22812 ( .B1(n20721), .B2(n20496), .A(n20719), .ZN(P1_U2805) );
  INV_X1 U22813 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22814 ( .B1(n19879), .B2(n19878), .A(n19877), .ZN(P1_U2806) );
  NOR4_X1 U22815 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19883) );
  NOR4_X1 U22816 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19882) );
  NOR4_X1 U22817 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19881) );
  NOR4_X1 U22818 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19880) );
  NAND4_X1 U22819 ( .A1(n19883), .A2(n19882), .A3(n19881), .A4(n19880), .ZN(
        n19889) );
  NOR4_X1 U22820 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19887) );
  AOI211_X1 U22821 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_17__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19886) );
  NOR4_X1 U22822 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19885) );
  NOR4_X1 U22823 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19884) );
  NAND4_X1 U22824 ( .A1(n19887), .A2(n19886), .A3(n19885), .A4(n19884), .ZN(
        n19888) );
  NOR2_X1 U22825 ( .A1(n19889), .A2(n19888), .ZN(n20736) );
  INV_X1 U22826 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20714) );
  NOR3_X1 U22827 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19891) );
  OAI21_X1 U22828 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19891), .A(n20736), .ZN(
        n19890) );
  OAI21_X1 U22829 ( .B1(n20736), .B2(n20714), .A(n19890), .ZN(P1_U2807) );
  INV_X1 U22830 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20720) );
  AOI21_X1 U22831 ( .B1(n20729), .B2(n20720), .A(n19891), .ZN(n19892) );
  INV_X1 U22832 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20711) );
  INV_X1 U22833 ( .A(n20736), .ZN(n20731) );
  AOI22_X1 U22834 ( .A1(n20736), .A2(n19892), .B1(n20711), .B2(n20731), .ZN(
        P1_U2808) );
  OAI22_X1 U22835 ( .A1(n19969), .A2(n19924), .B1(n19965), .B2(n19893), .ZN(
        n19894) );
  INV_X1 U22836 ( .A(n19894), .ZN(n19901) );
  INV_X1 U22837 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20668) );
  AOI22_X1 U22838 ( .A1(n19895), .A2(n19936), .B1(n19955), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19896) );
  OAI211_X1 U22839 ( .C1(n19919), .C2(n14119), .A(n19896), .B(n19933), .ZN(
        n19897) );
  AOI221_X1 U22840 ( .B1(n19899), .B2(n20668), .C1(n19898), .C2(
        P1_REIP_REG_9__SCAN_IN), .A(n19897), .ZN(n19900) );
  NAND2_X1 U22841 ( .A1(n19901), .A2(n19900), .ZN(P1_U2831) );
  NAND2_X1 U22842 ( .A1(n19903), .A2(n19902), .ZN(n19915) );
  NOR2_X1 U22843 ( .A1(n19905), .A2(n19904), .ZN(n19928) );
  AOI22_X1 U22844 ( .A1(n19936), .A2(n19906), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19928), .ZN(n19914) );
  NAND2_X1 U22845 ( .A1(n19953), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19911) );
  INV_X1 U22846 ( .A(n19907), .ZN(n19908) );
  NAND2_X1 U22847 ( .A1(n19909), .A2(n19908), .ZN(n19910) );
  NAND3_X1 U22848 ( .A1(n19911), .A2(n19910), .A3(n19933), .ZN(n19912) );
  AOI21_X1 U22849 ( .B1(n19955), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19912), .ZN(
        n19913) );
  AND3_X1 U22850 ( .A1(n19915), .A2(n19914), .A3(n19913), .ZN(n19916) );
  OAI21_X1 U22851 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n19917), .A(n19916), .ZN(
        P1_U2833) );
  OAI21_X1 U22852 ( .B1(n19919), .B2(n19918), .A(n19933), .ZN(n19922) );
  NOR2_X1 U22853 ( .A1(n19920), .A2(n19948), .ZN(n19921) );
  AOI211_X1 U22854 ( .C1(n19955), .C2(P1_EBX_REG_6__SCAN_IN), .A(n19922), .B(
        n19921), .ZN(n19930) );
  OAI22_X1 U22855 ( .A1(n19925), .A2(n19924), .B1(n19923), .B2(n19965), .ZN(
        n19926) );
  AOI221_X1 U22856 ( .B1(n19928), .B2(P1_REIP_REG_6__SCAN_IN), .C1(n19927), 
        .C2(n20663), .A(n19926), .ZN(n19929) );
  NAND2_X1 U22857 ( .A1(n19930), .A2(n19929), .ZN(P1_U2834) );
  NAND2_X1 U22858 ( .A1(n19932), .A2(n19931), .ZN(n19961) );
  NAND2_X1 U22859 ( .A1(n19953), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19934) );
  NAND2_X1 U22860 ( .A1(n19934), .A2(n19933), .ZN(n19935) );
  AOI21_X1 U22861 ( .B1(n19955), .B2(P1_EBX_REG_5__SCAN_IN), .A(n19935), .ZN(
        n19939) );
  NAND2_X1 U22862 ( .A1(n19937), .A2(n19936), .ZN(n19938) );
  OAI211_X1 U22863 ( .C1(n19940), .C2(P1_REIP_REG_5__SCAN_IN), .A(n19939), .B(
        n19938), .ZN(n19941) );
  INV_X1 U22864 ( .A(n19941), .ZN(n19944) );
  NAND2_X1 U22865 ( .A1(n19942), .A2(n19958), .ZN(n19943) );
  OAI211_X1 U22866 ( .C1(n19961), .C2(n20661), .A(n19944), .B(n19943), .ZN(
        n19945) );
  INV_X1 U22867 ( .A(n19945), .ZN(n19946) );
  OAI21_X1 U22868 ( .B1(n19947), .B2(n19965), .A(n19946), .ZN(P1_U2835) );
  OAI22_X1 U22869 ( .A1(n19950), .A2(n19949), .B1(n19948), .B2(n19994), .ZN(
        n19951) );
  AOI211_X1 U22870 ( .C1(n19953), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19952), .B(n19951), .ZN(n19964) );
  NOR2_X1 U22871 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19954), .ZN(n19956) );
  AOI22_X1 U22872 ( .A1(n19957), .A2(n19956), .B1(n19955), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19960) );
  NAND2_X1 U22873 ( .A1(n19979), .A2(n19958), .ZN(n19959) );
  OAI211_X1 U22874 ( .C1(n19961), .C2(n20659), .A(n19960), .B(n19959), .ZN(
        n19962) );
  INV_X1 U22875 ( .A(n19962), .ZN(n19963) );
  OAI211_X1 U22876 ( .C1(n19984), .C2(n19965), .A(n19964), .B(n19963), .ZN(
        P1_U2836) );
  OAI22_X1 U22877 ( .A1(n19969), .A2(n19968), .B1(n19967), .B2(n19966), .ZN(
        n19970) );
  INV_X1 U22878 ( .A(n19970), .ZN(n19971) );
  OAI21_X1 U22879 ( .B1(n14535), .B2(n19972), .A(n19971), .ZN(P1_U2863) );
  AOI22_X1 U22880 ( .A1(n19974), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19973), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19983) );
  OAI21_X1 U22881 ( .B1(n9613), .B2(n19976), .A(n19975), .ZN(n19978) );
  INV_X1 U22882 ( .A(n19978), .ZN(n19997) );
  AOI22_X1 U22883 ( .A1(n19997), .A2(n19981), .B1(n19980), .B2(n19979), .ZN(
        n19982) );
  OAI211_X1 U22884 ( .C1(n19985), .C2(n19984), .A(n19983), .B(n19982), .ZN(
        P1_U2995) );
  OAI21_X1 U22885 ( .B1(n19988), .B2(n19987), .A(n19986), .ZN(n19989) );
  AOI21_X1 U22886 ( .B1(n19990), .B2(n20015), .A(n19989), .ZN(n20008) );
  OAI211_X1 U22887 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19991), .B(n20003), .ZN(n19992) );
  INV_X1 U22888 ( .A(n19992), .ZN(n19996) );
  OAI22_X1 U22889 ( .A1(n19994), .A2(n19993), .B1(n20659), .B2(n19933), .ZN(
        n19995) );
  AOI211_X1 U22890 ( .C1(n19997), .C2(n20013), .A(n19996), .B(n19995), .ZN(
        n19998) );
  OAI21_X1 U22891 ( .B1(n20008), .B2(n19999), .A(n19998), .ZN(P1_U3027) );
  INV_X1 U22892 ( .A(n20000), .ZN(n20002) );
  AOI21_X1 U22893 ( .B1(n20002), .B2(n20021), .A(n20001), .ZN(n20006) );
  AOI22_X1 U22894 ( .A1(n20004), .A2(n20013), .B1(n20003), .B2(n20007), .ZN(
        n20005) );
  OAI211_X1 U22895 ( .C1(n20008), .C2(n20007), .A(n20006), .B(n20005), .ZN(
        P1_U3028) );
  NAND2_X1 U22896 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20009), .ZN(
        n20027) );
  AOI21_X1 U22897 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(n20025) );
  NAND3_X1 U22898 ( .A1(n20014), .A2(n13565), .A3(n20013), .ZN(n20023) );
  AND2_X1 U22899 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20016) );
  AOI21_X1 U22900 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20016), .A(
        n20015), .ZN(n20017) );
  INV_X1 U22901 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20656) );
  OAI22_X1 U22902 ( .A1(n20018), .A2(n20017), .B1(n20656), .B2(n19933), .ZN(
        n20019) );
  AOI21_X1 U22903 ( .B1(n20021), .B2(n20020), .A(n20019), .ZN(n20022) );
  AND2_X1 U22904 ( .A1(n20023), .A2(n20022), .ZN(n20024) );
  OAI221_X1 U22905 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20027), .C1(
        n20026), .C2(n20025), .A(n20024), .ZN(P1_U3029) );
  NOR2_X1 U22906 ( .A1(n20029), .A2(n20028), .ZN(P1_U3032) );
  INV_X1 U22907 ( .A(n20525), .ZN(n20578) );
  AOI22_X1 U22908 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9580), .B1(DATAI_24_), 
        .B2(n9579), .ZN(n20535) );
  NAND2_X1 U22909 ( .A1(n20084), .A2(n20037), .ZN(n20442) );
  NOR2_X1 U22910 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20158) );
  INV_X1 U22911 ( .A(n20158), .ZN(n20038) );
  NOR2_X1 U22912 ( .A1(n20038), .A2(n20441), .ZN(n20047) );
  INV_X1 U22913 ( .A(n20047), .ZN(n20085) );
  OAI22_X1 U22914 ( .A1(n20632), .A2(n20535), .B1(n20442), .B2(n20085), .ZN(
        n20039) );
  INV_X1 U22915 ( .A(n20039), .ZN(n20053) );
  NAND2_X1 U22916 ( .A1(n20049), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20521) );
  INV_X1 U22917 ( .A(n20632), .ZN(n20040) );
  NOR3_X1 U22918 ( .A1(n20111), .A2(n20040), .A3(n20574), .ZN(n20042) );
  NAND2_X1 U22919 ( .A1(n20499), .A2(n20496), .ZN(n20445) );
  INV_X1 U22920 ( .A(n20445), .ZN(n20041) );
  NOR2_X1 U22921 ( .A1(n20042), .A2(n20041), .ZN(n20051) );
  INV_X1 U22922 ( .A(n20051), .ZN(n20045) );
  NOR2_X1 U22923 ( .A1(n20319), .A2(n20043), .ZN(n20163) );
  NAND2_X1 U22924 ( .A1(n20163), .A2(n20449), .ZN(n20050) );
  INV_X1 U22925 ( .A(n20321), .ZN(n20044) );
  NAND2_X1 U22926 ( .A1(n20044), .A2(n20375), .ZN(n20199) );
  AOI22_X1 U22927 ( .A1(n20045), .A2(n20050), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20199), .ZN(n20046) );
  NOR2_X2 U22928 ( .A1(n20048), .A2(n20095), .ZN(n20577) );
  OR2_X1 U22929 ( .A1(n20049), .A2(n20638), .ZN(n20379) );
  OAI22_X1 U22930 ( .A1(n20051), .A2(n20050), .B1(n20379), .B2(n20199), .ZN(
        n20088) );
  AOI22_X1 U22931 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20089), .B1(
        n20577), .B2(n20088), .ZN(n20052) );
  OAI211_X1 U22932 ( .C1(n20586), .C2(n20120), .A(n20053), .B(n20052), .ZN(
        P1_U3033) );
  AOI22_X1 U22933 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9580), .B1(DATAI_25_), 
        .B2(n9579), .ZN(n20539) );
  NAND2_X1 U22934 ( .A1(n20084), .A2(n20054), .ZN(n20459) );
  OAI22_X1 U22935 ( .A1(n20632), .A2(n20539), .B1(n20459), .B2(n20085), .ZN(
        n20055) );
  INV_X1 U22936 ( .A(n20055), .ZN(n20058) );
  NOR2_X2 U22937 ( .A1(n20056), .A2(n20095), .ZN(n20588) );
  AOI22_X1 U22938 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20089), .B1(
        n20588), .B2(n20088), .ZN(n20057) );
  OAI211_X1 U22939 ( .C1(n20592), .C2(n20120), .A(n20058), .B(n20057), .ZN(
        P1_U3034) );
  AOI22_X1 U22940 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9580), .B1(DATAI_26_), 
        .B2(n9579), .ZN(n20543) );
  NAND2_X1 U22941 ( .A1(n20084), .A2(n20059), .ZN(n20463) );
  OAI22_X1 U22942 ( .A1(n20632), .A2(n20543), .B1(n20463), .B2(n20085), .ZN(
        n20060) );
  INV_X1 U22943 ( .A(n20060), .ZN(n20063) );
  NOR2_X2 U22944 ( .A1(n20061), .A2(n20095), .ZN(n20594) );
  AOI22_X1 U22945 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20089), .B1(
        n20594), .B2(n20088), .ZN(n20062) );
  OAI211_X1 U22946 ( .C1(n20598), .C2(n20120), .A(n20063), .B(n20062), .ZN(
        P1_U3035) );
  AOI22_X1 U22947 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9580), .B1(DATAI_27_), 
        .B2(n9579), .ZN(n20547) );
  NAND2_X1 U22948 ( .A1(n20084), .A2(n20064), .ZN(n20467) );
  OAI22_X1 U22949 ( .A1(n20632), .A2(n20547), .B1(n20467), .B2(n20085), .ZN(
        n20065) );
  INV_X1 U22950 ( .A(n20065), .ZN(n20068) );
  NOR2_X2 U22951 ( .A1(n20066), .A2(n20095), .ZN(n20600) );
  AOI22_X1 U22952 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20089), .B1(
        n20600), .B2(n20088), .ZN(n20067) );
  OAI211_X1 U22953 ( .C1(n20604), .C2(n20120), .A(n20068), .B(n20067), .ZN(
        P1_U3036) );
  AOI22_X1 U22954 ( .A1(DATAI_20_), .A2(n9579), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n9580), .ZN(n20610) );
  NAND2_X1 U22955 ( .A1(n20084), .A2(n11115), .ZN(n20471) );
  OAI22_X1 U22956 ( .A1(n20632), .A2(n20551), .B1(n20471), .B2(n20085), .ZN(
        n20069) );
  INV_X1 U22957 ( .A(n20069), .ZN(n20072) );
  NOR2_X2 U22958 ( .A1(n20070), .A2(n20095), .ZN(n20606) );
  AOI22_X1 U22959 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20089), .B1(
        n20606), .B2(n20088), .ZN(n20071) );
  OAI211_X1 U22960 ( .C1(n20610), .C2(n20120), .A(n20072), .B(n20071), .ZN(
        P1_U3037) );
  AOI22_X1 U22961 ( .A1(DATAI_21_), .A2(n9579), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n9580), .ZN(n20616) );
  NAND2_X1 U22962 ( .A1(n20084), .A2(n20073), .ZN(n20475) );
  OAI22_X1 U22963 ( .A1(n20632), .A2(n20555), .B1(n20475), .B2(n20085), .ZN(
        n20074) );
  INV_X1 U22964 ( .A(n20074), .ZN(n20077) );
  NOR2_X2 U22965 ( .A1(n20075), .A2(n20095), .ZN(n20612) );
  AOI22_X1 U22966 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20089), .B1(
        n20612), .B2(n20088), .ZN(n20076) );
  OAI211_X1 U22967 ( .C1(n20616), .C2(n20120), .A(n20077), .B(n20076), .ZN(
        P1_U3038) );
  AOI22_X1 U22968 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9580), .B1(DATAI_22_), 
        .B2(n9579), .ZN(n20622) );
  NAND2_X1 U22969 ( .A1(n20084), .A2(n20078), .ZN(n20479) );
  OAI22_X1 U22970 ( .A1(n20632), .A2(n20559), .B1(n20479), .B2(n20085), .ZN(
        n20079) );
  INV_X1 U22971 ( .A(n20079), .ZN(n20082) );
  NOR2_X2 U22972 ( .A1(n20080), .A2(n20095), .ZN(n20618) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20089), .B1(
        n20618), .B2(n20088), .ZN(n20081) );
  OAI211_X1 U22974 ( .C1(n20622), .C2(n20120), .A(n20082), .B(n20081), .ZN(
        P1_U3039) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n9580), .B1(DATAI_31_), 
        .B2(n9579), .ZN(n20567) );
  NAND2_X1 U22976 ( .A1(n20084), .A2(n9634), .ZN(n20484) );
  OAI22_X1 U22977 ( .A1(n20632), .A2(n20567), .B1(n20484), .B2(n20085), .ZN(
        n20086) );
  INV_X1 U22978 ( .A(n20086), .ZN(n20091) );
  NOR2_X2 U22979 ( .A1(n20087), .A2(n20095), .ZN(n20626) );
  AOI22_X1 U22980 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20089), .B1(
        n20626), .B2(n20088), .ZN(n20090) );
  OAI211_X1 U22981 ( .C1(n20633), .C2(n20120), .A(n20091), .B(n20090), .ZN(
        P1_U3040) );
  NAND2_X1 U22982 ( .A1(n20158), .A2(n20572), .ZN(n20094) );
  NOR2_X1 U22983 ( .A1(n20493), .A2(n20094), .ZN(n20114) );
  AOI21_X1 U22984 ( .B1(n20163), .B2(n9603), .A(n20114), .ZN(n20096) );
  OAI22_X1 U22985 ( .A1(n20096), .A2(n20574), .B1(n20094), .B2(n20638), .ZN(
        n20115) );
  AOI22_X1 U22986 ( .A1(n20577), .A2(n20115), .B1(n20576), .B2(n20114), .ZN(
        n20100) );
  INV_X1 U22987 ( .A(n20094), .ZN(n20098) );
  INV_X1 U22988 ( .A(n20156), .ZN(n20164) );
  OAI211_X1 U22989 ( .C1(n20164), .C2(n20496), .A(n20499), .B(n20096), .ZN(
        n20097) );
  OAI211_X1 U22990 ( .C1(n20499), .C2(n20098), .A(n20580), .B(n20097), .ZN(
        n20117) );
  INV_X1 U22991 ( .A(n20535), .ZN(n20583) );
  AOI22_X1 U22992 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20117), .B1(
        n20111), .B2(n20583), .ZN(n20099) );
  OAI211_X1 U22993 ( .C1(n20586), .C2(n20150), .A(n20100), .B(n20099), .ZN(
        P1_U3041) );
  AOI22_X1 U22994 ( .A1(n20588), .A2(n20115), .B1(n20587), .B2(n20114), .ZN(
        n20102) );
  INV_X1 U22995 ( .A(n20150), .ZN(n20116) );
  INV_X1 U22996 ( .A(n20592), .ZN(n20536) );
  AOI22_X1 U22997 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20536), .ZN(n20101) );
  OAI211_X1 U22998 ( .C1(n20539), .C2(n20120), .A(n20102), .B(n20101), .ZN(
        P1_U3042) );
  AOI22_X1 U22999 ( .A1(n20594), .A2(n20115), .B1(n20593), .B2(n20114), .ZN(
        n20104) );
  INV_X1 U23000 ( .A(n20543), .ZN(n20595) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20117), .B1(
        n20111), .B2(n20595), .ZN(n20103) );
  OAI211_X1 U23002 ( .C1(n20598), .C2(n20150), .A(n20104), .B(n20103), .ZN(
        P1_U3043) );
  AOI22_X1 U23003 ( .A1(n20600), .A2(n20115), .B1(n20599), .B2(n20114), .ZN(
        n20106) );
  INV_X1 U23004 ( .A(n20604), .ZN(n20544) );
  AOI22_X1 U23005 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20544), .ZN(n20105) );
  OAI211_X1 U23006 ( .C1(n20547), .C2(n20120), .A(n20106), .B(n20105), .ZN(
        P1_U3044) );
  AOI22_X1 U23007 ( .A1(n20606), .A2(n20115), .B1(n20605), .B2(n20114), .ZN(
        n20108) );
  INV_X1 U23008 ( .A(n20610), .ZN(n20548) );
  AOI22_X1 U23009 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20548), .ZN(n20107) );
  OAI211_X1 U23010 ( .C1(n20551), .C2(n20120), .A(n20108), .B(n20107), .ZN(
        P1_U3045) );
  AOI22_X1 U23011 ( .A1(n20612), .A2(n20115), .B1(n20611), .B2(n20114), .ZN(
        n20110) );
  INV_X1 U23012 ( .A(n20555), .ZN(n20613) );
  AOI22_X1 U23013 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20117), .B1(
        n20111), .B2(n20613), .ZN(n20109) );
  OAI211_X1 U23014 ( .C1(n20616), .C2(n20150), .A(n20110), .B(n20109), .ZN(
        P1_U3046) );
  AOI22_X1 U23015 ( .A1(n20618), .A2(n20115), .B1(n20617), .B2(n20114), .ZN(
        n20113) );
  INV_X1 U23016 ( .A(n20559), .ZN(n20619) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20117), .B1(
        n20111), .B2(n20619), .ZN(n20112) );
  OAI211_X1 U23018 ( .C1(n20622), .C2(n20150), .A(n20113), .B(n20112), .ZN(
        P1_U3047) );
  AOI22_X1 U23019 ( .A1(n20626), .A2(n20115), .B1(n20624), .B2(n20114), .ZN(
        n20119) );
  INV_X1 U23020 ( .A(n20633), .ZN(n20562) );
  AOI22_X1 U23021 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20117), .B1(
        n20116), .B2(n20562), .ZN(n20118) );
  OAI211_X1 U23022 ( .C1(n20567), .C2(n20120), .A(n20119), .B(n20118), .ZN(
        P1_U3048) );
  NAND2_X1 U23023 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20158), .ZN(
        n20167) );
  OR2_X1 U23024 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20167), .ZN(
        n20149) );
  OAI22_X1 U23025 ( .A1(n20150), .A2(n20535), .B1(n20442), .B2(n20149), .ZN(
        n20121) );
  INV_X1 U23026 ( .A(n20121), .ZN(n20130) );
  NAND2_X1 U23027 ( .A1(n20150), .A2(n20191), .ZN(n20122) );
  AOI21_X1 U23028 ( .B1(n20122), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20574), 
        .ZN(n20124) );
  NAND2_X1 U23029 ( .A1(n20163), .A2(n20520), .ZN(n20127) );
  AOI22_X1 U23030 ( .A1(n20124), .A2(n20127), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20149), .ZN(n20123) );
  OAI21_X1 U23031 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20375), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20254) );
  NAND3_X1 U23032 ( .A1(n20377), .A2(n20123), .A3(n20254), .ZN(n20153) );
  INV_X1 U23033 ( .A(n20124), .ZN(n20128) );
  NAND2_X1 U23034 ( .A1(n20126), .A2(n20125), .ZN(n20257) );
  OAI22_X1 U23035 ( .A1(n20128), .A2(n20127), .B1(n20379), .B2(n20257), .ZN(
        n20152) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20153), .B1(
        n20577), .B2(n20152), .ZN(n20129) );
  OAI211_X1 U23037 ( .C1(n20586), .C2(n20191), .A(n20130), .B(n20129), .ZN(
        P1_U3049) );
  OAI22_X1 U23038 ( .A1(n20150), .A2(n20539), .B1(n20149), .B2(n20459), .ZN(
        n20131) );
  INV_X1 U23039 ( .A(n20131), .ZN(n20133) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20153), .B1(
        n20588), .B2(n20152), .ZN(n20132) );
  OAI211_X1 U23041 ( .C1(n20592), .C2(n20191), .A(n20133), .B(n20132), .ZN(
        P1_U3050) );
  OAI22_X1 U23042 ( .A1(n20191), .A2(n20598), .B1(n20149), .B2(n20463), .ZN(
        n20134) );
  INV_X1 U23043 ( .A(n20134), .ZN(n20136) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20153), .B1(
        n20594), .B2(n20152), .ZN(n20135) );
  OAI211_X1 U23045 ( .C1(n20543), .C2(n20150), .A(n20136), .B(n20135), .ZN(
        P1_U3051) );
  OAI22_X1 U23046 ( .A1(n20150), .A2(n20547), .B1(n20149), .B2(n20467), .ZN(
        n20137) );
  INV_X1 U23047 ( .A(n20137), .ZN(n20139) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20153), .B1(
        n20600), .B2(n20152), .ZN(n20138) );
  OAI211_X1 U23049 ( .C1(n20604), .C2(n20191), .A(n20139), .B(n20138), .ZN(
        P1_U3052) );
  OAI22_X1 U23050 ( .A1(n20191), .A2(n20610), .B1(n20149), .B2(n20471), .ZN(
        n20140) );
  INV_X1 U23051 ( .A(n20140), .ZN(n20142) );
  AOI22_X1 U23052 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20153), .B1(
        n20606), .B2(n20152), .ZN(n20141) );
  OAI211_X1 U23053 ( .C1(n20551), .C2(n20150), .A(n20142), .B(n20141), .ZN(
        P1_U3053) );
  OAI22_X1 U23054 ( .A1(n20150), .A2(n20555), .B1(n20149), .B2(n20475), .ZN(
        n20143) );
  INV_X1 U23055 ( .A(n20143), .ZN(n20145) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20153), .B1(
        n20612), .B2(n20152), .ZN(n20144) );
  OAI211_X1 U23057 ( .C1(n20616), .C2(n20191), .A(n20145), .B(n20144), .ZN(
        P1_U3054) );
  OAI22_X1 U23058 ( .A1(n20191), .A2(n20622), .B1(n20149), .B2(n20479), .ZN(
        n20146) );
  INV_X1 U23059 ( .A(n20146), .ZN(n20148) );
  AOI22_X1 U23060 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20153), .B1(
        n20618), .B2(n20152), .ZN(n20147) );
  OAI211_X1 U23061 ( .C1(n20559), .C2(n20150), .A(n20148), .B(n20147), .ZN(
        P1_U3055) );
  OAI22_X1 U23062 ( .A1(n20150), .A2(n20567), .B1(n20149), .B2(n20484), .ZN(
        n20151) );
  INV_X1 U23063 ( .A(n20151), .ZN(n20155) );
  AOI22_X1 U23064 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20153), .B1(
        n20626), .B2(n20152), .ZN(n20154) );
  OAI211_X1 U23065 ( .C1(n20633), .C2(n20191), .A(n20155), .B(n20154), .ZN(
        P1_U3056) );
  NAND2_X1 U23066 ( .A1(n20158), .A2(n20157), .ZN(n20190) );
  OAI22_X1 U23067 ( .A1(n20191), .A2(n20535), .B1(n20442), .B2(n20190), .ZN(
        n20159) );
  INV_X1 U23068 ( .A(n20159), .ZN(n20171) );
  AND2_X1 U23069 ( .A1(n20161), .A2(n20160), .ZN(n20569) );
  INV_X1 U23070 ( .A(n20190), .ZN(n20162) );
  AOI21_X1 U23071 ( .B1(n20163), .B2(n20569), .A(n20162), .ZN(n20168) );
  AOI21_X1 U23072 ( .B1(n20164), .B2(n20499), .A(n20415), .ZN(n20169) );
  INV_X1 U23073 ( .A(n20169), .ZN(n20165) );
  AOI22_X1 U23074 ( .A1(n20168), .A2(n20165), .B1(n20574), .B2(n20167), .ZN(
        n20166) );
  NAND2_X1 U23075 ( .A1(n20580), .A2(n20166), .ZN(n20194) );
  OAI22_X1 U23076 ( .A1(n20169), .A2(n20168), .B1(n20638), .B2(n20167), .ZN(
        n20193) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20194), .B1(
        n20577), .B2(n20193), .ZN(n20170) );
  OAI211_X1 U23078 ( .C1(n20586), .C2(n20218), .A(n20171), .B(n20170), .ZN(
        P1_U3057) );
  OAI22_X1 U23079 ( .A1(n20218), .A2(n20592), .B1(n20459), .B2(n20190), .ZN(
        n20172) );
  INV_X1 U23080 ( .A(n20172), .ZN(n20174) );
  AOI22_X1 U23081 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20194), .B1(
        n20588), .B2(n20193), .ZN(n20173) );
  OAI211_X1 U23082 ( .C1(n20539), .C2(n20191), .A(n20174), .B(n20173), .ZN(
        P1_U3058) );
  OAI22_X1 U23083 ( .A1(n20218), .A2(n20598), .B1(n20463), .B2(n20190), .ZN(
        n20175) );
  INV_X1 U23084 ( .A(n20175), .ZN(n20177) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20194), .B1(
        n20594), .B2(n20193), .ZN(n20176) );
  OAI211_X1 U23086 ( .C1(n20543), .C2(n20191), .A(n20177), .B(n20176), .ZN(
        P1_U3059) );
  OAI22_X1 U23087 ( .A1(n20218), .A2(n20604), .B1(n20467), .B2(n20190), .ZN(
        n20178) );
  INV_X1 U23088 ( .A(n20178), .ZN(n20180) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20194), .B1(
        n20600), .B2(n20193), .ZN(n20179) );
  OAI211_X1 U23090 ( .C1(n20547), .C2(n20191), .A(n20180), .B(n20179), .ZN(
        P1_U3060) );
  OAI22_X1 U23091 ( .A1(n20218), .A2(n20610), .B1(n20471), .B2(n20190), .ZN(
        n20181) );
  INV_X1 U23092 ( .A(n20181), .ZN(n20183) );
  AOI22_X1 U23093 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20194), .B1(
        n20606), .B2(n20193), .ZN(n20182) );
  OAI211_X1 U23094 ( .C1(n20551), .C2(n20191), .A(n20183), .B(n20182), .ZN(
        P1_U3061) );
  OAI22_X1 U23095 ( .A1(n20218), .A2(n20616), .B1(n20475), .B2(n20190), .ZN(
        n20184) );
  INV_X1 U23096 ( .A(n20184), .ZN(n20186) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20194), .B1(
        n20612), .B2(n20193), .ZN(n20185) );
  OAI211_X1 U23098 ( .C1(n20555), .C2(n20191), .A(n20186), .B(n20185), .ZN(
        P1_U3062) );
  OAI22_X1 U23099 ( .A1(n20218), .A2(n20622), .B1(n20479), .B2(n20190), .ZN(
        n20187) );
  INV_X1 U23100 ( .A(n20187), .ZN(n20189) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20194), .B1(
        n20618), .B2(n20193), .ZN(n20188) );
  OAI211_X1 U23102 ( .C1(n20559), .C2(n20191), .A(n20189), .B(n20188), .ZN(
        P1_U3063) );
  OAI22_X1 U23103 ( .A1(n20191), .A2(n20567), .B1(n20484), .B2(n20190), .ZN(
        n20192) );
  INV_X1 U23104 ( .A(n20192), .ZN(n20196) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20194), .B1(
        n20626), .B2(n20193), .ZN(n20195) );
  OAI211_X1 U23106 ( .C1(n20633), .C2(n20218), .A(n20196), .B(n20195), .ZN(
        P1_U3064) );
  NAND3_X1 U23107 ( .A1(n9880), .A2(n20499), .A3(n20449), .ZN(n20198) );
  OAI21_X1 U23108 ( .B1(n20521), .B2(n20199), .A(n20198), .ZN(n20219) );
  AOI22_X1 U23109 ( .A1(n20577), .A2(n20219), .B1(n20576), .B2(n9875), .ZN(
        n20205) );
  AOI21_X1 U23110 ( .B1(n20244), .B2(n20218), .A(n20496), .ZN(n20200) );
  AOI21_X1 U23111 ( .B1(n9880), .B2(n20449), .A(n20200), .ZN(n20201) );
  NOR2_X1 U23112 ( .A1(n20201), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20203) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20221), .B1(
        n20220), .B2(n20583), .ZN(n20204) );
  OAI211_X1 U23114 ( .C1(n20586), .C2(n20244), .A(n20205), .B(n20204), .ZN(
        P1_U3065) );
  AOI22_X1 U23115 ( .A1(n20588), .A2(n20219), .B1(n20587), .B2(n9875), .ZN(
        n20207) );
  INV_X1 U23116 ( .A(n20539), .ZN(n20589) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20221), .B1(
        n20220), .B2(n20589), .ZN(n20206) );
  OAI211_X1 U23118 ( .C1(n20592), .C2(n20244), .A(n20207), .B(n20206), .ZN(
        P1_U3066) );
  AOI22_X1 U23119 ( .A1(n20594), .A2(n20219), .B1(n20593), .B2(n9875), .ZN(
        n20209) );
  INV_X1 U23120 ( .A(n20598), .ZN(n20540) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20221), .B1(
        n20247), .B2(n20540), .ZN(n20208) );
  OAI211_X1 U23122 ( .C1(n20543), .C2(n20218), .A(n20209), .B(n20208), .ZN(
        P1_U3067) );
  AOI22_X1 U23123 ( .A1(n20600), .A2(n20219), .B1(n20599), .B2(n9875), .ZN(
        n20211) );
  INV_X1 U23124 ( .A(n20547), .ZN(n20601) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20221), .B1(
        n20220), .B2(n20601), .ZN(n20210) );
  OAI211_X1 U23126 ( .C1(n20604), .C2(n20244), .A(n20211), .B(n20210), .ZN(
        P1_U3068) );
  AOI22_X1 U23127 ( .A1(n20606), .A2(n20219), .B1(n20605), .B2(n9875), .ZN(
        n20213) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20221), .B1(
        n20247), .B2(n20548), .ZN(n20212) );
  OAI211_X1 U23129 ( .C1(n20551), .C2(n20218), .A(n20213), .B(n20212), .ZN(
        P1_U3069) );
  AOI22_X1 U23130 ( .A1(n20612), .A2(n20219), .B1(n20611), .B2(n9875), .ZN(
        n20215) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20221), .B1(
        n20220), .B2(n20613), .ZN(n20214) );
  OAI211_X1 U23132 ( .C1(n20616), .C2(n20244), .A(n20215), .B(n20214), .ZN(
        P1_U3070) );
  AOI22_X1 U23133 ( .A1(n20618), .A2(n20219), .B1(n20617), .B2(n9875), .ZN(
        n20217) );
  INV_X1 U23134 ( .A(n20622), .ZN(n20556) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20221), .B1(
        n20247), .B2(n20556), .ZN(n20216) );
  OAI211_X1 U23136 ( .C1(n20559), .C2(n20218), .A(n20217), .B(n20216), .ZN(
        P1_U3071) );
  AOI22_X1 U23137 ( .A1(n20626), .A2(n20219), .B1(n20624), .B2(n9875), .ZN(
        n20223) );
  INV_X1 U23138 ( .A(n20567), .ZN(n20627) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20221), .B1(
        n20220), .B2(n20627), .ZN(n20222) );
  OAI211_X1 U23140 ( .C1(n20633), .C2(n20244), .A(n20223), .B(n20222), .ZN(
        P1_U3072) );
  NOR2_X1 U23141 ( .A1(n20251), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20227) );
  INV_X1 U23142 ( .A(n20227), .ZN(n20224) );
  NOR2_X1 U23143 ( .A1(n20493), .A2(n20224), .ZN(n20245) );
  AOI21_X1 U23144 ( .B1(n9880), .B2(n9603), .A(n20245), .ZN(n20225) );
  OAI22_X1 U23145 ( .A1(n20225), .A2(n20574), .B1(n20224), .B2(n20638), .ZN(
        n20246) );
  AOI22_X1 U23146 ( .A1(n20577), .A2(n20246), .B1(n20576), .B2(n20245), .ZN(
        n20230) );
  OAI211_X1 U23147 ( .C1(n20290), .C2(n20496), .A(n20499), .B(n20225), .ZN(
        n20226) );
  OAI211_X1 U23148 ( .C1(n20499), .C2(n20227), .A(n20580), .B(n20226), .ZN(
        n20248) );
  INV_X1 U23149 ( .A(n20286), .ZN(n20241) );
  INV_X1 U23150 ( .A(n20586), .ZN(n20532) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20248), .B1(
        n20241), .B2(n20532), .ZN(n20229) );
  OAI211_X1 U23152 ( .C1(n20535), .C2(n20244), .A(n20230), .B(n20229), .ZN(
        P1_U3073) );
  AOI22_X1 U23153 ( .A1(n20588), .A2(n20246), .B1(n20587), .B2(n20245), .ZN(
        n20232) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20248), .B1(
        n20247), .B2(n20589), .ZN(n20231) );
  OAI211_X1 U23155 ( .C1(n20592), .C2(n20286), .A(n20232), .B(n20231), .ZN(
        P1_U3074) );
  AOI22_X1 U23156 ( .A1(n20594), .A2(n20246), .B1(n20593), .B2(n20245), .ZN(
        n20234) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20248), .B1(
        n20247), .B2(n20595), .ZN(n20233) );
  OAI211_X1 U23158 ( .C1(n20598), .C2(n20286), .A(n20234), .B(n20233), .ZN(
        P1_U3075) );
  AOI22_X1 U23159 ( .A1(n20600), .A2(n20246), .B1(n20599), .B2(n20245), .ZN(
        n20236) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20248), .B1(
        n20247), .B2(n20601), .ZN(n20235) );
  OAI211_X1 U23161 ( .C1(n20604), .C2(n20286), .A(n20236), .B(n20235), .ZN(
        P1_U3076) );
  AOI22_X1 U23162 ( .A1(n20606), .A2(n20246), .B1(n20605), .B2(n20245), .ZN(
        n20238) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20248), .B1(
        n20241), .B2(n20548), .ZN(n20237) );
  OAI211_X1 U23164 ( .C1(n20551), .C2(n20244), .A(n20238), .B(n20237), .ZN(
        P1_U3077) );
  AOI22_X1 U23165 ( .A1(n20612), .A2(n20246), .B1(n20611), .B2(n20245), .ZN(
        n20240) );
  INV_X1 U23166 ( .A(n20616), .ZN(n20552) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20248), .B1(
        n20241), .B2(n20552), .ZN(n20239) );
  OAI211_X1 U23168 ( .C1(n20555), .C2(n20244), .A(n20240), .B(n20239), .ZN(
        P1_U3078) );
  AOI22_X1 U23169 ( .A1(n20618), .A2(n20246), .B1(n20617), .B2(n20245), .ZN(
        n20243) );
  AOI22_X1 U23170 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20248), .B1(
        n20241), .B2(n20556), .ZN(n20242) );
  OAI211_X1 U23171 ( .C1(n20559), .C2(n20244), .A(n20243), .B(n20242), .ZN(
        P1_U3079) );
  AOI22_X1 U23172 ( .A1(n20626), .A2(n20246), .B1(n20624), .B2(n20245), .ZN(
        n20250) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20248), .B1(
        n20247), .B2(n20627), .ZN(n20249) );
  OAI211_X1 U23174 ( .C1(n20633), .C2(n20286), .A(n20250), .B(n20249), .ZN(
        P1_U3080) );
  NOR2_X1 U23175 ( .A1(n20572), .A2(n20251), .ZN(n20295) );
  INV_X1 U23176 ( .A(n20295), .ZN(n20289) );
  OR2_X1 U23177 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20289), .ZN(
        n20280) );
  OAI22_X1 U23178 ( .A1(n20317), .A2(n20586), .B1(n20442), .B2(n20280), .ZN(
        n20252) );
  INV_X1 U23179 ( .A(n20252), .ZN(n20261) );
  NAND3_X1 U23180 ( .A1(n20317), .A2(n20286), .A3(n20499), .ZN(n20253) );
  NAND2_X1 U23181 ( .A1(n20253), .A2(n20445), .ZN(n20256) );
  NAND2_X1 U23182 ( .A1(n9880), .A2(n20520), .ZN(n20258) );
  AOI22_X1 U23183 ( .A1(n20256), .A2(n20258), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20280), .ZN(n20255) );
  NAND3_X1 U23184 ( .A1(n20530), .A2(n20255), .A3(n20254), .ZN(n20283) );
  INV_X1 U23185 ( .A(n20256), .ZN(n20259) );
  OAI22_X1 U23186 ( .A1(n20259), .A2(n20258), .B1(n20257), .B2(n20521), .ZN(
        n20282) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20283), .B1(
        n20577), .B2(n20282), .ZN(n20260) );
  OAI211_X1 U23188 ( .C1(n20535), .C2(n20286), .A(n20261), .B(n20260), .ZN(
        P1_U3081) );
  OAI22_X1 U23189 ( .A1(n20286), .A2(n20539), .B1(n20459), .B2(n20280), .ZN(
        n20262) );
  INV_X1 U23190 ( .A(n20262), .ZN(n20264) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20283), .B1(
        n20588), .B2(n20282), .ZN(n20263) );
  OAI211_X1 U23192 ( .C1(n20592), .C2(n20317), .A(n20264), .B(n20263), .ZN(
        P1_U3082) );
  OAI22_X1 U23193 ( .A1(n20317), .A2(n20598), .B1(n20463), .B2(n20280), .ZN(
        n20265) );
  INV_X1 U23194 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20283), .B1(
        n20594), .B2(n20282), .ZN(n20266) );
  OAI211_X1 U23196 ( .C1(n20543), .C2(n20286), .A(n20267), .B(n20266), .ZN(
        P1_U3083) );
  OAI22_X1 U23197 ( .A1(n20317), .A2(n20604), .B1(n20467), .B2(n20280), .ZN(
        n20268) );
  INV_X1 U23198 ( .A(n20268), .ZN(n20270) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20283), .B1(
        n20600), .B2(n20282), .ZN(n20269) );
  OAI211_X1 U23200 ( .C1(n20547), .C2(n20286), .A(n20270), .B(n20269), .ZN(
        P1_U3084) );
  OAI22_X1 U23201 ( .A1(n20317), .A2(n20610), .B1(n20471), .B2(n20280), .ZN(
        n20271) );
  INV_X1 U23202 ( .A(n20271), .ZN(n20273) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20283), .B1(
        n20606), .B2(n20282), .ZN(n20272) );
  OAI211_X1 U23204 ( .C1(n20551), .C2(n20286), .A(n20273), .B(n20272), .ZN(
        P1_U3085) );
  OAI22_X1 U23205 ( .A1(n20317), .A2(n20616), .B1(n20475), .B2(n20280), .ZN(
        n20274) );
  INV_X1 U23206 ( .A(n20274), .ZN(n20276) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20283), .B1(
        n20612), .B2(n20282), .ZN(n20275) );
  OAI211_X1 U23208 ( .C1(n20555), .C2(n20286), .A(n20276), .B(n20275), .ZN(
        P1_U3086) );
  OAI22_X1 U23209 ( .A1(n20317), .A2(n20622), .B1(n20479), .B2(n20280), .ZN(
        n20277) );
  INV_X1 U23210 ( .A(n20277), .ZN(n20279) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20283), .B1(
        n20618), .B2(n20282), .ZN(n20278) );
  OAI211_X1 U23212 ( .C1(n20559), .C2(n20286), .A(n20279), .B(n20278), .ZN(
        P1_U3087) );
  OAI22_X1 U23213 ( .A1(n20317), .A2(n20633), .B1(n20484), .B2(n20280), .ZN(
        n20281) );
  INV_X1 U23214 ( .A(n20281), .ZN(n20285) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20283), .B1(
        n20626), .B2(n20282), .ZN(n20284) );
  OAI211_X1 U23216 ( .C1(n20567), .C2(n20286), .A(n20285), .B(n20284), .ZN(
        P1_U3088) );
  NAND2_X1 U23217 ( .A1(n20287), .A2(n20491), .ZN(n20307) );
  INV_X1 U23218 ( .A(n20288), .ZN(n20312) );
  AOI21_X1 U23219 ( .B1(n9880), .B2(n20569), .A(n20312), .ZN(n20292) );
  OAI22_X1 U23220 ( .A1(n20292), .A2(n20574), .B1(n20289), .B2(n20638), .ZN(
        n20313) );
  AOI22_X1 U23221 ( .A1(n20577), .A2(n20313), .B1(n20312), .B2(n20576), .ZN(
        n20297) );
  INV_X1 U23222 ( .A(n20290), .ZN(n20291) );
  NOR2_X1 U23223 ( .A1(n20291), .A2(n20574), .ZN(n20293) );
  OAI21_X1 U23224 ( .B1(n20293), .B2(n20415), .A(n20292), .ZN(n20294) );
  OAI211_X1 U23225 ( .C1(n20499), .C2(n20295), .A(n20580), .B(n20294), .ZN(
        n20314) );
  INV_X1 U23226 ( .A(n20317), .ZN(n20304) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20314), .B1(
        n20304), .B2(n20583), .ZN(n20296) );
  OAI211_X1 U23228 ( .C1(n20586), .C2(n20307), .A(n20297), .B(n20296), .ZN(
        P1_U3089) );
  AOI22_X1 U23229 ( .A1(n20588), .A2(n20313), .B1(n20312), .B2(n20587), .ZN(
        n20299) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20314), .B1(
        n20304), .B2(n20589), .ZN(n20298) );
  OAI211_X1 U23231 ( .C1(n20592), .C2(n20307), .A(n20299), .B(n20298), .ZN(
        P1_U3090) );
  AOI22_X1 U23232 ( .A1(n20594), .A2(n20313), .B1(n20312), .B2(n20593), .ZN(
        n20301) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20314), .B1(
        n20304), .B2(n20595), .ZN(n20300) );
  OAI211_X1 U23234 ( .C1(n20598), .C2(n20307), .A(n20301), .B(n20300), .ZN(
        P1_U3091) );
  AOI22_X1 U23235 ( .A1(n20600), .A2(n20313), .B1(n20312), .B2(n20599), .ZN(
        n20303) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20314), .B1(
        n20341), .B2(n20544), .ZN(n20302) );
  OAI211_X1 U23237 ( .C1(n20547), .C2(n20317), .A(n20303), .B(n20302), .ZN(
        P1_U3092) );
  AOI22_X1 U23238 ( .A1(n20606), .A2(n20313), .B1(n20312), .B2(n20605), .ZN(
        n20306) );
  INV_X1 U23239 ( .A(n20551), .ZN(n20607) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20314), .B1(
        n20304), .B2(n20607), .ZN(n20305) );
  OAI211_X1 U23241 ( .C1(n20610), .C2(n20307), .A(n20306), .B(n20305), .ZN(
        P1_U3093) );
  AOI22_X1 U23242 ( .A1(n20612), .A2(n20313), .B1(n20312), .B2(n20611), .ZN(
        n20309) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20314), .B1(
        n20341), .B2(n20552), .ZN(n20308) );
  OAI211_X1 U23244 ( .C1(n20555), .C2(n20317), .A(n20309), .B(n20308), .ZN(
        P1_U3094) );
  AOI22_X1 U23245 ( .A1(n20618), .A2(n20313), .B1(n20312), .B2(n20617), .ZN(
        n20311) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20314), .B1(
        n20341), .B2(n20556), .ZN(n20310) );
  OAI211_X1 U23247 ( .C1(n20559), .C2(n20317), .A(n20311), .B(n20310), .ZN(
        P1_U3095) );
  AOI22_X1 U23248 ( .A1(n20626), .A2(n20313), .B1(n20312), .B2(n20624), .ZN(
        n20316) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20314), .B1(
        n20341), .B2(n20562), .ZN(n20315) );
  OAI211_X1 U23250 ( .C1(n20567), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        P1_U3096) );
  NAND2_X1 U23251 ( .A1(n20413), .A2(n20318), .ZN(n20350) );
  NAND2_X1 U23252 ( .A1(n20319), .A2(n20448), .ZN(n20374) );
  INV_X1 U23253 ( .A(n20374), .ZN(n20411) );
  NAND2_X1 U23254 ( .A1(n20320), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20410) );
  AOI21_X1 U23255 ( .B1(n20411), .B2(n20449), .A(n9879), .ZN(n20323) );
  NAND2_X1 U23256 ( .A1(n20321), .A2(n20375), .ZN(n20454) );
  OAI22_X1 U23257 ( .A1(n20323), .A2(n20574), .B1(n20379), .B2(n20454), .ZN(
        n20340) );
  AOI22_X1 U23258 ( .A1(n20577), .A2(n20340), .B1(n9879), .B2(n20576), .ZN(
        n20327) );
  INV_X1 U23259 ( .A(n20371), .ZN(n20322) );
  OAI21_X1 U23260 ( .B1(n20322), .B2(n20341), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20324) );
  NAND2_X1 U23261 ( .A1(n20324), .A2(n20323), .ZN(n20325) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20583), .ZN(n20326) );
  OAI211_X1 U23263 ( .C1(n20586), .C2(n20371), .A(n20327), .B(n20326), .ZN(
        P1_U3097) );
  AOI22_X1 U23264 ( .A1(n20588), .A2(n20340), .B1(n9879), .B2(n20587), .ZN(
        n20329) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20589), .ZN(n20328) );
  OAI211_X1 U23266 ( .C1(n20592), .C2(n20371), .A(n20329), .B(n20328), .ZN(
        P1_U3098) );
  AOI22_X1 U23267 ( .A1(n20594), .A2(n20340), .B1(n9879), .B2(n20593), .ZN(
        n20331) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20595), .ZN(n20330) );
  OAI211_X1 U23269 ( .C1(n20598), .C2(n20371), .A(n20331), .B(n20330), .ZN(
        P1_U3099) );
  AOI22_X1 U23270 ( .A1(n20600), .A2(n20340), .B1(n9879), .B2(n20599), .ZN(
        n20333) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20601), .ZN(n20332) );
  OAI211_X1 U23272 ( .C1(n20604), .C2(n20371), .A(n20333), .B(n20332), .ZN(
        P1_U3100) );
  AOI22_X1 U23273 ( .A1(n20606), .A2(n20340), .B1(n9879), .B2(n20605), .ZN(
        n20335) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20607), .ZN(n20334) );
  OAI211_X1 U23275 ( .C1(n20610), .C2(n20371), .A(n20335), .B(n20334), .ZN(
        P1_U3101) );
  AOI22_X1 U23276 ( .A1(n20612), .A2(n20340), .B1(n9879), .B2(n20611), .ZN(
        n20337) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20613), .ZN(n20336) );
  OAI211_X1 U23278 ( .C1(n20616), .C2(n20371), .A(n20337), .B(n20336), .ZN(
        P1_U3102) );
  AOI22_X1 U23279 ( .A1(n20618), .A2(n20340), .B1(n9879), .B2(n20617), .ZN(
        n20339) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20619), .ZN(n20338) );
  OAI211_X1 U23281 ( .C1(n20622), .C2(n20371), .A(n20339), .B(n20338), .ZN(
        P1_U3103) );
  AOI22_X1 U23282 ( .A1(n20626), .A2(n20340), .B1(n9879), .B2(n20624), .ZN(
        n20344) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20342), .B1(
        n20341), .B2(n20627), .ZN(n20343) );
  OAI211_X1 U23284 ( .C1(n20633), .C2(n20371), .A(n20344), .B(n20343), .ZN(
        P1_U3104) );
  NOR2_X1 U23285 ( .A1(n20410), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20349) );
  INV_X1 U23286 ( .A(n20349), .ZN(n20345) );
  NOR2_X1 U23287 ( .A1(n20493), .A2(n20345), .ZN(n20365) );
  AOI21_X1 U23288 ( .B1(n20411), .B2(n9603), .A(n20365), .ZN(n20346) );
  OAI22_X1 U23289 ( .A1(n20346), .A2(n20574), .B1(n20345), .B2(n20638), .ZN(
        n20366) );
  AOI22_X1 U23290 ( .A1(n20577), .A2(n20366), .B1(n20576), .B2(n20365), .ZN(
        n20352) );
  INV_X1 U23291 ( .A(n20413), .ZN(n20347) );
  OAI211_X1 U23292 ( .C1(n20347), .C2(n20496), .A(n20499), .B(n20346), .ZN(
        n20348) );
  OAI211_X1 U23293 ( .C1(n20499), .C2(n20349), .A(n20580), .B(n20348), .ZN(
        n20368) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20532), .ZN(n20351) );
  OAI211_X1 U23295 ( .C1(n20535), .C2(n20371), .A(n20352), .B(n20351), .ZN(
        P1_U3105) );
  AOI22_X1 U23296 ( .A1(n20588), .A2(n20366), .B1(n20587), .B2(n20365), .ZN(
        n20354) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20536), .ZN(n20353) );
  OAI211_X1 U23298 ( .C1(n20539), .C2(n20371), .A(n20354), .B(n20353), .ZN(
        P1_U3106) );
  AOI22_X1 U23299 ( .A1(n20594), .A2(n20366), .B1(n20593), .B2(n20365), .ZN(
        n20356) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20540), .ZN(n20355) );
  OAI211_X1 U23301 ( .C1(n20543), .C2(n20371), .A(n20356), .B(n20355), .ZN(
        P1_U3107) );
  AOI22_X1 U23302 ( .A1(n20600), .A2(n20366), .B1(n20599), .B2(n20365), .ZN(
        n20358) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20544), .ZN(n20357) );
  OAI211_X1 U23304 ( .C1(n20547), .C2(n20371), .A(n20358), .B(n20357), .ZN(
        P1_U3108) );
  AOI22_X1 U23305 ( .A1(n20606), .A2(n20366), .B1(n20605), .B2(n20365), .ZN(
        n20360) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20548), .ZN(n20359) );
  OAI211_X1 U23307 ( .C1(n20551), .C2(n20371), .A(n20360), .B(n20359), .ZN(
        P1_U3109) );
  AOI22_X1 U23308 ( .A1(n20612), .A2(n20366), .B1(n20611), .B2(n20365), .ZN(
        n20362) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20552), .ZN(n20361) );
  OAI211_X1 U23310 ( .C1(n20555), .C2(n20371), .A(n20362), .B(n20361), .ZN(
        P1_U3110) );
  AOI22_X1 U23311 ( .A1(n20618), .A2(n20366), .B1(n20617), .B2(n20365), .ZN(
        n20364) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20556), .ZN(n20363) );
  OAI211_X1 U23313 ( .C1(n20559), .C2(n20371), .A(n20364), .B(n20363), .ZN(
        P1_U3111) );
  AOI22_X1 U23314 ( .A1(n20626), .A2(n20366), .B1(n20624), .B2(n20365), .ZN(
        n20370) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20368), .B1(
        n20367), .B2(n20562), .ZN(n20369) );
  OAI211_X1 U23316 ( .C1(n20567), .C2(n20371), .A(n20370), .B(n20369), .ZN(
        P1_U3112) );
  NOR2_X1 U23317 ( .A1(n20572), .A2(n20410), .ZN(n20418) );
  INV_X1 U23318 ( .A(n20418), .ZN(n20412) );
  OR2_X1 U23319 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20412), .ZN(
        n20402) );
  OAI22_X1 U23320 ( .A1(n20408), .A2(n20535), .B1(n20442), .B2(n20402), .ZN(
        n20372) );
  INV_X1 U23321 ( .A(n20372), .ZN(n20383) );
  NAND3_X1 U23322 ( .A1(n20408), .A2(n20499), .A3(n20432), .ZN(n20373) );
  NAND2_X1 U23323 ( .A1(n20373), .A2(n20445), .ZN(n20378) );
  OR2_X1 U23324 ( .A1(n20374), .A2(n20449), .ZN(n20380) );
  AOI22_X1 U23325 ( .A1(n20378), .A2(n20380), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20402), .ZN(n20376) );
  OR2_X1 U23326 ( .A1(n20375), .A2(n20125), .ZN(n20522) );
  NAND2_X1 U23327 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20522), .ZN(n20529) );
  NAND3_X1 U23328 ( .A1(n20377), .A2(n20376), .A3(n20529), .ZN(n20405) );
  INV_X1 U23329 ( .A(n20378), .ZN(n20381) );
  OAI22_X1 U23330 ( .A1(n20381), .A2(n20380), .B1(n20379), .B2(n20522), .ZN(
        n20404) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20405), .B1(
        n20577), .B2(n20404), .ZN(n20382) );
  OAI211_X1 U23332 ( .C1(n20586), .C2(n20432), .A(n20383), .B(n20382), .ZN(
        P1_U3113) );
  OAI22_X1 U23333 ( .A1(n20432), .A2(n20592), .B1(n20459), .B2(n20402), .ZN(
        n20384) );
  INV_X1 U23334 ( .A(n20384), .ZN(n20386) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20405), .B1(
        n20588), .B2(n20404), .ZN(n20385) );
  OAI211_X1 U23336 ( .C1(n20539), .C2(n20408), .A(n20386), .B(n20385), .ZN(
        P1_U3114) );
  OAI22_X1 U23337 ( .A1(n20408), .A2(n20543), .B1(n20402), .B2(n20463), .ZN(
        n20387) );
  INV_X1 U23338 ( .A(n20387), .ZN(n20389) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20405), .B1(
        n20594), .B2(n20404), .ZN(n20388) );
  OAI211_X1 U23340 ( .C1(n20598), .C2(n20432), .A(n20389), .B(n20388), .ZN(
        P1_U3115) );
  OAI22_X1 U23341 ( .A1(n20432), .A2(n20604), .B1(n20467), .B2(n20402), .ZN(
        n20390) );
  INV_X1 U23342 ( .A(n20390), .ZN(n20392) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20405), .B1(
        n20600), .B2(n20404), .ZN(n20391) );
  OAI211_X1 U23344 ( .C1(n20547), .C2(n20408), .A(n20392), .B(n20391), .ZN(
        P1_U3116) );
  OAI22_X1 U23345 ( .A1(n20408), .A2(n20551), .B1(n20402), .B2(n20471), .ZN(
        n20393) );
  INV_X1 U23346 ( .A(n20393), .ZN(n20395) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20405), .B1(
        n20606), .B2(n20404), .ZN(n20394) );
  OAI211_X1 U23348 ( .C1(n20610), .C2(n20432), .A(n20395), .B(n20394), .ZN(
        P1_U3117) );
  OAI22_X1 U23349 ( .A1(n20408), .A2(n20555), .B1(n20475), .B2(n20402), .ZN(
        n20396) );
  INV_X1 U23350 ( .A(n20396), .ZN(n20398) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20405), .B1(
        n20612), .B2(n20404), .ZN(n20397) );
  OAI211_X1 U23352 ( .C1(n20616), .C2(n20432), .A(n20398), .B(n20397), .ZN(
        P1_U3118) );
  OAI22_X1 U23353 ( .A1(n20432), .A2(n20622), .B1(n20402), .B2(n20479), .ZN(
        n20399) );
  INV_X1 U23354 ( .A(n20399), .ZN(n20401) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20405), .B1(
        n20618), .B2(n20404), .ZN(n20400) );
  OAI211_X1 U23356 ( .C1(n20559), .C2(n20408), .A(n20401), .B(n20400), .ZN(
        P1_U3119) );
  OAI22_X1 U23357 ( .A1(n20432), .A2(n20633), .B1(n20484), .B2(n20402), .ZN(
        n20403) );
  INV_X1 U23358 ( .A(n20403), .ZN(n20407) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20405), .B1(
        n20626), .B2(n20404), .ZN(n20406) );
  OAI211_X1 U23360 ( .C1(n20567), .C2(n20408), .A(n20407), .B(n20406), .ZN(
        P1_U3120) );
  NOR2_X1 U23361 ( .A1(n20568), .A2(n20410), .ZN(n20435) );
  AOI21_X1 U23362 ( .B1(n20411), .B2(n20569), .A(n20435), .ZN(n20414) );
  OAI22_X1 U23363 ( .A1(n20414), .A2(n20574), .B1(n20412), .B2(n20638), .ZN(
        n20436) );
  AOI22_X1 U23364 ( .A1(n20577), .A2(n20436), .B1(n20576), .B2(n20435), .ZN(
        n20420) );
  NOR2_X1 U23365 ( .A1(n20413), .A2(n20574), .ZN(n20416) );
  OAI21_X1 U23366 ( .B1(n20416), .B2(n20415), .A(n20414), .ZN(n20417) );
  OAI211_X1 U23367 ( .C1(n20499), .C2(n20418), .A(n20580), .B(n20417), .ZN(
        n20438) );
  INV_X1 U23368 ( .A(n20432), .ZN(n20437) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20583), .ZN(n20419) );
  OAI211_X1 U23370 ( .C1(n20586), .C2(n20490), .A(n20420), .B(n20419), .ZN(
        P1_U3121) );
  AOI22_X1 U23371 ( .A1(n20588), .A2(n20436), .B1(n20587), .B2(n20435), .ZN(
        n20422) );
  INV_X1 U23372 ( .A(n20490), .ZN(n20429) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20438), .B1(
        n20429), .B2(n20536), .ZN(n20421) );
  OAI211_X1 U23374 ( .C1(n20539), .C2(n20432), .A(n20422), .B(n20421), .ZN(
        P1_U3122) );
  AOI22_X1 U23375 ( .A1(n20594), .A2(n20436), .B1(n20593), .B2(n20435), .ZN(
        n20424) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20438), .B1(
        n20429), .B2(n20540), .ZN(n20423) );
  OAI211_X1 U23377 ( .C1(n20543), .C2(n20432), .A(n20424), .B(n20423), .ZN(
        P1_U3123) );
  AOI22_X1 U23378 ( .A1(n20600), .A2(n20436), .B1(n20599), .B2(n20435), .ZN(
        n20426) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20601), .ZN(n20425) );
  OAI211_X1 U23380 ( .C1(n20604), .C2(n20490), .A(n20426), .B(n20425), .ZN(
        P1_U3124) );
  AOI22_X1 U23381 ( .A1(n20606), .A2(n20436), .B1(n20605), .B2(n20435), .ZN(
        n20428) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20438), .B1(
        n20429), .B2(n20548), .ZN(n20427) );
  OAI211_X1 U23383 ( .C1(n20551), .C2(n20432), .A(n20428), .B(n20427), .ZN(
        P1_U3125) );
  AOI22_X1 U23384 ( .A1(n20612), .A2(n20436), .B1(n20611), .B2(n20435), .ZN(
        n20431) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20438), .B1(
        n20429), .B2(n20552), .ZN(n20430) );
  OAI211_X1 U23386 ( .C1(n20555), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P1_U3126) );
  AOI22_X1 U23387 ( .A1(n20618), .A2(n20436), .B1(n20617), .B2(n20435), .ZN(
        n20434) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20619), .ZN(n20433) );
  OAI211_X1 U23389 ( .C1(n20622), .C2(n20490), .A(n20434), .B(n20433), .ZN(
        P1_U3127) );
  AOI22_X1 U23390 ( .A1(n20626), .A2(n20436), .B1(n20624), .B2(n20435), .ZN(
        n20440) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20438), .B1(
        n20437), .B2(n20627), .ZN(n20439) );
  OAI211_X1 U23392 ( .C1(n20633), .C2(n20490), .A(n20440), .B(n20439), .ZN(
        P1_U3128) );
  NAND2_X1 U23393 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20571) );
  OR2_X1 U23394 ( .A1(n20441), .A2(n20571), .ZN(n20483) );
  NOR2_X1 U23395 ( .A1(n20442), .A2(n20483), .ZN(n20443) );
  AOI21_X1 U23396 ( .B1(n20516), .B2(n20532), .A(n20443), .ZN(n20458) );
  INV_X1 U23397 ( .A(n20483), .ZN(n20452) );
  INV_X1 U23398 ( .A(n20516), .ZN(n20444) );
  NAND3_X1 U23399 ( .A1(n20444), .A2(n20499), .A3(n20490), .ZN(n20446) );
  NAND2_X1 U23400 ( .A1(n20446), .A2(n20445), .ZN(n20453) );
  NOR2_X1 U23401 ( .A1(n20448), .A2(n20447), .ZN(n20570) );
  NAND2_X1 U23402 ( .A1(n20570), .A2(n20449), .ZN(n20455) );
  AOI22_X1 U23403 ( .A1(n20453), .A2(n20455), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20454), .ZN(n20450) );
  OAI211_X1 U23404 ( .C1(n20452), .C2(n20451), .A(n20530), .B(n20450), .ZN(
        n20487) );
  INV_X1 U23405 ( .A(n20453), .ZN(n20456) );
  OAI22_X1 U23406 ( .A1(n20456), .A2(n20455), .B1(n20454), .B2(n20521), .ZN(
        n20486) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20487), .B1(
        n20577), .B2(n20486), .ZN(n20457) );
  OAI211_X1 U23408 ( .C1(n20535), .C2(n20490), .A(n20458), .B(n20457), .ZN(
        P1_U3129) );
  NOR2_X1 U23409 ( .A1(n20459), .A2(n20483), .ZN(n20460) );
  AOI21_X1 U23410 ( .B1(n20516), .B2(n20536), .A(n20460), .ZN(n20462) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20487), .B1(
        n20588), .B2(n20486), .ZN(n20461) );
  OAI211_X1 U23412 ( .C1(n20539), .C2(n20490), .A(n20462), .B(n20461), .ZN(
        P1_U3130) );
  NOR2_X1 U23413 ( .A1(n20463), .A2(n20483), .ZN(n20464) );
  AOI21_X1 U23414 ( .B1(n20516), .B2(n20540), .A(n20464), .ZN(n20466) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20487), .B1(
        n20594), .B2(n20486), .ZN(n20465) );
  OAI211_X1 U23416 ( .C1(n20543), .C2(n20490), .A(n20466), .B(n20465), .ZN(
        P1_U3131) );
  NOR2_X1 U23417 ( .A1(n20467), .A2(n20483), .ZN(n20468) );
  AOI21_X1 U23418 ( .B1(n20516), .B2(n20544), .A(n20468), .ZN(n20470) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20487), .B1(
        n20600), .B2(n20486), .ZN(n20469) );
  OAI211_X1 U23420 ( .C1(n20547), .C2(n20490), .A(n20470), .B(n20469), .ZN(
        P1_U3132) );
  NOR2_X1 U23421 ( .A1(n20471), .A2(n20483), .ZN(n20472) );
  AOI21_X1 U23422 ( .B1(n20516), .B2(n20548), .A(n20472), .ZN(n20474) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20487), .B1(
        n20606), .B2(n20486), .ZN(n20473) );
  OAI211_X1 U23424 ( .C1(n20551), .C2(n20490), .A(n20474), .B(n20473), .ZN(
        P1_U3133) );
  NOR2_X1 U23425 ( .A1(n20475), .A2(n20483), .ZN(n20476) );
  AOI21_X1 U23426 ( .B1(n20516), .B2(n20552), .A(n20476), .ZN(n20478) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20487), .B1(
        n20612), .B2(n20486), .ZN(n20477) );
  OAI211_X1 U23428 ( .C1(n20555), .C2(n20490), .A(n20478), .B(n20477), .ZN(
        P1_U3134) );
  NOR2_X1 U23429 ( .A1(n20479), .A2(n20483), .ZN(n20480) );
  AOI21_X1 U23430 ( .B1(n20516), .B2(n20556), .A(n20480), .ZN(n20482) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20487), .B1(
        n20618), .B2(n20486), .ZN(n20481) );
  OAI211_X1 U23432 ( .C1(n20559), .C2(n20490), .A(n20482), .B(n20481), .ZN(
        P1_U3135) );
  NOR2_X1 U23433 ( .A1(n20484), .A2(n20483), .ZN(n20485) );
  AOI21_X1 U23434 ( .B1(n20516), .B2(n20562), .A(n20485), .ZN(n20489) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20487), .B1(
        n20626), .B2(n20486), .ZN(n20488) );
  OAI211_X1 U23436 ( .C1(n20567), .C2(n20490), .A(n20489), .B(n20488), .ZN(
        P1_U3136) );
  AOI21_X1 U23437 ( .B1(n20570), .B2(n9603), .A(n20514), .ZN(n20495) );
  NOR2_X1 U23438 ( .A1(n20571), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20498) );
  INV_X1 U23439 ( .A(n20498), .ZN(n20494) );
  OAI22_X1 U23440 ( .A1(n20495), .A2(n20574), .B1(n20494), .B2(n20638), .ZN(
        n20515) );
  AOI22_X1 U23441 ( .A1(n20577), .A2(n20515), .B1(n20576), .B2(n20514), .ZN(
        n20501) );
  OAI21_X1 U23442 ( .B1(n20525), .B2(n20496), .A(n20495), .ZN(n20497) );
  OAI221_X1 U23443 ( .B1(n20499), .B2(n20498), .C1(n20574), .C2(n20497), .A(
        n20580), .ZN(n20517) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20583), .ZN(n20500) );
  OAI211_X1 U23445 ( .C1(n20586), .C2(n20566), .A(n20501), .B(n20500), .ZN(
        P1_U3137) );
  AOI22_X1 U23446 ( .A1(n20588), .A2(n20515), .B1(n20587), .B2(n20514), .ZN(
        n20503) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20589), .ZN(n20502) );
  OAI211_X1 U23448 ( .C1(n20592), .C2(n20566), .A(n20503), .B(n20502), .ZN(
        P1_U3138) );
  AOI22_X1 U23449 ( .A1(n20594), .A2(n20515), .B1(n20593), .B2(n20514), .ZN(
        n20505) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20595), .ZN(n20504) );
  OAI211_X1 U23451 ( .C1(n20598), .C2(n20566), .A(n20505), .B(n20504), .ZN(
        P1_U3139) );
  AOI22_X1 U23452 ( .A1(n20600), .A2(n20515), .B1(n20599), .B2(n20514), .ZN(
        n20507) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20601), .ZN(n20506) );
  OAI211_X1 U23454 ( .C1(n20604), .C2(n20566), .A(n20507), .B(n20506), .ZN(
        P1_U3140) );
  AOI22_X1 U23455 ( .A1(n20606), .A2(n20515), .B1(n20605), .B2(n20514), .ZN(
        n20509) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20607), .ZN(n20508) );
  OAI211_X1 U23457 ( .C1(n20610), .C2(n20566), .A(n20509), .B(n20508), .ZN(
        P1_U3141) );
  AOI22_X1 U23458 ( .A1(n20612), .A2(n20515), .B1(n20611), .B2(n20514), .ZN(
        n20511) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20613), .ZN(n20510) );
  OAI211_X1 U23460 ( .C1(n20616), .C2(n20566), .A(n20511), .B(n20510), .ZN(
        P1_U3142) );
  AOI22_X1 U23461 ( .A1(n20618), .A2(n20515), .B1(n20617), .B2(n20514), .ZN(
        n20513) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20619), .ZN(n20512) );
  OAI211_X1 U23463 ( .C1(n20622), .C2(n20566), .A(n20513), .B(n20512), .ZN(
        P1_U3143) );
  AOI22_X1 U23464 ( .A1(n20626), .A2(n20515), .B1(n20624), .B2(n20514), .ZN(
        n20519) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20517), .B1(
        n20516), .B2(n20627), .ZN(n20518) );
  OAI211_X1 U23466 ( .C1(n20633), .C2(n20566), .A(n20519), .B(n20518), .ZN(
        P1_U3144) );
  NAND2_X1 U23467 ( .A1(n20570), .A2(n20520), .ZN(n20527) );
  OAI22_X1 U23468 ( .A1(n20527), .A2(n20574), .B1(n20522), .B2(n20521), .ZN(
        n20561) );
  NOR3_X2 U23469 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20572), .A3(
        n20571), .ZN(n20560) );
  AOI22_X1 U23470 ( .A1(n20577), .A2(n20561), .B1(n20576), .B2(n20560), .ZN(
        n20534) );
  INV_X1 U23471 ( .A(n20566), .ZN(n20526) );
  INV_X1 U23472 ( .A(n20523), .ZN(n20524) );
  NOR2_X2 U23473 ( .A1(n20525), .A2(n20524), .ZN(n20628) );
  OAI21_X1 U23474 ( .B1(n20526), .B2(n20628), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20528) );
  AOI21_X1 U23475 ( .B1(n20528), .B2(n20527), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20531) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20532), .ZN(n20533) );
  OAI211_X1 U23477 ( .C1(n20535), .C2(n20566), .A(n20534), .B(n20533), .ZN(
        P1_U3145) );
  AOI22_X1 U23478 ( .A1(n20588), .A2(n20561), .B1(n20587), .B2(n20560), .ZN(
        n20538) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20536), .ZN(n20537) );
  OAI211_X1 U23480 ( .C1(n20539), .C2(n20566), .A(n20538), .B(n20537), .ZN(
        P1_U3146) );
  AOI22_X1 U23481 ( .A1(n20594), .A2(n20561), .B1(n20593), .B2(n20560), .ZN(
        n20542) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20540), .ZN(n20541) );
  OAI211_X1 U23483 ( .C1(n20543), .C2(n20566), .A(n20542), .B(n20541), .ZN(
        P1_U3147) );
  AOI22_X1 U23484 ( .A1(n20600), .A2(n20561), .B1(n20599), .B2(n20560), .ZN(
        n20546) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20544), .ZN(n20545) );
  OAI211_X1 U23486 ( .C1(n20547), .C2(n20566), .A(n20546), .B(n20545), .ZN(
        P1_U3148) );
  AOI22_X1 U23487 ( .A1(n20606), .A2(n20561), .B1(n20605), .B2(n20560), .ZN(
        n20550) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20548), .ZN(n20549) );
  OAI211_X1 U23489 ( .C1(n20551), .C2(n20566), .A(n20550), .B(n20549), .ZN(
        P1_U3149) );
  AOI22_X1 U23490 ( .A1(n20612), .A2(n20561), .B1(n20611), .B2(n20560), .ZN(
        n20554) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20552), .ZN(n20553) );
  OAI211_X1 U23492 ( .C1(n20555), .C2(n20566), .A(n20554), .B(n20553), .ZN(
        P1_U3150) );
  AOI22_X1 U23493 ( .A1(n20618), .A2(n20561), .B1(n20617), .B2(n20560), .ZN(
        n20558) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20556), .ZN(n20557) );
  OAI211_X1 U23495 ( .C1(n20559), .C2(n20566), .A(n20558), .B(n20557), .ZN(
        P1_U3151) );
  AOI22_X1 U23496 ( .A1(n20626), .A2(n20561), .B1(n20624), .B2(n20560), .ZN(
        n20565) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20563), .B1(
        n20628), .B2(n20562), .ZN(n20564) );
  OAI211_X1 U23498 ( .C1(n20567), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P1_U3152) );
  NOR2_X1 U23499 ( .A1(n20568), .A2(n20571), .ZN(n20623) );
  AOI21_X1 U23500 ( .B1(n20570), .B2(n20569), .A(n20623), .ZN(n20575) );
  NOR2_X1 U23501 ( .A1(n20572), .A2(n20571), .ZN(n20581) );
  INV_X1 U23502 ( .A(n20581), .ZN(n20573) );
  OAI22_X1 U23503 ( .A1(n20575), .A2(n20574), .B1(n20573), .B2(n20638), .ZN(
        n20625) );
  AOI22_X1 U23504 ( .A1(n20577), .A2(n20625), .B1(n20576), .B2(n20623), .ZN(
        n20585) );
  AND2_X1 U23505 ( .A1(n20579), .A2(n20578), .ZN(n20582) );
  OAI21_X1 U23506 ( .B1(n20582), .B2(n20581), .A(n20580), .ZN(n20629) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20583), .ZN(n20584) );
  OAI211_X1 U23508 ( .C1(n20586), .C2(n20632), .A(n20585), .B(n20584), .ZN(
        P1_U3153) );
  AOI22_X1 U23509 ( .A1(n20588), .A2(n20625), .B1(n20587), .B2(n20623), .ZN(
        n20591) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20589), .ZN(n20590) );
  OAI211_X1 U23511 ( .C1(n20592), .C2(n20632), .A(n20591), .B(n20590), .ZN(
        P1_U3154) );
  AOI22_X1 U23512 ( .A1(n20594), .A2(n20625), .B1(n20593), .B2(n20623), .ZN(
        n20597) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20595), .ZN(n20596) );
  OAI211_X1 U23514 ( .C1(n20598), .C2(n20632), .A(n20597), .B(n20596), .ZN(
        P1_U3155) );
  AOI22_X1 U23515 ( .A1(n20600), .A2(n20625), .B1(n20599), .B2(n20623), .ZN(
        n20603) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20601), .ZN(n20602) );
  OAI211_X1 U23517 ( .C1(n20604), .C2(n20632), .A(n20603), .B(n20602), .ZN(
        P1_U3156) );
  AOI22_X1 U23518 ( .A1(n20606), .A2(n20625), .B1(n20605), .B2(n20623), .ZN(
        n20609) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20607), .ZN(n20608) );
  OAI211_X1 U23520 ( .C1(n20610), .C2(n20632), .A(n20609), .B(n20608), .ZN(
        P1_U3157) );
  AOI22_X1 U23521 ( .A1(n20612), .A2(n20625), .B1(n20611), .B2(n20623), .ZN(
        n20615) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20613), .ZN(n20614) );
  OAI211_X1 U23523 ( .C1(n20616), .C2(n20632), .A(n20615), .B(n20614), .ZN(
        P1_U3158) );
  AOI22_X1 U23524 ( .A1(n20618), .A2(n20625), .B1(n20617), .B2(n20623), .ZN(
        n20621) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20619), .ZN(n20620) );
  OAI211_X1 U23526 ( .C1(n20622), .C2(n20632), .A(n20621), .B(n20620), .ZN(
        P1_U3159) );
  AOI22_X1 U23527 ( .A1(n20626), .A2(n20625), .B1(n20624), .B2(n20623), .ZN(
        n20631) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20627), .ZN(n20630) );
  OAI211_X1 U23529 ( .C1(n20633), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P1_U3160) );
  NOR2_X1 U23530 ( .A1(n20635), .A2(n20634), .ZN(n20639) );
  INV_X1 U23531 ( .A(n20636), .ZN(n20637) );
  OAI21_X1 U23532 ( .B1(n20639), .B2(n20638), .A(n20637), .ZN(P1_U3163) );
  AND2_X1 U23533 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20717), .ZN(
        P1_U3164) );
  AND2_X1 U23534 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20717), .ZN(
        P1_U3165) );
  AND2_X1 U23535 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20717), .ZN(
        P1_U3166) );
  AND2_X1 U23536 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20717), .ZN(
        P1_U3167) );
  AND2_X1 U23537 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20717), .ZN(
        P1_U3168) );
  AND2_X1 U23538 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20717), .ZN(
        P1_U3169) );
  AND2_X1 U23539 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20717), .ZN(
        P1_U3170) );
  AND2_X1 U23540 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20717), .ZN(
        P1_U3171) );
  AND2_X1 U23541 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20717), .ZN(
        P1_U3172) );
  AND2_X1 U23542 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20717), .ZN(
        P1_U3173) );
  AND2_X1 U23543 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20717), .ZN(
        P1_U3174) );
  AND2_X1 U23544 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20717), .ZN(
        P1_U3175) );
  AND2_X1 U23545 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20717), .ZN(
        P1_U3176) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20717), .ZN(
        P1_U3177) );
  AND2_X1 U23547 ( .A1(n20717), .A2(P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(
        P1_U3178) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20717), .ZN(
        P1_U3179) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20717), .ZN(
        P1_U3180) );
  AND2_X1 U23550 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20717), .ZN(
        P1_U3181) );
  AND2_X1 U23551 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20717), .ZN(
        P1_U3182) );
  AND2_X1 U23552 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20717), .ZN(
        P1_U3183) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20717), .ZN(
        P1_U3184) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20717), .ZN(
        P1_U3185) );
  AND2_X1 U23555 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20717), .ZN(P1_U3186) );
  AND2_X1 U23556 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20717), .ZN(P1_U3187) );
  AND2_X1 U23557 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20717), .ZN(P1_U3188) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20717), .ZN(P1_U3189) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20717), .ZN(P1_U3190) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20717), .ZN(P1_U3191) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20717), .ZN(P1_U3192) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20717), .ZN(P1_U3193) );
  AND2_X1 U23563 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20640), .ZN(n20652) );
  OAI21_X1 U23564 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20646), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20641) );
  AOI211_X1 U23565 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20642), .B(
        n20641), .ZN(n20643) );
  OAI22_X1 U23566 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20652), .B1(n20750), 
        .B2(n20643), .ZN(P1_U3194) );
  NAND2_X1 U23567 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20644) );
  OAI21_X1 U23568 ( .B1(NA), .B2(n20644), .A(n20653), .ZN(n20645) );
  OAI21_X1 U23569 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20646), .A(n20645), 
        .ZN(n20651) );
  INV_X1 U23570 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20648) );
  OAI211_X1 U23571 ( .C1(NA), .C2(n20741), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20653), .ZN(n20647) );
  OAI211_X1 U23572 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20648), .A(HOLD), .B(
        n20647), .ZN(n20649) );
  OAI22_X1 U23573 ( .A1(n20652), .A2(n20651), .B1(n20650), .B2(n20649), .ZN(
        P1_U3196) );
  NAND2_X1 U23574 ( .A1(n20750), .A2(n20653), .ZN(n20701) );
  INV_X1 U23575 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20654) );
  NAND2_X1 U23576 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20750), .ZN(n20705) );
  OAI222_X1 U23577 ( .A1(n20701), .A2(n20656), .B1(n20654), .B2(n20750), .C1(
        n20729), .C2(n20705), .ZN(P1_U3197) );
  INV_X1 U23578 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20655) );
  OAI222_X1 U23579 ( .A1(n20705), .A2(n20656), .B1(n20655), .B2(n20750), .C1(
        n13826), .C2(n20701), .ZN(P1_U3198) );
  OAI222_X1 U23580 ( .A1(n20705), .A2(n13826), .B1(n20657), .B2(n20750), .C1(
        n20659), .C2(n20701), .ZN(P1_U3199) );
  INV_X1 U23581 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20658) );
  OAI222_X1 U23582 ( .A1(n20705), .A2(n20659), .B1(n20658), .B2(n20750), .C1(
        n20661), .C2(n20701), .ZN(P1_U3200) );
  INV_X1 U23583 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20660) );
  OAI222_X1 U23584 ( .A1(n20705), .A2(n20661), .B1(n20660), .B2(n20750), .C1(
        n20663), .C2(n20701), .ZN(P1_U3201) );
  INV_X1 U23585 ( .A(n20701), .ZN(n20707) );
  AOI22_X1 U23586 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20707), .ZN(n20662) );
  OAI21_X1 U23587 ( .B1(n20663), .B2(n20705), .A(n20662), .ZN(P1_U3202) );
  INV_X1 U23588 ( .A(n20705), .ZN(n20708) );
  AOI22_X1 U23589 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20708), .ZN(n20664) );
  OAI21_X1 U23590 ( .B1(n20665), .B2(n20701), .A(n20664), .ZN(P1_U3203) );
  INV_X1 U23591 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20666) );
  OAI222_X1 U23592 ( .A1(n20701), .A2(n20668), .B1(n20666), .B2(n20750), .C1(
        n20665), .C2(n20705), .ZN(P1_U3204) );
  INV_X1 U23593 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20667) );
  OAI222_X1 U23594 ( .A1(n20705), .A2(n20668), .B1(n20667), .B2(n20750), .C1(
        n20671), .C2(n20701), .ZN(P1_U3205) );
  INV_X1 U23595 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20670) );
  OAI222_X1 U23596 ( .A1(n20705), .A2(n20671), .B1(n20670), .B2(n20750), .C1(
        n20669), .C2(n20701), .ZN(P1_U3206) );
  AOI222_X1 U23597 ( .A1(n20708), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20737), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20707), .ZN(n20672) );
  INV_X1 U23598 ( .A(n20672), .ZN(P1_U3207) );
  AOI222_X1 U23599 ( .A1(n20708), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20737), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20707), .ZN(n20673) );
  INV_X1 U23600 ( .A(n20673), .ZN(P1_U3208) );
  INV_X1 U23601 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20674) );
  OAI222_X1 U23602 ( .A1(n20705), .A2(n20675), .B1(n20674), .B2(n20750), .C1(
        n20677), .C2(n20701), .ZN(P1_U3209) );
  INV_X1 U23603 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20676) );
  OAI222_X1 U23604 ( .A1(n20705), .A2(n20677), .B1(n20676), .B2(n20750), .C1(
        n20678), .C2(n20701), .ZN(P1_U3210) );
  INV_X1 U23605 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20681) );
  INV_X1 U23606 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U23607 ( .A1(n20701), .A2(n20681), .B1(n20679), .B2(n20750), .C1(
        n20678), .C2(n20705), .ZN(P1_U3211) );
  AOI22_X1 U23608 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20707), .ZN(n20680) );
  OAI21_X1 U23609 ( .B1(n20681), .B2(n20705), .A(n20680), .ZN(P1_U3212) );
  INV_X1 U23610 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20684) );
  AOI22_X1 U23611 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20708), .ZN(n20682) );
  OAI21_X1 U23612 ( .B1(n20684), .B2(n20701), .A(n20682), .ZN(P1_U3213) );
  AOI22_X1 U23613 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20707), .ZN(n20683) );
  OAI21_X1 U23614 ( .B1(n20684), .B2(n20705), .A(n20683), .ZN(P1_U3214) );
  INV_X1 U23615 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20686) );
  AOI22_X1 U23616 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20708), .ZN(n20685) );
  OAI21_X1 U23617 ( .B1(n20686), .B2(n20701), .A(n20685), .ZN(P1_U3215) );
  INV_X1 U23618 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20687) );
  OAI222_X1 U23619 ( .A1(n20701), .A2(n20689), .B1(n20687), .B2(n20750), .C1(
        n20686), .C2(n20705), .ZN(P1_U3216) );
  AOI22_X1 U23620 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20707), .ZN(n20688) );
  OAI21_X1 U23621 ( .B1(n20689), .B2(n20705), .A(n20688), .ZN(P1_U3217) );
  AOI22_X1 U23622 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20737), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20708), .ZN(n20690) );
  OAI21_X1 U23623 ( .B1(n20692), .B2(n20701), .A(n20690), .ZN(P1_U3218) );
  INV_X1 U23624 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20691) );
  OAI222_X1 U23625 ( .A1(n20705), .A2(n20692), .B1(n20691), .B2(n20750), .C1(
        n20694), .C2(n20701), .ZN(P1_U3219) );
  INV_X1 U23626 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20693) );
  OAI222_X1 U23627 ( .A1(n20705), .A2(n20694), .B1(n20693), .B2(n20750), .C1(
        n20696), .C2(n20701), .ZN(P1_U3220) );
  INV_X1 U23628 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20695) );
  OAI222_X1 U23629 ( .A1(n20705), .A2(n20696), .B1(n20695), .B2(n20750), .C1(
        n20698), .C2(n20701), .ZN(P1_U3221) );
  INV_X1 U23630 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20697) );
  OAI222_X1 U23631 ( .A1(n20705), .A2(n20698), .B1(n20697), .B2(n20750), .C1(
        n20700), .C2(n20701), .ZN(P1_U3222) );
  INV_X1 U23632 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20699) );
  OAI222_X1 U23633 ( .A1(n20705), .A2(n20700), .B1(n20699), .B2(n20750), .C1(
        n20704), .C2(n20701), .ZN(P1_U3223) );
  INV_X1 U23634 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20703) );
  OAI222_X1 U23635 ( .A1(n20705), .A2(n20704), .B1(n20703), .B2(n20750), .C1(
        n20702), .C2(n20701), .ZN(P1_U3224) );
  AOI222_X1 U23636 ( .A1(n20707), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20737), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20708), .ZN(n20706) );
  INV_X1 U23637 ( .A(n20706), .ZN(P1_U3225) );
  AOI222_X1 U23638 ( .A1(n20708), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20737), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20707), .ZN(n20709) );
  INV_X1 U23639 ( .A(n20709), .ZN(P1_U3226) );
  INV_X1 U23640 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20710) );
  AOI22_X1 U23641 ( .A1(n20750), .A2(n20711), .B1(n20710), .B2(n20737), .ZN(
        P1_U3458) );
  INV_X1 U23642 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20732) );
  INV_X1 U23643 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20712) );
  AOI22_X1 U23644 ( .A1(n20750), .A2(n20732), .B1(n20712), .B2(n20737), .ZN(
        P1_U3459) );
  INV_X1 U23645 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20713) );
  AOI22_X1 U23646 ( .A1(n20750), .A2(n20714), .B1(n20713), .B2(n20737), .ZN(
        P1_U3460) );
  INV_X1 U23647 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20735) );
  INV_X1 U23648 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20715) );
  AOI22_X1 U23649 ( .A1(n20750), .A2(n20735), .B1(n20715), .B2(n20737), .ZN(
        P1_U3461) );
  INV_X1 U23650 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20718) );
  INV_X1 U23651 ( .A(n20719), .ZN(n20716) );
  AOI21_X1 U23652 ( .B1(n20718), .B2(n20717), .A(n20716), .ZN(P1_U3464) );
  OAI21_X1 U23653 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(P1_U3465) );
  AOI22_X1 U23654 ( .A1(n20725), .A2(n20724), .B1(n20723), .B2(n20722), .ZN(
        n20726) );
  INV_X1 U23655 ( .A(n20726), .ZN(n20728) );
  MUX2_X1 U23656 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20728), .S(
        n20727), .Z(P1_U3469) );
  AOI21_X1 U23657 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20730) );
  AOI22_X1 U23658 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20730), .B2(n20729), .ZN(n20733) );
  AOI22_X1 U23659 ( .A1(n20736), .A2(n20733), .B1(n20732), .B2(n20731), .ZN(
        P1_U3481) );
  OAI21_X1 U23660 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20736), .ZN(n20734) );
  OAI21_X1 U23661 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(P1_U3482) );
  AOI22_X1 U23662 ( .A1(n20750), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20738), 
        .B2(n20737), .ZN(P1_U3483) );
  AOI211_X1 U23663 ( .C1(n20742), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        n20749) );
  OAI211_X1 U23664 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20744), .A(n20743), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20746) );
  AOI21_X1 U23665 ( .B1(n20746), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20745), 
        .ZN(n20748) );
  NAND2_X1 U23666 ( .A1(n20749), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20747) );
  OAI21_X1 U23667 ( .B1(n20749), .B2(n20748), .A(n20747), .ZN(P1_U3485) );
  MUX2_X1 U23668 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20750), .Z(P1_U3486) );
  NOR4_X1 U23669 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__4__SCAN_IN), .A3(P3_INSTQUEUE_REG_4__4__SCAN_IN), 
        .A4(n20880), .ZN(n20755) );
  INV_X1 U23670 ( .A(DATAI_6_), .ZN(n20862) );
  NOR3_X1 U23671 ( .A1(DATAI_19_), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n20862), 
        .ZN(n20754) );
  INV_X1 U23672 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20833) );
  NAND4_X1 U23673 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20851), .A3(
        n20791), .A4(n20833), .ZN(n20752) );
  NAND4_X1 U23674 ( .A1(n10964), .A2(P2_LWORD_REG_15__SCAN_IN), .A3(n20805), 
        .A4(n20794), .ZN(n20751) );
  NOR2_X1 U23675 ( .A1(n20752), .A2(n20751), .ZN(n20753) );
  NAND3_X1 U23676 ( .A1(n20755), .A2(n20754), .A3(n20753), .ZN(n20773) );
  INV_X1 U23677 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20870) );
  NAND4_X1 U23678 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(n20870), .A4(n13826), .ZN(n20772)
         );
  NOR3_X1 U23679 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(
        n20758) );
  NOR4_X1 U23680 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .A3(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A4(n20854), .ZN(n20757) );
  NOR4_X1 U23681 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n20756) );
  NAND4_X1 U23682 ( .A1(P3_ADDRESS_REG_20__SCAN_IN), .A2(n20758), .A3(n20757), 
        .A4(n20756), .ZN(n20771) );
  NOR4_X1 U23683 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(DATAI_13_), .A3(
        P3_DATAO_REG_29__SCAN_IN), .A4(n20759), .ZN(n20769) );
  INV_X1 U23684 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20787) );
  NAND4_X1 U23685 ( .A1(P2_BYTEENABLE_REG_3__SCAN_IN), .A2(n20788), .A3(n20806), .A4(n20787), .ZN(n20762) );
  NAND3_X1 U23686 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), 
        .ZN(n20761) );
  INV_X1 U23687 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20837) );
  NAND4_X1 U23688 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_UWORD_REG_0__SCAN_IN), .A3(n20837), .A4(n12009), .ZN(n20760) );
  NOR4_X1 U23689 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n20762), .A3(n20761), 
        .A4(n20760), .ZN(n20768) );
  NOR4_X1 U23690 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_15__SCAN_IN), .A3(n20893), .A4(n20898), .ZN(n20767) );
  NAND4_X1 U23691 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(P2_EBX_REG_22__SCAN_IN), 
        .A3(DATAI_1_), .A4(P3_BE_N_REG_1__SCAN_IN), .ZN(n20765) );
  NAND3_X1 U23692 ( .A1(P3_UWORD_REG_4__SCAN_IN), .A2(
        P3_ADDRESS_REG_24__SCAN_IN), .A3(P3_UWORD_REG_11__SCAN_IN), .ZN(n20764) );
  NAND4_X1 U23693 ( .A1(BUF2_REG_20__SCAN_IN), .A2(P2_ADDRESS_REG_26__SCAN_IN), 
        .A3(P3_UWORD_REG_3__SCAN_IN), .A4(n20885), .ZN(n20763) );
  NOR4_X1 U23694 ( .A1(P3_LWORD_REG_3__SCAN_IN), .A2(n20765), .A3(n20764), 
        .A4(n20763), .ZN(n20766) );
  NAND4_X1 U23695 ( .A1(n20769), .A2(n20768), .A3(n20767), .A4(n20766), .ZN(
        n20770) );
  NOR4_X1 U23696 ( .A1(n20773), .A2(n20772), .A3(n20771), .A4(n20770), .ZN(
        n20782) );
  INV_X1 U23697 ( .A(n20774), .ZN(n20779) );
  AOI21_X1 U23698 ( .B1(n20777), .B2(n20776), .A(n20775), .ZN(n20778) );
  AOI22_X1 U23699 ( .A1(n20780), .A2(n20779), .B1(n20778), .B2(n17258), .ZN(
        n20781) );
  XNOR2_X1 U23700 ( .A(n20782), .B(n20781), .ZN(n20912) );
  AOI22_X1 U23701 ( .A1(n20785), .A2(keyinput12), .B1(keyinput34), .B2(n20784), 
        .ZN(n20783) );
  OAI221_X1 U23702 ( .B1(n20785), .B2(keyinput12), .C1(n20784), .C2(keyinput34), .A(n20783), .ZN(n20798) );
  AOI22_X1 U23703 ( .A1(n20788), .A2(keyinput24), .B1(keyinput1), .B2(n20787), 
        .ZN(n20786) );
  OAI221_X1 U23704 ( .B1(n20788), .B2(keyinput24), .C1(n20787), .C2(keyinput1), 
        .A(n20786), .ZN(n20797) );
  INV_X1 U23705 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n20790) );
  AOI22_X1 U23706 ( .A1(n20791), .A2(keyinput55), .B1(keyinput33), .B2(n20790), 
        .ZN(n20789) );
  OAI221_X1 U23707 ( .B1(n20791), .B2(keyinput55), .C1(n20790), .C2(keyinput33), .A(n20789), .ZN(n20796) );
  INV_X1 U23708 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U23709 ( .A1(n20794), .A2(keyinput44), .B1(n20793), .B2(keyinput50), 
        .ZN(n20792) );
  OAI221_X1 U23710 ( .B1(n20794), .B2(keyinput44), .C1(n20793), .C2(keyinput50), .A(n20792), .ZN(n20795) );
  NOR4_X1 U23711 ( .A1(n20798), .A2(n20797), .A3(n20796), .A4(n20795), .ZN(
        n20910) );
  AOI22_X1 U23712 ( .A1(n10783), .A2(keyinput46), .B1(keyinput32), .B2(n20800), 
        .ZN(n20799) );
  OAI221_X1 U23713 ( .B1(n10783), .B2(keyinput46), .C1(n20800), .C2(keyinput32), .A(n20799), .ZN(n20803) );
  XNOR2_X1 U23714 ( .A(n20801), .B(keyinput19), .ZN(n20802) );
  NOR2_X1 U23715 ( .A1(n20803), .A2(n20802), .ZN(n20814) );
  AOI22_X1 U23716 ( .A1(n20806), .A2(keyinput28), .B1(keyinput61), .B2(n20805), 
        .ZN(n20804) );
  OAI221_X1 U23717 ( .B1(n20806), .B2(keyinput28), .C1(n20805), .C2(keyinput61), .A(n20804), .ZN(n20807) );
  INV_X1 U23718 ( .A(n20807), .ZN(n20813) );
  AOI22_X1 U23719 ( .A1(n12395), .A2(keyinput11), .B1(keyinput30), .B2(n20809), 
        .ZN(n20808) );
  OAI221_X1 U23720 ( .B1(n12395), .B2(keyinput11), .C1(n20809), .C2(keyinput30), .A(n20808), .ZN(n20810) );
  INV_X1 U23721 ( .A(n20810), .ZN(n20812) );
  XNOR2_X1 U23722 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput62), .ZN(
        n20811) );
  AND4_X1 U23723 ( .A1(n20814), .A2(n20813), .A3(n20812), .A4(n20811), .ZN(
        n20909) );
  INV_X1 U23724 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20817) );
  INV_X1 U23725 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U23726 ( .A1(n20817), .A2(keyinput22), .B1(n20816), .B2(keyinput0), 
        .ZN(n20815) );
  OAI221_X1 U23727 ( .B1(n20817), .B2(keyinput22), .C1(n20816), .C2(keyinput0), 
        .A(n20815), .ZN(n20823) );
  XNOR2_X1 U23728 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput14), .ZN(
        n20821) );
  XNOR2_X1 U23729 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(keyinput27), 
        .ZN(n20820) );
  XNOR2_X1 U23730 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput18), 
        .ZN(n20819) );
  XNOR2_X1 U23731 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput58), 
        .ZN(n20818) );
  NAND4_X1 U23732 ( .A1(n20821), .A2(n20820), .A3(n20819), .A4(n20818), .ZN(
        n20822) );
  NOR2_X1 U23733 ( .A1(n20823), .A2(n20822), .ZN(n20831) );
  INV_X1 U23734 ( .A(DATAI_1_), .ZN(n20824) );
  XNOR2_X1 U23735 ( .A(n20824), .B(keyinput15), .ZN(n20829) );
  XOR2_X1 U23736 ( .A(keyinput43), .B(P3_BE_N_REG_1__SCAN_IN), .Z(n20828) );
  XNOR2_X1 U23737 ( .A(keyinput36), .B(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n20826) );
  XNOR2_X1 U23738 ( .A(keyinput9), .B(P1_EBX_REG_23__SCAN_IN), .ZN(n20825) );
  NAND2_X1 U23739 ( .A1(n20826), .A2(n20825), .ZN(n20827) );
  NOR3_X1 U23740 ( .A1(n20829), .A2(n20828), .A3(n20827), .ZN(n20830) );
  AND2_X1 U23741 ( .A1(n20831), .A2(n20830), .ZN(n20843) );
  OAI22_X1 U23742 ( .A1(n20834), .A2(keyinput21), .B1(n20833), .B2(keyinput41), 
        .ZN(n20832) );
  AOI221_X1 U23743 ( .B1(n20834), .B2(keyinput21), .C1(keyinput41), .C2(n20833), .A(n20832), .ZN(n20842) );
  INV_X1 U23744 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n20836) );
  OAI22_X1 U23745 ( .A1(n20837), .A2(keyinput38), .B1(n20836), .B2(keyinput6), 
        .ZN(n20835) );
  AOI221_X1 U23746 ( .B1(n20837), .B2(keyinput38), .C1(keyinput6), .C2(n20836), 
        .A(n20835), .ZN(n20841) );
  INV_X1 U23747 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n20839) );
  OAI22_X1 U23748 ( .A1(n13765), .A2(keyinput53), .B1(n20839), .B2(keyinput63), 
        .ZN(n20838) );
  AOI221_X1 U23749 ( .B1(n13765), .B2(keyinput53), .C1(keyinput63), .C2(n20839), .A(n20838), .ZN(n20840) );
  AND4_X1 U23750 ( .A1(n20843), .A2(n20842), .A3(n20841), .A4(n20840), .ZN(
        n20908) );
  INV_X1 U23751 ( .A(keyinput45), .ZN(n20845) );
  OAI22_X1 U23752 ( .A1(keyinput59), .A2(n20846), .B1(n20845), .B2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20844) );
  AOI221_X1 U23753 ( .B1(n20846), .B2(keyinput59), .C1(n20845), .C2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .A(n20844), .ZN(n20859) );
  INV_X1 U23754 ( .A(keyinput51), .ZN(n20848) );
  OAI22_X1 U23755 ( .A1(keyinput60), .A2(n20849), .B1(n20848), .B2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20847) );
  AOI221_X1 U23756 ( .B1(n20849), .B2(keyinput60), .C1(n20848), .C2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A(n20847), .ZN(n20858) );
  OAI22_X1 U23757 ( .A1(n20852), .A2(keyinput56), .B1(n20851), .B2(keyinput49), 
        .ZN(n20850) );
  AOI221_X1 U23758 ( .B1(n20852), .B2(keyinput56), .C1(keyinput49), .C2(n20851), .A(n20850), .ZN(n20857) );
  INV_X1 U23759 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20855) );
  OAI22_X1 U23760 ( .A1(n20855), .A2(keyinput47), .B1(n20854), .B2(keyinput8), 
        .ZN(n20853) );
  AOI221_X1 U23761 ( .B1(n20855), .B2(keyinput47), .C1(keyinput8), .C2(n20854), 
        .A(n20853), .ZN(n20856) );
  NAND4_X1 U23762 ( .A1(n20859), .A2(n20858), .A3(n20857), .A4(n20856), .ZN(
        n20906) );
  OAI22_X1 U23763 ( .A1(n20862), .A2(keyinput42), .B1(n20861), .B2(keyinput57), 
        .ZN(n20860) );
  AOI221_X1 U23764 ( .B1(n20862), .B2(keyinput42), .C1(keyinput57), .C2(n20861), .A(n20860), .ZN(n20874) );
  INV_X1 U23765 ( .A(DATAI_19_), .ZN(n20865) );
  INV_X1 U23766 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20864) );
  OAI22_X1 U23767 ( .A1(n20865), .A2(keyinput26), .B1(n20864), .B2(keyinput31), 
        .ZN(n20863) );
  AOI221_X1 U23768 ( .B1(n20865), .B2(keyinput26), .C1(keyinput31), .C2(n20864), .A(n20863), .ZN(n20873) );
  OAI22_X1 U23769 ( .A1(n20868), .A2(keyinput16), .B1(n20867), .B2(keyinput7), 
        .ZN(n20866) );
  AOI221_X1 U23770 ( .B1(n20868), .B2(keyinput16), .C1(keyinput7), .C2(n20867), 
        .A(n20866), .ZN(n20872) );
  OAI22_X1 U23771 ( .A1(n20870), .A2(keyinput23), .B1(n13826), .B2(keyinput4), 
        .ZN(n20869) );
  AOI221_X1 U23772 ( .B1(n20870), .B2(keyinput23), .C1(keyinput4), .C2(n13826), 
        .A(n20869), .ZN(n20871) );
  NAND4_X1 U23773 ( .A1(n20874), .A2(n20873), .A3(n20872), .A4(n20871), .ZN(
        n20905) );
  INV_X1 U23774 ( .A(keyinput2), .ZN(n20876) );
  OAI22_X1 U23775 ( .A1(keyinput52), .A2(n20877), .B1(n20876), .B2(
        P3_UWORD_REG_11__SCAN_IN), .ZN(n20875) );
  AOI221_X1 U23776 ( .B1(n20877), .B2(keyinput52), .C1(n20876), .C2(
        P3_UWORD_REG_11__SCAN_IN), .A(n20875), .ZN(n20890) );
  INV_X1 U23777 ( .A(P3_UWORD_REG_4__SCAN_IN), .ZN(n20879) );
  OAI22_X1 U23778 ( .A1(n20880), .A2(keyinput48), .B1(n20879), .B2(keyinput29), 
        .ZN(n20878) );
  AOI221_X1 U23779 ( .B1(n20880), .B2(keyinput48), .C1(keyinput29), .C2(n20879), .A(n20878), .ZN(n20889) );
  OAI22_X1 U23780 ( .A1(n20883), .A2(keyinput25), .B1(n20882), .B2(keyinput37), 
        .ZN(n20881) );
  AOI221_X1 U23781 ( .B1(n20883), .B2(keyinput25), .C1(keyinput37), .C2(n20882), .A(n20881), .ZN(n20888) );
  OAI22_X1 U23782 ( .A1(n20886), .A2(keyinput54), .B1(n20885), .B2(keyinput5), 
        .ZN(n20884) );
  AOI221_X1 U23783 ( .B1(n20886), .B2(keyinput54), .C1(keyinput5), .C2(n20885), 
        .A(n20884), .ZN(n20887) );
  NAND4_X1 U23784 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n20904) );
  OAI22_X1 U23785 ( .A1(n20893), .A2(keyinput35), .B1(n20892), .B2(keyinput17), 
        .ZN(n20891) );
  AOI221_X1 U23786 ( .B1(n20893), .B2(keyinput35), .C1(keyinput17), .C2(n20892), .A(n20891), .ZN(n20902) );
  OAI22_X1 U23787 ( .A1(n10767), .A2(keyinput3), .B1(n15115), .B2(keyinput20), 
        .ZN(n20894) );
  AOI221_X1 U23788 ( .B1(n10767), .B2(keyinput3), .C1(keyinput20), .C2(n15115), 
        .A(n20894), .ZN(n20901) );
  INV_X1 U23789 ( .A(keyinput40), .ZN(n20896) );
  OAI22_X1 U23790 ( .A1(n11840), .A2(keyinput13), .B1(n20896), .B2(
        P3_LWORD_REG_3__SCAN_IN), .ZN(n20895) );
  AOI221_X1 U23791 ( .B1(n11840), .B2(keyinput13), .C1(P3_LWORD_REG_3__SCAN_IN), .C2(n20896), .A(n20895), .ZN(n20900) );
  OAI22_X1 U23792 ( .A1(n20898), .A2(keyinput39), .B1(n13658), .B2(keyinput10), 
        .ZN(n20897) );
  AOI221_X1 U23793 ( .B1(n20898), .B2(keyinput39), .C1(keyinput10), .C2(n13658), .A(n20897), .ZN(n20899) );
  NAND4_X1 U23794 ( .A1(n20902), .A2(n20901), .A3(n20900), .A4(n20899), .ZN(
        n20903) );
  NOR4_X1 U23795 ( .A1(n20906), .A2(n20905), .A3(n20904), .A4(n20903), .ZN(
        n20907) );
  NAND4_X1 U23796 ( .A1(n20910), .A2(n20909), .A3(n20908), .A4(n20907), .ZN(
        n20911) );
  XNOR2_X1 U23797 ( .A(n20912), .B(n20911), .ZN(P3_U2684) );
  AND2_X1 U11203 ( .A1(n10958), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10969) );
  INV_X1 U11045 ( .A(n15717), .ZN(n10914) );
  BUF_X2 U12418 ( .A(n12871), .Z(n16971) );
  AND2_X1 U11131 ( .A1(n11151), .A2(n11116), .ZN(n13373) );
  BUF_X2 U11026 ( .A(n12176), .Z(n14380) );
  CLKBUF_X1 U11037 ( .A(n11021), .Z(n12028) );
  CLKBUF_X1 U11051 ( .A(n11919), .Z(n12100) );
  CLKBUF_X2 U11061 ( .A(n11332), .Z(n11944) );
  NOR2_X1 U11063 ( .A1(n11288), .A2(n20635), .ZN(n11498) );
  CLKBUF_X1 U11064 ( .A(n10066), .Z(n10067) );
  CLKBUF_X1 U11065 ( .A(n11165), .Z(n9614) );
  CLKBUF_X1 U11071 ( .A(n14708), .Z(n16053) );
  CLKBUF_X1 U11083 ( .A(n10097), .Z(n9606) );
  CLKBUF_X1 U11089 ( .A(n10355), .Z(n10369) );
  INV_X1 U11094 ( .A(n12173), .ZN(n12156) );
  CLKBUF_X1 U11104 ( .A(n11470), .Z(n9604) );
  NOR2_X1 U11105 ( .A1(n15025), .A2(n15012), .ZN(n14990) );
  AND2_X1 U11116 ( .A1(n10408), .A2(n10407), .ZN(n10404) );
  OR2_X1 U11118 ( .A1(n11170), .A2(n11169), .ZN(n11171) );
  CLKBUF_X1 U11154 ( .A(n11107), .Z(n9635) );
  CLKBUF_X1 U11175 ( .A(n13703), .Z(n9631) );
  CLKBUF_X1 U11193 ( .A(n9779), .Z(n9627) );
  NAND2_X2 U11206 ( .A1(n19203), .A2(n10559), .ZN(n12350) );
  CLKBUF_X1 U11209 ( .A(n10404), .Z(n10410) );
  CLKBUF_X1 U11210 ( .A(n10090), .Z(n10091) );
  CLKBUF_X1 U11326 ( .A(n11536), .Z(n9632) );
  NAND2_X1 U11337 ( .A1(n10028), .A2(n12350), .ZN(n13107) );
  CLKBUF_X1 U11383 ( .A(n19165), .Z(n19860) );
  INV_X1 U11403 ( .A(n12980), .ZN(n17432) );
  CLKBUF_X1 U11410 ( .A(n16521), .Z(n16527) );
  AND2_X1 U11437 ( .A1(n17266), .A2(n18274), .ZN(n20913) );
  AND3_X4 U11466 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20914) );
  OR2_X1 U11479 ( .A1(n10744), .A2(n10544), .ZN(n20915) );
  NAND2_X2 U11527 ( .A1(n13161), .A2(n16367), .ZN(n19046) );
  AND2_X2 U11542 ( .A1(n13112), .A2(n10566), .ZN(n13161) );
endmodule

