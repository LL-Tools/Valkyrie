

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123;

  INV_X1 U3541 ( .A(n5697), .ZN(n4499) );
  NAND2_X1 U3543 ( .A1(n5336), .A2(n5788), .ZN(n5787) );
  INV_X1 U3544 ( .A(n3905), .ZN(n3547) );
  AND2_X1 U3545 ( .A1(n4187), .A2(n4758), .ZN(n4320) );
  CLKBUF_X2 U3546 ( .A(n3344), .Z(n3884) );
  BUF_X1 U3547 ( .A(n3427), .Z(n4753) );
  CLKBUF_X2 U3548 ( .A(n4097), .Z(n3970) );
  CLKBUF_X2 U3549 ( .A(n3315), .Z(n4044) );
  CLKBUF_X2 U3550 ( .A(n4067), .Z(n4090) );
  CLKBUF_X2 U3551 ( .A(n3339), .Z(n4025) );
  CLKBUF_X2 U3552 ( .A(n3392), .Z(n3925) );
  BUF_X2 U3553 ( .A(n3096), .Z(n4068) );
  CLKBUF_X2 U3554 ( .A(n3456), .Z(n4074) );
  NAND2_X1 U3555 ( .A1(n3313), .A2(n3312), .ZN(n3401) );
  AND4_X1 U3556 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3367)
         );
  AND3_X1 U3557 ( .A1(n3294), .A2(n3293), .A3(n3292), .ZN(n3303) );
  INV_X2 U3558 ( .A(n3473), .ZN(n4099) );
  AND2_X2 U3559 ( .A1(n3297), .A2(n4777), .ZN(n4100) );
  AND2_X1 U3560 ( .A1(n3510), .A2(n7027), .ZN(n3454) );
  CLKBUF_X2 U3561 ( .A(n3461), .Z(n4050) );
  NAND2_X1 U3562 ( .A1(n4612), .A2(n5383), .ZN(n4279) );
  AND2_X1 U3563 ( .A1(n4952), .A2(n5067), .ZN(n5066) );
  CLKBUF_X2 U3564 ( .A(n3401), .Z(n3810) );
  NOR2_X1 U3566 ( .A1(n6807), .A2(n4996), .ZN(n5295) );
  NOR2_X1 U3567 ( .A1(n4669), .A2(n4670), .ZN(n6407) );
  NOR3_X1 U3569 ( .A1(n5425), .A2(n3248), .A3(n3247), .ZN(n5402) );
  AND2_X1 U3570 ( .A1(n4437), .A2(n4436), .ZN(n3285) );
  AND2_X1 U3571 ( .A1(n6022), .A2(n4463), .ZN(n6011) );
  INV_X1 U3572 ( .A(n6334), .ZN(n6365) );
  INV_X1 U3573 ( .A(n6259), .ZN(n6247) );
  BUF_X1 U3574 ( .A(n3418), .Z(n4173) );
  BUF_X2 U3575 ( .A(n3338), .Z(n3644) );
  AND2_X2 U3576 ( .A1(n5480), .A2(n4302), .ZN(n5450) );
  NAND2_X2 U3577 ( .A1(n3579), .A2(n4724), .ZN(n3578) );
  NAND2_X2 U3578 ( .A1(n5787), .A2(n3203), .ZN(n5783) );
  XNOR2_X2 U3579 ( .A(n5796), .B(n4526), .ZN(n5973) );
  INV_X1 U3580 ( .A(n3185), .ZN(n4813) );
  NOR2_X2 U3581 ( .A1(n5951), .A2(n4476), .ZN(n5936) );
  AOI211_X2 U3582 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6250), .A(n5352), .B(n5351), 
        .ZN(n5353) );
  OAI22_X2 U3583 ( .A1(n4123), .A2(n4124), .B1(n4121), .B2(n4139), .ZN(n4129)
         );
  AND2_X1 U3584 ( .A1(n6098), .A2(n4466), .ZN(n6022) );
  NAND2_X1 U3585 ( .A1(n4461), .A2(n6038), .ZN(n6098) );
  OR3_X2 U3586 ( .A1(n6792), .A2(n6377), .A3(n4184), .ZN(n6183) );
  AND2_X1 U3587 ( .A1(n3497), .A2(n4489), .ZN(n4128) );
  NAND2_X2 U3588 ( .A1(n3542), .A2(n3541), .ZN(n4164) );
  CLKBUF_X3 U3589 ( .A(n4198), .Z(n3098) );
  INV_X1 U3590 ( .A(n3571), .ZN(n4082) );
  CLKBUF_X1 U3591 ( .A(n3570), .Z(n4488) );
  AND2_X1 U3592 ( .A1(n3810), .A2(n4602), .ZN(n4388) );
  BUF_X2 U3593 ( .A(n3355), .Z(n4489) );
  NAND4_X4 U3594 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n4187)
         );
  AND4_X1 U3595 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3384)
         );
  AND4_X1 U3596 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3387)
         );
  AND4_X1 U3597 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3335)
         );
  AND4_X1 U3598 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3386)
         );
  BUF_X2 U3599 ( .A(n3338), .Z(n3461) );
  INV_X4 U3600 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5334) );
  INV_X2 U3601 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3287) );
  NOR2_X1 U3602 ( .A1(n4545), .A2(n4544), .ZN(n4546) );
  NAND2_X1 U3603 ( .A1(n3231), .A2(n3118), .ZN(n3234) );
  XNOR2_X1 U3604 ( .A(n5372), .B(n5371), .ZN(n5758) );
  AOI211_X1 U3605 ( .C1(n5346), .C2(n6365), .A(n5345), .B(n5344), .ZN(n5347)
         );
  AOI211_X1 U3606 ( .C1(n6350), .C2(n5802), .A(n5801), .B(n5800), .ZN(n5803)
         );
  INV_X1 U3607 ( .A(n5424), .ZN(n5794) );
  NOR2_X1 U3608 ( .A1(n5820), .A2(n3144), .ZN(n5821) );
  OR2_X1 U3609 ( .A1(n4412), .A2(n3223), .ZN(n5884) );
  AOI21_X1 U3610 ( .B1(n4500), .B2(n4499), .A(n4498), .ZN(n4501) );
  NOR2_X1 U3611 ( .A1(n4311), .A2(n3172), .ZN(n3171) );
  OR2_X1 U3612 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  NAND2_X1 U3613 ( .A1(n4406), .A2(n4405), .ZN(n5909) );
  OR2_X1 U3614 ( .A1(n5402), .A2(n5401), .ZN(n5932) );
  AND2_X1 U3615 ( .A1(n3158), .A2(n3136), .ZN(n3154) );
  OR2_X1 U3616 ( .A1(n3183), .A2(n3182), .ZN(n3181) );
  AND2_X1 U3617 ( .A1(n4951), .A2(n3205), .ZN(n3158) );
  NAND2_X1 U3618 ( .A1(n3217), .A2(n4380), .ZN(n3216) );
  NAND2_X1 U3619 ( .A1(n3260), .A2(n5831), .ZN(n3259) );
  OR2_X1 U3620 ( .A1(n3262), .A2(n4420), .ZN(n3261) );
  OR2_X1 U3621 ( .A1(n5823), .A2(n5830), .ZN(n3144) );
  NAND2_X1 U3622 ( .A1(n3184), .A2(n3119), .ZN(n3183) );
  NAND2_X1 U3623 ( .A1(n3665), .A2(n3664), .ZN(n4951) );
  AND2_X1 U3624 ( .A1(n5870), .A2(n4418), .ZN(n4419) );
  AND2_X1 U3625 ( .A1(n3212), .A2(n6360), .ZN(n4691) );
  OR2_X1 U3626 ( .A1(n4407), .A2(n6383), .ZN(n5898) );
  AND2_X1 U3627 ( .A1(n4460), .A2(n5295), .ZN(n6054) );
  AND2_X1 U3628 ( .A1(n6392), .A2(n4464), .ZN(n6080) );
  OR2_X1 U3629 ( .A1(n6395), .A2(n6055), .ZN(n6059) );
  OR2_X1 U3630 ( .A1(n6416), .A2(n6055), .ZN(n6037) );
  CLKBUF_X1 U3631 ( .A(n5358), .Z(n5733) );
  OR2_X1 U3632 ( .A1(n5004), .A2(n5299), .ZN(n4996) );
  NAND2_X1 U3633 ( .A1(n4467), .A2(n4569), .ZN(n5004) );
  AND2_X1 U3634 ( .A1(n4467), .A2(n6117), .ZN(n6416) );
  CLKBUF_X2 U3635 ( .A(n4725), .Z(n3097) );
  AND2_X2 U3636 ( .A1(n4330), .A2(n6154), .ZN(n4467) );
  NAND2_X2 U3637 ( .A1(n5696), .A2(n4842), .ZN(n5694) );
  INV_X1 U3638 ( .A(n5608), .ZN(n3093) );
  CLKBUF_X1 U3639 ( .A(n4713), .Z(n5625) );
  NAND2_X1 U3640 ( .A1(n4604), .A2(n4565), .ZN(n6792) );
  NAND2_X1 U3641 ( .A1(n3166), .A2(n3164), .ZN(n4618) );
  NAND2_X1 U3642 ( .A1(n3540), .A2(n3539), .ZN(n6495) );
  AOI21_X1 U3643 ( .B1(n3535), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3515), 
        .ZN(n3532) );
  INV_X1 U3644 ( .A(n5137), .ZN(n6473) );
  NAND2_X1 U3645 ( .A1(n3502), .A2(n4334), .ZN(n3594) );
  AND2_X1 U3646 ( .A1(n3221), .A2(n3220), .ZN(n5137) );
  NAND2_X1 U3647 ( .A1(n4192), .A2(n4193), .ZN(n3244) );
  AOI21_X2 U3648 ( .B1(n4319), .B2(n4320), .A(n3400), .ZN(n3425) );
  OAI211_X1 U3649 ( .C1(n4157), .C2(n3508), .A(n3507), .B(n3506), .ZN(n3593)
         );
  AND3_X1 U3650 ( .A1(n4445), .A2(n4793), .A3(n3422), .ZN(n3423) );
  NAND2_X1 U3651 ( .A1(n4194), .A2(n5383), .ZN(n4665) );
  OR2_X1 U3652 ( .A1(n3501), .A2(n7027), .ZN(n4334) );
  INV_X1 U3653 ( .A(n3098), .ZN(n4612) );
  OR2_X1 U3654 ( .A1(n4843), .A2(n4489), .ZN(n3353) );
  OR2_X1 U3655 ( .A1(n3468), .A2(n3467), .ZN(n4348) );
  OR2_X1 U3656 ( .A1(n3483), .A2(n3482), .ZN(n4399) );
  OR2_X1 U3657 ( .A1(n3494), .A2(n3493), .ZN(n4355) );
  NAND4_X1 U3658 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3355)
         );
  NAND2_X1 U3659 ( .A1(n3412), .A2(n3411), .ZN(n4443) );
  OR2_X2 U3660 ( .A1(n3351), .A2(n3350), .ZN(n4842) );
  AND4_X1 U3661 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3411)
         );
  AND4_X1 U3662 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  AND4_X1 U3663 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3336)
         );
  AND4_X1 U3664 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3412)
         );
  NOR2_X1 U3665 ( .A1(n6334), .A2(n4762), .ZN(n6686) );
  AND4_X1 U3666 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3366)
         );
  NOR2_X1 U3667 ( .A1(n6334), .A2(n4737), .ZN(n6707) );
  AND4_X1 U3668 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3333)
         );
  INV_X2 U3669 ( .A(n3455), .ZN(n4098) );
  AND4_X1 U3670 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3313)
         );
  AND4_X1 U3671 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3334)
         );
  OR2_X2 U3672 ( .A1(n6717), .A2(n6651), .ZN(n6334) );
  BUF_X2 U3673 ( .A(n4100), .Z(n4049) );
  BUF_X2 U3674 ( .A(n3345), .Z(n4030) );
  AND2_X2 U3675 ( .A1(n3295), .A2(n4788), .ZN(n3314) );
  AND2_X2 U3676 ( .A1(n3288), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5321)
         );
  INV_X2 U3677 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3288) );
  NOR2_X2 U3678 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4788) );
  NAND2_X2 U3679 ( .A1(n3153), .A2(n3107), .ZN(n5568) );
  OR2_X2 U3680 ( .A1(n4675), .A2(n4674), .ZN(n4773) );
  OR2_X1 U3681 ( .A1(n3809), .A2(n3417), .ZN(n4793) );
  AND2_X1 U3682 ( .A1(n3417), .A2(n3427), .ZN(n4447) );
  NAND2_X1 U3683 ( .A1(n3534), .A2(n3533), .ZN(n4593) );
  OR2_X1 U3684 ( .A1(n5470), .A2(n3207), .ZN(n5438) );
  NAND2_X2 U3685 ( .A1(n4227), .A2(n4226), .ZN(n5587) );
  INV_X2 U3686 ( .A(n5232), .ZN(n4227) );
  AND2_X2 U3687 ( .A1(n3297), .A2(n3295), .ZN(n3484) );
  AND2_X1 U3688 ( .A1(n3295), .A2(n4789), .ZN(n3472) );
  AND2_X2 U3689 ( .A1(n3295), .A2(n3296), .ZN(n3344) );
  NOR2_X4 U3690 ( .A1(n5495), .A2(n5496), .ZN(n5484) );
  XNOR2_X2 U3691 ( .A(n4360), .B(n4339), .ZN(n4692) );
  BUF_X2 U3692 ( .A(n4185), .Z(n4186) );
  INV_X4 U3693 ( .A(n5503), .ZN(n5383) );
  INV_X2 U3694 ( .A(n4186), .ZN(n5503) );
  NAND4_X1 U3695 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3094)
         );
  NAND4_X2 U3696 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3095)
         );
  NOR2_X2 U3697 ( .A1(n3620), .A2(n4677), .ZN(n4703) );
  AND2_X4 U3698 ( .A1(n5334), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3297)
         );
  NAND2_X2 U3699 ( .A1(n5448), .A2(n5443), .ZN(n5425) );
  OAI21_X2 U3700 ( .B1(n5901), .B2(n3181), .A(n3222), .ZN(n4415) );
  NOR2_X4 U3701 ( .A1(n5470), .A2(n3209), .ZN(n5437) );
  NAND2_X2 U3702 ( .A1(n5484), .A2(n5485), .ZN(n5470) );
  AND2_X1 U3703 ( .A1(n3295), .A2(n4789), .ZN(n3096) );
  OAI21_X1 U3704 ( .B1(n5404), .B2(n5343), .A(n5381), .ZN(n5362) );
  NAND2_X2 U3705 ( .A1(n5342), .A2(n5343), .ZN(n5381) );
  NAND2_X1 U3706 ( .A1(n3530), .A2(n3529), .ZN(n3139) );
  XNOR2_X1 U3707 ( .A(n3596), .B(n3595), .ZN(n4725) );
  AOI21_X1 U3708 ( .B1(n4415), .B2(n3117), .A(n3255), .ZN(n5336) );
  OAI22_X2 U3709 ( .A1(n3592), .A2(n3509), .B1(n3593), .B2(n3594), .ZN(n3587)
         );
  NAND2_X1 U3710 ( .A1(n3419), .A2(n3094), .ZN(n4198) );
  XNOR2_X2 U3711 ( .A(n3268), .B(n5369), .ZN(n5365) );
  NOR2_X4 U3712 ( .A1(n5381), .A2(n5382), .ZN(n3268) );
  NAND2_X4 U3713 ( .A1(n4333), .A2(n4335), .ZN(n4407) );
  AND2_X1 U3714 ( .A1(n3432), .A2(n4842), .ZN(n3433) );
  NAND2_X1 U3715 ( .A1(n3421), .A2(n4842), .ZN(n3809) );
  NAND2_X1 U3716 ( .A1(n3169), .A2(n3168), .ZN(n3163) );
  NAND2_X1 U3717 ( .A1(n4159), .A2(n4158), .ZN(n3169) );
  NAND2_X1 U3718 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  NAND2_X1 U3719 ( .A1(n4128), .A2(n4388), .ZN(n4167) );
  AND2_X1 U3720 ( .A1(n3206), .A2(n5681), .ZN(n3205) );
  XNOR2_X1 U3721 ( .A(n4333), .B(n3667), .ZN(n4389) );
  INV_X1 U3722 ( .A(n4084), .ZN(n4110) );
  NAND2_X1 U3723 ( .A1(n3270), .A2(n5513), .ZN(n3269) );
  INV_X1 U3724 ( .A(n3271), .ZN(n3270) );
  NOR2_X1 U3725 ( .A1(n5315), .A2(n7027), .ZN(n4084) );
  NAND2_X1 U3726 ( .A1(n6592), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3967) );
  NOR2_X1 U3727 ( .A1(n4488), .A2(n6592), .ZN(n3800) );
  INV_X1 U3728 ( .A(n4419), .ZN(n3260) );
  AOI21_X1 U3729 ( .B1(n3223), .B2(n4413), .A(n3120), .ZN(n3222) );
  INV_X1 U3730 ( .A(n4413), .ZN(n3182) );
  NOR2_X1 U3731 ( .A1(n4656), .A2(n4455), .ZN(n4459) );
  AND2_X1 U3732 ( .A1(n4439), .A2(n5609), .ZN(n4577) );
  INV_X1 U3733 ( .A(n4714), .ZN(n3605) );
  INV_X1 U3734 ( .A(n4399), .ZN(n3503) );
  NAND2_X1 U3735 ( .A1(n4399), .A2(n4763), .ZN(n3501) );
  INV_X1 U3736 ( .A(n4128), .ZN(n4157) );
  NAND2_X1 U3737 ( .A1(n4169), .A2(n4175), .ZN(n4170) );
  INV_X1 U3738 ( .A(n3355), .ZN(n3426) );
  INV_X1 U3739 ( .A(n4600), .ZN(n6794) );
  NAND2_X1 U3740 ( .A1(n6183), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5608) );
  AOI22_X1 U3741 ( .A1(n3456), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3347) );
  CLKBUF_X1 U3742 ( .A(n4320), .Z(n4600) );
  OR2_X1 U3743 ( .A1(n4618), .A2(n4568), .ZN(n4604) );
  OR2_X1 U3744 ( .A1(n3965), .A2(n7044), .ZN(n4018) );
  INV_X1 U3745 ( .A(n3826), .ZN(n3827) );
  NOR2_X1 U3746 ( .A1(n3240), .A2(n5506), .ZN(n3239) );
  INV_X1 U3747 ( .A(n3241), .ZN(n3240) );
  NAND2_X1 U3748 ( .A1(n4722), .A2(n7027), .ZN(n5053) );
  INV_X1 U3749 ( .A(n6419), .ZN(n4900) );
  INV_X1 U3750 ( .A(n3484), .ZN(n3455) );
  NAND2_X1 U3751 ( .A1(n5321), .A2(n4788), .ZN(n3361) );
  INV_X1 U3752 ( .A(n3635), .ZN(n3140) );
  NAND2_X1 U3753 ( .A1(n3578), .A2(n3569), .ZN(n3148) );
  OR2_X1 U3754 ( .A1(n4489), .A2(n7027), .ZN(n3541) );
  INV_X1 U3755 ( .A(n4167), .ZN(n4169) );
  NAND2_X1 U3756 ( .A1(n3160), .A2(n4141), .ZN(n3159) );
  OAI21_X1 U3757 ( .B1(n4131), .B2(n4130), .A(n4137), .ZN(n3160) );
  NAND2_X1 U3758 ( .A1(n4788), .A2(n4776), .ZN(n3473) );
  AND2_X1 U3759 ( .A1(n4163), .A2(n4162), .ZN(n4175) );
  OR2_X1 U3760 ( .A1(n4161), .A2(n4160), .ZN(n4163) );
  AND2_X1 U3761 ( .A1(n6420), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4160)
         );
  NAND2_X1 U3762 ( .A1(n3113), .A2(n3158), .ZN(n3157) );
  NOR2_X1 U3763 ( .A1(n4020), .A2(n3193), .ZN(n3192) );
  NOR2_X1 U3764 ( .A1(n5462), .A2(n3197), .ZN(n3196) );
  INV_X1 U3765 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U3766 ( .A1(n3133), .A2(n3210), .ZN(n3209) );
  INV_X1 U3767 ( .A(n5472), .ZN(n3210) );
  INV_X1 U3768 ( .A(n5447), .ZN(n3211) );
  AND2_X1 U3769 ( .A1(n3276), .A2(n5229), .ZN(n3206) );
  AND2_X1 U3770 ( .A1(n3115), .A2(n3277), .ZN(n3276) );
  INV_X1 U3771 ( .A(n5686), .ZN(n3277) );
  AND2_X1 U3772 ( .A1(n4333), .A2(n3660), .ZN(n4381) );
  INV_X1 U3773 ( .A(n3800), .ZN(n3784) );
  OR3_X1 U3774 ( .A1(n3248), .A2(n3247), .A3(n3246), .ZN(n3245) );
  INV_X1 U3775 ( .A(n5348), .ZN(n3246) );
  INV_X1 U3776 ( .A(n5400), .ZN(n3247) );
  OR2_X1 U3777 ( .A1(n5427), .A2(n5416), .ZN(n3248) );
  OAI21_X1 U3778 ( .B1(n3259), .B2(n3256), .A(n3121), .ZN(n3255) );
  NAND2_X1 U3779 ( .A1(n3224), .A2(n5885), .ZN(n3223) );
  INV_X1 U3780 ( .A(n3284), .ZN(n3224) );
  NOR2_X1 U3781 ( .A1(n3101), .A2(n3238), .ZN(n3237) );
  INV_X1 U3782 ( .A(n5683), .ZN(n3238) );
  AND2_X1 U3783 ( .A1(n4447), .A2(n3337), .ZN(n3438) );
  NAND2_X1 U3784 ( .A1(n3444), .A2(n4753), .ZN(n3150) );
  NAND2_X1 U3785 ( .A1(n3513), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3267) );
  INV_X1 U3786 ( .A(n4119), .ZN(n3497) );
  INV_X1 U3787 ( .A(n3150), .ZN(n3149) );
  CLKBUF_X1 U3788 ( .A(n4313), .Z(n4654) );
  XNOR2_X1 U3789 ( .A(n4593), .B(n6495), .ZN(n4712) );
  AOI22_X1 U3790 ( .A1(n3456), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3299) );
  AND3_X1 U3791 ( .A1(n4446), .A2(n4447), .A3(n4324), .ZN(n4439) );
  NOR2_X1 U3792 ( .A1(n4758), .A2(n3095), .ZN(n5611) );
  NAND2_X1 U3793 ( .A1(n6155), .A2(n7027), .ZN(n4530) );
  NAND2_X1 U3794 ( .A1(n5490), .A2(n3137), .ZN(n5461) );
  INV_X1 U3795 ( .A(n5490), .ZN(n5464) );
  NAND2_X1 U3796 ( .A1(n3157), .A2(n3758), .ZN(n3759) );
  NAND2_X1 U3797 ( .A1(n3155), .A2(n3156), .ZN(n3772) );
  INV_X1 U3798 ( .A(n3157), .ZN(n3155) );
  NAND2_X1 U3799 ( .A1(n3719), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3720)
         );
  NAND2_X1 U3800 ( .A1(n3113), .A2(n3154), .ZN(n3153) );
  NAND2_X1 U3801 ( .A1(n4112), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4114)
         );
  INV_X1 U3802 ( .A(n3967), .ZN(n5370) );
  INV_X1 U3803 ( .A(n4086), .ZN(n4112) );
  INV_X1 U3804 ( .A(n4018), .ZN(n4019) );
  NAND2_X1 U3805 ( .A1(n4019), .A2(n3192), .ZN(n4042) );
  OAI21_X1 U3806 ( .B1(n5802), .B2(n3641), .A(n3985), .ZN(n5439) );
  NAND2_X1 U3807 ( .A1(n3935), .A2(n3196), .ZN(n3939) );
  INV_X1 U3808 ( .A(n3897), .ZN(n3935) );
  OR2_X1 U3809 ( .A1(n3894), .A2(n3893), .ZN(n3897) );
  NOR2_X1 U3810 ( .A1(n3201), .A2(n5547), .ZN(n3200) );
  NAND2_X1 U3811 ( .A1(n3827), .A2(n3199), .ZN(n3863) );
  AND2_X1 U3812 ( .A1(n3200), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3199)
         );
  OR2_X1 U3813 ( .A1(n3808), .A2(n3807), .ZN(n3826) );
  NOR2_X1 U3814 ( .A1(n6951), .A2(n3720), .ZN(n3753) );
  NOR2_X1 U3815 ( .A1(n5063), .A2(n3190), .ZN(n3189) );
  INV_X1 U3816 ( .A(n4951), .ZN(n3190) );
  NAND2_X1 U3817 ( .A1(n3116), .A2(n3104), .ZN(n3147) );
  INV_X1 U3818 ( .A(n3165), .ZN(n3164) );
  NAND2_X1 U3819 ( .A1(n4159), .A2(n3161), .ZN(n3166) );
  OAI21_X1 U3820 ( .B1(n3168), .B2(n3167), .A(n6154), .ZN(n3165) );
  AND2_X1 U3821 ( .A1(n3102), .A2(n4428), .ZN(n3263) );
  AND2_X2 U3822 ( .A1(n5384), .A2(n4285), .ZN(n4508) );
  INV_X1 U3823 ( .A(n3266), .ZN(n3203) );
  AND2_X1 U3824 ( .A1(n4407), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3204)
         );
  NOR2_X1 U3825 ( .A1(n5780), .A2(n3266), .ZN(n3264) );
  NOR2_X1 U3826 ( .A1(n5813), .A2(n3229), .ZN(n3228) );
  INV_X1 U3827 ( .A(n5795), .ZN(n3229) );
  INV_X1 U3828 ( .A(n5813), .ZN(n3230) );
  AND2_X1 U3829 ( .A1(n4257), .A2(n5504), .ZN(n5502) );
  NAND2_X1 U3830 ( .A1(n3254), .A2(n3259), .ZN(n5820) );
  AND2_X1 U3831 ( .A1(n4255), .A2(n4254), .ZN(n5506) );
  NAND2_X1 U3832 ( .A1(n4415), .A2(n4414), .ZN(n5840) );
  AND2_X1 U3833 ( .A1(n4247), .A2(n4246), .ZN(n5562) );
  OR2_X1 U3834 ( .A1(n4407), .A2(n6031), .ZN(n5870) );
  NOR2_X1 U3835 ( .A1(n3175), .A2(n3176), .ZN(n3174) );
  INV_X1 U3836 ( .A(n3213), .ZN(n3175) );
  NAND2_X1 U3837 ( .A1(n6362), .A2(n6359), .ZN(n3212) );
  NOR2_X1 U3838 ( .A1(n3151), .A2(n3150), .ZN(n4438) );
  NAND2_X1 U3839 ( .A1(n5609), .A2(n3152), .ZN(n3151) );
  NAND2_X1 U3840 ( .A1(n3219), .A2(n4357), .ZN(n4624) );
  NAND2_X1 U3841 ( .A1(n5137), .A2(n4388), .ZN(n3219) );
  OAI21_X1 U3842 ( .B1(n3501), .B2(n4355), .A(n3225), .ZN(n3495) );
  NOR2_X1 U3843 ( .A1(n4172), .A2(n4174), .ZN(n4573) );
  NAND2_X1 U3844 ( .A1(n3185), .A2(n3251), .ZN(n4960) );
  NOR2_X1 U3845 ( .A1(n3250), .A2(n3097), .ZN(n3251) );
  INV_X1 U3846 ( .A(n3250), .ZN(n6426) );
  AND2_X1 U3847 ( .A1(n3111), .A2(n5136), .ZN(n6474) );
  OR2_X1 U3848 ( .A1(n6596), .A2(n3097), .ZN(n5015) );
  INV_X2 U3849 ( .A(n3419), .ZN(n4758) );
  OR2_X1 U3850 ( .A1(n4906), .A2(n3097), .ZN(n4727) );
  INV_X1 U3851 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U3852 ( .A1(n4439), .A2(n3398), .ZN(n6133) );
  INV_X1 U3853 ( .A(n3641), .ZN(n4183) );
  INV_X1 U3854 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6592) );
  NOR2_X1 U3855 ( .A1(n5608), .A2(n5655), .ZN(n5635) );
  NAND2_X1 U3856 ( .A1(n4307), .A2(n3130), .ZN(n3172) );
  NOR2_X1 U3857 ( .A1(n6269), .A2(n4497), .ZN(n3173) );
  OR2_X1 U3858 ( .A1(n6232), .A2(n5571), .ZN(n5560) );
  NOR2_X1 U3859 ( .A1(n5754), .A2(n3202), .ZN(n6241) );
  INV_X1 U3860 ( .A(n4308), .ZN(n3202) );
  INV_X1 U3861 ( .A(n6252), .ZN(n6277) );
  AND2_X1 U3862 ( .A1(n5754), .A2(n4308), .ZN(n6259) );
  NAND2_X1 U3863 ( .A1(n4495), .A2(n4494), .ZN(n5696) );
  OR3_X1 U3864 ( .A1(n4652), .A2(n6152), .A3(n4781), .ZN(n4495) );
  INV_X1 U3865 ( .A(n4842), .ZN(n5698) );
  NAND2_X1 U3866 ( .A1(n6356), .A2(n4625), .ZN(n6370) );
  INV_X1 U3867 ( .A(n6370), .ZN(n6350) );
  OR2_X1 U3868 ( .A1(n4618), .A2(n6133), .ZN(n6339) );
  INV_X1 U3869 ( .A(n6356), .ZN(n6358) );
  INV_X1 U3870 ( .A(n6080), .ZN(n4461) );
  INV_X1 U3871 ( .A(n6651), .ZN(n6586) );
  OAI21_X1 U3872 ( .B1(n4812), .B2(n6714), .A(n5053), .ZN(n6419) );
  INV_X1 U3873 ( .A(n6115), .ZN(n5333) );
  INV_X1 U3874 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4816) );
  AND2_X1 U3875 ( .A1(n4591), .A2(n4590), .ZN(n4596) );
  NAND2_X1 U3876 ( .A1(n3140), .A2(n3633), .ZN(n3659) );
  INV_X1 U3877 ( .A(n4424), .ZN(n3256) );
  INV_X1 U3878 ( .A(n3634), .ZN(n3633) );
  OR2_X1 U3879 ( .A1(n3654), .A2(n3653), .ZN(n4391) );
  NOR2_X1 U3880 ( .A1(n3525), .A2(n3524), .ZN(n4342) );
  NAND2_X1 U3881 ( .A1(n3095), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4119) );
  AOI21_X1 U3882 ( .B1(n4173), .B2(n5611), .A(n3420), .ZN(n4445) );
  NAND2_X1 U3883 ( .A1(n3426), .A2(n3401), .ZN(n3418) );
  NAND2_X1 U3884 ( .A1(n3419), .A2(n3417), .ZN(n4185) );
  AOI22_X1 U3885 ( .A1(n4097), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U3886 ( .A1(n3484), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3307) );
  INV_X1 U3887 ( .A(n4323), .ZN(n4446) );
  AOI22_X1 U3888 ( .A1(n4100), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3346) );
  INV_X1 U3889 ( .A(n3279), .ZN(n3278) );
  AND2_X1 U3890 ( .A1(n5415), .A2(n3280), .ZN(n3279) );
  NOR2_X1 U3891 ( .A1(n5423), .A2(n3281), .ZN(n3280) );
  INV_X1 U3892 ( .A(n5439), .ZN(n3281) );
  NAND2_X1 U3893 ( .A1(n3275), .A2(n5539), .ZN(n3274) );
  INV_X1 U3894 ( .A(n5306), .ZN(n3142) );
  AND2_X1 U3895 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3574), .ZN(n3637)
         );
  NOR2_X1 U3896 ( .A1(n3589), .A2(n3187), .ZN(n3574) );
  INV_X1 U3897 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3187) );
  INV_X1 U3898 ( .A(n4170), .ZN(n3167) );
  NOR2_X1 U3899 ( .A1(n3167), .A2(n3162), .ZN(n3161) );
  INV_X1 U3900 ( .A(n4158), .ZN(n3162) );
  NOR2_X1 U3901 ( .A1(n3261), .A2(n3258), .ZN(n3257) );
  INV_X1 U3902 ( .A(n4414), .ZN(n3258) );
  INV_X1 U3903 ( .A(n5831), .ZN(n3262) );
  NOR2_X1 U3904 ( .A1(n5530), .A2(n3242), .ZN(n3241) );
  INV_X1 U3905 ( .A(n5543), .ZN(n3242) );
  INV_X1 U3906 ( .A(n5899), .ZN(n3184) );
  INV_X1 U3907 ( .A(n4380), .ZN(n3218) );
  NAND2_X1 U3908 ( .A1(n3112), .A2(n4388), .ZN(n4365) );
  INV_X1 U3909 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U3910 ( .A1(n3454), .A2(n3605), .ZN(n3470) );
  INV_X1 U3911 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3289) );
  INV_X1 U3912 ( .A(n4168), .ZN(n3168) );
  NAND2_X1 U3913 ( .A1(n3159), .A2(n4147), .ZN(n4150) );
  AND2_X1 U3914 ( .A1(n3536), .A2(n4911), .ZN(n5075) );
  INV_X1 U3915 ( .A(n4443), .ZN(n3427) );
  XNOR2_X1 U3916 ( .A(n7028), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5144)
         );
  INV_X1 U3917 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6827) );
  NOR2_X1 U3918 ( .A1(n5461), .A2(n4305), .ZN(n5429) );
  AND2_X1 U3919 ( .A1(n5497), .A2(n3138), .ZN(n5490) );
  AND2_X1 U3920 ( .A1(n6183), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4308) );
  INV_X1 U3921 ( .A(n5648), .ZN(n5615) );
  NAND2_X1 U3922 ( .A1(n4666), .A2(n4612), .ZN(n3243) );
  XNOR2_X1 U3923 ( .A(n3244), .B(n4666), .ZN(n4613) );
  CLKBUF_X1 U3924 ( .A(n5555), .Z(n5556) );
  INV_X1 U3925 ( .A(n5609), .ZN(n4836) );
  AOI21_X1 U3926 ( .B1(n4389), .B2(n3800), .A(n3673), .ZN(n5063) );
  NAND2_X1 U3927 ( .A1(n4019), .A2(n3108), .ZN(n4062) );
  OR2_X1 U3928 ( .A1(n4062), .A2(n5349), .ZN(n4086) );
  NAND2_X1 U3929 ( .A1(n3935), .A2(n3194), .ZN(n3965) );
  NOR2_X1 U3930 ( .A1(n3195), .A2(n3198), .ZN(n3194) );
  INV_X1 U3931 ( .A(n3196), .ZN(n3195) );
  NAND2_X1 U3932 ( .A1(n3208), .A2(n5439), .ZN(n3207) );
  INV_X1 U3933 ( .A(n3209), .ZN(n3208) );
  OAI21_X1 U3934 ( .B1(n5808), .B2(n3641), .A(n3963), .ZN(n5447) );
  OAI21_X1 U3935 ( .B1(n5816), .B2(n3641), .A(n3920), .ZN(n5472) );
  CLKBUF_X1 U3936 ( .A(n5470), .Z(n5471) );
  NAND2_X1 U3937 ( .A1(n3862), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3894)
         );
  INV_X1 U3938 ( .A(n3863), .ZN(n3862) );
  NAND2_X1 U3939 ( .A1(n3273), .A2(n3272), .ZN(n3271) );
  INV_X1 U3940 ( .A(n3274), .ZN(n3273) );
  INV_X1 U3941 ( .A(n5526), .ZN(n3272) );
  CLKBUF_X1 U3942 ( .A(n5495), .Z(n5512) );
  AND2_X1 U3943 ( .A1(n3753), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3754)
         );
  NAND2_X1 U3944 ( .A1(n3754), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3808)
         );
  NAND2_X1 U3945 ( .A1(n3752), .A2(n3751), .ZN(n5681) );
  AND2_X1 U3946 ( .A1(n3735), .A2(n3734), .ZN(n5686) );
  NAND3_X1 U3947 ( .A1(n3637), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n3106), 
        .ZN(n3688) );
  NOR2_X1 U3948 ( .A1(n6981), .A2(n3688), .ZN(n3719) );
  NAND2_X1 U3949 ( .A1(n3637), .A2(n3105), .ZN(n3668) );
  INV_X1 U3950 ( .A(n3663), .ZN(n3664) );
  AND2_X1 U3951 ( .A1(n3637), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3661)
         );
  NAND2_X1 U3952 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3589) );
  OAI21_X1 U3953 ( .B1(n5783), .B2(n3283), .A(n4432), .ZN(n4433) );
  NAND2_X1 U3954 ( .A1(n4512), .A2(n4511), .ZN(n5390) );
  NAND2_X1 U3955 ( .A1(n5388), .A2(n4510), .ZN(n4511) );
  AND2_X1 U3956 ( .A1(n4281), .A2(n4280), .ZN(n5400) );
  AND2_X1 U3957 ( .A1(n4278), .A2(n4277), .ZN(n5416) );
  NOR2_X1 U3958 ( .A1(n3233), .A2(n5797), .ZN(n3227) );
  AND2_X1 U3959 ( .A1(n4268), .A2(n4267), .ZN(n5458) );
  AND3_X1 U3960 ( .A1(n5995), .A2(n4470), .A3(n4469), .ZN(n5974) );
  INV_X1 U3961 ( .A(n5861), .ZN(n5852) );
  NAND2_X1 U3962 ( .A1(n5541), .A2(n5543), .ZN(n5542) );
  NAND2_X1 U3963 ( .A1(n5541), .A2(n3241), .ZN(n5528) );
  AND2_X1 U3964 ( .A1(n4245), .A2(n4244), .ZN(n5575) );
  INV_X1 U3965 ( .A(n5679), .ZN(n4241) );
  CLKBUF_X1 U3966 ( .A(n5677), .Z(n5682) );
  NOR2_X1 U3967 ( .A1(n5587), .A2(n3101), .ZN(n5688) );
  INV_X1 U3968 ( .A(n6054), .ZN(n6038) );
  NAND2_X1 U3969 ( .A1(n3236), .A2(n4232), .ZN(n5690) );
  CLKBUF_X1 U3970 ( .A(n4824), .Z(n4953) );
  NOR2_X2 U3971 ( .A1(n4773), .A2(n4774), .ZN(n4772) );
  AND2_X1 U3972 ( .A1(n4830), .A2(n4359), .ZN(n6362) );
  NAND2_X1 U3973 ( .A1(n4828), .A2(n4829), .ZN(n4830) );
  NAND2_X1 U3974 ( .A1(n4712), .A2(n7027), .ZN(n3555) );
  NAND2_X1 U3975 ( .A1(n3149), .A2(n5609), .ZN(n4653) );
  XNOR2_X1 U3976 ( .A(n4714), .B(n4716), .ZN(n5637) );
  INV_X1 U3977 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4804) );
  AND2_X1 U3979 ( .A1(n4589), .A2(n4588), .ZN(n6121) );
  OAI21_X1 U3980 ( .B1(n6468), .B2(n6467), .A(n6586), .ZN(n6504) );
  CLKBUF_X1 U3981 ( .A(n4813), .Z(n6432) );
  INV_X1 U3982 ( .A(n3417), .ZN(n4733) );
  AND2_X2 U3983 ( .A1(n3303), .A2(n3302), .ZN(n3421) );
  OR2_X1 U3984 ( .A1(n5053), .A2(n4816), .ZN(n4764) );
  AND2_X1 U3985 ( .A1(n4711), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4908)
         );
  NAND2_X1 U3986 ( .A1(n3250), .A2(n4724), .ZN(n4906) );
  AND2_X1 U3987 ( .A1(n6810), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4171) );
  NOR2_X1 U3988 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6795) );
  NAND2_X1 U3989 ( .A1(n3935), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3936)
         );
  NAND2_X1 U3990 ( .A1(n3134), .A2(n3772), .ZN(n5673) );
  AND2_X1 U3991 ( .A1(n6183), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6234) );
  INV_X1 U3992 ( .A(n6241), .ZN(n6207) );
  INV_X1 U3993 ( .A(n6264), .ZN(n6249) );
  OR2_X1 U3994 ( .A1(n5608), .A2(n4295), .ZN(n6269) );
  AND2_X1 U3995 ( .A1(n5635), .A2(n4292), .ZN(n6252) );
  INV_X1 U3996 ( .A(n5696), .ZN(n5684) );
  NOR2_X2 U3997 ( .A1(n5748), .A2(n5357), .ZN(n5732) );
  NOR2_X1 U3998 ( .A1(n5748), .A2(n4845), .ZN(n5749) );
  INV_X1 U3999 ( .A(n5748), .ZN(n5746) );
  OR3_X1 U4000 ( .A1(n4618), .A2(n4617), .A3(n4616), .ZN(n6302) );
  AND2_X2 U4001 ( .A1(n6302), .A2(n6306), .ZN(n6303) );
  INV_X1 U4002 ( .A(n6300), .ZN(n6306) );
  OR2_X1 U4003 ( .A1(n4604), .A2(n4603), .ZN(n4841) );
  INV_X1 U4004 ( .A(n4642), .ZN(n4681) );
  INV_X1 U4005 ( .A(n4681), .ZN(n6328) );
  INV_X1 U4006 ( .A(n4841), .ZN(n6327) );
  XNOR2_X1 U4007 ( .A(n4116), .B(n4115), .ZN(n5754) );
  OR2_X1 U4008 ( .A1(n4114), .A2(n6937), .ZN(n4116) );
  AOI22_X1 U4009 ( .A1(n3571), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5370), .ZN(n5371) );
  NAND2_X1 U4010 ( .A1(n3268), .A2(n5369), .ZN(n5372) );
  INV_X1 U4011 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U4012 ( .A1(n4019), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4021)
         );
  OAI21_X1 U4013 ( .B1(n5414), .B2(n5415), .A(n5403), .ZN(n5786) );
  INV_X1 U4014 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U4015 ( .A1(n3827), .A2(n3200), .ZN(n3846) );
  NAND2_X1 U4016 ( .A1(n3827), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3845)
         );
  NAND2_X1 U4017 ( .A1(n6339), .A2(n4531), .ZN(n6356) );
  NAND2_X1 U4018 ( .A1(n5787), .A2(n3263), .ZN(n3265) );
  NAND2_X1 U4019 ( .A1(n5787), .A2(n3102), .ZN(n5759) );
  INV_X1 U4020 ( .A(n5783), .ZN(n5761) );
  NAND2_X1 U4021 ( .A1(n5787), .A2(n3132), .ZN(n5340) );
  NAND2_X1 U4022 ( .A1(n3231), .A2(n3228), .ZN(n5805) );
  INV_X1 U4023 ( .A(n3235), .ZN(n5812) );
  AND2_X1 U4024 ( .A1(n5541), .A2(n3239), .ZN(n5486) );
  OAI21_X1 U4025 ( .B1(n5840), .B2(n4420), .A(n4419), .ZN(n5833) );
  XNOR2_X1 U4026 ( .A(n3178), .B(n7026), .ZN(n6029) );
  NAND2_X1 U4027 ( .A1(n3180), .A2(n3179), .ZN(n3178) );
  OAI21_X1 U4028 ( .B1(n5861), .B2(n5853), .A(n4407), .ZN(n3179) );
  NAND2_X1 U4029 ( .A1(n5854), .A2(n4524), .ZN(n3180) );
  NAND2_X1 U4030 ( .A1(n5884), .A2(n4413), .ZN(n5877) );
  INV_X1 U4031 ( .A(n6098), .ZN(n6084) );
  NAND2_X1 U4032 ( .A1(n5305), .A2(n5306), .ZN(n3177) );
  NAND2_X1 U4033 ( .A1(n4993), .A2(n4994), .ZN(n3215) );
  OR2_X1 U4034 ( .A1(n6416), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4457)
         );
  INV_X1 U4035 ( .A(n5004), .ZN(n6395) );
  OR2_X1 U4036 ( .A1(n6059), .A2(n6416), .ZN(n6415) );
  INV_X1 U4037 ( .A(n6101), .ZN(n6412) );
  AND2_X1 U4038 ( .A1(n4467), .A2(n4332), .ZN(n6410) );
  NAND2_X1 U4039 ( .A1(n4467), .A2(n4442), .ZN(n6101) );
  INV_X1 U4040 ( .A(n6496), .ZN(n6583) );
  NAND2_X1 U4041 ( .A1(n3613), .A2(n3614), .ZN(n3220) );
  NAND2_X1 U4042 ( .A1(n3612), .A2(n3615), .ZN(n3221) );
  AND2_X1 U4043 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4890) );
  INV_X1 U4044 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6462) );
  INV_X1 U4045 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U4046 ( .A1(n4652), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U4047 ( .A1(n4596), .A2(n4592), .ZN(n6115) );
  OAI21_X1 U4048 ( .B1(n5196), .B2(n5199), .A(n5195), .ZN(n5221) );
  NAND2_X1 U4049 ( .A1(n3185), .A2(n3252), .ZN(n6454) );
  NOR2_X1 U4050 ( .A1(n5189), .A2(n3250), .ZN(n3252) );
  NAND2_X1 U4051 ( .A1(n3185), .A2(n3253), .ZN(n6494) );
  NOR2_X1 U4052 ( .A1(n6595), .A2(n3250), .ZN(n3253) );
  INV_X1 U4053 ( .A(n6637), .ZN(n5287) );
  NOR2_X1 U4054 ( .A1(n4853), .A2(n5053), .ZN(n6649) );
  INV_X1 U4055 ( .A(n6507), .ZN(n6666) );
  NOR2_X1 U4056 ( .A1(n4846), .A2(n5053), .ZN(n6667) );
  NOR2_X1 U4057 ( .A1(n4852), .A2(n5053), .ZN(n6673) );
  NOR2_X1 U4058 ( .A1(n4644), .A2(n5053), .ZN(n6679) );
  INV_X1 U4059 ( .A(n6613), .ZN(n6684) );
  INV_X1 U4060 ( .A(n6523), .ZN(n6690) );
  NOR2_X1 U4061 ( .A1(n4847), .A2(n5053), .ZN(n6691) );
  NOR2_X1 U4062 ( .A1(n4956), .A2(n5053), .ZN(n6697) );
  INV_X1 U4063 ( .A(n6650), .ZN(n6706) );
  INV_X1 U4064 ( .A(n6633), .ZN(n6703) );
  NOR2_X1 U4065 ( .A1(n7079), .A2(n5053), .ZN(n6704) );
  OAI211_X1 U4066 ( .C1(n6586), .C2(n6647), .A(n4729), .B(n6585), .ZN(n4768)
         );
  INV_X1 U4067 ( .A(n4889), .ZN(n4767) );
  OR2_X1 U4068 ( .A1(n4764), .A2(n4748), .ZN(n6544) );
  OR2_X1 U4069 ( .A1(n4764), .A2(n4758), .ZN(n6507) );
  INV_X1 U4070 ( .A(n6667), .ZN(n6556) );
  OR2_X1 U4071 ( .A1(n4764), .A2(n4753), .ZN(n7112) );
  INV_X1 U4072 ( .A(n6673), .ZN(n7113) );
  OR2_X1 U4073 ( .A1(n4764), .A2(n4733), .ZN(n6606) );
  INV_X1 U4074 ( .A(n6679), .ZN(n6562) );
  OR2_X1 U4075 ( .A1(n4764), .A2(n4763), .ZN(n6613) );
  INV_X1 U4076 ( .A(n6685), .ZN(n6565) );
  INV_X1 U4077 ( .A(n6697), .ZN(n6574) );
  OR2_X1 U4078 ( .A1(n4764), .A2(n5698), .ZN(n6633) );
  INV_X1 U4079 ( .A(n6704), .ZN(n6580) );
  INV_X1 U4080 ( .A(n4932), .ZN(n4948) );
  OR2_X1 U4081 ( .A1(n4906), .A2(n6595), .ZN(n5127) );
  INV_X1 U4082 ( .A(n6154), .ZN(n6152) );
  AND2_X1 U4083 ( .A1(n4171), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6154) );
  NOR2_X1 U4084 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6155) );
  INV_X2 U4085 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7027) );
  AND2_X1 U4086 ( .A1(n4557), .A2(n6800), .ZN(n6778) );
  INV_X1 U4087 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4550) );
  NOR2_X1 U4088 ( .A1(n6800), .A2(STATE_REG_2__SCAN_IN), .ZN(n6765) );
  INV_X2 U4089 ( .A(n6789), .ZN(n6800) );
  NOR2_X1 U4090 ( .A1(n5696), .A2(n4497), .ZN(n4498) );
  NAND2_X1 U4091 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  OAI21_X1 U4092 ( .B1(n5718), .B2(n6334), .A(n4535), .ZN(n4536) );
  XNOR2_X1 U4093 ( .A(n6582), .B(n3250), .ZN(n4893) );
  NOR2_X1 U4094 ( .A1(n5470), .A2(n5472), .ZN(n3099) );
  NAND2_X1 U4095 ( .A1(n3191), .A2(n4951), .ZN(n4950) );
  INV_X1 U4096 ( .A(n4407), .ZN(n4524) );
  AND2_X1 U4097 ( .A1(n5064), .A2(n5229), .ZN(n3100) );
  NAND2_X1 U4098 ( .A1(n3099), .A2(n4528), .ZN(n4527) );
  OR2_X1 U4099 ( .A1(n5689), .A2(n5586), .ZN(n3101) );
  NAND2_X1 U4100 ( .A1(n3140), .A2(n3131), .ZN(n4333) );
  INV_X1 U4101 ( .A(n5357), .ZN(n3152) );
  AND2_X1 U4102 ( .A1(n3264), .A2(n4502), .ZN(n3102) );
  AND2_X1 U4103 ( .A1(n4398), .A2(n4387), .ZN(n3103) );
  OR2_X1 U4104 ( .A1(n3577), .A2(n3568), .ZN(n3104) );
  AND2_X1 U4105 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3105) );
  AND2_X1 U4106 ( .A1(n3105), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3106)
         );
  OR2_X1 U4107 ( .A1(n3758), .A2(n5675), .ZN(n3107) );
  AND2_X1 U4108 ( .A1(n3192), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3108)
         );
  NAND2_X2 U4109 ( .A1(n4733), .A2(n4187), .ZN(n4194) );
  NOR2_X2 U4110 ( .A1(n5015), .A2(n6473), .ZN(n3109) );
  OR2_X1 U4111 ( .A1(n5555), .A2(n3274), .ZN(n5525) );
  AND2_X1 U4112 ( .A1(n5064), .A2(n3206), .ZN(n3110) );
  NOR2_X1 U4113 ( .A1(n5425), .A2(n3248), .ZN(n5399) );
  NAND2_X1 U4114 ( .A1(n3100), .A2(n5247), .ZN(n5246) );
  AND2_X1 U4115 ( .A1(n4815), .A2(n3250), .ZN(n3111) );
  AND2_X1 U4116 ( .A1(n3189), .A2(n3191), .ZN(n5064) );
  AND2_X1 U4117 ( .A1(n3635), .A2(n3148), .ZN(n3112) );
  AND2_X1 U4118 ( .A1(n3188), .A2(n3191), .ZN(n3113) );
  NOR2_X1 U4119 ( .A1(n5390), .A2(n5389), .ZN(n3114) );
  AND2_X1 U4120 ( .A1(n5247), .A2(n3718), .ZN(n3115) );
  NAND2_X1 U4121 ( .A1(n3174), .A2(n3214), .ZN(n5305) );
  NAND2_X1 U4122 ( .A1(n3177), .A2(n4398), .ZN(n5293) );
  OR2_X1 U4123 ( .A1(n3577), .A2(n3800), .ZN(n3116) );
  NOR2_X1 U4124 ( .A1(n5555), .A2(n3271), .ZN(n5511) );
  NAND2_X1 U4125 ( .A1(n3772), .A2(n3759), .ZN(n5674) );
  AND2_X1 U4126 ( .A1(n3257), .A2(n4424), .ZN(n3117) );
  AND2_X1 U4127 ( .A1(n3228), .A2(n5967), .ZN(n3118) );
  AND2_X1 U4128 ( .A1(n6090), .A2(n5890), .ZN(n3119) );
  INV_X1 U4129 ( .A(n4387), .ZN(n3176) );
  NAND2_X1 U4130 ( .A1(n3429), .A2(n4842), .ZN(n4319) );
  NOR2_X1 U4131 ( .A1(n4407), .A2(n6062), .ZN(n3120) );
  INV_X1 U4132 ( .A(n3249), .ZN(n5426) );
  NOR2_X1 U4133 ( .A1(n5425), .A2(n5427), .ZN(n3249) );
  OR2_X1 U4134 ( .A1(n4407), .A2(n4423), .ZN(n3121) );
  NAND2_X1 U4135 ( .A1(n3100), .A2(n3115), .ZN(n5583) );
  AND2_X1 U4136 ( .A1(n5437), .A2(n3280), .ZN(n5414) );
  NAND2_X1 U4137 ( .A1(n3267), .A2(n3496), .ZN(n3601) );
  INV_X1 U4138 ( .A(n5586), .ZN(n4232) );
  AND2_X1 U4139 ( .A1(n4231), .A2(n4230), .ZN(n5586) );
  NAND2_X1 U4140 ( .A1(n5787), .A2(n3264), .ZN(n3122) );
  AND2_X2 U4141 ( .A1(n4788), .A2(n4777), .ZN(n3339) );
  OR2_X1 U4142 ( .A1(n5901), .A2(n5899), .ZN(n3123) );
  AND2_X1 U4143 ( .A1(n3239), .A2(n4261), .ZN(n3124) );
  AND2_X1 U4144 ( .A1(n3567), .A2(n3566), .ZN(n3569) );
  INV_X1 U4145 ( .A(n3569), .ZN(n3568) );
  AND2_X1 U4146 ( .A1(n4753), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3125) );
  AND2_X1 U4147 ( .A1(n3424), .A2(n3423), .ZN(n3126) );
  AND2_X1 U4148 ( .A1(n4407), .A2(n5999), .ZN(n3127) );
  NOR2_X1 U4149 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4023) );
  INV_X1 U4150 ( .A(n4023), .ZN(n3641) );
  NAND2_X1 U4151 ( .A1(n3106), .A2(n3637), .ZN(n3128) );
  AND3_X1 U4152 ( .A1(n4314), .A2(n4187), .A3(n4296), .ZN(n3129) );
  NAND2_X1 U4153 ( .A1(n3215), .A2(n4380), .ZN(n5183) );
  NOR2_X1 U4154 ( .A1(n4310), .A2(n3173), .ZN(n3130) );
  AND2_X1 U4155 ( .A1(n3633), .A2(n3657), .ZN(n3131) );
  AND2_X1 U4156 ( .A1(n3203), .A2(n3204), .ZN(n3132) );
  INV_X1 U4157 ( .A(n3233), .ZN(n3232) );
  NOR2_X1 U4158 ( .A1(n4524), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3233)
         );
  INV_X1 U4159 ( .A(n5675), .ZN(n3771) );
  AND2_X1 U4160 ( .A1(n3211), .A2(n4528), .ZN(n3133) );
  AND2_X1 U4161 ( .A1(n3759), .A2(n3771), .ZN(n3134) );
  NOR2_X1 U4162 ( .A1(n5405), .A2(n3278), .ZN(n3135) );
  OR2_X1 U4163 ( .A1(n3156), .A2(n3771), .ZN(n3136) );
  NAND2_X1 U4164 ( .A1(n4613), .A2(n4612), .ZN(n4611) );
  INV_X1 U4165 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3193) );
  AND2_X1 U4166 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n3137) );
  AND2_X1 U4167 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n3138) );
  NOR4_X2 U4168 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n6785)
         );
  AND2_X2 U4169 ( .A1(n3139), .A2(n3531), .ZN(n3579) );
  XNOR2_X1 U4170 ( .A(n3587), .B(n3139), .ZN(n4340) );
  AND2_X2 U4171 ( .A1(n4748), .A2(n4758), .ZN(n5609) );
  AND2_X4 U4172 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4777) );
  NAND3_X1 U4173 ( .A1(n3143), .A2(n3141), .A3(n5294), .ZN(n4406) );
  NAND2_X1 U4174 ( .A1(n3142), .A2(n4398), .ZN(n3141) );
  XNOR2_X1 U4175 ( .A(n4397), .B(n4396), .ZN(n5306) );
  NAND3_X1 U4176 ( .A1(n3214), .A2(n3213), .A3(n3103), .ZN(n3143) );
  OR2_X2 U4177 ( .A1(n5821), .A2(n3127), .ZN(n3231) );
  OAI21_X1 U4178 ( .B1(n3635), .B2(n3577), .A(n3145), .ZN(n4702) );
  NAND2_X1 U4179 ( .A1(n3146), .A2(n3147), .ZN(n3145) );
  NAND3_X1 U4180 ( .A1(n3579), .A2(n3116), .A3(n4724), .ZN(n3146) );
  NAND4_X1 U4181 ( .A1(n5609), .A2(n3444), .A3(n3125), .A4(n3152), .ZN(n3445)
         );
  NAND2_X2 U4182 ( .A1(n5568), .A2(n5569), .ZN(n5555) );
  INV_X1 U4183 ( .A(n3758), .ZN(n3156) );
  NAND2_X2 U4184 ( .A1(n3163), .A2(n4170), .ZN(n4652) );
  NAND3_X1 U4185 ( .A1(n4306), .A2(n3171), .A3(n3170), .ZN(U2797) );
  INV_X2 U4187 ( .A(n4187), .ZN(n4748) );
  INV_X2 U4188 ( .A(n6232), .ZN(n6263) );
  NAND2_X4 U4189 ( .A1(n3093), .A2(n3129), .ZN(n6232) );
  NOR2_X1 U4190 ( .A1(n5901), .A2(n3183), .ZN(n4412) );
  OAI21_X2 U4191 ( .B1(n3579), .B2(n4724), .A(n3578), .ZN(n3185) );
  NAND2_X2 U4192 ( .A1(n3555), .A2(n3554), .ZN(n4724) );
  NAND2_X1 U4193 ( .A1(n3186), .A2(n3618), .ZN(n3617) );
  NAND2_X1 U4194 ( .A1(n3588), .A2(n3967), .ZN(n3186) );
  OR2_X1 U4195 ( .A1(n3186), .A2(n3618), .ZN(n4679) );
  OR2_X2 U4196 ( .A1(n5555), .A2(n3269), .ZN(n5495) );
  INV_X1 U4197 ( .A(n5063), .ZN(n3188) );
  INV_X1 U4198 ( .A(n4821), .ZN(n3191) );
  INV_X1 U4199 ( .A(n4042), .ZN(n4061) );
  INV_X1 U4200 ( .A(n3939), .ZN(n3964) );
  INV_X1 U4201 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3198) );
  INV_X1 U4202 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3201) );
  NAND3_X1 U4203 ( .A1(n4333), .A2(n3660), .A3(n4388), .ZN(n4384) );
  NAND3_X1 U4204 ( .A1(n4993), .A2(n5184), .A3(n3216), .ZN(n3214) );
  NAND3_X1 U4205 ( .A1(n3216), .A2(n5184), .A3(n3218), .ZN(n3213) );
  INV_X1 U4206 ( .A(n4994), .ZN(n3217) );
  NOR2_X1 U4207 ( .A1(n4412), .A2(n3284), .ZN(n5886) );
  NAND3_X1 U4208 ( .A1(n3503), .A2(n4763), .A3(n4355), .ZN(n3225) );
  NAND2_X1 U4209 ( .A1(n3231), .A2(n3230), .ZN(n3235) );
  INV_X1 U4210 ( .A(n3231), .ZN(n5814) );
  NAND2_X1 U4211 ( .A1(n3235), .A2(n3227), .ZN(n3226) );
  NAND2_X1 U4212 ( .A1(n3235), .A2(n3232), .ZN(n5796) );
  NAND2_X1 U4213 ( .A1(n3234), .A2(n3226), .ZN(n5798) );
  INV_X1 U4214 ( .A(n5587), .ZN(n3236) );
  NAND2_X1 U4215 ( .A1(n3236), .A2(n3237), .ZN(n5677) );
  NAND2_X1 U4216 ( .A1(n5541), .A2(n3124), .ZN(n5476) );
  NAND2_X1 U4217 ( .A1(n3244), .A2(n3243), .ZN(n4675) );
  NOR2_X2 U4218 ( .A1(n5425), .A2(n3245), .ZN(n4285) );
  NAND2_X1 U4219 ( .A1(n4340), .A2(n4388), .ZN(n4345) );
  CLKBUF_X1 U4220 ( .A(n4340), .Z(n3250) );
  NAND2_X1 U4221 ( .A1(n4415), .A2(n3257), .ZN(n3254) );
  NAND2_X1 U4222 ( .A1(n4505), .A2(n3265), .ZN(n4507) );
  NOR2_X1 U4223 ( .A1(n4524), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3266)
         );
  AND2_X2 U4224 ( .A1(n3601), .A2(n3602), .ZN(n4714) );
  NAND4_X1 U4225 ( .A1(n3425), .A2(n3126), .A3(n3437), .A4(n4451), .ZN(n3602)
         );
  OAI21_X2 U4226 ( .B1(n5909), .B2(n4408), .A(n4409), .ZN(n5901) );
  AOI21_X1 U4227 ( .B1(n5381), .B2(n5382), .A(n3268), .ZN(n5767) );
  NAND3_X1 U4228 ( .A1(n3579), .A2(n4724), .A3(n3568), .ZN(n3635) );
  NOR2_X1 U4229 ( .A1(n5555), .A2(n5557), .ZN(n5538) );
  INV_X1 U4230 ( .A(n5557), .ZN(n3275) );
  NAND2_X1 U4231 ( .A1(n5437), .A2(n3279), .ZN(n5403) );
  AND2_X2 U4232 ( .A1(n5437), .A2(n3135), .ZN(n5342) );
  NAND2_X1 U4233 ( .A1(n4213), .A2(n4212), .ZN(n4824) );
  INV_X1 U4234 ( .A(n4705), .ZN(n4213) );
  NAND2_X1 U4235 ( .A1(n4242), .A2(n4241), .ZN(n5574) );
  INV_X1 U4236 ( .A(n5677), .ZN(n4242) );
  OR2_X4 U4237 ( .A1(n5473), .A2(n5458), .ZN(n5460) );
  AND2_X2 U4238 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4789) );
  AND2_X2 U4239 ( .A1(n3289), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3296)
         );
  INV_X4 U4240 ( .A(n4284), .ZN(n4199) );
  AOI22_X1 U4241 ( .A1(n3472), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3357) );
  INV_X1 U4242 ( .A(n4319), .ZN(n3439) );
  AOI22_X1 U4243 ( .A1(n3096), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3290) );
  OAI21_X1 U4244 ( .B1(n4291), .B2(n4513), .A(n4290), .ZN(n4496) );
  CLKBUF_X1 U4245 ( .A(n5342), .Z(n5404) );
  OR2_X2 U4246 ( .A1(n5748), .A2(n4844), .ZN(n5747) );
  AND2_X2 U4247 ( .A1(n4841), .A2(n4840), .ZN(n5748) );
  INV_X1 U4248 ( .A(READY_N), .ZN(n4601) );
  AND2_X1 U4249 ( .A1(n4890), .A2(n7027), .ZN(n6300) );
  AND4_X1 U4250 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3282)
         );
  INV_X1 U4251 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U4252 ( .A1(n5696), .A2(n5698), .ZN(n5697) );
  INV_X1 U4253 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6981) );
  INV_X1 U4254 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5462) );
  INV_X1 U4255 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6951) );
  INV_X1 U4256 ( .A(n6377), .ZN(n6396) );
  AND2_X1 U4257 ( .A1(n4425), .A2(n4430), .ZN(n3283) );
  NAND2_X1 U4258 ( .A1(n4365), .A2(n4364), .ZN(n4367) );
  NAND2_X1 U4259 ( .A1(n5898), .A2(n4411), .ZN(n3284) );
  AND4_X1 U4260 ( .A1(n3398), .A2(STATE2_REG_0__SCAN_IN), .A3(n4748), .A4(
        n4758), .ZN(n3286) );
  AND2_X1 U4261 ( .A1(n4187), .A2(n4443), .ZN(n3420) );
  AOI22_X1 U4262 ( .A1(n4100), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3393) );
  OR2_X1 U4263 ( .A1(n3452), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3453)
         );
  OR2_X1 U4264 ( .A1(n3361), .A2(n3324), .ZN(n3327) );
  AND2_X1 U4265 ( .A1(n7028), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4132)
         );
  OR2_X1 U4266 ( .A1(n3565), .A2(n3564), .ZN(n4370) );
  NAND2_X1 U4267 ( .A1(n4067), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3369) );
  INV_X1 U4268 ( .A(n5585), .ZN(n3718) );
  AND2_X1 U4269 ( .A1(n3997), .A2(n3996), .ZN(n4013) );
  AND2_X1 U4270 ( .A1(n3632), .A2(n3631), .ZN(n3634) );
  AND2_X2 U4271 ( .A1(n3287), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3295)
         );
  OR3_X1 U4272 ( .A1(n4161), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6420), 
        .ZN(n4176) );
  OR2_X1 U4273 ( .A1(n3981), .A2(n3980), .ZN(n3997) );
  INV_X1 U4274 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3893) );
  NOR2_X1 U4275 ( .A1(n4334), .A2(n4376), .ZN(n4335) );
  OR2_X1 U4276 ( .A1(n3630), .A2(n3629), .ZN(n4373) );
  OR2_X1 U4277 ( .A1(n3553), .A2(n3552), .ZN(n4336) );
  OR2_X1 U4278 ( .A1(n3809), .A2(n3811), .ZN(n5315) );
  INV_X1 U4279 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5517) );
  INV_X1 U4280 ( .A(n5249), .ZN(n4226) );
  NAND2_X1 U4281 ( .A1(n4580), .A2(n4579), .ZN(n4839) );
  NAND2_X1 U4282 ( .A1(n5783), .A2(n4435), .ZN(n4436) );
  AND2_X1 U4283 ( .A1(n4524), .A2(n5339), .ZN(n5779) );
  INV_X1 U4284 ( .A(n4388), .ZN(n4376) );
  AND2_X1 U4285 ( .A1(n4467), .A2(n4456), .ZN(n6055) );
  OR2_X1 U4286 ( .A1(n4727), .A2(n6467), .ZN(n4814) );
  NAND2_X1 U4287 ( .A1(n3495), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3612) );
  OR2_X1 U4288 ( .A1(n6651), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4564) );
  AND2_X1 U4289 ( .A1(n6259), .A2(n4539), .ZN(n4310) );
  NAND2_X1 U4290 ( .A1(n4772), .A2(n4706), .ZN(n4705) );
  AOI21_X1 U4291 ( .B1(n4839), .B2(n6154), .A(n4838), .ZN(n4840) );
  INV_X1 U4292 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4506) );
  OR2_X1 U4293 ( .A1(n4346), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6360)
         );
  AND2_X1 U4294 ( .A1(n4573), .A2(n4758), .ZN(n4595) );
  NAND2_X1 U4295 ( .A1(n6145), .A2(n4721), .ZN(n4722) );
  NAND2_X1 U4296 ( .A1(n4961), .A2(n6473), .ZN(n5131) );
  AND2_X1 U4297 ( .A1(n5140), .A2(n5139), .ZN(n5195) );
  OR2_X1 U4298 ( .A1(n4957), .A2(n5625), .ZN(n5057) );
  OR2_X1 U4299 ( .A1(n6651), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5190) );
  AOI21_X1 U4300 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7028), .A(n5053), .ZN(
        n6585) );
  INV_X1 U4301 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6461) );
  OR2_X1 U4302 ( .A1(n4764), .A2(n3421), .ZN(n6625) );
  OR2_X1 U4303 ( .A1(n4906), .A2(n5189), .ZN(n4932) );
  OR2_X1 U4304 ( .A1(n4559), .A2(n6152), .ZN(n4565) );
  OR2_X1 U4305 ( .A1(n5580), .A2(n4298), .ZN(n5527) );
  INV_X1 U4306 ( .A(n6330), .ZN(n6324) );
  OR2_X1 U4307 ( .A1(n4654), .A2(n6794), .ZN(n4615) );
  AND2_X1 U4308 ( .A1(n5673), .A2(n5676), .ZN(n6189) );
  NAND2_X1 U4309 ( .A1(n6592), .A2(n4816), .ZN(n6651) );
  INV_X1 U4310 ( .A(n6339), .ZN(n6366) );
  AOI21_X1 U4311 ( .B1(n4484), .B2(n4483), .A(n4482), .ZN(n4485) );
  INV_X1 U4312 ( .A(n5637), .ZN(n4957) );
  AND2_X1 U4313 ( .A1(n4573), .A2(n4602), .ZN(n6117) );
  OR2_X1 U4314 ( .A1(n6121), .A2(n6152), .ZN(n4591) );
  OAI211_X1 U4315 ( .C1(n4966), .C2(n4965), .A(n6585), .B(n4964), .ZN(n4989)
         );
  INV_X1 U4316 ( .A(n6454), .ZN(n5225) );
  INV_X1 U4317 ( .A(n6494), .ZN(n6456) );
  OAI21_X1 U4318 ( .B1(n6504), .B2(n6472), .A(n6471), .ZN(n6491) );
  AND2_X1 U4319 ( .A1(n6474), .A2(n6473), .ZN(n6534) );
  NAND4_X1 U4320 ( .A1(n5143), .A2(n5195), .A3(n5142), .A4(n5141), .ZN(n5175)
         );
  AND2_X1 U4321 ( .A1(n3111), .A2(n5254), .ZN(n6576) );
  INV_X1 U4322 ( .A(n6570), .ZN(n7116) );
  OAI211_X1 U4323 ( .C1(n5020), .C2(n5019), .A(n6585), .B(n5018), .ZN(n5043)
         );
  OAI21_X1 U4324 ( .B1(n5263), .B2(n6584), .A(n5262), .ZN(n5289) );
  INV_X1 U4325 ( .A(n6711), .ZN(n6652) );
  AND2_X1 U4326 ( .A1(n5255), .A2(n5254), .ZN(n6637) );
  INV_X1 U4327 ( .A(n7112), .ZN(n6672) );
  NAND2_X1 U4328 ( .A1(n6432), .A2(n6426), .ZN(n6596) );
  NOR2_X1 U4329 ( .A1(n4849), .A2(n5053), .ZN(n6685) );
  OAI21_X1 U4330 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n4883) );
  AND2_X1 U4331 ( .A1(n7027), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4529) );
  INV_X1 U4332 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6943) );
  INV_X1 U4333 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6467) );
  INV_X1 U4334 ( .A(n6234), .ZN(n6266) );
  INV_X1 U4335 ( .A(n5858), .ZN(n5731) );
  INV_X1 U4336 ( .A(n5896), .ZN(n6195) );
  INV_X1 U4337 ( .A(n5749), .ZN(n5744) );
  INV_X1 U4338 ( .A(n6303), .ZN(n6299) );
  OR2_X1 U4339 ( .A1(n4618), .A2(n4615), .ZN(n6330) );
  INV_X1 U4340 ( .A(n6189), .ZN(n5889) );
  INV_X1 U4341 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U4342 ( .B1(n3285), .B2(n6101), .A(n4485), .ZN(n4486) );
  NAND2_X1 U4343 ( .A1(n5973), .A2(n6412), .ZN(n5980) );
  INV_X1 U4344 ( .A(n6410), .ZN(n6398) );
  INV_X1 U4345 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6420) );
  INV_X1 U4346 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U4347 ( .A1(n4963), .A2(n4965), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4959), .ZN(n4992) );
  INV_X1 U4348 ( .A(n5191), .ZN(n5228) );
  AOI21_X1 U4349 ( .B1(n6499), .B2(n6503), .A(n6498), .ZN(n6539) );
  INV_X1 U4350 ( .A(n6533), .ZN(n5182) );
  OR2_X1 U4351 ( .A1(n5015), .A2(n5137), .ZN(n7121) );
  AOI22_X1 U4352 ( .A1(n5017), .A2(n5019), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5014), .ZN(n5046) );
  AOI22_X1 U4353 ( .A1(n5259), .A2(n6584), .B1(n6658), .B2(n5258), .ZN(n5292)
         );
  AOI21_X1 U4354 ( .B1(n6588), .B2(n6593), .A(n6587), .ZN(n6641) );
  OR2_X1 U4355 ( .A1(n6596), .A2(n6595), .ZN(n6711) );
  INV_X1 U4356 ( .A(n6649), .ZN(n6553) );
  INV_X1 U4357 ( .A(n6691), .ZN(n6568) );
  INV_X1 U4358 ( .A(n6609), .ZN(n6683) );
  OR2_X1 U4359 ( .A1(n4727), .A2(n6473), .ZN(n4889) );
  INV_X1 U4360 ( .A(n6778), .ZN(n6718) );
  AND2_X1 U4361 ( .A1(n6943), .A2(STATE_REG_1__SCAN_IN), .ZN(n6789) );
  INV_X1 U4362 ( .A(n6765), .ZN(n6773) );
  OAI21_X1 U4363 ( .B1(n5365), .B2(n6334), .A(n4546), .ZN(U2956) );
  AND2_X2 U4364 ( .A1(n5321), .A2(n3296), .ZN(n4067) );
  AOI22_X1 U4365 ( .A1(n3484), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3294) );
  AND2_X2 U4366 ( .A1(n5321), .A2(n4789), .ZN(n3315) );
  AOI22_X1 U4367 ( .A1(n3314), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3291) );
  NOR2_X4 U4368 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4776) );
  AND2_X2 U4369 ( .A1(n3297), .A2(n4776), .ZN(n3338) );
  AND2_X1 U4370 ( .A1(n3291), .A2(n3290), .ZN(n3293) );
  AOI22_X1 U4371 ( .A1(n4099), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3292) );
  AND2_X4 U4372 ( .A1(n3297), .A2(n5321), .ZN(n4073) );
  NAND2_X2 U4373 ( .A1(n3296), .A2(n4777), .ZN(n3462) );
  INV_X2 U4374 ( .A(n3462), .ZN(n3402) );
  AOI22_X1 U4375 ( .A1(n4073), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3301) );
  AND2_X2 U4376 ( .A1(n3296), .A2(n4776), .ZN(n3903) );
  AOI22_X1 U4377 ( .A1(n3344), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3300) );
  INV_X2 U4378 ( .A(n3361), .ZN(n3456) );
  AND2_X2 U4379 ( .A1(n4777), .A2(n4789), .ZN(n3392) );
  AND2_X2 U4380 ( .A1(n4776), .A2(n4789), .ZN(n3345) );
  AOI22_X1 U4381 ( .A1(n4100), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4382 ( .A1(n3472), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4383 ( .A1(n4099), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4384 ( .A1(n3344), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4385 ( .A1(n3456), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4386 ( .A1(n3461), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4387 ( .A1(n4073), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4388 ( .A1(n4100), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3308) );
  AND4_X2 U4389 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3312)
         );
  NAND2_X1 U4390 ( .A1(n3421), .A2(n3401), .ZN(n4843) );
  BUF_X4 U4391 ( .A(n3314), .Z(n4097) );
  NAND2_X1 U4392 ( .A1(n4097), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4393 ( .A1(n3315), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4394 ( .A1(n4099), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4395 ( .A1(n3339), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4396 ( .A1(n3484), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4397 ( .A1(n3472), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3322)
         );
  NAND2_X1 U4398 ( .A1(n3644), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4399 ( .A1(n4067), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4400 ( .A1(n4100), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3328)
         );
  INV_X1 U4401 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4402 ( .A1(n3392), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4403 ( .A1(n3345), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3325)
         );
  NAND2_X1 U4404 ( .A1(n3344), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4405 ( .A1(n4073), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4406 ( .A1(n3903), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4407 ( .A1(n3402), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3329) );
  INV_X1 U4408 ( .A(n3401), .ZN(n3337) );
  NAND2_X1 U4409 ( .A1(n3337), .A2(n3570), .ZN(n3356) );
  AOI22_X1 U4410 ( .A1(n3484), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4411 ( .A1(n3096), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4412 ( .A1(n4097), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4413 ( .A1(n4099), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3340) );
  NAND4_X1 U4414 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3351)
         );
  AOI22_X1 U4415 ( .A1(n3344), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4416 ( .A1(n4073), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3348) );
  NAND4_X1 U4417 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3350)
         );
  AND2_X1 U4418 ( .A1(n3356), .A2(n4842), .ZN(n3352) );
  NAND2_X1 U4419 ( .A1(n3353), .A2(n3352), .ZN(n4323) );
  AND2_X1 U4420 ( .A1(n4843), .A2(n4489), .ZN(n3354) );
  NOR2_X1 U4421 ( .A1(n4323), .A2(n3354), .ZN(n3435) );
  AND2_X2 U4422 ( .A1(n3356), .A2(n3426), .ZN(n3429) );
  AOI22_X1 U4423 ( .A1(n4099), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4424 ( .A1(n3484), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4425 ( .A1(n4100), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4426 ( .A1(n4073), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4427 ( .A1(n3344), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4428 ( .A1(n3456), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3362) );
  NAND2_X2 U4429 ( .A1(n3367), .A2(n3366), .ZN(n3419) );
  NAND2_X1 U4430 ( .A1(n4097), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4431 ( .A1(n3484), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4432 ( .A1(n3339), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U4433 ( .A1(n4100), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3375)
         );
  NAND2_X1 U4434 ( .A1(n3472), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3374)
         );
  NAND2_X1 U4435 ( .A1(n4073), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4436 ( .A1(n3903), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4437 ( .A1(n3315), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3379)
         );
  NAND2_X1 U4438 ( .A1(n3644), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U4439 ( .A1(n3456), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U4440 ( .A1(n4099), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3376) );
  AND4_X2 U4441 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3385)
         );
  NAND2_X1 U4442 ( .A1(n3344), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4443 ( .A1(n3402), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4444 ( .A1(n3345), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3381)
         );
  NAND2_X1 U4445 ( .A1(n3392), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3380)
         );
  AOI22_X1 U4446 ( .A1(n3484), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4447 ( .A1(n3472), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3644), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4448 ( .A1(n4097), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4449 ( .A1(n4099), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3388) );
  AND4_X2 U4450 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3397)
         );
  AOI22_X1 U4451 ( .A1(n3344), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4452 ( .A1(n4073), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4453 ( .A1(n3456), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3394) );
  NAND2_X2 U4454 ( .A1(n3397), .A2(n3282), .ZN(n3417) );
  INV_X1 U4455 ( .A(n4185), .ZN(n3399) );
  INV_X1 U4456 ( .A(n3418), .ZN(n3398) );
  NAND2_X2 U4457 ( .A1(n3399), .A2(n3398), .ZN(n4454) );
  INV_X1 U4458 ( .A(n4454), .ZN(n3400) );
  XNOR2_X1 U4459 ( .A(n4550), .B(STATE_REG_1__SCAN_IN), .ZN(n4293) );
  NOR2_X1 U4460 ( .A1(n3419), .A2(n4293), .ZN(n3441) );
  AOI22_X1 U4461 ( .A1(n3903), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4462 ( .A1(n3472), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3456), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4463 ( .A1(n3484), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4464 ( .A1(n3314), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4465 ( .A1(n3344), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4073), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4466 ( .A1(n4099), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4467 ( .A1(n4100), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4468 ( .A1(n3461), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3407) );
  OAI211_X1 U4469 ( .C1(n3441), .C2(n3810), .A(n4447), .B(n3095), .ZN(n3414)
         );
  INV_X1 U4470 ( .A(n4843), .ZN(n4321) );
  NAND3_X1 U4471 ( .A1(n4447), .A2(n4321), .A3(n4758), .ZN(n3413) );
  NAND2_X1 U4472 ( .A1(n3414), .A2(n3413), .ZN(n3415) );
  NAND3_X1 U4473 ( .A1(n3435), .A2(n3425), .A3(n3415), .ZN(n3416) );
  NAND2_X1 U4474 ( .A1(n3416), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3448) );
  INV_X1 U4475 ( .A(n3448), .ZN(n3513) );
  MUX2_X1 U4476 ( .A(n4171), .B(n4530), .S(n7028), .Z(n3496) );
  NAND2_X1 U4477 ( .A1(n4843), .A2(n3417), .ZN(n3432) );
  NAND2_X1 U4478 ( .A1(n3432), .A2(n4320), .ZN(n3424) );
  INV_X1 U4479 ( .A(n6155), .ZN(n6113) );
  NOR2_X1 U4480 ( .A1(n6113), .A2(n7027), .ZN(n3422) );
  INV_X2 U4481 ( .A(n3421), .ZN(n3570) );
  OAI21_X1 U4482 ( .B1(n4763), .B2(n3570), .A(n3810), .ZN(n3428) );
  NAND2_X1 U4483 ( .A1(n3428), .A2(n4753), .ZN(n3431) );
  NAND3_X1 U4484 ( .A1(n3809), .A2(n4443), .A3(n3429), .ZN(n3430) );
  NAND2_X1 U4485 ( .A1(n3431), .A2(n3430), .ZN(n3434) );
  NAND2_X1 U4486 ( .A1(n3434), .A2(n3433), .ZN(n4172) );
  NAND2_X1 U4487 ( .A1(n4172), .A2(n5609), .ZN(n4451) );
  INV_X1 U4488 ( .A(n3435), .ZN(n3436) );
  OAI21_X1 U4489 ( .B1(n3436), .B2(n4733), .A(n4602), .ZN(n3437) );
  NAND2_X1 U4490 ( .A1(n3439), .A2(n3438), .ZN(n4313) );
  INV_X1 U4491 ( .A(n4313), .ZN(n3440) );
  NAND2_X2 U4492 ( .A1(n3440), .A2(n4187), .ZN(n4568) );
  INV_X1 U4493 ( .A(n3441), .ZN(n3442) );
  NAND2_X1 U4494 ( .A1(n3442), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3447) );
  INV_X1 U4495 ( .A(n4172), .ZN(n3443) );
  NAND2_X1 U4496 ( .A1(n3443), .A2(n3286), .ZN(n3446) );
  NOR2_X1 U4497 ( .A1(n3810), .A2(n3417), .ZN(n3444) );
  NAND2_X1 U4498 ( .A1(n3570), .A2(n4842), .ZN(n5357) );
  OAI211_X2 U4499 ( .C1(n4568), .C2(n3447), .A(n3446), .B(n3445), .ZN(n3450)
         );
  INV_X1 U4500 ( .A(n4530), .ZN(n3538) );
  INV_X1 U4501 ( .A(n4171), .ZN(n3537) );
  AOI22_X1 U4502 ( .A1(n3538), .A2(n5144), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3537), .ZN(n3451) );
  OAI21_X1 U4503 ( .B1(n3448), .B2(n3287), .A(n3451), .ZN(n3449) );
  OR2_X2 U4504 ( .A1(n3450), .A2(n3449), .ZN(n3510) );
  INV_X1 U4505 ( .A(n3451), .ZN(n3452) );
  NAND2_X1 U4506 ( .A1(n3450), .A2(n3453), .ZN(n3511) );
  NAND2_X1 U4507 ( .A1(n3510), .A2(n3511), .ZN(n4715) );
  NAND3_X1 U4508 ( .A1(n4714), .A2(n4715), .A3(n7027), .ZN(n3471) );
  INV_X1 U4509 ( .A(n3541), .ZN(n3504) );
  AOI22_X1 U4510 ( .A1(n4098), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4511 ( .A1(n3884), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4073), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4512 ( .A1(n4068), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4513 ( .A1(n4074), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3457) );
  NAND4_X1 U4514 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n3468)
         );
  AOI22_X1 U4515 ( .A1(n4050), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3466) );
  INV_X2 U4516 ( .A(n3462), .ZN(n4091) );
  AOI22_X1 U4517 ( .A1(n3547), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4518 ( .A1(n3971), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4519 ( .A1(n4049), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4520 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3467)
         );
  NAND2_X1 U4521 ( .A1(n3504), .A2(n4348), .ZN(n3469) );
  NAND3_X1 U4522 ( .A1(n3471), .A2(n3470), .A3(n3469), .ZN(n3592) );
  AOI22_X1 U4523 ( .A1(n4098), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4524 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4068), .B1(n4050), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4525 ( .A1(n3970), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3475) );
  INV_X2 U4526 ( .A(n3473), .ZN(n3971) );
  AOI22_X1 U4527 ( .A1(n3971), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3474) );
  NAND4_X1 U4528 ( .A1(n3477), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3483)
         );
  AOI22_X1 U4529 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n3344), .B1(n3903), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3481) );
  INV_X1 U4530 ( .A(n4073), .ZN(n3910) );
  INV_X2 U4531 ( .A(n3910), .ZN(n4092) );
  AOI22_X1 U4532 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4092), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4533 ( .A1(n4074), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4534 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n4049), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3478) );
  NAND4_X1 U4535 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(n3482)
         );
  AOI22_X1 U4536 ( .A1(n3484), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4537 ( .A1(n4049), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4073), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4538 ( .A1(n4068), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4539 ( .A1(n3971), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3485) );
  NAND4_X1 U4540 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3494)
         );
  AOI22_X1 U4541 ( .A1(n3970), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4542 ( .A1(n3884), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4543 ( .A1(n4090), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4544 ( .A1(n3903), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3489) );
  NAND4_X1 U4545 ( .A1(n3492), .A2(n3491), .A3(n3490), .A4(n3489), .ZN(n3493)
         );
  NAND2_X1 U4546 ( .A1(n3496), .A2(n7027), .ZN(n3611) );
  NAND2_X1 U4547 ( .A1(n3612), .A2(n3611), .ZN(n3500) );
  INV_X1 U4548 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3499) );
  AOI21_X1 U4549 ( .B1(n4748), .B2(n4355), .A(n7027), .ZN(n3498) );
  OAI211_X1 U4550 ( .C1(n4157), .C2(n3499), .A(n3498), .B(n3501), .ZN(n3614)
         );
  NAND2_X1 U4551 ( .A1(n3500), .A2(n3614), .ZN(n3502) );
  NAND2_X1 U4552 ( .A1(n3504), .A2(n3503), .ZN(n3507) );
  NAND2_X2 U4553 ( .A1(n4748), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3542) );
  INV_X1 U4554 ( .A(n3542), .ZN(n3505) );
  NAND2_X1 U4555 ( .A1(n3505), .A2(n4348), .ZN(n3506) );
  AND2_X1 U4556 ( .A1(n3594), .A2(n3593), .ZN(n3509) );
  INV_X1 U4557 ( .A(n3587), .ZN(n3531) );
  NAND2_X1 U4558 ( .A1(n4714), .A2(n3510), .ZN(n3512) );
  NAND2_X1 U4559 ( .A1(n3512), .A2(n3511), .ZN(n3534) );
  NAND2_X1 U4561 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3514) );
  XNOR2_X1 U4562 ( .A(n6827), .B(n3514), .ZN(n4860) );
  OAI22_X1 U4563 ( .A1(n4860), .A2(n4530), .B1(n4171), .B2(n6827), .ZN(n3515)
         );
  XNOR2_X1 U4564 ( .A(n3534), .B(n3532), .ZN(n4713) );
  NAND2_X1 U4565 ( .A1(n4713), .A2(n7027), .ZN(n3530) );
  INV_X1 U4566 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4567 ( .A1(n4098), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4568 ( .A1(n4068), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4569 ( .A1(n3970), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4570 ( .A1(n4099), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4571 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3525)
         );
  AOI22_X1 U4572 ( .A1(n3884), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4573 ( .A1(n4073), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4574 ( .A1(n4074), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4575 ( .A1(n4100), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4576 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  OAI22_X1 U4577 ( .A1(n4157), .A2(n3526), .B1(n3542), .B2(n4342), .ZN(n3528)
         );
  NOR2_X1 U4578 ( .A1(n4342), .A2(n3541), .ZN(n3527) );
  XNOR2_X1 U4579 ( .A(n3528), .B(n3527), .ZN(n3529) );
  INV_X1 U4580 ( .A(n3532), .ZN(n3533) );
  NAND2_X1 U4581 ( .A1(n3535), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3540) );
  AND3_X1 U4582 ( .A1(n6462), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U4583 ( .A1(n6550), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U4584 ( .A1(n6569), .A2(n6462), .ZN(n3536) );
  AND2_X1 U4585 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U4586 ( .A1(n4908), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U4587 ( .A1(n5075), .A2(n3538), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3537), .ZN(n3539) );
  AOI22_X1 U4588 ( .A1(n4098), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4589 ( .A1(n4068), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4590 ( .A1(n3970), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4591 ( .A1(n3971), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4592 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3553)
         );
  AOI22_X1 U4593 ( .A1(n3884), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4594 ( .A1(n4092), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4595 ( .A1(n4074), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4596 ( .A1(n4049), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4597 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3552)
         );
  AOI22_X1 U4598 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n4128), .B1(n4164), 
        .B2(n4336), .ZN(n3554) );
  AOI22_X1 U4599 ( .A1(n4098), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4600 ( .A1(n4068), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4601 ( .A1(n3970), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4602 ( .A1(n3971), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4603 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3565)
         );
  AOI22_X1 U4604 ( .A1(n3884), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4605 ( .A1(n4092), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4606 ( .A1(n4074), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4607 ( .A1(n4049), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4608 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3564)
         );
  NAND2_X1 U4609 ( .A1(n4164), .A2(n4370), .ZN(n3567) );
  NAND2_X1 U4610 ( .A1(n4128), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3566) );
  NAND2_X1 U4611 ( .A1(n3152), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3597) );
  NOR2_X2 U4612 ( .A1(n4842), .A2(n6592), .ZN(n3571) );
  INV_X1 U4613 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6297) );
  INV_X1 U4614 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6864) );
  OAI22_X1 U4615 ( .A1(n4082), .A2(n6297), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6864), .ZN(n3572) );
  INV_X1 U4616 ( .A(n3572), .ZN(n3573) );
  OAI21_X1 U4617 ( .B1(n3597), .B2(n4598), .A(n3573), .ZN(n3576) );
  INV_X1 U4618 ( .A(n3637), .ZN(n3638) );
  INV_X1 U4619 ( .A(n3574), .ZN(n3580) );
  NAND2_X1 U4620 ( .A1(n6864), .A2(n3580), .ZN(n3575) );
  NAND2_X1 U4621 ( .A1(n3638), .A2(n3575), .ZN(n6257) );
  MUX2_X1 U4622 ( .A(n3576), .B(n6257), .S(n4023), .Z(n3577) );
  INV_X1 U4623 ( .A(n4702), .ZN(n3586) );
  INV_X1 U4624 ( .A(n3589), .ZN(n3581) );
  OAI21_X1 U4625 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3581), .A(n3580), 
        .ZN(n5624) );
  AOI22_X1 U4626 ( .A1(n4023), .A2(n5624), .B1(n5370), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3583) );
  NAND2_X1 U4627 ( .A1(n3571), .A2(EAX_REG_3__SCAN_IN), .ZN(n3582) );
  OAI211_X1 U4628 ( .C1(n3597), .C2(n4804), .A(n3583), .B(n3582), .ZN(n3584)
         );
  AOI21_X1 U4629 ( .B1(n4813), .B2(n3800), .A(n3584), .ZN(n4693) );
  INV_X1 U4630 ( .A(n4693), .ZN(n3585) );
  NAND2_X1 U4631 ( .A1(n3586), .A2(n3585), .ZN(n3620) );
  NAND2_X1 U4632 ( .A1(n4340), .A2(n3800), .ZN(n3588) );
  OAI21_X1 U4633 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3589), .ZN(n6369) );
  AOI22_X1 U4634 ( .A1(n5370), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4023), 
        .B2(n6369), .ZN(n3591) );
  NAND2_X1 U4635 ( .A1(n3571), .A2(EAX_REG_2__SCAN_IN), .ZN(n3590) );
  OAI211_X1 U4636 ( .C1(n3597), .C2(n5334), .A(n3591), .B(n3590), .ZN(n3618)
         );
  BUF_X1 U4637 ( .A(n3592), .Z(n3596) );
  XNOR2_X1 U4638 ( .A(n3594), .B(n3593), .ZN(n3595) );
  NAND2_X1 U4639 ( .A1(n4725), .A2(n3800), .ZN(n3600) );
  INV_X1 U4640 ( .A(n3597), .ZN(n3608) );
  INV_X1 U4641 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4648) );
  INV_X1 U4642 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4833) );
  OAI22_X1 U4643 ( .A1(n4082), .A2(n4648), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4833), .ZN(n3598) );
  AOI21_X1 U4644 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3608), .A(n3598), 
        .ZN(n3599) );
  NAND2_X1 U4645 ( .A1(n3600), .A2(n3599), .ZN(n4610) );
  INV_X1 U4646 ( .A(n3601), .ZN(n3604) );
  INV_X1 U4647 ( .A(n3602), .ZN(n3603) );
  NAND2_X1 U4648 ( .A1(n3604), .A2(n3603), .ZN(n3606) );
  NAND2_X1 U4649 ( .A1(n3606), .A2(n3605), .ZN(n6496) );
  OR2_X1 U4650 ( .A1(n6496), .A2(n3784), .ZN(n3610) );
  INV_X1 U4651 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4854) );
  INV_X1 U4652 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5643) );
  OAI22_X1 U4653 ( .A1(n4082), .A2(n4854), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5643), .ZN(n3607) );
  AOI21_X1 U4654 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3608), .A(n3607), 
        .ZN(n3609) );
  NAND2_X1 U4655 ( .A1(n3610), .A2(n3609), .ZN(n4627) );
  NAND2_X1 U4656 ( .A1(n3614), .A2(n3611), .ZN(n3615) );
  INV_X1 U4657 ( .A(n3612), .ZN(n3613) );
  INV_X1 U4658 ( .A(n3809), .ZN(n3616) );
  AOI21_X1 U4659 ( .B1(n6473), .B2(n3616), .A(n6592), .ZN(n4626) );
  NAND2_X1 U4660 ( .A1(n4627), .A2(n4626), .ZN(n4628) );
  OAI21_X1 U4661 ( .B1(n4627), .B2(n3641), .A(n4628), .ZN(n4609) );
  NAND2_X1 U4662 ( .A1(n4610), .A2(n4609), .ZN(n4608) );
  NAND2_X1 U4663 ( .A1(n3617), .A2(n4608), .ZN(n3619) );
  NAND2_X1 U4664 ( .A1(n3619), .A2(n4679), .ZN(n4677) );
  AOI22_X1 U4665 ( .A1(n4098), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4666 ( .A1(n4068), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4667 ( .A1(n3970), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4668 ( .A1(n3971), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4669 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3630)
         );
  AOI22_X1 U4670 ( .A1(n3884), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4671 ( .A1(n4092), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4672 ( .A1(n4074), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4673 ( .A1(n4049), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4674 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3629)
         );
  NAND2_X1 U4675 ( .A1(n4164), .A2(n4373), .ZN(n3632) );
  NAND2_X1 U4676 ( .A1(n4128), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3631) );
  NAND2_X1 U4677 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  NAND2_X1 U4678 ( .A1(n3659), .A2(n3636), .ZN(n4377) );
  INV_X1 U4679 ( .A(n3661), .ZN(n3640) );
  INV_X1 U4680 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U4681 ( .A1(n3638), .A2(n6357), .ZN(n3639) );
  NAND2_X1 U4682 ( .A1(n3640), .A2(n3639), .ZN(n6349) );
  AOI22_X1 U4683 ( .A1(n6349), .A2(n4183), .B1(n5370), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3643) );
  NAND2_X1 U4684 ( .A1(n3571), .A2(EAX_REG_5__SCAN_IN), .ZN(n3642) );
  OAI211_X1 U4685 ( .C1(n4377), .C2(n3784), .A(n3643), .B(n3642), .ZN(n4822)
         );
  NAND2_X1 U4686 ( .A1(n4703), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U4687 ( .A1(n4128), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4688 ( .A1(n4098), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4689 ( .A1(n4068), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4690 ( .A1(n3970), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4691 ( .A1(n3971), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3645) );
  NAND4_X1 U4692 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(n3654)
         );
  AOI22_X1 U4693 ( .A1(n3884), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4694 ( .A1(n4092), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4695 ( .A1(n4074), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3650) );
  INV_X1 U4696 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6922) );
  AOI22_X1 U4697 ( .A1(n4049), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4698 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3653)
         );
  NAND2_X1 U4699 ( .A1(n4164), .A2(n4391), .ZN(n3655) );
  INV_X1 U4700 ( .A(n3657), .ZN(n3658) );
  NAND2_X1 U4701 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  NAND2_X1 U4702 ( .A1(n4381), .A2(n3800), .ZN(n3665) );
  INV_X1 U4703 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4650) );
  OAI21_X1 U4704 ( .B1(n3661), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3668), 
        .ZN(n5599) );
  AOI22_X1 U4705 ( .A1(n5599), .A2(n4183), .B1(n5370), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3662) );
  OAI21_X1 U4706 ( .B1(n4082), .B2(n4650), .A(n3662), .ZN(n3663) );
  INV_X1 U4707 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U4708 ( .A1(n4164), .A2(n4399), .ZN(n3666) );
  OAI21_X1 U4709 ( .B1(n4157), .B2(n6802), .A(n3666), .ZN(n3667) );
  INV_X1 U4710 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4711 ( .A1(n3668), .A2(n6347), .ZN(n3669) );
  NAND2_X1 U4712 ( .A1(n3669), .A2(n3128), .ZN(n6341) );
  NOR2_X1 U4713 ( .A1(n3967), .A2(n6347), .ZN(n3670) );
  AOI21_X1 U4714 ( .B1(n6341), .B2(n4183), .A(n3670), .ZN(n3671) );
  OAI21_X1 U4715 ( .B1(n4082), .B2(n3672), .A(n3671), .ZN(n3673) );
  AOI22_X1 U4716 ( .A1(n4068), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4717 ( .A1(n3884), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4718 ( .A1(n4092), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4719 ( .A1(n4050), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3674) );
  NAND4_X1 U4720 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3683)
         );
  AOI22_X1 U4721 ( .A1(n4098), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4722 ( .A1(n3970), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4723 ( .A1(n4049), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4724 ( .A1(n4090), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4725 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3682)
         );
  NOR2_X1 U4726 ( .A1(n3683), .A2(n3682), .ZN(n3687) );
  NAND2_X1 U4727 ( .A1(n3571), .A2(EAX_REG_8__SCAN_IN), .ZN(n3686) );
  XNOR2_X1 U4728 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3128), .ZN(n6221) );
  INV_X1 U4729 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5310) );
  OAI22_X1 U4730 ( .A1(n6221), .A2(n3641), .B1(n3967), .B2(n5310), .ZN(n3684)
         );
  INV_X1 U4731 ( .A(n3684), .ZN(n3685) );
  OAI211_X1 U4732 ( .C1(n3687), .C2(n3784), .A(n3686), .B(n3685), .ZN(n5229)
         );
  AOI21_X1 U4733 ( .B1(n6981), .B2(n3688), .A(n3719), .ZN(n6212) );
  OR2_X1 U4734 ( .A1(n6212), .A2(n3641), .ZN(n3703) );
  AOI22_X1 U4735 ( .A1(n4090), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4736 ( .A1(n4068), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4737 ( .A1(n3884), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4738 ( .A1(n3970), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4739 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3698)
         );
  AOI22_X1 U4740 ( .A1(n4092), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4741 ( .A1(n4098), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4742 ( .A1(n3547), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4743 ( .A1(n4049), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4744 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3697)
         );
  NOR2_X1 U4745 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  OAI22_X1 U4746 ( .A1(n3784), .A2(n3699), .B1(n3967), .B2(n6981), .ZN(n3701)
         );
  INV_X1 U4747 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5253) );
  NOR2_X1 U4748 ( .A1(n4082), .A2(n5253), .ZN(n3700) );
  NOR2_X1 U4749 ( .A1(n3701), .A2(n3700), .ZN(n3702) );
  NAND2_X1 U4750 ( .A1(n3703), .A2(n3702), .ZN(n5247) );
  XNOR2_X1 U4751 ( .A(n3719), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5904)
         );
  AOI22_X1 U4752 ( .A1(n4050), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4753 ( .A1(n3884), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4754 ( .A1(n4092), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4755 ( .A1(n4090), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4756 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3713)
         );
  AOI22_X1 U4757 ( .A1(n4098), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4758 ( .A1(n3970), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4759 ( .A1(n4049), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4760 ( .A1(n4068), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4761 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3712)
         );
  OAI21_X1 U4762 ( .B1(n3713), .B2(n3712), .A(n3800), .ZN(n3716) );
  NAND2_X1 U4763 ( .A1(n3571), .A2(EAX_REG_10__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4764 ( .A1(n5370), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3714)
         );
  NAND3_X1 U4765 ( .A1(n3716), .A2(n3715), .A3(n3714), .ZN(n3717) );
  AOI21_X1 U4766 ( .B1(n5904), .B2(n4183), .A(n3717), .ZN(n5585) );
  AOI21_X1 U4767 ( .B1(n6951), .B2(n3720), .A(n3753), .ZN(n6332) );
  OR2_X1 U4768 ( .A1(n6332), .A2(n3641), .ZN(n3735) );
  AOI22_X1 U4769 ( .A1(n3970), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4770 ( .A1(n4050), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4771 ( .A1(n4092), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4772 ( .A1(n4049), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4773 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3730)
         );
  AOI22_X1 U4774 ( .A1(n4098), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4775 ( .A1(n3884), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4776 ( .A1(n3971), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4777 ( .A1(n4068), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4778 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  NOR2_X1 U4779 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  OAI22_X1 U4780 ( .A1(n3784), .A2(n3731), .B1(n3967), .B2(n6951), .ZN(n3733)
         );
  INV_X1 U4781 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5745) );
  NOR2_X1 U4782 ( .A1(n4082), .A2(n5745), .ZN(n3732) );
  NOR2_X1 U4783 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  INV_X1 U4784 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3736) );
  XNOR2_X1 U4785 ( .A(n3753), .B(n3736), .ZN(n6198) );
  NAND2_X1 U4786 ( .A1(n6198), .A2(n4183), .ZN(n3740) );
  INV_X1 U4787 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5742) );
  AOI21_X1 U4788 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3736), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3737) );
  INV_X1 U4789 ( .A(n3737), .ZN(n3738) );
  OAI21_X1 U4790 ( .B1(n4082), .B2(n5742), .A(n3738), .ZN(n3739) );
  NAND2_X1 U4791 ( .A1(n3740), .A2(n3739), .ZN(n3752) );
  AOI22_X1 U4792 ( .A1(n4098), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4793 ( .A1(n3547), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4794 ( .A1(n4044), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4795 ( .A1(n4074), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4796 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3750)
         );
  AOI22_X1 U4797 ( .A1(n4068), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4798 ( .A1(n3884), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4073), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4799 ( .A1(n3970), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4800 ( .A1(n4049), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4801 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  OAI21_X1 U4802 ( .B1(n3750), .B2(n3749), .A(n3800), .ZN(n3751) );
  INV_X1 U4803 ( .A(n3754), .ZN(n3755) );
  INV_X1 U4804 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U4805 ( .A1(n3755), .A2(n6192), .ZN(n3756) );
  NAND2_X1 U4806 ( .A1(n3808), .A2(n3756), .ZN(n6187) );
  INV_X1 U4807 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5741) );
  OAI22_X1 U4808 ( .A1(n4082), .A2(n5741), .B1(n3967), .B2(n6192), .ZN(n3757)
         );
  AOI21_X1 U4809 ( .B1(n6187), .B2(n4183), .A(n3757), .ZN(n3758) );
  AOI22_X1 U4810 ( .A1(n4050), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4811 ( .A1(n4068), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4049), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4812 ( .A1(n4092), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4813 ( .A1(n3970), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4814 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4815 ( .A1(n4090), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4816 ( .A1(n3884), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4817 ( .A1(n4098), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4818 ( .A1(n4030), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4819 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  OR2_X1 U4820 ( .A1(n3769), .A2(n3768), .ZN(n3770) );
  NAND2_X1 U4821 ( .A1(n3800), .A2(n3770), .ZN(n5675) );
  INV_X1 U4822 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3789) );
  XNOR2_X1 U4823 ( .A(n3808), .B(n3789), .ZN(n5879) );
  NAND2_X1 U4824 ( .A1(n5879), .A2(n4183), .ZN(n3788) );
  AOI22_X1 U4825 ( .A1(n4098), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4826 ( .A1(n4092), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4827 ( .A1(n3970), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4828 ( .A1(n4074), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4829 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3782)
         );
  AOI22_X1 U4830 ( .A1(n4068), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4831 ( .A1(n3884), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4832 ( .A1(n4090), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4833 ( .A1(n4049), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4834 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  NOR2_X1 U4835 ( .A1(n3782), .A2(n3781), .ZN(n3783) );
  OAI22_X1 U4836 ( .A1(n3784), .A2(n3783), .B1(n3967), .B2(n3789), .ZN(n3786)
         );
  INV_X1 U4837 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5738) );
  NOR2_X1 U4838 ( .A1(n4082), .A2(n5738), .ZN(n3785) );
  NOR2_X1 U4839 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  NAND2_X1 U4840 ( .A1(n3788), .A2(n3787), .ZN(n5569) );
  OR2_X1 U4841 ( .A1(n3808), .A2(n3789), .ZN(n3791) );
  INV_X1 U4842 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3790) );
  XNOR2_X1 U4843 ( .A(n3791), .B(n3790), .ZN(n5867) );
  AOI22_X1 U4844 ( .A1(n3884), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4845 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n4044), .B1(n4025), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4846 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n3547), .B1(n4030), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4847 ( .A1(n4068), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4848 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3802)
         );
  AOI22_X1 U4849 ( .A1(n4098), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4850 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4049), .B1(n4073), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4851 ( .A1(n4050), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4852 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3970), .B1(n3971), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4853 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3801)
         );
  OAI21_X1 U4854 ( .B1(n3802), .B2(n3801), .A(n3800), .ZN(n3805) );
  NAND2_X1 U4855 ( .A1(n3571), .A2(EAX_REG_15__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4856 ( .A1(n5370), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3803)
         );
  NAND3_X1 U4857 ( .A1(n3805), .A2(n3804), .A3(n3803), .ZN(n3806) );
  AOI21_X1 U4858 ( .B1(n5867), .B2(n4183), .A(n3806), .ZN(n5557) );
  NAND2_X1 U4859 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3807) );
  INV_X1 U4860 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5547) );
  XNOR2_X1 U4861 ( .A(n3826), .B(n5547), .ZN(n5862) );
  NAND2_X1 U4862 ( .A1(n5862), .A2(n4183), .ZN(n3825) );
  NAND2_X1 U4863 ( .A1(n3810), .A2(n4489), .ZN(n3811) );
  AOI22_X1 U4864 ( .A1(n4068), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4865 ( .A1(n3884), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4866 ( .A1(n4092), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4867 ( .A1(n4074), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4868 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3821)
         );
  AOI22_X1 U4869 ( .A1(n4098), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3970), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4870 ( .A1(n4050), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4871 ( .A1(n3971), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4872 ( .A1(n4049), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4873 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  OR2_X1 U4874 ( .A1(n3821), .A2(n3820), .ZN(n3823) );
  INV_X1 U4875 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4645) );
  OAI22_X1 U4876 ( .A1(n4082), .A2(n4645), .B1(n3967), .B2(n5547), .ZN(n3822)
         );
  AOI21_X1 U4877 ( .B1(n4084), .B2(n3823), .A(n3822), .ZN(n3824) );
  NAND2_X1 U4878 ( .A1(n3825), .A2(n3824), .ZN(n5539) );
  XNOR2_X1 U4879 ( .A(n3845), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5855)
         );
  NAND2_X1 U4880 ( .A1(n5855), .A2(n4183), .ZN(n3844) );
  AOI22_X1 U4881 ( .A1(n4049), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4882 ( .A1(n3970), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4883 ( .A1(n4092), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4884 ( .A1(n4025), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4885 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3839)
         );
  NAND2_X1 U4886 ( .A1(n4091), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3833)
         );
  NAND2_X1 U4887 ( .A1(n4044), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3832) );
  AND3_X1 U4888 ( .A1(n3833), .A2(n3832), .A3(n3641), .ZN(n3837) );
  AOI22_X1 U4889 ( .A1(n4068), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4890 ( .A1(n4098), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4891 ( .A1(n4050), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4892 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  NAND2_X1 U4893 ( .A1(n4110), .A2(n3641), .ZN(n3898) );
  OAI21_X1 U4894 ( .B1(n3839), .B2(n3838), .A(n3898), .ZN(n3842) );
  NAND2_X1 U4895 ( .A1(n3571), .A2(EAX_REG_17__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4896 ( .A1(n6592), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3840)
         );
  NAND3_X1 U4897 ( .A1(n3842), .A2(n3841), .A3(n3840), .ZN(n3843) );
  NAND2_X1 U4898 ( .A1(n3844), .A2(n3843), .ZN(n5526) );
  NAND2_X1 U4899 ( .A1(n3846), .A2(n5517), .ZN(n3847) );
  NAND2_X1 U4900 ( .A1(n3863), .A2(n3847), .ZN(n5848) );
  AOI22_X1 U4901 ( .A1(n4050), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4902 ( .A1(n3884), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4903 ( .A1(n4090), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4904 ( .A1(n4049), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4905 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AOI22_X1 U4906 ( .A1(n4098), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4907 ( .A1(n4092), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4908 ( .A1(n3970), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4909 ( .A1(n4068), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4910 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  NOR2_X1 U4911 ( .A1(n3857), .A2(n3856), .ZN(n3860) );
  INV_X1 U4912 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6906) );
  OAI22_X1 U4913 ( .A1(n4082), .A2(n6906), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5517), .ZN(n3858) );
  INV_X1 U4914 ( .A(n3858), .ZN(n3859) );
  OAI21_X1 U4915 ( .B1(n4110), .B2(n3860), .A(n3859), .ZN(n3861) );
  MUX2_X1 U4916 ( .A(n5848), .B(n3861), .S(n3641), .Z(n5513) );
  INV_X1 U4917 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U4918 ( .A1(n3863), .A2(n6967), .ZN(n3864) );
  NAND2_X1 U4919 ( .A1(n3894), .A2(n3864), .ZN(n5836) );
  AOI22_X1 U4920 ( .A1(n4049), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4921 ( .A1(n4068), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4922 ( .A1(n4098), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4923 ( .A1(n4044), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4924 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3876)
         );
  INV_X1 U4925 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3869) );
  NOR2_X1 U4926 ( .A1(n3462), .A2(n3869), .ZN(n3870) );
  AOI211_X1 U4927 ( .C1(n4097), .C2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n4183), 
        .B(n3870), .ZN(n3874) );
  AOI22_X1 U4928 ( .A1(n4074), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4929 ( .A1(n4050), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3884), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4930 ( .A1(n4092), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4931 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3875)
         );
  OAI21_X1 U4932 ( .B1(n3876), .B2(n3875), .A(n3898), .ZN(n3878) );
  NAND2_X1 U4933 ( .A1(n3571), .A2(EAX_REG_19__SCAN_IN), .ZN(n3877) );
  OAI211_X1 U4934 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6967), .A(n3878), .B(
        n3877), .ZN(n3879) );
  OAI21_X1 U4935 ( .B1(n5836), .B2(n3641), .A(n3879), .ZN(n5496) );
  AOI22_X1 U4936 ( .A1(n4050), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4937 ( .A1(n4044), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4938 ( .A1(n4091), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4939 ( .A1(n4049), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4940 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3890)
         );
  AOI22_X1 U4941 ( .A1(n4098), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4942 ( .A1(n3884), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4092), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4943 ( .A1(n4074), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4944 ( .A1(n3970), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4945 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3889)
         );
  OAI21_X1 U4946 ( .B1(n3890), .B2(n3889), .A(n4084), .ZN(n3892) );
  AOI22_X1 U4947 ( .A1(n3571), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6592), .ZN(n3891) );
  NAND2_X1 U4948 ( .A1(n3892), .A2(n3891), .ZN(n3896) );
  NAND2_X1 U4949 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  NAND2_X1 U4950 ( .A1(n3897), .A2(n3895), .ZN(n5826) );
  MUX2_X1 U4951 ( .A(n3896), .B(n5826), .S(n4023), .Z(n5485) );
  XNOR2_X1 U4952 ( .A(n3935), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5816)
         );
  INV_X1 U4953 ( .A(n3898), .ZN(n3919) );
  AOI22_X1 U4954 ( .A1(n4049), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4955 ( .A1(n4068), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4956 ( .A1(n4050), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4957 ( .A1(n4044), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4958 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3916)
         );
  INV_X1 U4959 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3906) );
  INV_X1 U4960 ( .A(n3903), .ZN(n3905) );
  INV_X1 U4961 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3904) );
  OAI22_X1 U4962 ( .A1(n3455), .A2(n3906), .B1(n3905), .B2(n3904), .ZN(n3915)
         );
  INV_X1 U4963 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4964 ( .A1(n3884), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3908) );
  AOI21_X1 U4965 ( .B1(n4097), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n4183), 
        .ZN(n3907) );
  OAI211_X1 U4966 ( .C1(n3910), .C2(n3909), .A(n3908), .B(n3907), .ZN(n3914)
         );
  INV_X1 U4967 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3912) );
  INV_X1 U4968 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3911) );
  OAI22_X1 U4969 ( .A1(n3361), .A2(n3912), .B1(n3473), .B2(n3911), .ZN(n3913)
         );
  NOR4_X1 U4970 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3918)
         );
  AOI22_X1 U4971 ( .A1(n3571), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6592), .ZN(n3917) );
  OAI21_X1 U4972 ( .B1(n3919), .B2(n3918), .A(n3917), .ZN(n3920) );
  AOI22_X1 U4973 ( .A1(n3970), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4974 ( .A1(n4068), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4975 ( .A1(n4100), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4976 ( .A1(n3884), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4977 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3931)
         );
  AOI22_X1 U4978 ( .A1(n4098), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4979 ( .A1(n4092), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4980 ( .A1(n3971), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4981 ( .A1(n4030), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4982 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NOR2_X1 U4983 ( .A1(n3931), .A2(n3930), .ZN(n3934) );
  INV_X1 U4984 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7014) );
  OAI22_X1 U4985 ( .A1(n4082), .A2(n7014), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5462), .ZN(n3932) );
  INV_X1 U4986 ( .A(n3932), .ZN(n3933) );
  OAI21_X1 U4987 ( .B1(n4110), .B2(n3934), .A(n3933), .ZN(n3938) );
  NAND2_X1 U4988 ( .A1(n3936), .A2(n5462), .ZN(n3937) );
  NAND2_X1 U4989 ( .A1(n3939), .A2(n3937), .ZN(n5457) );
  MUX2_X1 U4990 ( .A(n3938), .B(n5457), .S(n4023), .Z(n4528) );
  XNOR2_X1 U4991 ( .A(n3964), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5808)
         );
  AOI22_X1 U4992 ( .A1(n4098), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4993 ( .A1(n4068), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3942) );
  INV_X1 U4994 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U4995 ( .A1(n3970), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4996 ( .A1(n3971), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4997 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3949)
         );
  AOI22_X1 U4998 ( .A1(n3884), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4999 ( .A1(n4073), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U5000 ( .A1(n4074), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U5001 ( .A1(n4049), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U5002 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  NOR2_X1 U5003 ( .A1(n3949), .A2(n3948), .ZN(n3969) );
  AOI22_X1 U5004 ( .A1(n4098), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U5005 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n4068), .B1(n4050), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U5006 ( .A1(n3970), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U5007 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3971), .B1(n4025), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U5008 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3959)
         );
  AOI22_X1 U5009 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n3884), .B1(n3547), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U5010 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4092), .B1(n4091), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U5011 ( .A1(n4074), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U5012 ( .A1(n4049), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U5013 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3958)
         );
  NOR2_X1 U5014 ( .A1(n3959), .A2(n3958), .ZN(n3968) );
  XNOR2_X1 U5015 ( .A(n3969), .B(n3968), .ZN(n3962) );
  NAND2_X1 U5016 ( .A1(n3571), .A2(EAX_REG_23__SCAN_IN), .ZN(n3961) );
  OAI21_X1 U5017 ( .B1(n6467), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6592), 
        .ZN(n3960) );
  OAI211_X1 U5018 ( .C1(n4110), .C2(n3962), .A(n3961), .B(n3960), .ZN(n3963)
         );
  NAND2_X1 U5019 ( .A1(n3965), .A2(n7044), .ZN(n3966) );
  AND2_X1 U5020 ( .A1(n4018), .A2(n3966), .ZN(n5802) );
  NOR2_X1 U5021 ( .A1(n3967), .A2(n7044), .ZN(n3984) );
  NOR2_X1 U5022 ( .A1(n3969), .A2(n3968), .ZN(n3996) );
  AOI22_X1 U5023 ( .A1(n4098), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5024 ( .A1(n4068), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5025 ( .A1(n3970), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5026 ( .A1(n3971), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U5027 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U5028 ( .A1(n3884), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U5029 ( .A1(n4092), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5030 ( .A1(n4074), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5031 ( .A1(n4049), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U5032 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  NOR2_X1 U5033 ( .A1(n3996), .A2(n3997), .ZN(n3982) );
  AOI211_X1 U5034 ( .C1(n3996), .C2(n3997), .A(n3982), .B(n4110), .ZN(n3983)
         );
  AOI211_X1 U5035 ( .C1(n3571), .C2(EAX_REG_24__SCAN_IN), .A(n3984), .B(n3983), 
        .ZN(n3985) );
  AOI22_X1 U5036 ( .A1(n4098), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U5037 ( .A1(n4068), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U5038 ( .A1(n3970), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U5039 ( .A1(n4099), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U5040 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3995)
         );
  AOI22_X1 U5041 ( .A1(n3884), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5042 ( .A1(n4073), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U5043 ( .A1(n4074), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5044 ( .A1(n4049), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U5045 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  OR2_X1 U5046 ( .A1(n3995), .A2(n3994), .ZN(n4012) );
  XOR2_X1 U5047 ( .A(n4012), .B(n4013), .Z(n4000) );
  INV_X1 U5048 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3998) );
  OAI22_X1 U5049 ( .A1(n4082), .A2(n3998), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3193), .ZN(n3999) );
  AOI21_X1 U5050 ( .B1(n4084), .B2(n4000), .A(n3999), .ZN(n4001) );
  XNOR2_X1 U5051 ( .A(n4018), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5790)
         );
  MUX2_X1 U5052 ( .A(n4001), .B(n5790), .S(n4023), .Z(n5423) );
  AOI22_X1 U5053 ( .A1(n4098), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4068), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U5054 ( .A1(n3884), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5055 ( .A1(n4044), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5056 ( .A1(n4049), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3925), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U5057 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4011)
         );
  AOI22_X1 U5058 ( .A1(n4050), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4090), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5059 ( .A1(n4073), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5060 ( .A1(n3970), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5061 ( .A1(n4074), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U5062 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  NOR2_X1 U5063 ( .A1(n4011), .A2(n4010), .ZN(n4038) );
  NAND2_X1 U5064 ( .A1(n4013), .A2(n4012), .ZN(n4037) );
  XNOR2_X1 U5065 ( .A(n4038), .B(n4037), .ZN(n4017) );
  INV_X1 U5066 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4014) );
  OAI22_X1 U5067 ( .A1(n4082), .A2(n4014), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4020), .ZN(n4015) );
  INV_X1 U5068 ( .A(n4015), .ZN(n4016) );
  OAI21_X1 U5069 ( .B1(n4017), .B2(n4110), .A(n4016), .ZN(n4024) );
  NAND2_X1 U5070 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  NAND2_X1 U5071 ( .A1(n4042), .A2(n4022), .ZN(n5777) );
  MUX2_X1 U5072 ( .A(n4024), .B(n5777), .S(n4023), .Z(n5415) );
  AOI22_X1 U5073 ( .A1(n4098), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5074 ( .A1(n4068), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4050), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5075 ( .A1(n3970), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5076 ( .A1(n3971), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4025), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U5077 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4036)
         );
  AOI22_X1 U5078 ( .A1(n3884), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3547), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5079 ( .A1(n4073), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5080 ( .A1(n4074), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5081 ( .A1(n4049), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4030), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U5082 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4035)
         );
  OR2_X1 U5083 ( .A1(n4036), .A2(n4035), .ZN(n4057) );
  NOR2_X1 U5084 ( .A1(n4038), .A2(n4037), .ZN(n4058) );
  XOR2_X1 U5085 ( .A(n4057), .B(n4058), .Z(n4041) );
  INV_X1 U5086 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4039) );
  INV_X1 U5087 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5773) );
  OAI22_X1 U5088 ( .A1(n4082), .A2(n4039), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5773), .ZN(n4040) );
  AOI21_X1 U5089 ( .B1(n4041), .B2(n4084), .A(n4040), .ZN(n4043) );
  XOR2_X1 U5090 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n4061), .Z(n5771) );
  MUX2_X1 U5091 ( .A(n4043), .B(n5771), .S(n4183), .Z(n5405) );
  AOI22_X1 U5092 ( .A1(n4090), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5093 ( .A1(n4068), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4074), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5094 ( .A1(n3971), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5095 ( .A1(n3884), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5096 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4056)
         );
  AOI22_X1 U5097 ( .A1(n4098), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5098 ( .A1(n4050), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4049), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5099 ( .A1(n4073), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U5100 ( .A1(n3903), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U5101 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4055)
         );
  NOR2_X1 U5102 ( .A1(n4056), .A2(n4055), .ZN(n4066) );
  NAND2_X1 U5103 ( .A1(n4058), .A2(n4057), .ZN(n4065) );
  XNOR2_X1 U5104 ( .A(n4066), .B(n4065), .ZN(n4060) );
  AOI22_X1 U5105 ( .A1(n3571), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6592), .ZN(n4059) );
  OAI21_X1 U5106 ( .B1(n4060), .B2(n4110), .A(n4059), .ZN(n4064) );
  NAND2_X1 U5107 ( .A1(n4062), .A2(n5349), .ZN(n4063) );
  NAND2_X1 U5108 ( .A1(n4086), .A2(n4063), .ZN(n5354) );
  MUX2_X1 U5109 ( .A(n4064), .B(n5354), .S(n4183), .Z(n5343) );
  NOR2_X1 U5110 ( .A1(n4066), .A2(n4065), .ZN(n4089) );
  AOI22_X1 U5111 ( .A1(n4098), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4067), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5112 ( .A1(n4068), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5113 ( .A1(n4097), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5114 ( .A1(n4099), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U5115 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4080)
         );
  AOI22_X1 U5116 ( .A1(n3884), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5117 ( .A1(n4073), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5118 ( .A1(n4074), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5119 ( .A1(n4100), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5120 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  OR2_X1 U5121 ( .A1(n4080), .A2(n4079), .ZN(n4088) );
  XOR2_X1 U5122 ( .A(n4089), .B(n4088), .Z(n4085) );
  INV_X1 U5123 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4081) );
  INV_X1 U5124 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5765) );
  OAI22_X1 U5125 ( .A1(n4082), .A2(n4081), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5765), .ZN(n4083) );
  AOI21_X1 U5126 ( .B1(n4085), .B2(n4084), .A(n4083), .ZN(n4087) );
  XOR2_X1 U5127 ( .A(n4112), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .Z(n5763) );
  MUX2_X1 U5128 ( .A(n4087), .B(n5763), .S(n4183), .Z(n5382) );
  NAND2_X1 U5129 ( .A1(n4089), .A2(n4088), .ZN(n4108) );
  AOI22_X1 U5130 ( .A1(n4090), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4044), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5131 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n3884), .B1(n3903), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5132 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4092), .B1(n4091), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5133 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n4074), .B1(n3345), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U5134 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4106)
         );
  AOI22_X1 U5135 ( .A1(n4098), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5136 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4068), .B1(n3338), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5137 ( .A1(n4099), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5138 ( .A1(n4100), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5139 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  NOR2_X1 U5140 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  XNOR2_X1 U5141 ( .A(n4108), .B(n4107), .ZN(n4111) );
  AOI22_X1 U5142 ( .A1(n3571), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6592), .ZN(n4109) );
  OAI21_X1 U5143 ( .B1(n4111), .B2(n4110), .A(n4109), .ZN(n4113) );
  XOR2_X1 U5144 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4114), .Z(n4309) );
  MUX2_X1 U5145 ( .A(n4113), .B(n4309), .S(n4183), .Z(n5369) );
  INV_X1 U5146 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6937) );
  INV_X1 U5147 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4115) );
  NAND2_X1 U5148 ( .A1(n4164), .A2(n4602), .ZN(n4117) );
  NAND2_X1 U5149 ( .A1(n4117), .A2(n3810), .ZN(n4123) );
  INV_X1 U5150 ( .A(n4132), .ZN(n4118) );
  XNOR2_X1 U5151 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4133) );
  XNOR2_X1 U5152 ( .A(n4118), .B(n4133), .ZN(n4178) );
  AND2_X1 U5153 ( .A1(n4178), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4124) );
  XNOR2_X1 U5154 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4122) );
  AOI21_X1 U5155 ( .B1(n4173), .B2(n4122), .A(n4119), .ZN(n4121) );
  NAND2_X1 U5156 ( .A1(n4758), .A2(n3810), .ZN(n4120) );
  NAND2_X1 U5157 ( .A1(n4836), .A2(n4120), .ZN(n4139) );
  NAND2_X1 U5158 ( .A1(n4164), .A2(n4122), .ZN(n4127) );
  INV_X1 U5159 ( .A(n4123), .ZN(n4126) );
  INV_X1 U5160 ( .A(n4124), .ZN(n4125) );
  OAI22_X1 U5161 ( .A1(n4129), .A2(n4127), .B1(n4126), .B2(n4125), .ZN(n4131)
         );
  AOI21_X1 U5162 ( .B1(n4129), .B2(n4178), .A(n4167), .ZN(n4130) );
  NAND2_X1 U5163 ( .A1(n4133), .A2(n4132), .ZN(n4135) );
  NAND2_X1 U5164 ( .A1(n6461), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4134) );
  NAND2_X1 U5165 ( .A1(n4135), .A2(n4134), .ZN(n4144) );
  XNOR2_X1 U5166 ( .A(n6827), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4142)
         );
  XNOR2_X1 U5167 ( .A(n4144), .B(n4142), .ZN(n4177) );
  NAND2_X1 U5168 ( .A1(n4164), .A2(n4177), .ZN(n4138) );
  INV_X1 U5169 ( .A(n4139), .ZN(n4136) );
  OAI211_X1 U5170 ( .C1(n4177), .C2(n4157), .A(n4138), .B(n4136), .ZN(n4137)
         );
  INV_X1 U5171 ( .A(n4138), .ZN(n4140) );
  NAND2_X1 U5172 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  INV_X1 U5173 ( .A(n4142), .ZN(n4143) );
  NAND2_X1 U5174 ( .A1(n4144), .A2(n4143), .ZN(n4146) );
  NAND2_X1 U5175 ( .A1(n6827), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U5176 ( .A1(n4146), .A2(n4145), .ZN(n4153) );
  XNOR2_X1 U5177 ( .A(n4804), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4151)
         );
  XNOR2_X1 U5178 ( .A(n4153), .B(n4151), .ZN(n4179) );
  INV_X1 U5179 ( .A(n4179), .ZN(n4148) );
  NAND2_X1 U5180 ( .A1(n4157), .A2(n4148), .ZN(n4147) );
  NAND2_X1 U5181 ( .A1(n4169), .A2(n4148), .ZN(n4149) );
  NAND2_X1 U5182 ( .A1(n4150), .A2(n4149), .ZN(n4159) );
  INV_X1 U5183 ( .A(n4151), .ZN(n4152) );
  NAND2_X1 U5184 ( .A1(n4153), .A2(n4152), .ZN(n4155) );
  NAND2_X1 U5185 ( .A1(n6462), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5186 ( .A1(n4155), .A2(n4154), .ZN(n4161) );
  INV_X1 U5187 ( .A(n4176), .ZN(n4156) );
  NAND2_X1 U5188 ( .A1(n4157), .A2(n4156), .ZN(n4158) );
  NAND2_X1 U5189 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4598), .ZN(n4162) );
  NAND2_X1 U5190 ( .A1(n4164), .A2(n4175), .ZN(n4166) );
  NAND2_X1 U5191 ( .A1(n7027), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4165) );
  OAI211_X1 U5192 ( .C1(n4167), .C2(n4176), .A(n4166), .B(n4165), .ZN(n4168)
         );
  OR2_X1 U5193 ( .A1(n4173), .A2(n3095), .ZN(n4174) );
  INV_X1 U5194 ( .A(n4175), .ZN(n4181) );
  NAND4_X1 U5195 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  NAND2_X1 U5196 ( .A1(n4181), .A2(n4180), .ZN(n4572) );
  INV_X1 U5197 ( .A(n4572), .ZN(n4182) );
  NAND2_X1 U5198 ( .A1(n4573), .A2(n4182), .ZN(n4559) );
  NOR2_X4 U5199 ( .A1(n4564), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U5200 ( .A1(n4183), .A2(n4529), .ZN(n6159) );
  NAND3_X1 U5201 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), 
        .A3(n6795), .ZN(n6147) );
  NAND2_X1 U5202 ( .A1(n6159), .A2(n6147), .ZN(n4184) );
  INV_X1 U5203 ( .A(n4665), .ZN(n4448) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4479) );
  NOR2_X1 U5205 ( .A1(n3098), .A2(EBX_REG_29__SCAN_IN), .ZN(n4188) );
  AOI21_X1 U5206 ( .B1(n4448), .B2(n4479), .A(n4188), .ZN(n5384) );
  INV_X1 U5207 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4189) );
  NAND2_X1 U5208 ( .A1(n4194), .A2(n4189), .ZN(n4190) );
  OAI211_X1 U5209 ( .C1(n3098), .C2(EBX_REG_1__SCAN_IN), .A(n4190), .B(n4186), 
        .ZN(n4193) );
  OR2_X2 U5210 ( .A1(n4198), .A2(n4186), .ZN(n4284) );
  INV_X1 U5211 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U5212 ( .A1(n4199), .A2(n4191), .ZN(n4192) );
  NAND2_X1 U5213 ( .A1(n4194), .A2(EBX_REG_0__SCAN_IN), .ZN(n4197) );
  INV_X1 U5214 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U5215 ( .A1(n4186), .A2(n4195), .ZN(n4196) );
  NAND2_X1 U5216 ( .A1(n4197), .A2(n4196), .ZN(n4666) );
  INV_X1 U5217 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5218 ( .A1(n4199), .A2(n4680), .ZN(n4203) );
  NAND2_X1 U5219 ( .A1(n4186), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4200)
         );
  NAND2_X1 U5220 ( .A1(n4194), .A2(n4200), .ZN(n4201) );
  OAI21_X1 U5221 ( .B1(EBX_REG_2__SCAN_IN), .B2(n3098), .A(n4201), .ZN(n4202)
         );
  AND2_X1 U5222 ( .A1(n4203), .A2(n4202), .ZN(n4674) );
  OR2_X1 U5223 ( .A1(n4279), .A2(EBX_REG_3__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5224 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4204)
         );
  OAI211_X1 U5225 ( .C1(n3098), .C2(EBX_REG_3__SCAN_IN), .A(n4194), .B(n4204), 
        .ZN(n4205) );
  NAND2_X1 U5226 ( .A1(n4206), .A2(n4205), .ZN(n4774) );
  INV_X1 U5227 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U5228 ( .A1(n4199), .A2(n6925), .ZN(n4209) );
  INV_X1 U5229 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U5230 ( .A1(n4194), .A2(n4366), .ZN(n4207) );
  OAI211_X1 U5231 ( .C1(n3098), .C2(EBX_REG_4__SCAN_IN), .A(n4207), .B(n5383), 
        .ZN(n4208) );
  NAND2_X1 U5232 ( .A1(n4209), .A2(n4208), .ZN(n4706) );
  MUX2_X1 U5233 ( .A(n4279), .B(n5383), .S(EBX_REG_5__SCAN_IN), .Z(n4211) );
  OR2_X1 U5234 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4210)
         );
  NAND2_X1 U5235 ( .A1(n4211), .A2(n4210), .ZN(n4826) );
  INV_X1 U5236 ( .A(n4826), .ZN(n4212) );
  INV_X1 U5237 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4214) );
  NAND2_X1 U5238 ( .A1(n4199), .A2(n4214), .ZN(n4217) );
  INV_X1 U5239 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U5240 ( .A1(n4194), .A2(n4385), .ZN(n4215) );
  OAI211_X1 U5241 ( .C1(n3098), .C2(EBX_REG_6__SCAN_IN), .A(n4215), .B(n5383), 
        .ZN(n4216) );
  AND2_X1 U5242 ( .A1(n4217), .A2(n4216), .ZN(n4954) );
  NOR2_X2 U5243 ( .A1(n4824), .A2(n4954), .ZN(n4952) );
  OR2_X1 U5244 ( .A1(n4279), .A2(EBX_REG_7__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U5245 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4218)
         );
  OAI211_X1 U5246 ( .C1(n3098), .C2(EBX_REG_7__SCAN_IN), .A(n4194), .B(n4218), 
        .ZN(n4219) );
  AND2_X1 U5247 ( .A1(n4220), .A2(n4219), .ZN(n5067) );
  INV_X1 U5248 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U5249 ( .A1(n4612), .A2(n6891), .ZN(n4223) );
  NAND2_X1 U5250 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4221)
         );
  NAND2_X1 U5251 ( .A1(n4194), .A2(n4221), .ZN(n4222) );
  NAND2_X1 U5252 ( .A1(n4223), .A2(n4222), .ZN(n4224) );
  OAI21_X1 U5253 ( .B1(EBX_REG_8__SCAN_IN), .B2(n4284), .A(n4224), .ZN(n5231)
         );
  NAND2_X1 U5254 ( .A1(n5066), .A2(n5231), .ZN(n5232) );
  MUX2_X1 U5255 ( .A(n4279), .B(n5383), .S(EBX_REG_9__SCAN_IN), .Z(n4225) );
  OAI21_X1 U5256 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4665), .A(n4225), 
        .ZN(n5249) );
  NAND2_X1 U5257 ( .A1(n4199), .A2(n5695), .ZN(n4231) );
  NAND2_X1 U5258 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4228) );
  NAND2_X1 U5259 ( .A1(n4194), .A2(n4228), .ZN(n4229) );
  OAI21_X1 U5260 ( .B1(EBX_REG_10__SCAN_IN), .B2(n3098), .A(n4229), .ZN(n4230)
         );
  MUX2_X1 U5261 ( .A(n4279), .B(n5383), .S(EBX_REG_11__SCAN_IN), .Z(n4234) );
  OR2_X1 U5262 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4233)
         );
  NAND2_X1 U5263 ( .A1(n4234), .A2(n4233), .ZN(n5689) );
  INV_X1 U5264 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U5265 ( .A1(n4199), .A2(n4235), .ZN(n4238) );
  INV_X1 U5266 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U5267 ( .A1(n4194), .A2(n6082), .ZN(n4236) );
  OAI211_X1 U5268 ( .C1(n3098), .C2(EBX_REG_12__SCAN_IN), .A(n4236), .B(n5383), 
        .ZN(n4237) );
  NAND2_X1 U5269 ( .A1(n4238), .A2(n4237), .ZN(n5683) );
  MUX2_X1 U5270 ( .A(n4279), .B(n5383), .S(EBX_REG_13__SCAN_IN), .Z(n4240) );
  OR2_X1 U5271 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4239)
         );
  NAND2_X1 U5272 ( .A1(n4240), .A2(n4239), .ZN(n5679) );
  INV_X1 U5273 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U5274 ( .A1(n4199), .A2(n5672), .ZN(n4245) );
  INV_X1 U5275 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U5276 ( .A1(n4194), .A2(n6062), .ZN(n4243) );
  OAI211_X1 U5277 ( .C1(EBX_REG_14__SCAN_IN), .C2(n3098), .A(n4243), .B(n5383), 
        .ZN(n4244) );
  NOR2_X2 U5278 ( .A1(n5574), .A2(n5575), .ZN(n5561) );
  MUX2_X1 U5279 ( .A(n4279), .B(n5383), .S(EBX_REG_15__SCAN_IN), .Z(n4247) );
  OR2_X1 U5280 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4246)
         );
  AND2_X2 U5281 ( .A1(n5561), .A2(n5562), .ZN(n5541) );
  INV_X1 U5282 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U5283 ( .A1(n4194), .A2(n5853), .ZN(n4248) );
  OAI211_X1 U5284 ( .C1(EBX_REG_16__SCAN_IN), .C2(n3098), .A(n4248), .B(n5383), 
        .ZN(n4249) );
  OAI21_X1 U5285 ( .B1(EBX_REG_16__SCAN_IN), .B2(n4284), .A(n4249), .ZN(n5543)
         );
  OR2_X1 U5286 ( .A1(n4279), .A2(EBX_REG_17__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U5287 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4250) );
  OAI211_X1 U5288 ( .C1(n3098), .C2(EBX_REG_17__SCAN_IN), .A(n4194), .B(n4250), 
        .ZN(n4251) );
  NAND2_X1 U5289 ( .A1(n4252), .A2(n4251), .ZN(n5530) );
  INV_X1 U5290 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U5291 ( .A1(n4199), .A2(n5665), .ZN(n4255) );
  INV_X1 U5292 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U5293 ( .A1(n4194), .A2(n6010), .ZN(n4253) );
  OAI211_X1 U5294 ( .C1(EBX_REG_19__SCAN_IN), .C2(n3098), .A(n4253), .B(n5383), 
        .ZN(n4254) );
  OR2_X1 U5295 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4257)
         );
  INV_X1 U5296 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U5297 ( .A1(n4612), .A2(n4256), .ZN(n5504) );
  OAI22_X1 U5298 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n3098), .ZN(n5487) );
  NAND2_X1 U5299 ( .A1(n5502), .A2(n5487), .ZN(n4259) );
  NAND2_X1 U5300 ( .A1(n5503), .A2(EBX_REG_20__SCAN_IN), .ZN(n4258) );
  OAI211_X1 U5301 ( .C1(n5502), .C2(n5503), .A(n4259), .B(n4258), .ZN(n4260)
         );
  INV_X1 U5302 ( .A(n4260), .ZN(n4261) );
  OR2_X1 U5303 ( .A1(n4279), .A2(EBX_REG_21__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U5304 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4262) );
  OAI211_X1 U5305 ( .C1(n3098), .C2(EBX_REG_21__SCAN_IN), .A(n4194), .B(n4262), 
        .ZN(n4263) );
  NAND2_X1 U5306 ( .A1(n4264), .A2(n4263), .ZN(n5475) );
  OR2_X2 U5307 ( .A1(n5476), .A2(n5475), .ZN(n5473) );
  INV_X1 U5308 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U5309 ( .A1(n4199), .A2(n5662), .ZN(n4268) );
  NAND2_X1 U5310 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U5311 ( .A1(n4194), .A2(n4265), .ZN(n4266) );
  OAI21_X1 U5312 ( .B1(EBX_REG_22__SCAN_IN), .B2(n3098), .A(n4266), .ZN(n4267)
         );
  MUX2_X1 U5313 ( .A(n4279), .B(n5383), .S(EBX_REG_23__SCAN_IN), .Z(n4270) );
  OR2_X1 U5314 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4269)
         );
  NAND2_X1 U5315 ( .A1(n4270), .A2(n4269), .ZN(n5449) );
  NOR2_X4 U5316 ( .A1(n5460), .A2(n5449), .ZN(n5448) );
  INV_X1 U5317 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5318 ( .A1(n4194), .A2(n4422), .ZN(n4271) );
  OAI211_X1 U5319 ( .C1(EBX_REG_24__SCAN_IN), .C2(n3098), .A(n4271), .B(n5383), 
        .ZN(n4272) );
  OAI21_X1 U5320 ( .B1(EBX_REG_24__SCAN_IN), .B2(n4284), .A(n4272), .ZN(n5443)
         );
  MUX2_X1 U5321 ( .A(n4279), .B(n5383), .S(EBX_REG_25__SCAN_IN), .Z(n4274) );
  OR2_X1 U5322 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4273)
         );
  NAND2_X1 U5323 ( .A1(n4274), .A2(n4273), .ZN(n5427) );
  INV_X1 U5324 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U5325 ( .A1(n4199), .A2(n4275), .ZN(n4278) );
  INV_X1 U5326 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U5327 ( .A1(n4194), .A2(n5339), .ZN(n4276) );
  OAI211_X1 U5328 ( .C1(EBX_REG_26__SCAN_IN), .C2(n3098), .A(n4276), .B(n5383), 
        .ZN(n4277) );
  MUX2_X1 U5329 ( .A(n4279), .B(n5383), .S(EBX_REG_27__SCAN_IN), .Z(n4281) );
  OR2_X1 U5330 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4280)
         );
  INV_X1 U5331 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U5332 ( .A1(n4194), .A2(n5925), .ZN(n4282) );
  OAI211_X1 U5333 ( .C1(EBX_REG_28__SCAN_IN), .C2(n3098), .A(n4282), .B(n5383), 
        .ZN(n4283) );
  OAI21_X1 U5334 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4284), .A(n4283), .ZN(n5348)
         );
  INV_X1 U5335 ( .A(n5388), .ZN(n4288) );
  AND2_X1 U5336 ( .A1(n3098), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4286)
         );
  AOI21_X1 U5337 ( .B1(n4665), .B2(EBX_REG_30__SCAN_IN), .A(n4286), .ZN(n4514)
         );
  INV_X1 U5338 ( .A(n4514), .ZN(n4287) );
  OAI21_X1 U5339 ( .B1(n4508), .B2(n4288), .A(n4287), .ZN(n4291) );
  NOR2_X1 U5340 ( .A1(n4508), .A2(n5503), .ZN(n4513) );
  INV_X1 U5341 ( .A(n4508), .ZN(n4289) );
  OAI211_X1 U5342 ( .C1(n5388), .C2(n5383), .A(n4289), .B(n4514), .ZN(n4290)
         );
  INV_X1 U5343 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U5344 ( .A1(n4601), .A2(n6467), .ZN(n5634) );
  INV_X1 U5345 ( .A(n5634), .ZN(n4296) );
  NOR2_X1 U5346 ( .A1(n3098), .A2(n4296), .ZN(n4292) );
  NOR2_X1 U5347 ( .A1(n4496), .A2(n6277), .ZN(n4311) );
  INV_X1 U5348 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U5349 ( .A1(n4293), .A2(n6943), .ZN(n4616) );
  OR2_X1 U5350 ( .A1(n4616), .A2(n5634), .ZN(n6140) );
  NAND2_X1 U5351 ( .A1(n4600), .A2(n6140), .ZN(n5377) );
  NAND3_X1 U5352 ( .A1(n3095), .A2(n5634), .A3(n5655), .ZN(n4294) );
  AND2_X1 U5353 ( .A1(n5377), .A2(n4294), .ZN(n4295) );
  NAND2_X1 U5354 ( .A1(n4758), .A2(n4616), .ZN(n4314) );
  NAND2_X1 U5355 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n4303) );
  AND2_X1 U5356 ( .A1(n6232), .A2(n6183), .ZN(n5648) );
  NAND2_X1 U5357 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5428) );
  INV_X1 U5358 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7062) );
  NOR2_X1 U5359 ( .A1(n5428), .A2(n7062), .ZN(n5406) );
  INV_X1 U5360 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6746) );
  INV_X1 U5361 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6741) );
  INV_X1 U5362 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6737) );
  INV_X1 U5363 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6969) );
  INV_X1 U5364 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6730) );
  INV_X1 U5365 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6869) );
  INV_X1 U5366 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6782) );
  INV_X1 U5367 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6728) );
  NOR3_X1 U5368 ( .A1(n6869), .A2(n6782), .A3(n6728), .ZN(n6262) );
  NAND2_X1 U5369 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6262), .ZN(n6245) );
  NOR2_X1 U5370 ( .A1(n6730), .A2(n6245), .ZN(n5602) );
  NAND2_X1 U5371 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5602), .ZN(n6231) );
  NOR2_X1 U5372 ( .A1(n6969), .A2(n6231), .ZN(n6223) );
  NAND2_X1 U5373 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6223), .ZN(n5594) );
  NOR2_X1 U5374 ( .A1(n6737), .A2(n5594), .ZN(n5589) );
  NAND2_X1 U5375 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5589), .ZN(n6204) );
  NOR2_X1 U5376 ( .A1(n6741), .A2(n6204), .ZN(n6181) );
  NAND2_X1 U5377 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6181), .ZN(n6179) );
  NOR2_X1 U5378 ( .A1(n6746), .A2(n6179), .ZN(n5570) );
  NAND2_X1 U5379 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5570), .ZN(n5571) );
  NAND2_X1 U5380 ( .A1(n6263), .A2(n5571), .ZN(n4297) );
  NAND2_X1 U5381 ( .A1(n4297), .A2(n6183), .ZN(n5580) );
  AND2_X1 U5382 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5544) );
  NAND2_X1 U5383 ( .A1(n5544), .A2(REIP_REG_17__SCAN_IN), .ZN(n4304) );
  AND2_X1 U5384 ( .A1(n6263), .A2(n4304), .ZN(n4298) );
  INV_X1 U5385 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6752) );
  INV_X1 U5386 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U5387 ( .A1(n6752), .A2(n6753), .ZN(n4299) );
  NAND2_X1 U5388 ( .A1(n4299), .A2(REIP_REG_20__SCAN_IN), .ZN(n4300) );
  AND2_X1 U5389 ( .A1(n6263), .A2(n4300), .ZN(n4301) );
  NOR2_X1 U5390 ( .A1(n5527), .A2(n4301), .ZN(n5480) );
  NAND2_X1 U5391 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .ZN(
        n4305) );
  INV_X1 U5392 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6756) );
  OAI21_X1 U5393 ( .B1(n4305), .B2(n6756), .A(n6263), .ZN(n4302) );
  OAI21_X1 U5394 ( .B1(n5648), .B2(n5406), .A(n5450), .ZN(n5417) );
  AOI21_X1 U5395 ( .B1(n6263), .B2(n4303), .A(n5417), .ZN(n5350) );
  NAND2_X1 U5396 ( .A1(n5350), .A2(REIP_REG_29__SCAN_IN), .ZN(n5392) );
  NAND3_X1 U5397 ( .A1(n5392), .A2(REIP_REG_30__SCAN_IN), .A3(n5615), .ZN(
        n4307) );
  NOR2_X1 U5398 ( .A1(n5560), .A2(n4304), .ZN(n5497) );
  NAND3_X1 U5399 ( .A1(n5429), .A2(REIP_REG_27__SCAN_IN), .A3(n5406), .ZN(
        n5391) );
  INV_X1 U5400 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7075) );
  INV_X1 U5401 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6768) );
  NOR3_X1 U5402 ( .A1(n5391), .A2(n7075), .A3(n6768), .ZN(n5374) );
  INV_X1 U5403 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U5404 ( .A1(n6234), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(n5374), 
        .B2(n6770), .ZN(n4306) );
  INV_X1 U5405 ( .A(n4309), .ZN(n4539) );
  NAND2_X1 U5406 ( .A1(n4602), .A2(n4616), .ZN(n4312) );
  NOR2_X1 U5407 ( .A1(READY_N), .A2(n4572), .ZN(n4578) );
  NAND2_X1 U5408 ( .A1(n4312), .A2(n4578), .ZN(n4318) );
  NAND2_X1 U5409 ( .A1(n4314), .A2(n4601), .ZN(n4315) );
  OAI211_X1 U5410 ( .C1(n4654), .C2(n4315), .A(n4187), .B(n5357), .ZN(n4316)
         );
  NAND2_X1 U5411 ( .A1(n4652), .A2(n4316), .ZN(n4317) );
  MUX2_X1 U5412 ( .A(n4318), .B(n4317), .S(n4753), .Z(n4329) );
  INV_X1 U5413 ( .A(n4573), .ZN(n4326) );
  NAND2_X1 U5414 ( .A1(n4319), .A2(n3095), .ZN(n4322) );
  MUX2_X1 U5415 ( .A(n4322), .B(n6794), .S(n4321), .Z(n4453) );
  NAND2_X1 U5416 ( .A1(n5315), .A2(n4748), .ZN(n4324) );
  NAND2_X1 U5417 ( .A1(n4453), .A2(n4439), .ZN(n4325) );
  NAND2_X1 U5418 ( .A1(n4326), .A2(n4325), .ZN(n4582) );
  NOR2_X1 U5419 ( .A1(n5315), .A2(n4758), .ZN(n4458) );
  INV_X1 U5420 ( .A(n4458), .ZN(n4327) );
  OR2_X1 U5421 ( .A1(n4652), .A2(n4327), .ZN(n4328) );
  NAND3_X1 U5422 ( .A1(n4329), .A2(n4582), .A3(n4328), .ZN(n4330) );
  NAND2_X1 U5423 ( .A1(n4438), .A2(n4763), .ZN(n4331) );
  NAND2_X1 U5424 ( .A1(n4615), .A2(n4331), .ZN(n4332) );
  NOR2_X1 U5425 ( .A1(n4496), .A2(n6398), .ZN(n4487) );
  NAND2_X1 U5426 ( .A1(n4813), .A2(n4388), .ZN(n4338) );
  NAND2_X1 U5427 ( .A1(n4348), .A2(n4355), .ZN(n4347) );
  NAND2_X1 U5428 ( .A1(n4347), .A2(n4342), .ZN(n4341) );
  NAND2_X1 U5429 ( .A1(n4341), .A2(n4336), .ZN(n4372) );
  OAI211_X1 U5430 ( .C1(n4336), .C2(n4341), .A(n4372), .B(n4600), .ZN(n4337)
         );
  NAND2_X1 U5431 ( .A1(n4338), .A2(n4337), .ZN(n4360) );
  INV_X1 U5432 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4339) );
  OAI21_X1 U5433 ( .B1(n4342), .B2(n4347), .A(n4341), .ZN(n4343) );
  AND2_X1 U5434 ( .A1(n4748), .A2(n3417), .ZN(n4353) );
  AOI21_X1 U5435 ( .B1(n4343), .B2(n4600), .A(n4353), .ZN(n4344) );
  NAND2_X1 U5436 ( .A1(n4345), .A2(n4344), .ZN(n4346) );
  NAND2_X1 U5437 ( .A1(n4346), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6359)
         );
  NAND2_X1 U5438 ( .A1(n3097), .A2(n4388), .ZN(n4352) );
  OAI21_X1 U5439 ( .B1(n4355), .B2(n4348), .A(n4347), .ZN(n4349) );
  OAI211_X1 U5440 ( .C1(n4349), .C2(n6794), .A(n4447), .B(n3810), .ZN(n4350)
         );
  INV_X1 U5441 ( .A(n4350), .ZN(n4351) );
  NAND2_X1 U5442 ( .A1(n4352), .A2(n4351), .ZN(n4829) );
  INV_X1 U5443 ( .A(n4353), .ZN(n4354) );
  OAI21_X1 U5444 ( .B1(n6794), .B2(n4355), .A(n4354), .ZN(n4356) );
  INV_X1 U5445 ( .A(n4356), .ZN(n4357) );
  NAND2_X1 U5446 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4623)
         );
  XNOR2_X1 U5447 ( .A(n4623), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4828)
         );
  INV_X1 U5448 ( .A(n4623), .ZN(n4358) );
  NAND2_X1 U5449 ( .A1(n4358), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4359)
         );
  NAND2_X1 U5450 ( .A1(n4692), .A2(n4691), .ZN(n4362) );
  NAND2_X1 U5451 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4361)
         );
  NAND2_X1 U5452 ( .A1(n4362), .A2(n4361), .ZN(n5047) );
  XNOR2_X1 U5453 ( .A(n4372), .B(n4370), .ZN(n4363) );
  NAND2_X1 U5454 ( .A1(n4363), .A2(n4600), .ZN(n4364) );
  XNOR2_X1 U5455 ( .A(n4367), .B(n4366), .ZN(n5048) );
  NAND2_X1 U5456 ( .A1(n5047), .A2(n5048), .ZN(n4369) );
  NAND2_X1 U5457 ( .A1(n4367), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4368)
         );
  NAND2_X1 U5458 ( .A1(n4369), .A2(n4368), .ZN(n4993) );
  INV_X1 U5459 ( .A(n4370), .ZN(n4371) );
  NOR2_X1 U5460 ( .A1(n4372), .A2(n4371), .ZN(n4374) );
  NAND2_X1 U5461 ( .A1(n4374), .A2(n4373), .ZN(n4390) );
  OAI211_X1 U5462 ( .C1(n4374), .C2(n4373), .A(n4390), .B(n4600), .ZN(n4375)
         );
  OAI21_X1 U5463 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(n4379) );
  INV_X1 U5464 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4378) );
  XNOR2_X1 U5465 ( .A(n4379), .B(n4378), .ZN(n4994) );
  NAND2_X1 U5466 ( .A1(n4379), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4380)
         );
  XNOR2_X1 U5467 ( .A(n4390), .B(n4391), .ZN(n4382) );
  NAND2_X1 U5468 ( .A1(n4382), .A2(n4600), .ZN(n4383) );
  NAND2_X1 U5469 ( .A1(n4384), .A2(n4383), .ZN(n4386) );
  XNOR2_X1 U5470 ( .A(n4386), .B(n4385), .ZN(n5184) );
  NAND2_X1 U5471 ( .A1(n4386), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4387)
         );
  NAND2_X1 U5472 ( .A1(n4389), .A2(n4388), .ZN(n4395) );
  INV_X1 U5473 ( .A(n4390), .ZN(n4392) );
  NAND2_X1 U5474 ( .A1(n4392), .A2(n4391), .ZN(n4401) );
  XNOR2_X1 U5475 ( .A(n4401), .B(n4399), .ZN(n4393) );
  NAND2_X1 U5476 ( .A1(n4393), .A2(n4600), .ZN(n4394) );
  NAND2_X1 U5477 ( .A1(n4395), .A2(n4394), .ZN(n4397) );
  INV_X1 U5478 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5479 ( .A1(n4397), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4398)
         );
  NAND2_X1 U5480 ( .A1(n4600), .A2(n4399), .ZN(n4400) );
  OR2_X1 U5481 ( .A1(n4401), .A2(n4400), .ZN(n4402) );
  NAND2_X1 U5482 ( .A1(n4407), .A2(n4402), .ZN(n4404) );
  INV_X1 U5483 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4403) );
  XNOR2_X1 U5484 ( .A(n4404), .B(n4403), .ZN(n5294) );
  NAND2_X1 U5485 ( .A1(n4404), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4405)
         );
  INV_X1 U5486 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7064) );
  NOR2_X1 U5487 ( .A1(n4407), .A2(n7064), .ZN(n4408) );
  NAND2_X1 U5488 ( .A1(n4407), .A2(n7064), .ZN(n4409) );
  INV_X1 U5489 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6383) );
  AND2_X1 U5490 ( .A1(n4407), .A2(n6383), .ZN(n5899) );
  INV_X1 U5491 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U5492 ( .A1(n4407), .A2(n6099), .ZN(n6090) );
  NAND2_X1 U5493 ( .A1(n4407), .A2(n6082), .ZN(n5890) );
  NOR2_X1 U5494 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4410) );
  OR2_X1 U5495 ( .A1(n4407), .A2(n4410), .ZN(n4411) );
  XNOR2_X1 U5496 ( .A(n4407), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5885)
         );
  INV_X1 U5497 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U5498 ( .A1(n4407), .A2(n6072), .ZN(n4413) );
  NAND2_X1 U5499 ( .A1(n4407), .A2(n6062), .ZN(n4414) );
  AND2_X1 U5500 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4462) );
  AND2_X1 U5501 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5502 ( .A1(n4462), .A2(n4463), .ZN(n4416) );
  AND2_X1 U5503 ( .A1(n4407), .A2(n4416), .ZN(n4420) );
  INV_X1 U5504 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6031) );
  INV_X1 U5505 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U5506 ( .A1(n7026), .A2(n5853), .ZN(n5842) );
  NOR2_X1 U5507 ( .A1(n5842), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4417)
         );
  OR2_X1 U5508 ( .A1(n4407), .A2(n4417), .ZN(n4418) );
  NAND2_X1 U5509 ( .A1(n4407), .A2(n6010), .ZN(n5831) );
  AND2_X1 U5510 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5976) );
  AND2_X1 U5511 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4473) );
  NAND3_X1 U5512 ( .A1(n5976), .A2(n4473), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U5513 ( .A1(n4407), .A2(n4421), .ZN(n4424) );
  NOR2_X1 U5514 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5991) );
  NOR2_X1 U5515 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5975) );
  INV_X1 U5516 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5967) );
  AND4_X1 U5517 ( .A1(n5991), .A2(n5975), .A3(n4422), .A4(n5967), .ZN(n4423)
         );
  XNOR2_X1 U5518 ( .A(n4407), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5788)
         );
  AND2_X1 U5519 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4502) );
  INV_X1 U5520 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4480) );
  AND2_X1 U5521 ( .A1(n4480), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4483)
         );
  NAND4_X1 U5522 ( .A1(n4407), .A2(n4502), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n4483), .ZN(n4425) );
  NAND2_X1 U5523 ( .A1(n4479), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5524 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4517) );
  INV_X1 U5525 ( .A(n4517), .ZN(n4428) );
  AOI21_X1 U5526 ( .B1(n4502), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n4517), 
        .ZN(n4427) );
  NOR2_X1 U5527 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5920) );
  NOR2_X1 U5528 ( .A1(n5920), .A2(n4430), .ZN(n4426) );
  AOI211_X1 U5529 ( .C1(n4524), .C2(n4428), .A(n4427), .B(n4426), .ZN(n4429)
         );
  OAI21_X1 U5530 ( .B1(n5779), .B2(n4430), .A(n4429), .ZN(n4431) );
  INV_X1 U5531 ( .A(n4431), .ZN(n4432) );
  INV_X1 U5532 ( .A(n4433), .ZN(n4437) );
  NAND2_X1 U5533 ( .A1(n5779), .A2(n5920), .ZN(n5760) );
  NOR2_X1 U5534 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4503) );
  INV_X1 U5535 ( .A(n4503), .ZN(n4434) );
  OAI21_X1 U5536 ( .B1(n5760), .B2(n4434), .A(n4517), .ZN(n4435) );
  INV_X1 U5537 ( .A(n4577), .ZN(n4780) );
  AOI22_X1 U5538 ( .A1(n3440), .A2(n4612), .B1(n4438), .B2(n4489), .ZN(n4440)
         );
  NAND3_X1 U5539 ( .A1(n4780), .A2(n4440), .A3(n6133), .ZN(n4441) );
  OR2_X1 U5540 ( .A1(n4441), .A2(n4595), .ZN(n4442) );
  NAND2_X1 U5541 ( .A1(n5357), .A2(n4443), .ZN(n4444) );
  OAI211_X1 U5542 ( .C1(n4446), .C2(n5383), .A(n4445), .B(n4444), .ZN(n4450)
         );
  NAND2_X1 U5543 ( .A1(n5611), .A2(n4753), .ZN(n4581) );
  AOI21_X1 U5544 ( .B1(n4448), .B2(n4581), .A(n4447), .ZN(n4449) );
  NOR2_X1 U5545 ( .A1(n4450), .A2(n4449), .ZN(n4452) );
  NAND3_X1 U5546 ( .A1(n4453), .A2(n4452), .A3(n4451), .ZN(n4656) );
  OAI21_X1 U5547 ( .B1(n4454), .B2(n3095), .A(n4793), .ZN(n4455) );
  INV_X1 U5548 ( .A(n4459), .ZN(n4456) );
  AND2_X2 U5549 ( .A1(n6037), .A2(n4457), .ZN(n6392) );
  NAND2_X1 U5550 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6807) );
  NAND4_X1 U5551 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4998) );
  NOR2_X1 U5552 ( .A1(n6807), .A2(n4998), .ZN(n5297) );
  NAND2_X1 U5553 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6373) );
  NOR3_X1 U5554 ( .A1(n7064), .A2(n6383), .A3(n6373), .ZN(n4460) );
  NAND2_X1 U5555 ( .A1(n5297), .A2(n4460), .ZN(n6036) );
  INV_X1 U5556 ( .A(n6036), .ZN(n4464) );
  NAND2_X1 U5557 ( .A1(n4459), .A2(n4458), .ZN(n4781) );
  INV_X1 U5558 ( .A(n4781), .ZN(n4569) );
  INV_X1 U5559 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U5560 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U5561 ( .A1(n6404), .A2(n6805), .ZN(n6393) );
  NAND3_X1 U5562 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6393), .ZN(n5299) );
  NAND2_X1 U5563 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6060) );
  NOR2_X1 U5564 ( .A1(n6060), .A2(n6072), .ZN(n6063) );
  AND2_X1 U5565 ( .A1(n6063), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6042)
         );
  AND2_X1 U5566 ( .A1(n6042), .A2(n4462), .ZN(n4466) );
  AND2_X1 U5567 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U5568 ( .A1(n6011), .A2(n5990), .ZN(n5985) );
  INV_X1 U5569 ( .A(n5976), .ZN(n4471) );
  NOR2_X2 U5570 ( .A1(n5985), .A2(n4471), .ZN(n5964) );
  NAND2_X1 U5571 ( .A1(n5964), .A2(n4473), .ZN(n5951) );
  NAND2_X1 U5572 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5573 ( .A1(n5936), .A2(n4502), .ZN(n5916) );
  INV_X1 U5574 ( .A(n5916), .ZN(n4484) );
  NAND2_X1 U5575 ( .A1(n4464), .A2(n4466), .ZN(n4465) );
  NAND2_X1 U5576 ( .A1(n6037), .A2(n4465), .ZN(n5995) );
  NAND4_X1 U5577 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U5578 ( .A1(n6037), .A2(n4468), .ZN(n4470) );
  NAND2_X1 U5579 ( .A1(n6054), .A2(n4466), .ZN(n5993) );
  INV_X1 U5580 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7047) );
  AND2_X1 U5581 ( .A1(n7047), .A2(n6059), .ZN(n4669) );
  NOR2_X1 U5582 ( .A1(n4467), .A2(n6377), .ZN(n4670) );
  NAND2_X1 U5583 ( .A1(n5004), .A2(n6407), .ZN(n6039) );
  OAI21_X1 U5584 ( .B1(n4468), .B2(n5993), .A(n6039), .ZN(n4469) );
  NAND2_X1 U5585 ( .A1(n6415), .A2(n4471), .ZN(n4472) );
  AND2_X1 U5586 ( .A1(n5974), .A2(n4472), .ZN(n5968) );
  INV_X1 U5587 ( .A(n4473), .ZN(n4474) );
  OAI21_X1 U5588 ( .B1(n6392), .B2(n6395), .A(n4474), .ZN(n4475) );
  AND2_X2 U5589 ( .A1(n5968), .A2(n4475), .ZN(n5958) );
  NAND2_X1 U5590 ( .A1(n6415), .A2(n4476), .ZN(n4477) );
  AND2_X2 U5591 ( .A1(n5958), .A2(n4477), .ZN(n5931) );
  INV_X1 U5592 ( .A(n4502), .ZN(n5921) );
  NAND2_X1 U5593 ( .A1(n6415), .A2(n5921), .ZN(n4478) );
  NAND2_X1 U5594 ( .A1(n5931), .A2(n4478), .ZN(n5913) );
  AOI21_X1 U5595 ( .B1(n4479), .B2(n6415), .A(n5913), .ZN(n4481) );
  NAND2_X1 U5596 ( .A1(n6377), .A2(REIP_REG_30__SCAN_IN), .ZN(n4540) );
  OAI21_X1 U5597 ( .B1(n4481), .B2(n4480), .A(n4540), .ZN(n4482) );
  OR2_X1 U5598 ( .A1(n4487), .A2(n4486), .ZN(U2988) );
  AND2_X1 U5599 ( .A1(n4733), .A2(n4488), .ZN(n4492) );
  NOR2_X1 U5600 ( .A1(n3810), .A2(n6152), .ZN(n4491) );
  NOR2_X1 U5601 ( .A1(n4842), .A2(n4489), .ZN(n4490) );
  NAND4_X1 U5602 ( .A1(n4492), .A2(n4753), .A3(n4491), .A4(n4490), .ZN(n4837)
         );
  INV_X1 U5603 ( .A(n4837), .ZN(n4493) );
  NAND2_X1 U5604 ( .A1(n4493), .A2(n4612), .ZN(n4494) );
  INV_X1 U5605 ( .A(n4496), .ZN(n4500) );
  OAI21_X1 U5606 ( .B1(n5365), .B2(n5694), .A(n4501), .ZN(U2829) );
  NAND2_X1 U5607 ( .A1(n4407), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5780) );
  NAND3_X1 U5608 ( .A1(n5779), .A2(n4503), .A3(n5920), .ZN(n4504) );
  OR2_X1 U5609 ( .A1(n5787), .A2(n4504), .ZN(n4505) );
  XNOR2_X1 U5610 ( .A(n4507), .B(n4506), .ZN(n5756) );
  INV_X1 U5611 ( .A(n5756), .ZN(n4523) );
  NAND2_X1 U5612 ( .A1(n4508), .A2(n5383), .ZN(n4512) );
  INV_X1 U5613 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U5614 ( .A1(n4199), .A2(n4509), .ZN(n5385) );
  INV_X1 U5615 ( .A(n5385), .ZN(n4510) );
  AOI21_X1 U5616 ( .B1(n4514), .B2(n5390), .A(n4513), .ZN(n4516) );
  AOI22_X1 U5617 ( .A1(n4665), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3098), .ZN(n4515) );
  XNOR2_X1 U5618 ( .A(n4516), .B(n4515), .ZN(n5654) );
  NOR3_X1 U5619 ( .A1(n5916), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4517), 
        .ZN(n4520) );
  AOI21_X1 U5620 ( .B1(n4517), .B2(n6415), .A(n5913), .ZN(n4518) );
  NAND2_X1 U5621 ( .A1(n6377), .A2(REIP_REG_31__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U5622 ( .B1(n4518), .B2(n4506), .A(n5753), .ZN(n4519) );
  AOI21_X1 U5623 ( .B1(n5654), .B2(n6410), .A(n4521), .ZN(n4522) );
  OAI21_X1 U5624 ( .B1(n4523), .B2(n6101), .A(n4522), .ZN(U2987) );
  INV_X1 U5625 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5999) );
  AND2_X1 U5626 ( .A1(n4524), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5830)
         );
  XNOR2_X1 U5627 ( .A(n4407), .B(n5999), .ZN(n5823) );
  XNOR2_X1 U5628 ( .A(n4524), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5813)
         );
  NOR2_X1 U5629 ( .A1(n4407), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5795)
         );
  AOI21_X1 U5630 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4407), .A(n5795), 
        .ZN(n4525) );
  INV_X1 U5631 ( .A(n4525), .ZN(n4526) );
  NAND2_X1 U5632 ( .A1(n5973), .A2(n6366), .ZN(n4538) );
  OAI21_X1 U5633 ( .B1(n3099), .B2(n4528), .A(n4527), .ZN(n5718) );
  NAND2_X1 U5634 ( .A1(n4529), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6717) );
  NAND2_X1 U5635 ( .A1(n4530), .A2(n6651), .ZN(n6790) );
  NAND2_X1 U5636 ( .A1(n6790), .A2(n7027), .ZN(n4531) );
  INV_X1 U5637 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6758) );
  NOR2_X1 U5638 ( .A1(n6396), .A2(n6758), .ZN(n5978) );
  NAND2_X1 U5639 ( .A1(n6467), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U5640 ( .A1(n7027), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4532) );
  NAND2_X1 U5641 ( .A1(n4533), .A2(n4532), .ZN(n4625) );
  NOR2_X1 U5642 ( .A1(n5457), .A2(n6370), .ZN(n4534) );
  AOI211_X1 U5643 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5978), 
        .B(n4534), .ZN(n4535) );
  INV_X1 U5644 ( .A(n4536), .ZN(n4537) );
  NAND2_X1 U5645 ( .A1(n4538), .A2(n4537), .ZN(U2964) );
  NOR2_X1 U5646 ( .A1(n3285), .A2(n6339), .ZN(n4545) );
  NAND2_X1 U5647 ( .A1(n4539), .A2(n6350), .ZN(n4543) );
  OAI21_X1 U5648 ( .B1(n6356), .B2(n6937), .A(n4540), .ZN(n4541) );
  INV_X1 U5649 ( .A(n4541), .ZN(n4542) );
  INV_X1 U5650 ( .A(HOLD), .ZN(n7001) );
  INV_X1 U5651 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4556) );
  NOR2_X1 U5652 ( .A1(n7001), .A2(n4556), .ZN(n4552) );
  INV_X1 U5653 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4551) );
  NOR2_X1 U5654 ( .A1(n6943), .A2(n4551), .ZN(n6719) );
  NOR2_X1 U5655 ( .A1(n4552), .A2(n6719), .ZN(n4548) );
  NOR2_X1 U5656 ( .A1(n7001), .A2(n4550), .ZN(n4549) );
  NAND2_X1 U5657 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n4547) );
  OAI211_X1 U5658 ( .C1(n4548), .C2(n4549), .A(n4547), .B(n4616), .ZN(U3182)
         );
  AOI21_X1 U5659 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n4549), .ZN(
        n6724) );
  NOR2_X1 U5660 ( .A1(n4556), .A2(n4550), .ZN(n4555) );
  INV_X1 U5661 ( .A(NA_N), .ZN(n6965) );
  AOI221_X1 U5662 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6965), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6721) );
  INV_X1 U5663 ( .A(n6721), .ZN(n4554) );
  OAI21_X1 U5664 ( .B1(n4552), .B2(n4551), .A(n6800), .ZN(n4553) );
  OAI211_X1 U5665 ( .C1(n6724), .C2(n4555), .A(n4554), .B(n4553), .ZN(U3181)
         );
  INV_X1 U5666 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4558) );
  OAI21_X1 U5667 ( .B1(n4556), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4557) );
  OAI21_X1 U5668 ( .B1(n6789), .B2(n4558), .A(n6718), .ZN(U2789) );
  OR2_X1 U5669 ( .A1(n4652), .A2(n5609), .ZN(n4561) );
  NAND2_X1 U5670 ( .A1(n4559), .A2(n4568), .ZN(n4560) );
  NAND2_X1 U5671 ( .A1(n4561), .A2(n4560), .ZN(n4567) );
  OAI21_X1 U5672 ( .B1(n4567), .B2(n6152), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4563) );
  NAND3_X1 U5673 ( .A1(n6155), .A2(STATE2_REG_0__SCAN_IN), .A3(n6592), .ZN(
        n4562) );
  NAND2_X1 U5674 ( .A1(n4563), .A2(n4562), .ZN(U2790) );
  INV_X1 U5675 ( .A(n4564), .ZN(n5498) );
  INV_X1 U5676 ( .A(n4604), .ZN(n4599) );
  AOI211_X1 U5677 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4565), .A(n5498), .B(
        n4599), .ZN(n4566) );
  INV_X1 U5678 ( .A(n4566), .ZN(U2788) );
  OR2_X1 U5679 ( .A1(n4600), .A2(n5611), .ZN(n5366) );
  AOI21_X1 U5680 ( .B1(n5366), .B2(n4616), .A(READY_N), .ZN(n6793) );
  NOR2_X1 U5681 ( .A1(n4567), .A2(n6793), .ZN(n6131) );
  OR2_X1 U5682 ( .A1(n6131), .A2(n6152), .ZN(n4574) );
  INV_X1 U5683 ( .A(n4574), .ZN(n6165) );
  INV_X1 U5684 ( .A(MORE_REG_SCAN_IN), .ZN(n4576) );
  NAND3_X1 U5685 ( .A1(n4780), .A2(n4568), .A3(n6133), .ZN(n4570) );
  MUX2_X1 U5686 ( .A(n4570), .B(n4569), .S(n4652), .Z(n4571) );
  AOI21_X1 U5687 ( .B1(n4573), .B2(n4572), .A(n4571), .ZN(n6134) );
  OR2_X1 U5688 ( .A1(n6134), .A2(n4574), .ZN(n4575) );
  OAI21_X1 U5689 ( .B1(n6165), .B2(n4576), .A(n4575), .ZN(U3471) );
  NAND2_X1 U5690 ( .A1(n4652), .A2(n4577), .ZN(n4580) );
  NAND2_X1 U5691 ( .A1(n4595), .A2(n4578), .ZN(n4579) );
  NAND2_X1 U5692 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  NOR2_X1 U5693 ( .A1(n4839), .A2(n4583), .ZN(n4589) );
  INV_X1 U5694 ( .A(n4616), .ZN(n4585) );
  NAND2_X1 U5695 ( .A1(n3098), .A2(n4616), .ZN(n4584) );
  AOI22_X1 U5696 ( .A1(n6117), .A2(n4585), .B1(n3440), .B2(n4584), .ZN(n4586)
         );
  OR2_X1 U5697 ( .A1(n4586), .A2(READY_N), .ZN(n4587) );
  MUX2_X1 U5698 ( .A(n4781), .B(n4587), .S(n4652), .Z(n4588) );
  AND2_X1 U5699 ( .A1(n4890), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U5700 ( .A1(n6779), .A2(FLUSH_REG_SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5701 ( .A1(n7027), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4592) );
  INV_X1 U5702 ( .A(n6495), .ZN(n6654) );
  NOR2_X1 U5703 ( .A1(n4593), .A2(n6654), .ZN(n4594) );
  XNOR2_X1 U5704 ( .A(n4594), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6268)
         );
  INV_X1 U5705 ( .A(n4595), .ZN(n4658) );
  NOR3_X1 U5706 ( .A1(n6268), .A2(STATE2_REG_1__SCAN_IN), .A3(n4658), .ZN(
        n4808) );
  NAND2_X1 U5707 ( .A1(n4808), .A2(n4816), .ZN(n4597) );
  OAI22_X1 U5708 ( .A1(n4598), .A2(n6115), .B1(n4597), .B2(n4596), .ZN(U3455)
         );
  OAI21_X1 U5709 ( .B1(n4600), .B2(n4601), .A(n4599), .ZN(n4642) );
  AOI22_X1 U5710 ( .A1(n4642), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n6324), .ZN(n4605) );
  NAND2_X1 U5711 ( .A1(n4602), .A2(n4601), .ZN(n4603) );
  NAND2_X1 U5712 ( .A1(n6327), .A2(DATAI_11_), .ZN(n4682) );
  NAND2_X1 U5713 ( .A1(n4605), .A2(n4682), .ZN(U2935) );
  AOI22_X1 U5714 ( .A1(n4642), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6324), .ZN(n4606) );
  NAND2_X1 U5715 ( .A1(n6327), .A2(DATAI_8_), .ZN(n4689) );
  NAND2_X1 U5716 ( .A1(n4606), .A2(n4689), .ZN(U2932) );
  AOI22_X1 U5717 ( .A1(n4642), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6324), .ZN(n4607) );
  NAND2_X1 U5718 ( .A1(n6327), .A2(DATAI_7_), .ZN(n4685) );
  NAND2_X1 U5719 ( .A1(n4607), .A2(n4685), .ZN(U2931) );
  OAI21_X1 U5720 ( .B1(n4610), .B2(n4609), .A(n4608), .ZN(n5642) );
  OAI21_X1 U5721 ( .B1(n4613), .B2(n4612), .A(n4611), .ZN(n6409) );
  AOI22_X1 U5722 ( .A1(n4499), .A2(n6409), .B1(n5684), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4614) );
  OAI21_X1 U5723 ( .B1(n5642), .B2(n5694), .A(n4614), .ZN(U2858) );
  INV_X1 U5724 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4622) );
  INV_X1 U5725 ( .A(n4615), .ZN(n6143) );
  NOR2_X1 U5726 ( .A1(n6117), .A2(n6143), .ZN(n4617) );
  NOR2_X2 U5727 ( .A1(n6302), .A2(n4748), .ZN(n6282) );
  INV_X1 U5728 ( .A(n6282), .ZN(n4621) );
  INV_X1 U5729 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4620) );
  INV_X1 U5730 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4619) );
  OAI222_X1 U5731 ( .A1(n4622), .A2(n6299), .B1(n4621), .B2(n4620), .C1(n6306), 
        .C2(n4619), .ZN(U2899) );
  OAI21_X1 U5732 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4624), .A(n4623), 
        .ZN(n4673) );
  OAI21_X1 U5733 ( .B1(n6358), .B2(n4625), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4632) );
  OR2_X1 U5734 ( .A1(n4627), .A2(n4626), .ZN(n4629) );
  NAND2_X1 U5735 ( .A1(n4629), .A2(n4628), .ZN(n5652) );
  INV_X1 U5736 ( .A(n5652), .ZN(n4630) );
  INV_X1 U5737 ( .A(REIP_REG_0__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U5738 ( .A1(n6396), .A2(n7077), .ZN(n4668) );
  AOI21_X1 U5739 ( .B1(n4630), .B2(n6365), .A(n4668), .ZN(n4631) );
  OAI211_X1 U5740 ( .C1(n4673), .C2(n6339), .A(n4632), .B(n4631), .ZN(U2986)
         );
  AOI222_X1 U5741 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_17__SCAN_IN), .C1(n6300), .C2(UWORD_REG_1__SCAN_IN), .ZN(
        n4633) );
  INV_X1 U5742 ( .A(n4633), .ZN(U2906) );
  AOI222_X1 U5743 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_20__SCAN_IN), .C1(n6300), .C2(UWORD_REG_4__SCAN_IN), .ZN(
        n4634) );
  INV_X1 U5744 ( .A(n4634), .ZN(U2903) );
  AOI222_X1 U5745 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_16__SCAN_IN), .C1(n6300), .C2(UWORD_REG_0__SCAN_IN), .ZN(
        n4635) );
  INV_X1 U5746 ( .A(n4635), .ZN(U2907) );
  AOI222_X1 U5747 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6300), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n4636) );
  INV_X1 U5748 ( .A(n4636), .ZN(U2902) );
  AOI222_X1 U5749 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_18__SCAN_IN), .C1(n6300), .C2(UWORD_REG_2__SCAN_IN), .ZN(
        n4637) );
  INV_X1 U5750 ( .A(n4637), .ZN(U2905) );
  AOI222_X1 U5751 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6300), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4638) );
  INV_X1 U5752 ( .A(n4638), .ZN(U2901) );
  AOI222_X1 U5753 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6300), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4639) );
  INV_X1 U5754 ( .A(n4639), .ZN(U2893) );
  AOI222_X1 U5755 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_25__SCAN_IN), .C1(n6300), .C2(UWORD_REG_9__SCAN_IN), .ZN(
        n4640) );
  INV_X1 U5756 ( .A(n4640), .ZN(U2898) );
  AOI222_X1 U5757 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6282), .B1(n6303), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6300), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n4641) );
  INV_X1 U5758 ( .A(n4641), .ZN(U2895) );
  INV_X1 U5759 ( .A(DATAI_3_), .ZN(n4644) );
  INV_X1 U5760 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n7000) );
  INV_X1 U5761 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4643) );
  OAI222_X1 U5762 ( .A1(n4644), .A2(n4841), .B1(n4681), .B2(n7000), .C1(n4643), 
        .C2(n6330), .ZN(U2927) );
  INV_X1 U5763 ( .A(DATAI_0_), .ZN(n4853) );
  INV_X1 U5764 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6998) );
  OAI222_X1 U5765 ( .A1(n4853), .A2(n4841), .B1(n4681), .B2(n6998), .C1(n4645), 
        .C2(n6330), .ZN(U2924) );
  INV_X1 U5766 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4646) );
  INV_X1 U5767 ( .A(DATAI_4_), .ZN(n4849) );
  OAI222_X1 U5768 ( .A1(n6330), .A2(n6297), .B1(n4646), .B2(n4681), .C1(n4841), 
        .C2(n4849), .ZN(U2943) );
  INV_X1 U5769 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4647) );
  INV_X1 U5770 ( .A(DATAI_1_), .ZN(n4846) );
  OAI222_X1 U5771 ( .A1(n6330), .A2(n4648), .B1(n4647), .B2(n4681), .C1(n4841), 
        .C2(n4846), .ZN(U2940) );
  INV_X1 U5772 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4649) );
  INV_X1 U5773 ( .A(DATAI_6_), .ZN(n4956) );
  OAI222_X1 U5774 ( .A1(n6330), .A2(n4650), .B1(n4649), .B2(n4681), .C1(n4841), 
        .C2(n4956), .ZN(U2945) );
  INV_X1 U5775 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4651) );
  OAI222_X1 U5776 ( .A1(n6330), .A2(n4854), .B1(n4651), .B2(n4681), .C1(n4841), 
        .C2(n4853), .ZN(U2939) );
  AOI21_X1 U5777 ( .B1(n6117), .B2(n6155), .A(n5333), .ZN(n4662) );
  INV_X1 U5778 ( .A(n6145), .ZN(n5325) );
  NAND3_X1 U5779 ( .A1(n4654), .A2(n4454), .A3(n4653), .ZN(n4655) );
  NOR2_X1 U5780 ( .A1(n4656), .A2(n4655), .ZN(n4657) );
  AND2_X1 U5781 ( .A1(n4658), .A2(n4657), .ZN(n5316) );
  INV_X1 U5782 ( .A(n5316), .ZN(n4802) );
  NOR2_X1 U5783 ( .A1(n5315), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4659)
         );
  AOI21_X1 U5784 ( .B1(n6583), .B2(n4802), .A(n4659), .ZN(n6119) );
  OAI22_X1 U5785 ( .A1(n6119), .A2(n6113), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6810), .ZN(n4660) );
  AOI21_X1 U5786 ( .B1(n5325), .B2(n3288), .A(n4660), .ZN(n4661) );
  OAI22_X1 U5787 ( .A1(n4662), .A2(n3288), .B1(n5333), .B2(n4661), .ZN(U3461)
         );
  INV_X1 U5788 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n7015) );
  OAI22_X1 U5789 ( .A1(n4681), .A2(n7015), .B1(n5742), .B2(n6330), .ZN(n4663)
         );
  INV_X1 U5790 ( .A(DATAI_12_), .ZN(n5743) );
  NOR2_X1 U5791 ( .A1(n4841), .A2(n5743), .ZN(n6317) );
  OR2_X1 U5792 ( .A1(n4663), .A2(n6317), .ZN(U2951) );
  INV_X1 U5793 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n7092) );
  OAI22_X1 U5794 ( .A1(n4681), .A2(n7092), .B1(n5253), .B2(n6330), .ZN(n4664)
         );
  INV_X1 U5795 ( .A(DATAI_9_), .ZN(n5252) );
  NOR2_X1 U5796 ( .A1(n4841), .A2(n5252), .ZN(n6314) );
  OR2_X1 U5797 ( .A1(n4664), .A2(n6314), .ZN(U2948) );
  OR2_X1 U5798 ( .A1(n4665), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4667)
         );
  AND2_X1 U5799 ( .A1(n4667), .A2(n4666), .ZN(n5645) );
  AOI211_X1 U5800 ( .C1(n6410), .C2(n5645), .A(n4669), .B(n4668), .ZN(n4672)
         );
  OAI21_X1 U5801 ( .B1(n6416), .B2(n4670), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4671) );
  OAI211_X1 U5802 ( .C1(n6101), .C2(n4673), .A(n4672), .B(n4671), .ZN(U3018)
         );
  NAND2_X1 U5803 ( .A1(n4675), .A2(n4674), .ZN(n4676) );
  NAND2_X1 U5804 ( .A1(n4773), .A2(n4676), .ZN(n6397) );
  INV_X1 U5805 ( .A(n4608), .ZN(n4678) );
  OAI21_X1 U5806 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n6363) );
  OAI222_X1 U5807 ( .A1(n6397), .A2(n5697), .B1(n4680), .B2(n5696), .C1(n6363), 
        .C2(n5694), .ZN(U2857) );
  AOI22_X1 U5808 ( .A1(n6328), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6324), .ZN(n4683) );
  NAND2_X1 U5809 ( .A1(n4683), .A2(n4682), .ZN(U2950) );
  AOI22_X1 U5810 ( .A1(n6328), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6324), .ZN(n4684) );
  NAND2_X1 U5811 ( .A1(n6327), .A2(DATAI_13_), .ZN(n4687) );
  NAND2_X1 U5812 ( .A1(n4684), .A2(n4687), .ZN(U2952) );
  AOI22_X1 U5813 ( .A1(n6328), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6324), .ZN(n4686) );
  NAND2_X1 U5814 ( .A1(n4686), .A2(n4685), .ZN(U2946) );
  AOI22_X1 U5815 ( .A1(n6328), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6324), .ZN(n4688) );
  NAND2_X1 U5816 ( .A1(n4688), .A2(n4687), .ZN(U2937) );
  AOI22_X1 U5817 ( .A1(n6328), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6324), .ZN(n4690) );
  NAND2_X1 U5818 ( .A1(n4690), .A2(n4689), .ZN(U2947) );
  XNOR2_X1 U5819 ( .A(n4692), .B(n4691), .ZN(n5010) );
  OR2_X1 U5820 ( .A1(n4677), .A2(n4693), .ZN(n4701) );
  INV_X1 U5821 ( .A(n4701), .ZN(n4694) );
  AOI21_X1 U5822 ( .B1(n4693), .B2(n4677), .A(n4694), .ZN(n5610) );
  AND2_X1 U5823 ( .A1(n6377), .A2(REIP_REG_3__SCAN_IN), .ZN(n5007) );
  AOI21_X1 U5824 ( .B1(n6358), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5007), 
        .ZN(n4695) );
  OAI21_X1 U5825 ( .B1(n5624), .B2(n6370), .A(n4695), .ZN(n4696) );
  AOI21_X1 U5826 ( .B1(n5610), .B2(n6365), .A(n4696), .ZN(n4697) );
  OAI21_X1 U5827 ( .B1(n5010), .B2(n6339), .A(n4697), .ZN(U2983) );
  INV_X1 U5828 ( .A(DATAI_2_), .ZN(n4852) );
  AOI22_X1 U5829 ( .A1(n6328), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6324), .ZN(n4698) );
  OAI21_X1 U5830 ( .B1(n4852), .B2(n4841), .A(n4698), .ZN(U2941) );
  INV_X1 U5831 ( .A(DATAI_5_), .ZN(n4847) );
  AOI22_X1 U5832 ( .A1(n6328), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6324), .ZN(n4699) );
  OAI21_X1 U5833 ( .B1(n4847), .B2(n4841), .A(n4699), .ZN(U2944) );
  AOI22_X1 U5834 ( .A1(n6328), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6324), .ZN(n4700) );
  OAI21_X1 U5835 ( .B1(n4644), .B2(n4841), .A(n4700), .ZN(U2942) );
  AND2_X1 U5836 ( .A1(n4702), .A2(n4701), .ZN(n4704) );
  OR2_X1 U5837 ( .A1(n4704), .A2(n4703), .ZN(n6261) );
  OR2_X1 U5838 ( .A1(n4772), .A2(n4706), .ZN(n4707) );
  NAND2_X1 U5839 ( .A1(n4705), .A2(n4707), .ZN(n6276) );
  INV_X1 U5840 ( .A(n6276), .ZN(n4708) );
  AOI22_X1 U5841 ( .A1(n4499), .A2(n4708), .B1(n5684), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4709) );
  OAI21_X1 U5842 ( .B1(n6261), .B2(n5694), .A(n4709), .ZN(U2855) );
  INV_X1 U5843 ( .A(n5645), .ZN(n4710) );
  OAI222_X1 U5844 ( .A1(n4710), .A2(n5697), .B1(n5696), .B2(n4195), .C1(n5652), 
        .C2(n5694), .ZN(U2859) );
  AND2_X1 U5845 ( .A1(n4711), .A2(n6461), .ZN(n6647) );
  NAND2_X1 U5846 ( .A1(n5612), .A2(n6583), .ZN(n5013) );
  INV_X1 U5847 ( .A(n5013), .ZN(n4719) );
  INV_X1 U5848 ( .A(n4715), .ZN(n4716) );
  NAND2_X1 U5849 ( .A1(n5625), .A2(n5637), .ZN(n6653) );
  INV_X1 U5850 ( .A(n6653), .ZN(n4718) );
  NAND2_X1 U5851 ( .A1(n6647), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4765) );
  INV_X1 U5852 ( .A(n4765), .ZN(n4717) );
  AOI21_X1 U5853 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4728) );
  NOR2_X1 U5854 ( .A1(n4728), .A2(n6651), .ZN(n4720) );
  AOI21_X1 U5855 ( .B1(n6647), .B2(STATE2_REG_2__SCAN_IN), .A(n4720), .ZN(
        n4771) );
  INV_X1 U5856 ( .A(n4890), .ZN(n6156) );
  INV_X1 U5857 ( .A(n6795), .ZN(n6713) );
  NAND2_X1 U5858 ( .A1(n6156), .A2(n6713), .ZN(n4721) );
  INV_X1 U5859 ( .A(DATAI_21_), .ZN(n4723) );
  NOR2_X2 U5860 ( .A1(n6334), .A2(n4723), .ZN(n6692) );
  OR2_X1 U5861 ( .A1(n4727), .A2(n5137), .ZN(n6650) );
  NAND2_X1 U5862 ( .A1(n6365), .A2(DATAI_29_), .ZN(n6695) );
  OR2_X1 U5863 ( .A1(n4764), .A2(n3337), .ZN(n6523) );
  OAI22_X1 U5864 ( .A1(n6650), .A2(n6695), .B1(n6523), .B2(n4765), .ZN(n4726)
         );
  AOI21_X1 U5865 ( .B1(n6692), .B2(n4767), .A(n4726), .ZN(n4731) );
  NAND3_X1 U5866 ( .A1(n4814), .A2(n6586), .A3(n4728), .ZN(n4729) );
  NAND2_X1 U5867 ( .A1(n4768), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4730)
         );
  OAI211_X1 U5868 ( .C1(n4771), .C2(n6568), .A(n4731), .B(n4730), .ZN(U3129)
         );
  INV_X1 U5869 ( .A(DATAI_19_), .ZN(n4732) );
  NOR2_X1 U5870 ( .A1(n6334), .A2(n4732), .ZN(n6680) );
  INV_X1 U5871 ( .A(DATAI_27_), .ZN(n6912) );
  NOR2_X1 U5872 ( .A1(n6334), .A2(n6912), .ZN(n6609) );
  OAI22_X1 U5873 ( .A1(n6650), .A2(n6683), .B1(n6606), .B2(n4765), .ZN(n4734)
         );
  AOI21_X1 U5874 ( .B1(n6680), .B2(n4767), .A(n4734), .ZN(n4736) );
  NAND2_X1 U5875 ( .A1(n4768), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4735)
         );
  OAI211_X1 U5876 ( .C1(n4771), .C2(n6562), .A(n4736), .B(n4735), .ZN(U3127)
         );
  INV_X1 U5877 ( .A(DATAI_7_), .ZN(n7079) );
  INV_X1 U5878 ( .A(DATAI_23_), .ZN(n4737) );
  NAND2_X1 U5879 ( .A1(n6365), .A2(DATAI_31_), .ZN(n6712) );
  OAI22_X1 U5880 ( .A1(n6650), .A2(n6712), .B1(n6633), .B2(n4765), .ZN(n4738)
         );
  AOI21_X1 U5881 ( .B1(n6707), .B2(n4767), .A(n4738), .ZN(n4740) );
  NAND2_X1 U5882 ( .A1(n4768), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4739)
         );
  OAI211_X1 U5883 ( .C1(n4771), .C2(n6580), .A(n4740), .B(n4739), .ZN(U3131)
         );
  INV_X1 U5884 ( .A(DATAI_22_), .ZN(n4741) );
  NOR2_X1 U5885 ( .A1(n6334), .A2(n4741), .ZN(n6698) );
  INV_X1 U5886 ( .A(DATAI_30_), .ZN(n4742) );
  NOR2_X1 U5887 ( .A1(n6334), .A2(n4742), .ZN(n6628) );
  INV_X1 U5888 ( .A(n6628), .ZN(n6701) );
  OAI22_X1 U5889 ( .A1(n6650), .A2(n6701), .B1(n6625), .B2(n4765), .ZN(n4743)
         );
  AOI21_X1 U5890 ( .B1(n6698), .B2(n4767), .A(n4743), .ZN(n4745) );
  NAND2_X1 U5891 ( .A1(n4768), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4744)
         );
  OAI211_X1 U5892 ( .C1(n4771), .C2(n6574), .A(n4745), .B(n4744), .ZN(U3130)
         );
  INV_X1 U5893 ( .A(DATAI_16_), .ZN(n4746) );
  NOR2_X2 U5894 ( .A1(n6334), .A2(n4746), .ZN(n6662) );
  INV_X1 U5895 ( .A(DATAI_24_), .ZN(n4747) );
  NOR2_X1 U5896 ( .A1(n6334), .A2(n4747), .ZN(n6589) );
  INV_X1 U5897 ( .A(n6589), .ZN(n6665) );
  OAI22_X1 U5898 ( .A1(n6650), .A2(n6665), .B1(n6544), .B2(n4765), .ZN(n4749)
         );
  AOI21_X1 U5899 ( .B1(n6662), .B2(n4767), .A(n4749), .ZN(n4751) );
  NAND2_X1 U5900 ( .A1(n4768), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4750)
         );
  OAI211_X1 U5901 ( .C1(n4771), .C2(n6553), .A(n4751), .B(n4750), .ZN(U3124)
         );
  INV_X1 U5902 ( .A(DATAI_18_), .ZN(n4752) );
  NOR2_X2 U5903 ( .A1(n6334), .A2(n4752), .ZN(n6674) );
  NAND2_X1 U5904 ( .A1(n6365), .A2(DATAI_26_), .ZN(n6677) );
  OAI22_X1 U5905 ( .A1(n6650), .A2(n6677), .B1(n7112), .B2(n4765), .ZN(n4754)
         );
  AOI21_X1 U5906 ( .B1(n6674), .B2(n4767), .A(n4754), .ZN(n4756) );
  NAND2_X1 U5907 ( .A1(n4768), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4755)
         );
  OAI211_X1 U5908 ( .C1(n4771), .C2(n7113), .A(n4756), .B(n4755), .ZN(U3126)
         );
  INV_X1 U5909 ( .A(DATAI_17_), .ZN(n4757) );
  NOR2_X2 U5910 ( .A1(n6334), .A2(n4757), .ZN(n6668) );
  NAND2_X1 U5911 ( .A1(n6365), .A2(DATAI_25_), .ZN(n6671) );
  OAI22_X1 U5912 ( .A1(n6650), .A2(n6671), .B1(n6507), .B2(n4765), .ZN(n4759)
         );
  AOI21_X1 U5913 ( .B1(n6668), .B2(n4767), .A(n4759), .ZN(n4761) );
  NAND2_X1 U5914 ( .A1(n4768), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4760)
         );
  OAI211_X1 U5915 ( .C1(n4771), .C2(n6556), .A(n4761), .B(n4760), .ZN(U3125)
         );
  INV_X1 U5916 ( .A(DATAI_20_), .ZN(n4762) );
  NAND2_X1 U5917 ( .A1(n6365), .A2(DATAI_28_), .ZN(n6689) );
  OAI22_X1 U5918 ( .A1(n6650), .A2(n6689), .B1(n6613), .B2(n4765), .ZN(n4766)
         );
  AOI21_X1 U5919 ( .B1(n6686), .B2(n4767), .A(n4766), .ZN(n4770) );
  NAND2_X1 U5920 ( .A1(n4768), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4769)
         );
  OAI211_X1 U5921 ( .C1(n4771), .C2(n6565), .A(n4770), .B(n4769), .ZN(U3128)
         );
  AOI21_X1 U5922 ( .B1(n4774), .B2(n4773), .A(n4772), .ZN(n5621) );
  INV_X1 U5923 ( .A(n5621), .ZN(n4775) );
  INV_X1 U5924 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5614) );
  INV_X1 U5925 ( .A(n5610), .ZN(n4851) );
  OAI222_X1 U5926 ( .A1(n4775), .A2(n5697), .B1(n5614), .B2(n5696), .C1(n4851), 
        .C2(n5694), .ZN(U2856) );
  INV_X1 U5927 ( .A(n4776), .ZN(n4811) );
  INV_X1 U5928 ( .A(n6117), .ZN(n4799) );
  XNOR2_X1 U5929 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4779) );
  XNOR2_X1 U5930 ( .A(n4777), .B(n5334), .ZN(n4782) );
  INV_X1 U5931 ( .A(n4782), .ZN(n4778) );
  OAI22_X1 U5932 ( .A1(n4799), .A2(n4779), .B1(n4793), .B2(n4778), .ZN(n4784)
         );
  AND2_X1 U5933 ( .A1(n4781), .A2(n4780), .ZN(n4787) );
  NOR2_X1 U5934 ( .A1(n4787), .A2(n4782), .ZN(n4783) );
  AOI211_X1 U5935 ( .C1(n5625), .C2(n4802), .A(n4784), .B(n4783), .ZN(n5326)
         );
  MUX2_X1 U5936 ( .A(n5326), .B(n5334), .S(n6121), .Z(n6126) );
  INV_X1 U5937 ( .A(n6126), .ZN(n6128) );
  NAND2_X1 U5938 ( .A1(n6128), .A2(n6810), .ZN(n4807) );
  NAND2_X1 U5939 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4786) );
  INV_X1 U5940 ( .A(n4786), .ZN(n4785) );
  MUX2_X1 U5941 ( .A(n4786), .B(n4785), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4800) );
  INV_X1 U5942 ( .A(n4787), .ZN(n4792) );
  MUX2_X1 U5943 ( .A(n4788), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4777), 
        .Z(n4790) );
  NOR2_X1 U5944 ( .A1(n4790), .A2(n4789), .ZN(n4791) );
  NAND2_X1 U5945 ( .A1(n4792), .A2(n4791), .ZN(n4798) );
  INV_X1 U5946 ( .A(n4793), .ZN(n4796) );
  NOR2_X1 U5947 ( .A1(n4777), .A2(n4804), .ZN(n4794) );
  NOR2_X1 U5948 ( .A1(n4794), .A2(n3297), .ZN(n4795) );
  NAND2_X1 U5949 ( .A1(n3462), .A2(n4795), .ZN(n6111) );
  NAND2_X1 U5950 ( .A1(n4796), .A2(n6111), .ZN(n4797) );
  OAI211_X1 U5951 ( .C1(n4800), .C2(n4799), .A(n4798), .B(n4797), .ZN(n4801)
         );
  AOI21_X1 U5952 ( .B1(n5612), .B2(n4802), .A(n4801), .ZN(n6114) );
  INV_X1 U5953 ( .A(n6121), .ZN(n4803) );
  MUX2_X1 U5954 ( .A(n4804), .B(n6114), .S(n4803), .Z(n6130) );
  INV_X1 U5955 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6164) );
  NAND2_X1 U5956 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6164), .ZN(n4806) );
  INV_X1 U5957 ( .A(n4789), .ZN(n4805) );
  OAI22_X1 U5958 ( .A1(n4807), .A2(n6130), .B1(n4806), .B2(n4805), .ZN(n6137)
         );
  MUX2_X1 U5959 ( .A(n6164), .B(n6121), .S(n6810), .Z(n4809) );
  AOI21_X1 U5960 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4809), .A(n4808), 
        .ZN(n6135) );
  INV_X1 U5961 ( .A(n6135), .ZN(n4810) );
  AOI21_X1 U5962 ( .B1(n4811), .B2(n6137), .A(n4810), .ZN(n6149) );
  AND2_X1 U5963 ( .A1(n6149), .A2(n6164), .ZN(n4812) );
  INV_X1 U5964 ( .A(n6779), .ZN(n6714) );
  AND2_X1 U5965 ( .A1(n4814), .A2(n6596), .ZN(n6427) );
  INV_X1 U5966 ( .A(n4724), .ZN(n4815) );
  NAND2_X1 U5967 ( .A1(n3097), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6582) );
  INV_X1 U5968 ( .A(n6582), .ZN(n6425) );
  NAND2_X1 U5969 ( .A1(n3111), .A2(n6425), .ZN(n6548) );
  AOI21_X1 U5970 ( .B1(n6427), .B2(n6548), .A(n6651), .ZN(n4819) );
  INV_X1 U5971 ( .A(n5612), .ZN(n5192) );
  NAND2_X1 U5972 ( .A1(n4816), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4896) );
  INV_X1 U5973 ( .A(n4896), .ZN(n4817) );
  OAI22_X1 U5974 ( .A1(n3185), .A2(n5190), .B1(n5192), .B2(n4817), .ZN(n4818)
         );
  OAI21_X1 U5975 ( .B1(n4819), .B2(n4818), .A(n6419), .ZN(n4820) );
  OAI21_X1 U5976 ( .B1(n6419), .B2(n6462), .A(n4820), .ZN(U3462) );
  OR2_X1 U5977 ( .A1(n4703), .A2(n4822), .ZN(n4823) );
  AND2_X1 U5978 ( .A1(n4821), .A2(n4823), .ZN(n6352) );
  INV_X1 U5979 ( .A(n6352), .ZN(n4848) );
  INV_X1 U5980 ( .A(n4953), .ZN(n4825) );
  AOI21_X1 U5981 ( .B1(n4826), .B2(n4705), .A(n4825), .ZN(n6251) );
  AOI22_X1 U5982 ( .A1(n6251), .A2(n4499), .B1(EBX_REG_5__SCAN_IN), .B2(n5684), 
        .ZN(n4827) );
  OAI21_X1 U5983 ( .B1(n4848), .B2(n5694), .A(n4827), .ZN(U2854) );
  OR2_X1 U5984 ( .A1(n4829), .A2(n4828), .ZN(n4831) );
  AND2_X1 U5985 ( .A1(n4831), .A2(n4830), .ZN(n6411) );
  NAND2_X1 U5986 ( .A1(n6350), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5987 ( .A1(n6377), .A2(REIP_REG_1__SCAN_IN), .ZN(n6406) );
  OAI211_X1 U5988 ( .C1(n6356), .C2(n4833), .A(n4832), .B(n6406), .ZN(n4834)
         );
  AOI21_X1 U5989 ( .B1(n6366), .B2(n6411), .A(n4834), .ZN(n4835) );
  OAI21_X1 U5990 ( .B1(n6334), .B2(n5642), .A(n4835), .ZN(U2985) );
  NOR2_X1 U5991 ( .A1(n4837), .A2(n4836), .ZN(n4838) );
  AND2_X1 U5992 ( .A1(n4843), .A2(n4842), .ZN(n4844) );
  INV_X1 U5993 ( .A(n4844), .ZN(n4845) );
  OAI222_X1 U5994 ( .A1(n5642), .A2(n5747), .B1(n5744), .B2(n4846), .C1(n5746), 
        .C2(n4648), .ZN(U2890) );
  INV_X1 U5995 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6295) );
  OAI222_X1 U5996 ( .A1(n4848), .A2(n5747), .B1(n5744), .B2(n4847), .C1(n5746), 
        .C2(n6295), .ZN(U2886) );
  OAI222_X1 U5997 ( .A1(n6261), .A2(n5747), .B1(n5744), .B2(n4849), .C1(n6297), 
        .C2(n5746), .ZN(U2887) );
  INV_X1 U5998 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4850) );
  OAI222_X1 U5999 ( .A1(n4851), .A2(n5747), .B1(n5744), .B2(n4644), .C1(n5746), 
        .C2(n4850), .ZN(U2888) );
  INV_X1 U6000 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6952) );
  OAI222_X1 U6001 ( .A1(n6363), .A2(n5747), .B1(n5744), .B2(n4852), .C1(n5746), 
        .C2(n6952), .ZN(U2889) );
  OAI222_X1 U6002 ( .A1(n5652), .A2(n5747), .B1(n5746), .B2(n4854), .C1(n5744), 
        .C2(n4853), .ZN(U2891) );
  AND2_X1 U6003 ( .A1(n3097), .A2(n6473), .ZN(n5254) );
  INV_X1 U6004 ( .A(n5254), .ZN(n5189) );
  AOI21_X1 U6005 ( .B1(n4889), .B2(n4932), .A(n6467), .ZN(n4859) );
  NAND2_X1 U6006 ( .A1(n4957), .A2(n5625), .ZN(n5146) );
  OR2_X1 U6007 ( .A1(n5612), .A2(n6651), .ZN(n6466) );
  INV_X1 U6008 ( .A(n6466), .ZN(n5072) );
  AOI21_X1 U6009 ( .B1(n6586), .B2(n5146), .A(n5072), .ZN(n4858) );
  NAND2_X1 U6010 ( .A1(n4908), .A2(n7028), .ZN(n4884) );
  AND2_X1 U6011 ( .A1(n4860), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6658) );
  NOR2_X1 U6012 ( .A1(n5144), .A2(n6592), .ZN(n4855) );
  NOR2_X1 U6013 ( .A1(n5053), .A2(n4855), .ZN(n5140) );
  NAND2_X1 U6014 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6462), .ZN(n4856) );
  NAND2_X1 U6015 ( .A1(n5140), .A2(n4856), .ZN(n5261) );
  AOI211_X1 U6016 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4884), .A(n6658), .B(
        n5261), .ZN(n4857) );
  NAND2_X1 U6017 ( .A1(n4883), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4864)
         );
  NOR2_X1 U6018 ( .A1(n5192), .A2(n6651), .ZN(n6642) );
  INV_X1 U6019 ( .A(n5146), .ZN(n6542) );
  NOR2_X1 U6020 ( .A1(n4860), .A2(n6592), .ZN(n6463) );
  INV_X1 U6021 ( .A(n5144), .ZN(n4861) );
  NOR2_X1 U6022 ( .A1(n4861), .A2(n6462), .ZN(n5258) );
  AOI22_X1 U6023 ( .A1(n6642), .A2(n6542), .B1(n6463), .B2(n5258), .ZN(n4885)
         );
  OAI22_X1 U6024 ( .A1(n4885), .A2(n6562), .B1(n6606), .B2(n4884), .ZN(n4862)
         );
  AOI21_X1 U6025 ( .B1(n6680), .B2(n4948), .A(n4862), .ZN(n4863) );
  OAI211_X1 U6026 ( .C1(n4889), .C2(n6683), .A(n4864), .B(n4863), .ZN(U3135)
         );
  NAND2_X1 U6027 ( .A1(n4883), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4867)
         );
  OAI22_X1 U6028 ( .A1(n4885), .A2(n6574), .B1(n6625), .B2(n4884), .ZN(n4865)
         );
  AOI21_X1 U6029 ( .B1(n6698), .B2(n4948), .A(n4865), .ZN(n4866) );
  OAI211_X1 U6030 ( .C1(n4889), .C2(n6701), .A(n4867), .B(n4866), .ZN(U3138)
         );
  NAND2_X1 U6031 ( .A1(n4883), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4870)
         );
  OAI22_X1 U6032 ( .A1(n4885), .A2(n6580), .B1(n6633), .B2(n4884), .ZN(n4868)
         );
  AOI21_X1 U6033 ( .B1(n6707), .B2(n4948), .A(n4868), .ZN(n4869) );
  OAI211_X1 U6034 ( .C1(n4889), .C2(n6712), .A(n4870), .B(n4869), .ZN(U3139)
         );
  NAND2_X1 U6035 ( .A1(n4883), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4873)
         );
  OAI22_X1 U6036 ( .A1(n4885), .A2(n6565), .B1(n6613), .B2(n4884), .ZN(n4871)
         );
  AOI21_X1 U6037 ( .B1(n6686), .B2(n4948), .A(n4871), .ZN(n4872) );
  OAI211_X1 U6038 ( .C1(n4889), .C2(n6689), .A(n4873), .B(n4872), .ZN(U3136)
         );
  NAND2_X1 U6039 ( .A1(n4883), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4876)
         );
  OAI22_X1 U6040 ( .A1(n4885), .A2(n7113), .B1(n7112), .B2(n4884), .ZN(n4874)
         );
  AOI21_X1 U6041 ( .B1(n6674), .B2(n4948), .A(n4874), .ZN(n4875) );
  OAI211_X1 U6042 ( .C1(n4889), .C2(n6677), .A(n4876), .B(n4875), .ZN(U3134)
         );
  NAND2_X1 U6043 ( .A1(n4883), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4879)
         );
  OAI22_X1 U6044 ( .A1(n4885), .A2(n6568), .B1(n6523), .B2(n4884), .ZN(n4877)
         );
  AOI21_X1 U6045 ( .B1(n6692), .B2(n4948), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6046 ( .C1(n4889), .C2(n6695), .A(n4879), .B(n4878), .ZN(U3137)
         );
  NAND2_X1 U6047 ( .A1(n4883), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4882)
         );
  OAI22_X1 U6048 ( .A1(n4885), .A2(n6556), .B1(n6507), .B2(n4884), .ZN(n4880)
         );
  AOI21_X1 U6049 ( .B1(n6668), .B2(n4948), .A(n4880), .ZN(n4881) );
  OAI211_X1 U6050 ( .C1(n4889), .C2(n6671), .A(n4882), .B(n4881), .ZN(U3133)
         );
  NAND2_X1 U6051 ( .A1(n4883), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4888)
         );
  OAI22_X1 U6052 ( .A1(n4885), .A2(n6553), .B1(n6544), .B2(n4884), .ZN(n4886)
         );
  AOI21_X1 U6053 ( .B1(n6662), .B2(n4948), .A(n4886), .ZN(n4887) );
  OAI211_X1 U6054 ( .C1(n4889), .C2(n6665), .A(n4888), .B(n4887), .ZN(U3132)
         );
  AOI222_X1 U6055 ( .A1(n4896), .A2(n6583), .B1(n4890), .B2(n6149), .C1(n5137), 
        .C2(n6586), .ZN(n4892) );
  NAND2_X1 U6056 ( .A1(n4900), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4891) );
  OAI21_X1 U6057 ( .B1(n4892), .B2(n4900), .A(n4891), .ZN(U3465) );
  AOI22_X1 U6058 ( .A1(n4893), .A2(n6586), .B1(n5625), .B2(n4896), .ZN(n4895)
         );
  NAND2_X1 U6059 ( .A1(n4900), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4894) );
  OAI21_X1 U6060 ( .B1(n4900), .B2(n4895), .A(n4894), .ZN(U3463) );
  INV_X1 U6061 ( .A(n3097), .ZN(n5136) );
  AOI21_X1 U6062 ( .B1(n5136), .B2(n6467), .A(n6651), .ZN(n4897) );
  AOI22_X1 U6063 ( .A1(n4897), .A2(n6582), .B1(n4957), .B2(n4896), .ZN(n4899)
         );
  NAND2_X1 U6064 ( .A1(n4900), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4898) );
  OAI21_X1 U6065 ( .B1(n4900), .B2(n4899), .A(n4898), .ZN(U3464) );
  INV_X1 U6066 ( .A(n4908), .ZN(n4905) );
  INV_X1 U6067 ( .A(n6585), .ZN(n4904) );
  OAI21_X1 U6068 ( .B1(n4906), .B2(n5136), .A(n6365), .ZN(n4902) );
  OR2_X1 U6069 ( .A1(n5013), .A2(n5146), .ZN(n4901) );
  NAND2_X1 U6070 ( .A1(n4901), .A2(n4911), .ZN(n4907) );
  AOI21_X1 U6071 ( .B1(n4902), .B2(n5190), .A(n4907), .ZN(n4903) );
  AOI211_X1 U6072 ( .C1(n4905), .C2(n6651), .A(n4904), .B(n4903), .ZN(n4945)
         );
  INV_X1 U6073 ( .A(n4945), .ZN(n4936) );
  NOR2_X1 U6074 ( .A1(n4932), .A2(n6677), .ZN(n4914) );
  INV_X1 U6075 ( .A(n6674), .ZN(n7120) );
  NAND2_X1 U6076 ( .A1(n3097), .A2(n5137), .ZN(n6595) );
  NAND2_X1 U6077 ( .A1(n4907), .A2(n6586), .ZN(n4910) );
  NAND2_X1 U6078 ( .A1(n4908), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U6079 ( .A1(n4910), .A2(n4909), .ZN(n4943) );
  INV_X1 U6080 ( .A(n4911), .ZN(n4942) );
  AOI22_X1 U6081 ( .A1(n4943), .A2(n6673), .B1(n6672), .B2(n4942), .ZN(n4912)
         );
  OAI21_X1 U6082 ( .B1(n7120), .B2(n5127), .A(n4912), .ZN(n4913) );
  AOI211_X1 U6083 ( .C1(n4936), .C2(INSTQUEUE_REG_15__2__SCAN_IN), .A(n4914), 
        .B(n4913), .ZN(n4915) );
  INV_X1 U6084 ( .A(n4915), .ZN(U3142) );
  NOR2_X1 U6085 ( .A1(n4932), .A2(n6683), .ZN(n4918) );
  INV_X1 U6086 ( .A(n6680), .ZN(n6607) );
  INV_X1 U6087 ( .A(n6606), .ZN(n6678) );
  AOI22_X1 U6088 ( .A1(n4943), .A2(n6679), .B1(n6678), .B2(n4942), .ZN(n4916)
         );
  OAI21_X1 U6089 ( .B1(n6607), .B2(n5127), .A(n4916), .ZN(n4917) );
  AOI211_X1 U6090 ( .C1(n4936), .C2(INSTQUEUE_REG_15__3__SCAN_IN), .A(n4918), 
        .B(n4917), .ZN(n4919) );
  INV_X1 U6091 ( .A(n4919), .ZN(U3143) );
  NOR2_X1 U6092 ( .A1(n4932), .A2(n6712), .ZN(n4922) );
  INV_X1 U6093 ( .A(n6707), .ZN(n6634) );
  AOI22_X1 U6094 ( .A1(n4943), .A2(n6704), .B1(n6703), .B2(n4942), .ZN(n4920)
         );
  OAI21_X1 U6095 ( .B1(n6634), .B2(n5127), .A(n4920), .ZN(n4921) );
  AOI211_X1 U6096 ( .C1(n4936), .C2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4922), 
        .B(n4921), .ZN(n4923) );
  INV_X1 U6097 ( .A(n4923), .ZN(U3147) );
  NOR2_X1 U6098 ( .A1(n4932), .A2(n6695), .ZN(n4926) );
  INV_X1 U6099 ( .A(n6692), .ZN(n5266) );
  AOI22_X1 U6100 ( .A1(n4943), .A2(n6691), .B1(n6690), .B2(n4942), .ZN(n4924)
         );
  OAI21_X1 U6101 ( .B1(n5266), .B2(n5127), .A(n4924), .ZN(n4925) );
  AOI211_X1 U6102 ( .C1(n4936), .C2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4926), 
        .B(n4925), .ZN(n4927) );
  INV_X1 U6103 ( .A(n4927), .ZN(U3145) );
  NOR2_X1 U6104 ( .A1(n4932), .A2(n6689), .ZN(n4930) );
  INV_X1 U6105 ( .A(n6686), .ZN(n6614) );
  AOI22_X1 U6106 ( .A1(n4943), .A2(n6685), .B1(n6684), .B2(n4942), .ZN(n4928)
         );
  OAI21_X1 U6107 ( .B1(n6614), .B2(n5127), .A(n4928), .ZN(n4929) );
  AOI211_X1 U6108 ( .C1(n4936), .C2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n4930), 
        .B(n4929), .ZN(n4931) );
  INV_X1 U6109 ( .A(n4931), .ZN(U3144) );
  NOR2_X1 U6110 ( .A1(n4932), .A2(n6701), .ZN(n4935) );
  INV_X1 U6111 ( .A(n6698), .ZN(n6626) );
  INV_X1 U6112 ( .A(n6625), .ZN(n6696) );
  AOI22_X1 U6113 ( .A1(n4943), .A2(n6697), .B1(n6696), .B2(n4942), .ZN(n4933)
         );
  OAI21_X1 U6114 ( .B1(n6626), .B2(n5127), .A(n4933), .ZN(n4934) );
  AOI211_X1 U6115 ( .C1(n4936), .C2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4935), 
        .B(n4934), .ZN(n4937) );
  INV_X1 U6116 ( .A(n4937), .ZN(U3146) );
  INV_X1 U6117 ( .A(n6662), .ZN(n6545) );
  INV_X1 U6118 ( .A(n6544), .ZN(n6648) );
  AOI22_X1 U6119 ( .A1(n4943), .A2(n6649), .B1(n6648), .B2(n4942), .ZN(n4938)
         );
  OAI21_X1 U6120 ( .B1(n6545), .B2(n5127), .A(n4938), .ZN(n4940) );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n7091) );
  NOR2_X1 U6122 ( .A1(n4945), .A2(n7091), .ZN(n4939) );
  AOI211_X1 U6123 ( .C1(n4948), .C2(n6589), .A(n4940), .B(n4939), .ZN(n4941)
         );
  INV_X1 U6124 ( .A(n4941), .ZN(U3140) );
  INV_X1 U6125 ( .A(n6671), .ZN(n6599) );
  INV_X1 U6126 ( .A(n6668), .ZN(n5279) );
  AOI22_X1 U6127 ( .A1(n4943), .A2(n6667), .B1(n6666), .B2(n4942), .ZN(n4944)
         );
  OAI21_X1 U6128 ( .B1(n5279), .B2(n5127), .A(n4944), .ZN(n4947) );
  INV_X1 U6129 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U6130 ( .A1(n4945), .A2(n6876), .ZN(n4946) );
  AOI211_X1 U6131 ( .C1(n4948), .C2(n6599), .A(n4947), .B(n4946), .ZN(n4949)
         );
  INV_X1 U6132 ( .A(n4949), .ZN(U3141) );
  OAI21_X1 U6133 ( .B1(n3191), .B2(n4951), .A(n4950), .ZN(n5607) );
  AOI21_X1 U6134 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(n5601) );
  AOI22_X1 U6135 ( .A1(n5601), .A2(n4499), .B1(n5684), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4955) );
  OAI21_X1 U6136 ( .B1(n5607), .B2(n5694), .A(n4955), .ZN(U2853) );
  OAI222_X1 U6137 ( .A1(n5607), .A2(n5747), .B1(n5744), .B2(n4956), .C1(n5746), 
        .C2(n4650), .ZN(U2885) );
  INV_X1 U6138 ( .A(n4960), .ZN(n4961) );
  OAI21_X1 U6139 ( .B1(n4961), .B2(n6651), .A(n5190), .ZN(n4963) );
  OR2_X1 U6140 ( .A1(n5612), .A2(n6496), .ZN(n4958) );
  NOR2_X1 U6141 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6142 ( .A1(n5012), .A2(n6462), .ZN(n5052) );
  OR2_X1 U6143 ( .A1(n5052), .A2(n7028), .ZN(n4987) );
  OAI21_X1 U6144 ( .B1(n4958), .B2(n5057), .A(n4987), .ZN(n4965) );
  INV_X1 U6145 ( .A(n5052), .ZN(n4959) );
  NOR2_X1 U6146 ( .A1(n4960), .A2(n6473), .ZN(n5191) );
  OAI22_X1 U6147 ( .A1(n5131), .A2(n6712), .B1(n6633), .B2(n4987), .ZN(n4962)
         );
  AOI21_X1 U6148 ( .B1(n6707), .B2(n5191), .A(n4962), .ZN(n4968) );
  INV_X1 U6149 ( .A(n4963), .ZN(n4966) );
  NAND2_X1 U6150 ( .A1(n5052), .A2(n6651), .ZN(n4964) );
  NAND2_X1 U6151 ( .A1(n4989), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4967) );
  OAI211_X1 U6152 ( .C1(n4992), .C2(n6580), .A(n4968), .B(n4967), .ZN(U3035)
         );
  OAI22_X1 U6153 ( .A1(n5131), .A2(n6683), .B1(n6606), .B2(n4987), .ZN(n4969)
         );
  AOI21_X1 U6154 ( .B1(n6680), .B2(n5191), .A(n4969), .ZN(n4971) );
  NAND2_X1 U6155 ( .A1(n4989), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4970) );
  OAI211_X1 U6156 ( .C1(n4992), .C2(n6562), .A(n4971), .B(n4970), .ZN(U3031)
         );
  OAI22_X1 U6157 ( .A1(n5131), .A2(n6689), .B1(n6613), .B2(n4987), .ZN(n4972)
         );
  AOI21_X1 U6158 ( .B1(n6686), .B2(n5191), .A(n4972), .ZN(n4974) );
  NAND2_X1 U6159 ( .A1(n4989), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4973) );
  OAI211_X1 U6160 ( .C1(n4992), .C2(n6565), .A(n4974), .B(n4973), .ZN(U3032)
         );
  OAI22_X1 U6161 ( .A1(n5131), .A2(n6665), .B1(n6544), .B2(n4987), .ZN(n4975)
         );
  AOI21_X1 U6162 ( .B1(n6662), .B2(n5191), .A(n4975), .ZN(n4977) );
  NAND2_X1 U6163 ( .A1(n4989), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4976) );
  OAI211_X1 U6164 ( .C1(n4992), .C2(n6553), .A(n4977), .B(n4976), .ZN(U3028)
         );
  OAI22_X1 U6165 ( .A1(n5131), .A2(n6701), .B1(n6625), .B2(n4987), .ZN(n4978)
         );
  AOI21_X1 U6166 ( .B1(n6698), .B2(n5191), .A(n4978), .ZN(n4980) );
  NAND2_X1 U6167 ( .A1(n4989), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4979) );
  OAI211_X1 U6168 ( .C1(n4992), .C2(n6574), .A(n4980), .B(n4979), .ZN(U3034)
         );
  OAI22_X1 U6169 ( .A1(n5131), .A2(n6695), .B1(n6523), .B2(n4987), .ZN(n4981)
         );
  AOI21_X1 U6170 ( .B1(n6692), .B2(n5191), .A(n4981), .ZN(n4983) );
  NAND2_X1 U6171 ( .A1(n4989), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4982) );
  OAI211_X1 U6172 ( .C1(n4992), .C2(n6568), .A(n4983), .B(n4982), .ZN(U3033)
         );
  OAI22_X1 U6173 ( .A1(n5131), .A2(n6671), .B1(n6507), .B2(n4987), .ZN(n4984)
         );
  AOI21_X1 U6174 ( .B1(n6668), .B2(n5191), .A(n4984), .ZN(n4986) );
  NAND2_X1 U6175 ( .A1(n4989), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4985) );
  OAI211_X1 U6176 ( .C1(n4992), .C2(n6556), .A(n4986), .B(n4985), .ZN(U3029)
         );
  OAI22_X1 U6177 ( .A1(n5131), .A2(n6677), .B1(n7112), .B2(n4987), .ZN(n4988)
         );
  AOI21_X1 U6178 ( .B1(n6674), .B2(n5191), .A(n4988), .ZN(n4991) );
  NAND2_X1 U6179 ( .A1(n4989), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4990) );
  OAI211_X1 U6180 ( .C1(n4992), .C2(n7113), .A(n4991), .B(n4990), .ZN(U3030)
         );
  XNOR2_X1 U6181 ( .A(n4993), .B(n4994), .ZN(n6348) );
  INV_X1 U6182 ( .A(n6037), .ZN(n5298) );
  NOR2_X1 U6183 ( .A1(n6404), .A2(n4189), .ZN(n5005) );
  OAI22_X1 U6184 ( .A1(n5298), .A2(n5005), .B1(n6395), .B2(n6407), .ZN(n5003)
         );
  OR2_X1 U6185 ( .A1(n4378), .A2(n5299), .ZN(n5238) );
  AND2_X1 U6186 ( .A1(n6415), .A2(n5238), .ZN(n4995) );
  OR2_X1 U6187 ( .A1(n5003), .A2(n4995), .ZN(n5237) );
  INV_X1 U6188 ( .A(n6392), .ZN(n4997) );
  OAI211_X1 U6189 ( .C1(n4998), .C2(n4997), .A(n4996), .B(n4378), .ZN(n4999)
         );
  NAND2_X1 U6190 ( .A1(n5237), .A2(n4999), .ZN(n5002) );
  NAND2_X1 U6191 ( .A1(n6377), .A2(REIP_REG_5__SCAN_IN), .ZN(n6354) );
  INV_X1 U6192 ( .A(n6354), .ZN(n5000) );
  AOI21_X1 U6193 ( .B1(n6410), .B2(n6251), .A(n5000), .ZN(n5001) );
  OAI211_X1 U6194 ( .C1(n6101), .C2(n6348), .A(n5002), .B(n5001), .ZN(U3013)
         );
  INV_X1 U6195 ( .A(n5003), .ZN(n6403) );
  OAI21_X1 U6196 ( .B1(n5004), .B2(n6393), .A(n6403), .ZN(n6102) );
  INV_X1 U6197 ( .A(n6393), .ZN(n5006) );
  AOI21_X1 U6198 ( .B1(n5005), .B2(n6392), .A(n6395), .ZN(n5300) );
  NOR2_X1 U6199 ( .A1(n5006), .A2(n5300), .ZN(n6104) );
  AOI22_X1 U6200 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6102), .B1(n6104), 
        .B2(n4339), .ZN(n5009) );
  AOI21_X1 U6201 ( .B1(n6410), .B2(n5621), .A(n5007), .ZN(n5008) );
  OAI211_X1 U6202 ( .C1(n5010), .C2(n6101), .A(n5009), .B(n5008), .ZN(U3015)
         );
  INV_X1 U6203 ( .A(n5015), .ZN(n5011) );
  OAI21_X1 U6204 ( .B1(n5011), .B2(n6651), .A(n5190), .ZN(n5017) );
  NAND2_X1 U6205 ( .A1(n5012), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5073) );
  OR2_X1 U6206 ( .A1(n5073), .A2(n7028), .ZN(n5041) );
  OAI21_X1 U6207 ( .B1(n5013), .B2(n5057), .A(n5041), .ZN(n5019) );
  INV_X1 U6208 ( .A(n5073), .ZN(n5014) );
  OAI22_X1 U6209 ( .A1(n7121), .A2(n6695), .B1(n6523), .B2(n5041), .ZN(n5016)
         );
  AOI21_X1 U6210 ( .B1(n3109), .B2(n6692), .A(n5016), .ZN(n5022) );
  INV_X1 U6211 ( .A(n5017), .ZN(n5020) );
  NAND2_X1 U6212 ( .A1(n5073), .A2(n6651), .ZN(n5018) );
  NAND2_X1 U6213 ( .A1(n5043), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5021) );
  OAI211_X1 U6214 ( .C1(n5046), .C2(n6568), .A(n5022), .B(n5021), .ZN(U3097)
         );
  OAI22_X1 U6215 ( .A1(n7121), .A2(n6683), .B1(n6606), .B2(n5041), .ZN(n5023)
         );
  AOI21_X1 U6216 ( .B1(n3109), .B2(n6680), .A(n5023), .ZN(n5025) );
  NAND2_X1 U6217 ( .A1(n5043), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5024) );
  OAI211_X1 U6218 ( .C1(n5046), .C2(n6562), .A(n5025), .B(n5024), .ZN(U3095)
         );
  OAI22_X1 U6219 ( .A1(n7121), .A2(n6712), .B1(n6633), .B2(n5041), .ZN(n5026)
         );
  AOI21_X1 U6220 ( .B1(n3109), .B2(n6707), .A(n5026), .ZN(n5028) );
  NAND2_X1 U6221 ( .A1(n5043), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5027) );
  OAI211_X1 U6222 ( .C1(n5046), .C2(n6580), .A(n5028), .B(n5027), .ZN(U3099)
         );
  OAI22_X1 U6223 ( .A1(n7121), .A2(n6701), .B1(n6625), .B2(n5041), .ZN(n5029)
         );
  AOI21_X1 U6224 ( .B1(n3109), .B2(n6698), .A(n5029), .ZN(n5031) );
  NAND2_X1 U6225 ( .A1(n5043), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5030) );
  OAI211_X1 U6226 ( .C1(n5046), .C2(n6574), .A(n5031), .B(n5030), .ZN(U3098)
         );
  OAI22_X1 U6227 ( .A1(n7121), .A2(n6671), .B1(n6507), .B2(n5041), .ZN(n5032)
         );
  AOI21_X1 U6228 ( .B1(n3109), .B2(n6668), .A(n5032), .ZN(n5034) );
  NAND2_X1 U6229 ( .A1(n5043), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5033) );
  OAI211_X1 U6230 ( .C1(n5046), .C2(n6556), .A(n5034), .B(n5033), .ZN(U3093)
         );
  OAI22_X1 U6231 ( .A1(n7121), .A2(n6689), .B1(n6613), .B2(n5041), .ZN(n5035)
         );
  AOI21_X1 U6232 ( .B1(n3109), .B2(n6686), .A(n5035), .ZN(n5037) );
  NAND2_X1 U6233 ( .A1(n5043), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5036) );
  OAI211_X1 U6234 ( .C1(n5046), .C2(n6565), .A(n5037), .B(n5036), .ZN(U3096)
         );
  OAI22_X1 U6235 ( .A1(n7121), .A2(n6665), .B1(n6544), .B2(n5041), .ZN(n5038)
         );
  AOI21_X1 U6236 ( .B1(n3109), .B2(n6662), .A(n5038), .ZN(n5040) );
  NAND2_X1 U6237 ( .A1(n5043), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5039) );
  OAI211_X1 U6238 ( .C1(n5046), .C2(n6553), .A(n5040), .B(n5039), .ZN(U3092)
         );
  OAI22_X1 U6239 ( .A1(n7121), .A2(n6677), .B1(n7112), .B2(n5041), .ZN(n5042)
         );
  AOI21_X1 U6240 ( .B1(n3109), .B2(n6674), .A(n5042), .ZN(n5045) );
  NAND2_X1 U6241 ( .A1(n5043), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5044) );
  OAI211_X1 U6242 ( .C1(n5046), .C2(n7113), .A(n5045), .B(n5044), .ZN(U3094)
         );
  XOR2_X1 U6243 ( .A(n5047), .B(n5048), .Z(n6107) );
  NAND2_X1 U6244 ( .A1(n6107), .A2(n6366), .ZN(n5051) );
  INV_X1 U6245 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6727) );
  NOR2_X1 U6246 ( .A1(n6396), .A2(n6727), .ZN(n6106) );
  NOR2_X1 U6247 ( .A1(n6370), .A2(n6257), .ZN(n5049) );
  AOI211_X1 U6248 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6106), 
        .B(n5049), .ZN(n5050) );
  OAI211_X1 U6249 ( .C1(n6261), .C2(n6334), .A(n5051), .B(n5050), .ZN(U2982)
         );
  INV_X1 U6250 ( .A(n5057), .ZN(n5080) );
  NOR2_X1 U6251 ( .A1(n5080), .A2(n6651), .ZN(n5071) );
  OAI211_X1 U6252 ( .C1(n6642), .C2(n5071), .A(n5131), .B(n5127), .ZN(n5055)
         );
  INV_X1 U6253 ( .A(n5190), .ZN(n6655) );
  AOI21_X1 U6254 ( .B1(n5057), .B2(n6655), .A(n6463), .ZN(n5077) );
  OR2_X1 U6255 ( .A1(n5052), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5102)
         );
  INV_X1 U6256 ( .A(n5075), .ZN(n5079) );
  AOI21_X1 U6257 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5144), .A(n5053), .ZN(
        n5074) );
  OAI21_X1 U6258 ( .B1(n6592), .B2(n5079), .A(n5074), .ZN(n6469) );
  AOI21_X1 U6259 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5102), .A(n6469), .ZN(
        n5054) );
  NAND3_X1 U6260 ( .A1(n5055), .A2(n5077), .A3(n5054), .ZN(n5134) );
  NAND2_X1 U6261 ( .A1(n5134), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5062) );
  INV_X1 U6262 ( .A(n5131), .ZN(n5060) );
  NOR2_X1 U6263 ( .A1(n5075), .A2(n5144), .ZN(n6464) );
  NAND2_X1 U6264 ( .A1(n6464), .A2(n6658), .ZN(n5056) );
  OAI21_X1 U6265 ( .B1(n6466), .B2(n5057), .A(n5056), .ZN(n5128) );
  NAND2_X1 U6266 ( .A1(n5128), .A2(n6649), .ZN(n5058) );
  OAI21_X1 U6267 ( .B1(n5102), .B2(n6544), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6268 ( .B1(n5060), .B2(n6662), .A(n5059), .ZN(n5061) );
  OAI211_X1 U6269 ( .C1(n5127), .C2(n6665), .A(n5062), .B(n5061), .ZN(U3020)
         );
  AND2_X1 U6270 ( .A1(n4950), .A2(n5063), .ZN(n5065) );
  OR2_X1 U6271 ( .A1(n5065), .A2(n5064), .ZN(n6235) );
  INV_X1 U6272 ( .A(n5066), .ZN(n5233) );
  OAI21_X1 U6273 ( .B1(n5067), .B2(n4952), .A(n5233), .ZN(n6237) );
  INV_X1 U6274 ( .A(n6237), .ZN(n5068) );
  AOI22_X1 U6275 ( .A1(n5068), .A2(n4499), .B1(n5684), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5069) );
  OAI21_X1 U6276 ( .B1(n6235), .B2(n5694), .A(n5069), .ZN(U2852) );
  INV_X1 U6277 ( .A(n6595), .ZN(n5070) );
  NAND2_X1 U6278 ( .A1(n3111), .A2(n5070), .ZN(n6570) );
  OAI211_X1 U6279 ( .C1(n5072), .C2(n5071), .A(n7121), .B(n6570), .ZN(n5078)
         );
  OR2_X1 U6280 ( .A1(n5073), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7111)
         );
  OAI21_X1 U6281 ( .B1(n5075), .B2(n6592), .A(n5074), .ZN(n6657) );
  AOI21_X1 U6282 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7111), .A(n6657), .ZN(
        n5076) );
  NAND3_X1 U6283 ( .A1(n5078), .A2(n5077), .A3(n5076), .ZN(n7110) );
  NAND2_X1 U6284 ( .A1(n7110), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5083) );
  INV_X1 U6285 ( .A(n6712), .ZN(n6636) );
  NOR2_X1 U6286 ( .A1(n5079), .A2(n5144), .ZN(n6643) );
  AOI22_X1 U6287 ( .A1(n6642), .A2(n5080), .B1(n6658), .B2(n6643), .ZN(n7114)
         );
  OAI22_X1 U6288 ( .A1(n7114), .A2(n6580), .B1(n6633), .B2(n7111), .ZN(n5081)
         );
  AOI21_X1 U6289 ( .B1(n6636), .B2(n7116), .A(n5081), .ZN(n5082) );
  OAI211_X1 U6290 ( .C1(n7121), .C2(n6634), .A(n5083), .B(n5082), .ZN(U3091)
         );
  NAND2_X1 U6291 ( .A1(n7110), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5086) );
  OAI22_X1 U6292 ( .A1(n7114), .A2(n6574), .B1(n6625), .B2(n7111), .ZN(n5084)
         );
  AOI21_X1 U6293 ( .B1(n6628), .B2(n7116), .A(n5084), .ZN(n5085) );
  OAI211_X1 U6294 ( .C1(n7121), .C2(n6626), .A(n5086), .B(n5085), .ZN(U3090)
         );
  NAND2_X1 U6295 ( .A1(n7110), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5089) );
  OAI22_X1 U6296 ( .A1(n7114), .A2(n6553), .B1(n6544), .B2(n7111), .ZN(n5087)
         );
  AOI21_X1 U6297 ( .B1(n6589), .B2(n7116), .A(n5087), .ZN(n5088) );
  OAI211_X1 U6298 ( .C1(n7121), .C2(n6545), .A(n5089), .B(n5088), .ZN(U3084)
         );
  NAND2_X1 U6299 ( .A1(n7110), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U6300 ( .A1(n7114), .A2(n6562), .B1(n6606), .B2(n7111), .ZN(n5090)
         );
  AOI21_X1 U6301 ( .B1(n6609), .B2(n7116), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6302 ( .C1(n7121), .C2(n6607), .A(n5092), .B(n5091), .ZN(U3087)
         );
  NAND2_X1 U6303 ( .A1(n7110), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5095) );
  INV_X1 U6304 ( .A(n6689), .ZN(n6616) );
  OAI22_X1 U6305 ( .A1(n7114), .A2(n6565), .B1(n6613), .B2(n7111), .ZN(n5093)
         );
  AOI21_X1 U6306 ( .B1(n6616), .B2(n7116), .A(n5093), .ZN(n5094) );
  OAI211_X1 U6307 ( .C1(n7121), .C2(n6614), .A(n5095), .B(n5094), .ZN(U3088)
         );
  NAND2_X1 U6308 ( .A1(n7110), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U6309 ( .A1(n7114), .A2(n6556), .B1(n6507), .B2(n7111), .ZN(n5096)
         );
  AOI21_X1 U6310 ( .B1(n6599), .B2(n7116), .A(n5096), .ZN(n5097) );
  OAI211_X1 U6311 ( .C1(n7121), .C2(n5279), .A(n5098), .B(n5097), .ZN(U3085)
         );
  NAND2_X1 U6312 ( .A1(n7110), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5101) );
  INV_X1 U6313 ( .A(n6695), .ZN(n6621) );
  OAI22_X1 U6314 ( .A1(n7114), .A2(n6568), .B1(n6523), .B2(n7111), .ZN(n5099)
         );
  AOI21_X1 U6315 ( .B1(n6621), .B2(n7116), .A(n5099), .ZN(n5100) );
  OAI211_X1 U6316 ( .C1(n7121), .C2(n5266), .A(n5101), .B(n5100), .ZN(U3089)
         );
  OAI222_X1 U6317 ( .A1(n6235), .A2(n5747), .B1(n5744), .B2(n7079), .C1(n5746), 
        .C2(n3672), .ZN(U2884) );
  NOR2_X1 U6318 ( .A1(n5127), .A2(n6701), .ZN(n5105) );
  INV_X1 U6319 ( .A(n5102), .ZN(n5129) );
  AOI22_X1 U6320 ( .A1(n6696), .A2(n5129), .B1(n5128), .B2(n6697), .ZN(n5103)
         );
  OAI21_X1 U6321 ( .B1(n5131), .B2(n6626), .A(n5103), .ZN(n5104) );
  AOI211_X1 U6322 ( .C1(INSTQUEUE_REG_0__6__SCAN_IN), .C2(n5134), .A(n5105), 
        .B(n5104), .ZN(n5106) );
  INV_X1 U6323 ( .A(n5106), .ZN(U3026) );
  NOR2_X1 U6324 ( .A1(n5127), .A2(n6695), .ZN(n5109) );
  AOI22_X1 U6325 ( .A1(n6690), .A2(n5129), .B1(n5128), .B2(n6691), .ZN(n5107)
         );
  OAI21_X1 U6326 ( .B1(n5131), .B2(n5266), .A(n5107), .ZN(n5108) );
  AOI211_X1 U6327 ( .C1(INSTQUEUE_REG_0__5__SCAN_IN), .C2(n5134), .A(n5109), 
        .B(n5108), .ZN(n5110) );
  INV_X1 U6328 ( .A(n5110), .ZN(U3025) );
  NOR2_X1 U6329 ( .A1(n5127), .A2(n6689), .ZN(n5113) );
  AOI22_X1 U6330 ( .A1(n6684), .A2(n5129), .B1(n5128), .B2(n6685), .ZN(n5111)
         );
  OAI21_X1 U6331 ( .B1(n5131), .B2(n6614), .A(n5111), .ZN(n5112) );
  AOI211_X1 U6332 ( .C1(INSTQUEUE_REG_0__4__SCAN_IN), .C2(n5134), .A(n5113), 
        .B(n5112), .ZN(n5114) );
  INV_X1 U6333 ( .A(n5114), .ZN(U3024) );
  NOR2_X1 U6334 ( .A1(n5127), .A2(n6677), .ZN(n5117) );
  AOI22_X1 U6335 ( .A1(n6672), .A2(n5129), .B1(n5128), .B2(n6673), .ZN(n5115)
         );
  OAI21_X1 U6336 ( .B1(n5131), .B2(n7120), .A(n5115), .ZN(n5116) );
  AOI211_X1 U6337 ( .C1(INSTQUEUE_REG_0__2__SCAN_IN), .C2(n5134), .A(n5117), 
        .B(n5116), .ZN(n5118) );
  INV_X1 U6338 ( .A(n5118), .ZN(U3022) );
  NOR2_X1 U6339 ( .A1(n5127), .A2(n6683), .ZN(n5121) );
  AOI22_X1 U6340 ( .A1(n6678), .A2(n5129), .B1(n5128), .B2(n6679), .ZN(n5119)
         );
  OAI21_X1 U6341 ( .B1(n5131), .B2(n6607), .A(n5119), .ZN(n5120) );
  AOI211_X1 U6342 ( .C1(INSTQUEUE_REG_0__3__SCAN_IN), .C2(n5134), .A(n5121), 
        .B(n5120), .ZN(n5122) );
  INV_X1 U6343 ( .A(n5122), .ZN(U3023) );
  NOR2_X1 U6344 ( .A1(n5127), .A2(n6671), .ZN(n5125) );
  AOI22_X1 U6345 ( .A1(n6666), .A2(n5129), .B1(n5128), .B2(n6667), .ZN(n5123)
         );
  OAI21_X1 U6346 ( .B1(n5131), .B2(n5279), .A(n5123), .ZN(n5124) );
  AOI211_X1 U6347 ( .C1(INSTQUEUE_REG_0__1__SCAN_IN), .C2(n5134), .A(n5125), 
        .B(n5124), .ZN(n5126) );
  INV_X1 U6348 ( .A(n5126), .ZN(U3021) );
  NOR2_X1 U6349 ( .A1(n5127), .A2(n6712), .ZN(n5133) );
  AOI22_X1 U6350 ( .A1(n6703), .A2(n5129), .B1(n5128), .B2(n6704), .ZN(n5130)
         );
  OAI21_X1 U6351 ( .B1(n5131), .B2(n6634), .A(n5130), .ZN(n5132) );
  AOI211_X1 U6352 ( .C1(INSTQUEUE_REG_0__7__SCAN_IN), .C2(n5134), .A(n5133), 
        .B(n5132), .ZN(n5135) );
  INV_X1 U6353 ( .A(n5135), .ZN(U3027) );
  AND2_X1 U6354 ( .A1(n6474), .A2(n5137), .ZN(n6533) );
  NOR3_X1 U6355 ( .A1(n6533), .A2(n6576), .A3(n6651), .ZN(n5138) );
  OAI22_X1 U6356 ( .A1(n5138), .A2(n6655), .B1(n6495), .B2(n5146), .ZN(n5143)
         );
  NAND2_X1 U6357 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5139) );
  INV_X1 U6358 ( .A(n6658), .ZN(n5142) );
  NAND2_X1 U6359 ( .A1(n6550), .A2(n7028), .ZN(n5178) );
  NAND2_X1 U6360 ( .A1(n5178), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6361 ( .A1(n5175), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5150) );
  AND2_X1 U6362 ( .A1(n5144), .A2(n6462), .ZN(n5198) );
  NAND2_X1 U6363 ( .A1(n6463), .A2(n5198), .ZN(n5145) );
  OAI21_X1 U6364 ( .B1(n6466), .B2(n5146), .A(n5145), .ZN(n5176) );
  NAND2_X1 U6365 ( .A1(n5176), .A2(n6704), .ZN(n5147) );
  OAI21_X1 U6366 ( .B1(n5178), .B2(n6633), .A(n5147), .ZN(n5148) );
  AOI21_X1 U6367 ( .B1(n6576), .B2(n6707), .A(n5148), .ZN(n5149) );
  OAI211_X1 U6368 ( .C1(n5182), .C2(n6712), .A(n5150), .B(n5149), .ZN(U3075)
         );
  NAND2_X1 U6369 ( .A1(n5175), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6370 ( .A1(n5176), .A2(n6649), .ZN(n5151) );
  OAI21_X1 U6371 ( .B1(n5178), .B2(n6544), .A(n5151), .ZN(n5152) );
  AOI21_X1 U6372 ( .B1(n6576), .B2(n6662), .A(n5152), .ZN(n5153) );
  OAI211_X1 U6373 ( .C1(n5182), .C2(n6665), .A(n5154), .B(n5153), .ZN(U3068)
         );
  NAND2_X1 U6374 ( .A1(n5175), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6375 ( .A1(n5176), .A2(n6697), .ZN(n5155) );
  OAI21_X1 U6376 ( .B1(n5178), .B2(n6625), .A(n5155), .ZN(n5156) );
  AOI21_X1 U6377 ( .B1(n6576), .B2(n6698), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6378 ( .C1(n5182), .C2(n6701), .A(n5158), .B(n5157), .ZN(U3074)
         );
  NAND2_X1 U6379 ( .A1(n5175), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6380 ( .A1(n5176), .A2(n6667), .ZN(n5159) );
  OAI21_X1 U6381 ( .B1(n5178), .B2(n6507), .A(n5159), .ZN(n5160) );
  AOI21_X1 U6382 ( .B1(n6576), .B2(n6668), .A(n5160), .ZN(n5161) );
  OAI211_X1 U6383 ( .C1(n5182), .C2(n6671), .A(n5162), .B(n5161), .ZN(U3069)
         );
  NAND2_X1 U6384 ( .A1(n5175), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6385 ( .A1(n5176), .A2(n6685), .ZN(n5163) );
  OAI21_X1 U6386 ( .B1(n5178), .B2(n6613), .A(n5163), .ZN(n5164) );
  AOI21_X1 U6387 ( .B1(n6576), .B2(n6686), .A(n5164), .ZN(n5165) );
  OAI211_X1 U6388 ( .C1(n5182), .C2(n6689), .A(n5166), .B(n5165), .ZN(U3072)
         );
  NAND2_X1 U6389 ( .A1(n5175), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6390 ( .A1(n5176), .A2(n6679), .ZN(n5167) );
  OAI21_X1 U6391 ( .B1(n5178), .B2(n6606), .A(n5167), .ZN(n5168) );
  AOI21_X1 U6392 ( .B1(n6576), .B2(n6680), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6393 ( .C1(n5182), .C2(n6683), .A(n5170), .B(n5169), .ZN(U3071)
         );
  NAND2_X1 U6394 ( .A1(n5175), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6395 ( .A1(n5176), .A2(n6673), .ZN(n5171) );
  OAI21_X1 U6396 ( .B1(n5178), .B2(n7112), .A(n5171), .ZN(n5172) );
  AOI21_X1 U6397 ( .B1(n6576), .B2(n6674), .A(n5172), .ZN(n5173) );
  OAI211_X1 U6398 ( .C1(n5182), .C2(n6677), .A(n5174), .B(n5173), .ZN(U3070)
         );
  NAND2_X1 U6399 ( .A1(n5175), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6400 ( .A1(n5176), .A2(n6691), .ZN(n5177) );
  OAI21_X1 U6401 ( .B1(n5178), .B2(n6523), .A(n5177), .ZN(n5179) );
  AOI21_X1 U6402 ( .B1(n6576), .B2(n6692), .A(n5179), .ZN(n5180) );
  OAI211_X1 U6403 ( .C1(n5182), .C2(n6695), .A(n5181), .B(n5180), .ZN(U3073)
         );
  XNOR2_X1 U6404 ( .A(n5183), .B(n5184), .ZN(n5245) );
  INV_X1 U6405 ( .A(n5607), .ZN(n5187) );
  AND2_X1 U6406 ( .A1(n6377), .A2(REIP_REG_6__SCAN_IN), .ZN(n5242) );
  AOI21_X1 U6407 ( .B1(n6358), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5242), 
        .ZN(n5185) );
  OAI21_X1 U6408 ( .B1(n5599), .B2(n6370), .A(n5185), .ZN(n5186) );
  AOI21_X1 U6409 ( .B1(n5187), .B2(n6365), .A(n5186), .ZN(n5188) );
  OAI21_X1 U6410 ( .B1(n6339), .B2(n5245), .A(n5188), .ZN(U2980) );
  OAI21_X1 U6411 ( .B1(n5191), .B2(n5225), .A(n5190), .ZN(n5193) );
  NOR2_X1 U6412 ( .A1(n5625), .A2(n5637), .ZN(n5257) );
  NAND2_X1 U6413 ( .A1(n5257), .A2(n5192), .ZN(n5197) );
  AOI21_X1 U6414 ( .B1(n5193), .B2(n5197), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5196) );
  NOR2_X1 U6415 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5194) );
  AND2_X1 U6416 ( .A1(n5194), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6431)
         );
  AND2_X1 U6417 ( .A1(n6431), .A2(n7028), .ZN(n5199) );
  NAND2_X1 U6418 ( .A1(n5221), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5202) );
  INV_X1 U6419 ( .A(n5197), .ZN(n6421) );
  AOI22_X1 U6420 ( .A1(n6421), .A2(n6586), .B1(n6658), .B2(n5198), .ZN(n5223)
         );
  INV_X1 U6421 ( .A(n5199), .ZN(n5222) );
  OAI22_X1 U6422 ( .A1(n5223), .A2(n6568), .B1(n6523), .B2(n5222), .ZN(n5200)
         );
  AOI21_X1 U6423 ( .B1(n6692), .B2(n5225), .A(n5200), .ZN(n5201) );
  OAI211_X1 U6424 ( .C1(n5228), .C2(n6695), .A(n5202), .B(n5201), .ZN(U3041)
         );
  NAND2_X1 U6425 ( .A1(n5221), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5205) );
  OAI22_X1 U6426 ( .A1(n5223), .A2(n6562), .B1(n6606), .B2(n5222), .ZN(n5203)
         );
  AOI21_X1 U6427 ( .B1(n6680), .B2(n5225), .A(n5203), .ZN(n5204) );
  OAI211_X1 U6428 ( .C1(n5228), .C2(n6683), .A(n5205), .B(n5204), .ZN(U3039)
         );
  NAND2_X1 U6429 ( .A1(n5221), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5208) );
  OAI22_X1 U6430 ( .A1(n5223), .A2(n7113), .B1(n7112), .B2(n5222), .ZN(n5206)
         );
  AOI21_X1 U6431 ( .B1(n6674), .B2(n5225), .A(n5206), .ZN(n5207) );
  OAI211_X1 U6432 ( .C1(n5228), .C2(n6677), .A(n5208), .B(n5207), .ZN(U3038)
         );
  NAND2_X1 U6433 ( .A1(n5221), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5211) );
  OAI22_X1 U6434 ( .A1(n5223), .A2(n6556), .B1(n6507), .B2(n5222), .ZN(n5209)
         );
  AOI21_X1 U6435 ( .B1(n6668), .B2(n5225), .A(n5209), .ZN(n5210) );
  OAI211_X1 U6436 ( .C1(n5228), .C2(n6671), .A(n5211), .B(n5210), .ZN(U3037)
         );
  NAND2_X1 U6437 ( .A1(n5221), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5214) );
  OAI22_X1 U6438 ( .A1(n5223), .A2(n6565), .B1(n6613), .B2(n5222), .ZN(n5212)
         );
  AOI21_X1 U6439 ( .B1(n6686), .B2(n5225), .A(n5212), .ZN(n5213) );
  OAI211_X1 U6440 ( .C1(n5228), .C2(n6689), .A(n5214), .B(n5213), .ZN(U3040)
         );
  NAND2_X1 U6441 ( .A1(n5221), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5217) );
  OAI22_X1 U6442 ( .A1(n5223), .A2(n6580), .B1(n6633), .B2(n5222), .ZN(n5215)
         );
  AOI21_X1 U6443 ( .B1(n6707), .B2(n5225), .A(n5215), .ZN(n5216) );
  OAI211_X1 U6444 ( .C1(n5228), .C2(n6712), .A(n5217), .B(n5216), .ZN(U3043)
         );
  NAND2_X1 U6445 ( .A1(n5221), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5220) );
  OAI22_X1 U6446 ( .A1(n5223), .A2(n6553), .B1(n6544), .B2(n5222), .ZN(n5218)
         );
  AOI21_X1 U6447 ( .B1(n6662), .B2(n5225), .A(n5218), .ZN(n5219) );
  OAI211_X1 U6448 ( .C1(n5228), .C2(n6665), .A(n5220), .B(n5219), .ZN(U3036)
         );
  NAND2_X1 U6449 ( .A1(n5221), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5227) );
  OAI22_X1 U6450 ( .A1(n5223), .A2(n6574), .B1(n6625), .B2(n5222), .ZN(n5224)
         );
  AOI21_X1 U6451 ( .B1(n6698), .B2(n5225), .A(n5224), .ZN(n5226) );
  OAI211_X1 U6452 ( .C1(n5228), .C2(n6701), .A(n5227), .B(n5226), .ZN(U3042)
         );
  NOR2_X1 U6453 ( .A1(n5064), .A2(n5229), .ZN(n5230) );
  OR2_X1 U6454 ( .A1(n3100), .A2(n5230), .ZN(n6224) );
  INV_X1 U6455 ( .A(n5231), .ZN(n5234) );
  AOI21_X1 U6456 ( .B1(n5234), .B2(n5233), .A(n4227), .ZN(n6220) );
  AOI22_X1 U6457 ( .A1(n6220), .A2(n4499), .B1(n5684), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5235) );
  OAI21_X1 U6458 ( .B1(n6224), .B2(n5694), .A(n5235), .ZN(U2851) );
  AOI22_X1 U6459 ( .A1(n5749), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5748), .ZN(n5236) );
  OAI21_X1 U6460 ( .B1(n6224), .B2(n5747), .A(n5236), .ZN(U2883) );
  INV_X1 U6462 ( .A(n5237), .ZN(n5239) );
  OAI33_X1 U6463 ( .A1(1'b0), .A2(n5239), .A3(n4385), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n5300), .B3(n5238), .ZN(n5241) );
  INV_X1 U6464 ( .A(n5241), .ZN(n5244) );
  AOI21_X1 U6465 ( .B1(n6410), .B2(n5601), .A(n5242), .ZN(n5243) );
  OAI211_X1 U6466 ( .C1(n6101), .C2(n5245), .A(n5244), .B(n5243), .ZN(U3012)
         );
  OR2_X1 U6467 ( .A1(n3100), .A2(n5247), .ZN(n5248) );
  NAND2_X1 U6468 ( .A1(n5246), .A2(n5248), .ZN(n6215) );
  NAND2_X1 U6469 ( .A1(n5232), .A2(n5249), .ZN(n5250) );
  AND2_X1 U6470 ( .A1(n5587), .A2(n5250), .ZN(n6384) );
  AOI22_X1 U6471 ( .A1(n6384), .A2(n4499), .B1(EBX_REG_9__SCAN_IN), .B2(n5684), 
        .ZN(n5251) );
  OAI21_X1 U6472 ( .B1(n6215), .B2(n5694), .A(n5251), .ZN(U2850) );
  OAI222_X1 U6473 ( .A1(n6215), .A2(n5747), .B1(n5746), .B2(n5253), .C1(n5744), 
        .C2(n5252), .ZN(U2882) );
  INV_X1 U6474 ( .A(n6596), .ZN(n5255) );
  OAI21_X1 U6475 ( .B1(n3109), .B2(n6637), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5256) );
  NAND2_X1 U6476 ( .A1(n5256), .A2(n6586), .ZN(n5263) );
  INV_X1 U6477 ( .A(n5263), .ZN(n5259) );
  AND2_X1 U6478 ( .A1(n5257), .A2(n5612), .ZN(n6584) );
  AND3_X1 U6479 ( .A1(n6827), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U6480 ( .A1(n6590), .A2(n7028), .ZN(n5286) );
  OAI22_X1 U6481 ( .A1(n5287), .A2(n6634), .B1(n5286), .B2(n6633), .ZN(n5260)
         );
  AOI21_X1 U6482 ( .B1(n3109), .B2(n6636), .A(n5260), .ZN(n5265) );
  AOI211_X1 U6483 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5286), .A(n6463), .B(
        n5261), .ZN(n5262) );
  NAND2_X1 U6484 ( .A1(n5289), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5264)
         );
  OAI211_X1 U6485 ( .C1(n5292), .C2(n6580), .A(n5265), .B(n5264), .ZN(U3107)
         );
  OAI22_X1 U6486 ( .A1(n5287), .A2(n5266), .B1(n5286), .B2(n6523), .ZN(n5267)
         );
  AOI21_X1 U6487 ( .B1(n3109), .B2(n6621), .A(n5267), .ZN(n5269) );
  NAND2_X1 U6488 ( .A1(n5289), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5268)
         );
  OAI211_X1 U6489 ( .C1(n5292), .C2(n6568), .A(n5269), .B(n5268), .ZN(U3105)
         );
  INV_X1 U6490 ( .A(n6677), .ZN(n7117) );
  OAI22_X1 U6491 ( .A1(n5287), .A2(n7120), .B1(n5286), .B2(n7112), .ZN(n5270)
         );
  AOI21_X1 U6492 ( .B1(n3109), .B2(n7117), .A(n5270), .ZN(n5272) );
  NAND2_X1 U6493 ( .A1(n5289), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5271)
         );
  OAI211_X1 U6494 ( .C1(n5292), .C2(n7113), .A(n5272), .B(n5271), .ZN(U3102)
         );
  OAI22_X1 U6495 ( .A1(n5287), .A2(n6607), .B1(n5286), .B2(n6606), .ZN(n5273)
         );
  AOI21_X1 U6496 ( .B1(n3109), .B2(n6609), .A(n5273), .ZN(n5275) );
  NAND2_X1 U6497 ( .A1(n5289), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5274)
         );
  OAI211_X1 U6498 ( .C1(n5292), .C2(n6562), .A(n5275), .B(n5274), .ZN(U3103)
         );
  OAI22_X1 U6499 ( .A1(n5287), .A2(n6545), .B1(n5286), .B2(n6544), .ZN(n5276)
         );
  AOI21_X1 U6500 ( .B1(n3109), .B2(n6589), .A(n5276), .ZN(n5278) );
  NAND2_X1 U6501 ( .A1(n5289), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5277)
         );
  OAI211_X1 U6502 ( .C1(n5292), .C2(n6553), .A(n5278), .B(n5277), .ZN(U3100)
         );
  OAI22_X1 U6503 ( .A1(n5287), .A2(n5279), .B1(n5286), .B2(n6507), .ZN(n5280)
         );
  AOI21_X1 U6504 ( .B1(n3109), .B2(n6599), .A(n5280), .ZN(n5282) );
  NAND2_X1 U6505 ( .A1(n5289), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5281)
         );
  OAI211_X1 U6506 ( .C1(n5292), .C2(n6556), .A(n5282), .B(n5281), .ZN(U3101)
         );
  OAI22_X1 U6507 ( .A1(n5287), .A2(n6614), .B1(n5286), .B2(n6613), .ZN(n5283)
         );
  AOI21_X1 U6508 ( .B1(n3109), .B2(n6616), .A(n5283), .ZN(n5285) );
  NAND2_X1 U6509 ( .A1(n5289), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5284)
         );
  OAI211_X1 U6510 ( .C1(n5292), .C2(n6565), .A(n5285), .B(n5284), .ZN(U3104)
         );
  OAI22_X1 U6511 ( .A1(n5287), .A2(n6626), .B1(n5286), .B2(n6625), .ZN(n5288)
         );
  AOI21_X1 U6512 ( .B1(n3109), .B2(n6628), .A(n5288), .ZN(n5291) );
  NAND2_X1 U6513 ( .A1(n5289), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5290)
         );
  OAI211_X1 U6514 ( .C1(n5292), .C2(n6574), .A(n5291), .B(n5290), .ZN(U3106)
         );
  XNOR2_X1 U6515 ( .A(n5293), .B(n5294), .ZN(n5314) );
  INV_X1 U6516 ( .A(n6039), .ZN(n5296) );
  OAI22_X1 U6517 ( .A1(n5298), .A2(n5297), .B1(n5296), .B2(n5295), .ZN(n6371)
         );
  INV_X1 U6518 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6735) );
  NOR3_X1 U6519 ( .A1(n5300), .A2(n5299), .A3(n6807), .ZN(n6374) );
  OAI211_X1 U6520 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6374), .B(n6373), .ZN(n5302) );
  NAND2_X1 U6521 ( .A1(n6220), .A2(n6410), .ZN(n5301) );
  OAI211_X1 U6522 ( .C1(n6735), .C2(n6396), .A(n5302), .B(n5301), .ZN(n5303)
         );
  AOI21_X1 U6523 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n6371), .A(n5303), 
        .ZN(n5304) );
  OAI21_X1 U6524 ( .B1(n6101), .B2(n5314), .A(n5304), .ZN(U3010) );
  XOR2_X1 U6525 ( .A(n5305), .B(n5306), .Z(n6344) );
  AOI22_X1 U6526 ( .A1(n6374), .A2(n4396), .B1(n6412), .B2(n6344), .ZN(n5309)
         );
  NAND2_X1 U6527 ( .A1(n6377), .A2(REIP_REG_7__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U6528 ( .B1(n6398), .B2(n6237), .A(n6345), .ZN(n5307) );
  AOI21_X1 U6529 ( .B1(n6371), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5307), 
        .ZN(n5308) );
  NAND2_X1 U6530 ( .A1(n5309), .A2(n5308), .ZN(U3011) );
  OAI22_X1 U6531 ( .A1(n6356), .A2(n5310), .B1(n6396), .B2(n6735), .ZN(n5312)
         );
  NOR2_X1 U6532 ( .A1(n6224), .A2(n6334), .ZN(n5311) );
  AOI211_X1 U6533 ( .C1(n6350), .C2(n6221), .A(n5312), .B(n5311), .ZN(n5313)
         );
  OAI21_X1 U6534 ( .B1(n6339), .B2(n5314), .A(n5313), .ZN(U2978) );
  NAND2_X1 U6535 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5327) );
  AOI22_X1 U6536 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4506), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4189), .ZN(n5328) );
  INV_X1 U6537 ( .A(n5328), .ZN(n5320) );
  NOR3_X1 U6538 ( .A1(n5315), .A2(n4777), .A3(n4776), .ZN(n5318) );
  NOR2_X1 U6539 ( .A1(n5637), .A2(n5316), .ZN(n5317) );
  AOI211_X1 U6540 ( .C1(n6117), .C2(n3287), .A(n5318), .B(n5317), .ZN(n6120)
         );
  INV_X1 U6541 ( .A(n3295), .ZN(n5319) );
  OAI222_X1 U6542 ( .A1(n5327), .A2(n5320), .B1(n6113), .B2(n6120), .C1(n5319), 
        .C2(n6145), .ZN(n5322) );
  AOI22_X1 U6543 ( .A1(n5322), .A2(n6115), .B1(n5321), .B2(n5325), .ZN(n5323)
         );
  OAI21_X1 U6544 ( .B1(n3287), .B2(n6115), .A(n5323), .ZN(U3460) );
  INV_X1 U6545 ( .A(n4777), .ZN(n5324) );
  AOI21_X1 U6546 ( .B1(n5325), .B2(n5324), .A(n5333), .ZN(n5335) );
  INV_X1 U6547 ( .A(n5326), .ZN(n5331) );
  NAND2_X1 U6548 ( .A1(n4777), .A2(n5334), .ZN(n5329) );
  OAI22_X1 U6549 ( .A1(n6145), .A2(n5329), .B1(n5328), .B2(n5327), .ZN(n5330)
         );
  AOI21_X1 U6550 ( .B1(n5331), .B2(n6155), .A(n5330), .ZN(n5332) );
  OAI22_X1 U6551 ( .A1(n5335), .A2(n5334), .B1(n5333), .B2(n5332), .ZN(U3459)
         );
  CLKBUF_X1 U6552 ( .A(n5336), .Z(n5789) );
  INV_X1 U6553 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5337) );
  AND2_X1 U6554 ( .A1(n5779), .A2(n5337), .ZN(n5338) );
  NAND2_X1 U6555 ( .A1(n5789), .A2(n5338), .ZN(n5769) );
  AOI22_X1 U6556 ( .A1(n5340), .A2(n5769), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5339), .ZN(n5341) );
  XNOR2_X1 U6557 ( .A(n5341), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5929)
         );
  INV_X1 U6558 ( .A(n5362), .ZN(n5346) );
  NOR2_X1 U6559 ( .A1(n5354), .A2(n6370), .ZN(n5345) );
  NAND2_X1 U6560 ( .A1(n6377), .A2(REIP_REG_28__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6561 ( .B1(n6356), .B2(n5349), .A(n5923), .ZN(n5344) );
  OAI21_X1 U6562 ( .B1(n6339), .B2(n5929), .A(n5347), .ZN(U2958) );
  XNOR2_X1 U6563 ( .A(n5402), .B(n5348), .ZN(n5361) );
  INV_X1 U6564 ( .A(n5361), .ZN(n5927) );
  INV_X2 U6565 ( .A(n6269), .ZN(n6250) );
  OAI22_X1 U6566 ( .A1(n6266), .A2(n5349), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5391), .ZN(n5352) );
  NOR2_X1 U6567 ( .A1(n5350), .A2(n6768), .ZN(n5351) );
  OAI21_X1 U6568 ( .B1(n5354), .B2(n6247), .A(n5353), .ZN(n5355) );
  AOI21_X1 U6569 ( .B1(n5927), .B2(n6252), .A(n5355), .ZN(n5356) );
  OAI21_X1 U6570 ( .B1(n5362), .B2(n6207), .A(n5356), .ZN(U2799) );
  AOI22_X1 U6571 ( .A1(n5732), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5748), .ZN(n5360) );
  NOR3_X1 U6572 ( .A1(n5748), .A2(n5698), .A3(n3810), .ZN(n5358) );
  NAND2_X1 U6573 ( .A1(n5733), .A2(DATAI_12_), .ZN(n5359) );
  OAI211_X1 U6574 ( .C1(n5362), .C2(n5747), .A(n5360), .B(n5359), .ZN(U2863)
         );
  INV_X1 U6575 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6909) );
  OAI222_X1 U6576 ( .A1(n5362), .A2(n5694), .B1(n5697), .B2(n5361), .C1(n5696), 
        .C2(n6909), .ZN(U2831) );
  AOI22_X1 U6577 ( .A1(n5732), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5748), .ZN(n5364) );
  NAND2_X1 U6578 ( .A1(n5733), .A2(DATAI_14_), .ZN(n5363) );
  OAI211_X1 U6579 ( .C1(n5365), .C2(n5747), .A(n5364), .B(n5363), .ZN(U2861)
         );
  OR2_X1 U6580 ( .A1(n5498), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5368) );
  INV_X1 U6581 ( .A(n5366), .ZN(n5367) );
  MUX2_X1 U6582 ( .A(n5368), .B(n5367), .S(n6792), .Z(U3474) );
  INV_X1 U6583 ( .A(n5635), .ZN(n5378) );
  OAI211_X1 U6584 ( .C1(n5392), .C2(n6770), .A(REIP_REG_31__SCAN_IN), .B(n5615), .ZN(n5376) );
  NOR2_X1 U6585 ( .A1(n6770), .A2(REIP_REG_31__SCAN_IN), .ZN(n5373) );
  AOI22_X1 U6586 ( .A1(n6234), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n5374), 
        .B2(n5373), .ZN(n5375) );
  OAI211_X1 U6587 ( .C1(n5378), .C2(n5377), .A(n5376), .B(n5375), .ZN(n5379)
         );
  AOI21_X1 U6588 ( .B1(n5654), .B2(n6252), .A(n5379), .ZN(n5380) );
  OAI21_X1 U6589 ( .B1(n5758), .B2(n6207), .A(n5380), .ZN(U2796) );
  INV_X1 U6590 ( .A(n5767), .ZN(n5703) );
  NAND2_X1 U6591 ( .A1(n5384), .A2(n5383), .ZN(n5386) );
  NAND2_X1 U6592 ( .A1(n5386), .A2(n5385), .ZN(n5387) );
  NOR2_X1 U6593 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  INV_X1 U6594 ( .A(n5763), .ZN(n5396) );
  AOI22_X1 U6595 ( .A1(n6250), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6234), .ZN(n5395) );
  NOR2_X1 U6596 ( .A1(n5391), .A2(n6768), .ZN(n5393) );
  OAI21_X1 U6597 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5393), .A(n5392), .ZN(n5394) );
  OAI211_X1 U6598 ( .C1(n6247), .C2(n5396), .A(n5395), .B(n5394), .ZN(n5397)
         );
  AOI21_X1 U6599 ( .B1(n3114), .B2(n6252), .A(n5397), .ZN(n5398) );
  OAI21_X1 U6600 ( .B1(n5703), .B2(n6207), .A(n5398), .ZN(U2798) );
  NOR2_X1 U6601 ( .A1(n5399), .A2(n5400), .ZN(n5401) );
  AOI21_X1 U6602 ( .B1(n5405), .B2(n5403), .A(n5404), .ZN(n5775) );
  NAND2_X1 U6603 ( .A1(n5775), .A2(n6241), .ZN(n5413) );
  NAND2_X1 U6604 ( .A1(n6250), .A2(EBX_REG_27__SCAN_IN), .ZN(n5408) );
  INV_X1 U6605 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6764) );
  NAND3_X1 U6606 ( .A1(n5429), .A2(n5406), .A3(n6764), .ZN(n5407) );
  OAI211_X1 U6607 ( .C1(n6266), .C2(n5773), .A(n5408), .B(n5407), .ZN(n5411)
         );
  INV_X1 U6608 ( .A(n5771), .ZN(n5409) );
  NOR2_X1 U6609 ( .A1(n6247), .A2(n5409), .ZN(n5410) );
  AOI211_X1 U6610 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5417), .A(n5411), .B(n5410), .ZN(n5412) );
  OAI211_X1 U6611 ( .C1(n5932), .C2(n6277), .A(n5413), .B(n5412), .ZN(U2800)
         );
  AOI21_X1 U6612 ( .B1(n5416), .B2(n5426), .A(n5399), .ZN(n5939) );
  AOI22_X1 U6613 ( .A1(n6250), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6234), .ZN(n5420) );
  INV_X1 U6614 ( .A(n5429), .ZN(n5440) );
  NOR2_X1 U6615 ( .A1(n5440), .A2(n5428), .ZN(n5418) );
  OAI21_X1 U6616 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5418), .A(n5417), .ZN(n5419) );
  OAI211_X1 U6617 ( .C1(n6247), .C2(n5777), .A(n5420), .B(n5419), .ZN(n5421)
         );
  AOI21_X1 U6618 ( .B1(n5939), .B2(n6252), .A(n5421), .ZN(n5422) );
  OAI21_X1 U6619 ( .B1(n5786), .B2(n6207), .A(n5422), .ZN(U2801) );
  AOI21_X1 U6620 ( .B1(n5423), .B2(n5438), .A(n5414), .ZN(n5424) );
  AOI21_X1 U6621 ( .B1(n5427), .B2(n5425), .A(n3249), .ZN(n5953) );
  INV_X1 U6622 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6623 ( .A1(n6259), .A2(n5790), .ZN(n5433) );
  OAI211_X1 U6624 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5429), .B(n5428), .ZN(n5430) );
  OAI21_X1 U6625 ( .B1(n6266), .B2(n3193), .A(n5430), .ZN(n5431) );
  AOI21_X1 U6626 ( .B1(n6250), .B2(EBX_REG_25__SCAN_IN), .A(n5431), .ZN(n5432)
         );
  OAI211_X1 U6627 ( .C1(n5450), .C2(n5434), .A(n5433), .B(n5432), .ZN(n5435)
         );
  AOI21_X1 U6628 ( .B1(n5953), .B2(n6252), .A(n5435), .ZN(n5436) );
  OAI21_X1 U6629 ( .B1(n5794), .B2(n6207), .A(n5436), .ZN(U2802) );
  OAI21_X1 U6630 ( .B1(n5437), .B2(n5439), .A(n5438), .ZN(n5799) );
  INV_X1 U6631 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6761) );
  OAI22_X1 U6632 ( .A1(n6266), .A2(n7044), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5440), .ZN(n5441) );
  AOI21_X1 U6633 ( .B1(n6250), .B2(EBX_REG_24__SCAN_IN), .A(n5441), .ZN(n5442)
         );
  OAI21_X1 U6634 ( .B1(n5450), .B2(n6761), .A(n5442), .ZN(n5445) );
  OAI21_X1 U6635 ( .B1(n5448), .B2(n5443), .A(n5425), .ZN(n5956) );
  NOR2_X1 U6636 ( .A1(n5956), .A2(n6277), .ZN(n5444) );
  AOI211_X1 U6637 ( .C1(n6259), .C2(n5802), .A(n5445), .B(n5444), .ZN(n5446)
         );
  OAI21_X1 U6638 ( .B1(n5799), .B2(n6207), .A(n5446), .ZN(U2803) );
  AOI21_X1 U6639 ( .B1(n5447), .B2(n4527), .A(n5437), .ZN(n5810) );
  INV_X1 U6640 ( .A(n5810), .ZN(n5715) );
  AOI21_X1 U6641 ( .B1(n5449), .B2(n5460), .A(n5448), .ZN(n5970) );
  AOI22_X1 U6642 ( .A1(n6250), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6234), .ZN(n5454) );
  NOR2_X1 U6643 ( .A1(n5461), .A2(n6758), .ZN(n5452) );
  INV_X1 U6644 ( .A(n5450), .ZN(n5451) );
  OAI21_X1 U6645 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5452), .A(n5451), .ZN(n5453) );
  OAI211_X1 U6646 ( .C1(n6247), .C2(n5808), .A(n5454), .B(n5453), .ZN(n5455)
         );
  AOI21_X1 U6647 ( .B1(n5970), .B2(n6252), .A(n5455), .ZN(n5456) );
  OAI21_X1 U6648 ( .B1(n5715), .B2(n6207), .A(n5456), .ZN(U2804) );
  INV_X1 U6649 ( .A(n5457), .ZN(n5468) );
  NAND2_X1 U6650 ( .A1(n5473), .A2(n5458), .ZN(n5459) );
  NAND2_X1 U6651 ( .A1(n5460), .A2(n5459), .ZN(n5981) );
  OAI22_X1 U6652 ( .A1(n6266), .A2(n5462), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5461), .ZN(n5463) );
  AOI21_X1 U6653 ( .B1(n6250), .B2(EBX_REG_22__SCAN_IN), .A(n5463), .ZN(n5466)
         );
  INV_X1 U6654 ( .A(n5480), .ZN(n5489) );
  INV_X1 U6655 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6987) );
  NOR3_X1 U6656 ( .A1(n6987), .A2(REIP_REG_21__SCAN_IN), .A3(n5464), .ZN(n5477) );
  OAI21_X1 U6657 ( .B1(n5489), .B2(n5477), .A(REIP_REG_22__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U6658 ( .C1(n5981), .C2(n6277), .A(n5466), .B(n5465), .ZN(n5467)
         );
  AOI21_X1 U6659 ( .B1(n5468), .B2(n6259), .A(n5467), .ZN(n5469) );
  OAI21_X1 U6660 ( .B1(n5718), .B2(n6207), .A(n5469), .ZN(U2805) );
  XOR2_X1 U6661 ( .A(n5472), .B(n5471), .Z(n5818) );
  INV_X1 U6662 ( .A(n5818), .ZN(n5721) );
  INV_X1 U6663 ( .A(n5473), .ZN(n5474) );
  AOI21_X1 U6664 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5987) );
  AOI21_X1 U6665 ( .B1(n6234), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5477), 
        .ZN(n5479) );
  NAND2_X1 U6666 ( .A1(n6250), .A2(EBX_REG_21__SCAN_IN), .ZN(n5478) );
  OAI211_X1 U6667 ( .C1(n5480), .C2(n6756), .A(n5479), .B(n5478), .ZN(n5482)
         );
  NOR2_X1 U6668 ( .A1(n6247), .A2(n5816), .ZN(n5481) );
  AOI211_X1 U6669 ( .C1(n5987), .C2(n6252), .A(n5482), .B(n5481), .ZN(n5483)
         );
  OAI21_X1 U6670 ( .B1(n5721), .B2(n6207), .A(n5483), .ZN(U2806) );
  OAI21_X1 U6671 ( .B1(n5484), .B2(n5485), .A(n5471), .ZN(n5824) );
  MUX2_X1 U6672 ( .A(n5503), .B(n5502), .S(n5486), .Z(n5488) );
  XNOR2_X1 U6673 ( .A(n5488), .B(n5487), .ZN(n6002) );
  AOI22_X1 U6674 ( .A1(n6250), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6234), .ZN(n5492) );
  OAI21_X1 U6675 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5490), .A(n5489), .ZN(n5491) );
  OAI211_X1 U6676 ( .C1(n6247), .C2(n5826), .A(n5492), .B(n5491), .ZN(n5493)
         );
  AOI21_X1 U6677 ( .B1(n6252), .B2(n6002), .A(n5493), .ZN(n5494) );
  OAI21_X1 U6678 ( .B1(n5824), .B2(n6207), .A(n5494), .ZN(U2807) );
  AOI21_X1 U6679 ( .B1(n5496), .B2(n5512), .A(n5484), .ZN(n5838) );
  NAND2_X1 U6680 ( .A1(n5838), .A2(n6241), .ZN(n5510) );
  INV_X1 U6681 ( .A(n5497), .ZN(n5521) );
  XNOR2_X1 U6682 ( .A(REIP_REG_18__SCAN_IN), .B(REIP_REG_19__SCAN_IN), .ZN(
        n5501) );
  NAND2_X1 U6683 ( .A1(n6183), .A2(n5498), .ZN(n6264) );
  OAI21_X1 U6684 ( .B1(n6266), .B2(n6967), .A(n6264), .ZN(n5499) );
  AOI21_X1 U6685 ( .B1(n6250), .B2(EBX_REG_19__SCAN_IN), .A(n5499), .ZN(n5500)
         );
  OAI21_X1 U6686 ( .B1(n5521), .B2(n5501), .A(n5500), .ZN(n5508) );
  INV_X1 U6687 ( .A(n5502), .ZN(n5505) );
  MUX2_X1 U6688 ( .A(n5505), .B(n5504), .S(n5503), .Z(n5514) );
  NOR2_X1 U6689 ( .A1(n5528), .A2(n5514), .ZN(n5516) );
  XOR2_X1 U6690 ( .A(n5506), .B(n5516), .Z(n6007) );
  NOR2_X1 U6691 ( .A1(n6007), .A2(n6277), .ZN(n5507) );
  AOI211_X1 U6692 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5527), .A(n5508), .B(n5507), .ZN(n5509) );
  OAI211_X1 U6693 ( .C1(n6247), .C2(n5836), .A(n5510), .B(n5509), .ZN(U2808)
         );
  OAI21_X1 U6694 ( .B1(n5511), .B2(n5513), .A(n5512), .ZN(n5846) );
  AND2_X1 U6695 ( .A1(n5528), .A2(n5514), .ZN(n5515) );
  NOR2_X1 U6696 ( .A1(n5516), .A2(n5515), .ZN(n6019) );
  OAI21_X1 U6697 ( .B1(n6266), .B2(n5517), .A(n6264), .ZN(n5518) );
  AOI21_X1 U6698 ( .B1(n6250), .B2(EBX_REG_18__SCAN_IN), .A(n5518), .ZN(n5520)
         );
  NAND2_X1 U6699 ( .A1(n5527), .A2(REIP_REG_18__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U6700 ( .C1(n5521), .C2(REIP_REG_18__SCAN_IN), .A(n5520), .B(n5519), .ZN(n5523) );
  NOR2_X1 U6701 ( .A1(n6247), .A2(n5848), .ZN(n5522) );
  AOI211_X1 U6702 ( .C1(n6019), .C2(n6252), .A(n5523), .B(n5522), .ZN(n5524)
         );
  OAI21_X1 U6703 ( .B1(n5846), .B2(n6207), .A(n5524), .ZN(U2809) );
  XOR2_X1 U6704 ( .A(n5526), .B(n5525), .Z(n5858) );
  INV_X1 U6705 ( .A(n5527), .ZN(n5535) );
  INV_X1 U6706 ( .A(n5560), .ZN(n5546) );
  AOI21_X1 U6707 ( .B1(n5546), .B2(n5544), .A(REIP_REG_17__SCAN_IN), .ZN(n5534) );
  INV_X1 U6708 ( .A(n5528), .ZN(n5529) );
  AOI21_X1 U6709 ( .B1(n5530), .B2(n5542), .A(n5529), .ZN(n6027) );
  NAND2_X1 U6710 ( .A1(n6027), .A2(n6252), .ZN(n5533) );
  OAI21_X1 U6711 ( .B1(n6266), .B2(n3201), .A(n6264), .ZN(n5531) );
  AOI21_X1 U6712 ( .B1(n6250), .B2(EBX_REG_17__SCAN_IN), .A(n5531), .ZN(n5532)
         );
  OAI211_X1 U6713 ( .C1(n5535), .C2(n5534), .A(n5533), .B(n5532), .ZN(n5536)
         );
  AOI21_X1 U6714 ( .B1(n5855), .B2(n6259), .A(n5536), .ZN(n5537) );
  OAI21_X1 U6715 ( .B1(n5731), .B2(n6207), .A(n5537), .ZN(U2810) );
  OR2_X1 U6716 ( .A1(n5538), .A2(n5539), .ZN(n5540) );
  NAND2_X1 U6717 ( .A1(n5525), .A2(n5540), .ZN(n5866) );
  OAI21_X1 U6718 ( .B1(n5541), .B2(n5543), .A(n5542), .ZN(n5669) );
  INV_X1 U6719 ( .A(n5669), .ZN(n6034) );
  INV_X1 U6720 ( .A(n5580), .ZN(n5551) );
  INV_X1 U6721 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6750) );
  INV_X1 U6722 ( .A(n5544), .ZN(n5545) );
  OAI211_X1 U6723 ( .C1(REIP_REG_15__SCAN_IN), .C2(REIP_REG_16__SCAN_IN), .A(
        n5546), .B(n5545), .ZN(n5550) );
  OAI21_X1 U6724 ( .B1(n6266), .B2(n5547), .A(n6264), .ZN(n5548) );
  AOI21_X1 U6725 ( .B1(n6250), .B2(EBX_REG_16__SCAN_IN), .A(n5548), .ZN(n5549)
         );
  OAI211_X1 U6726 ( .C1(n5551), .C2(n6750), .A(n5550), .B(n5549), .ZN(n5553)
         );
  NOR2_X1 U6727 ( .A1(n6247), .A2(n5862), .ZN(n5552) );
  AOI211_X1 U6728 ( .C1(n6034), .C2(n6252), .A(n5553), .B(n5552), .ZN(n5554)
         );
  OAI21_X1 U6729 ( .B1(n5866), .B2(n6207), .A(n5554), .ZN(U2811) );
  AOI21_X1 U6730 ( .B1(n5557), .B2(n5556), .A(n5538), .ZN(n5670) );
  NAND2_X1 U6731 ( .A1(n5670), .A2(n6241), .ZN(n5567) );
  AOI21_X1 U6732 ( .B1(n6234), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6249), 
        .ZN(n5559) );
  NAND2_X1 U6733 ( .A1(n6250), .A2(EBX_REG_15__SCAN_IN), .ZN(n5558) );
  OAI211_X1 U6734 ( .C1(n5560), .C2(REIP_REG_15__SCAN_IN), .A(n5559), .B(n5558), .ZN(n5565) );
  NOR2_X1 U6735 ( .A1(n5561), .A2(n5562), .ZN(n5563) );
  OR2_X1 U6736 ( .A1(n5541), .A2(n5563), .ZN(n6053) );
  NOR2_X1 U6737 ( .A1(n6053), .A2(n6277), .ZN(n5564) );
  AOI211_X1 U6738 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5580), .A(n5565), .B(n5564), .ZN(n5566) );
  OAI211_X1 U6739 ( .C1(n6247), .C2(n5867), .A(n5567), .B(n5566), .ZN(U2812)
         );
  OAI21_X1 U6740 ( .B1(n5568), .B2(n5569), .A(n5556), .ZN(n5739) );
  INV_X1 U6741 ( .A(n5739), .ZN(n5881) );
  NAND2_X1 U6742 ( .A1(n5881), .A2(n6241), .ZN(n5582) );
  AOI21_X1 U6743 ( .B1(n6234), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6249), 
        .ZN(n5573) );
  NAND3_X1 U6744 ( .A1(n6263), .A2(n5571), .A3(n5570), .ZN(n5572) );
  OAI211_X1 U6745 ( .C1(n6269), .C2(n5672), .A(n5573), .B(n5572), .ZN(n5579)
         );
  INV_X1 U6746 ( .A(n5561), .ZN(n5577) );
  NAND2_X1 U6747 ( .A1(n5574), .A2(n5575), .ZN(n5576) );
  NAND2_X1 U6748 ( .A1(n5577), .A2(n5576), .ZN(n6066) );
  NOR2_X1 U6749 ( .A1(n6066), .A2(n6277), .ZN(n5578) );
  AOI211_X1 U6750 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5580), .A(n5579), .B(n5578), .ZN(n5581) );
  OAI211_X1 U6751 ( .C1(n6247), .C2(n5879), .A(n5582), .B(n5581), .ZN(U2813)
         );
  INV_X1 U6752 ( .A(n5583), .ZN(n5584) );
  AOI21_X1 U6753 ( .B1(n5585), .B2(n5246), .A(n5584), .ZN(n5906) );
  INV_X1 U6754 ( .A(n5906), .ZN(n5751) );
  NAND2_X1 U6755 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  NAND2_X1 U6756 ( .A1(n5690), .A2(n5588), .ZN(n6379) );
  OAI22_X1 U6757 ( .A1(n5904), .A2(n6247), .B1(n6277), .B2(n6379), .ZN(n5593)
         );
  INV_X1 U6758 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5591) );
  INV_X1 U6759 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6739) );
  NAND3_X1 U6760 ( .A1(n6263), .A2(n6739), .A3(n5589), .ZN(n5590) );
  OAI211_X1 U6761 ( .C1(n6266), .C2(n5591), .A(n6264), .B(n5590), .ZN(n5592)
         );
  AOI211_X1 U6762 ( .C1(n6250), .C2(EBX_REG_10__SCAN_IN), .A(n5593), .B(n5592), 
        .ZN(n5597) );
  NOR3_X1 U6763 ( .A1(n6232), .A2(REIP_REG_9__SCAN_IN), .A3(n5594), .ZN(n6214)
         );
  INV_X1 U6764 ( .A(n5594), .ZN(n5595) );
  NOR2_X1 U6765 ( .A1(n6232), .A2(n5595), .ZN(n6222) );
  INV_X1 U6766 ( .A(n6183), .ZN(n5616) );
  OR2_X1 U6767 ( .A1(n6222), .A2(n5616), .ZN(n6225) );
  OAI21_X1 U6768 ( .B1(n6214), .B2(n6225), .A(REIP_REG_10__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U6769 ( .C1(n5751), .C2(n6207), .A(n5597), .B(n5596), .ZN(U2817)
         );
  INV_X1 U6770 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6732) );
  INV_X1 U6771 ( .A(n5602), .ZN(n5598) );
  OAI21_X1 U6772 ( .B1(n5616), .B2(n5598), .A(n5615), .ZN(n6255) );
  OAI22_X1 U6773 ( .A1(n5599), .A2(n6247), .B1(n6732), .B2(n6255), .ZN(n5600)
         );
  AOI21_X1 U6774 ( .B1(n6252), .B2(n5601), .A(n5600), .ZN(n5606) );
  AOI22_X1 U6775 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6250), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6234), .ZN(n5604) );
  NAND3_X1 U6776 ( .A1(n6263), .A2(n5602), .A3(n6732), .ZN(n5603) );
  AND3_X1 U6777 ( .A1(n5604), .A2(n6264), .A3(n5603), .ZN(n5605) );
  OAI211_X1 U6778 ( .C1(n6207), .C2(n5607), .A(n5606), .B(n5605), .ZN(U2821)
         );
  AOI21_X1 U6779 ( .B1(n5609), .B2(n3093), .A(n6241), .ZN(n5653) );
  INV_X1 U6780 ( .A(n5653), .ZN(n6273) );
  NAND2_X1 U6781 ( .A1(n6273), .A2(n5610), .ZN(n5623) );
  NAND2_X1 U6782 ( .A1(n3093), .A2(n5611), .ZN(n6267) );
  INV_X1 U6783 ( .A(n6267), .ZN(n5644) );
  AOI22_X1 U6784 ( .A1(n5644), .A2(n5612), .B1(n6234), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5613) );
  OAI21_X1 U6785 ( .B1(n6269), .B2(n5614), .A(n5613), .ZN(n5620) );
  OAI21_X1 U6786 ( .B1(n5616), .B2(n6782), .A(n5615), .ZN(n5617) );
  NAND2_X1 U6787 ( .A1(n5617), .A2(REIP_REG_2__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U6788 ( .B1(n6232), .B2(n6262), .A(n6183), .ZN(n6258) );
  INV_X1 U6789 ( .A(n6258), .ZN(n5618) );
  AOI21_X1 U6790 ( .B1(n6728), .B2(n5631), .A(n5618), .ZN(n5619) );
  AOI211_X1 U6791 ( .C1(n5621), .C2(n6252), .A(n5620), .B(n5619), .ZN(n5622)
         );
  OAI211_X1 U6792 ( .C1(n6247), .C2(n5624), .A(n5623), .B(n5622), .ZN(U2824)
         );
  OAI21_X1 U6793 ( .B1(n6232), .B2(n6782), .A(n6869), .ZN(n5630) );
  AOI22_X1 U6794 ( .A1(n5644), .A2(n5625), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6234), .ZN(n5627) );
  NAND2_X1 U6795 ( .A1(n6250), .A2(EBX_REG_2__SCAN_IN), .ZN(n5626) );
  OAI211_X1 U6796 ( .C1(n6277), .C2(n6397), .A(n5627), .B(n5626), .ZN(n5629)
         );
  NOR2_X1 U6797 ( .A1(n6247), .A2(n6369), .ZN(n5628) );
  AOI211_X1 U6798 ( .C1(n5631), .C2(n5630), .A(n5629), .B(n5628), .ZN(n5632)
         );
  OAI21_X1 U6799 ( .B1(n5653), .B2(n6363), .A(n5632), .ZN(U2825) );
  INV_X1 U6800 ( .A(n4611), .ZN(n5633) );
  NAND3_X1 U6801 ( .A1(n5635), .A2(n5634), .A3(n5633), .ZN(n5636) );
  OAI21_X1 U6802 ( .B1(n6782), .B2(n6183), .A(n5636), .ZN(n5639) );
  OAI22_X1 U6803 ( .A1(n6232), .A2(REIP_REG_1__SCAN_IN), .B1(n5637), .B2(n6267), .ZN(n5638) );
  AOI211_X1 U6804 ( .C1(n6250), .C2(EBX_REG_1__SCAN_IN), .A(n5639), .B(n5638), 
        .ZN(n5641) );
  MUX2_X1 U6805 ( .A(n6247), .B(n6266), .S(PHYADDRPOINTER_REG_1__SCAN_IN), .Z(
        n5640) );
  OAI211_X1 U6806 ( .C1(n5653), .C2(n5642), .A(n5641), .B(n5640), .ZN(U2826)
         );
  AOI21_X1 U6807 ( .B1(n6247), .B2(n6266), .A(n5643), .ZN(n5650) );
  AOI22_X1 U6808 ( .A1(n5644), .A2(n6583), .B1(n6250), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5647) );
  NAND2_X1 U6809 ( .A1(n6252), .A2(n5645), .ZN(n5646) );
  OAI211_X1 U6810 ( .C1(n5648), .C2(n7077), .A(n5647), .B(n5646), .ZN(n5649)
         );
  NOR2_X1 U6811 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  OAI21_X1 U6812 ( .B1(n5653), .B2(n5652), .A(n5651), .ZN(U2827) );
  INV_X1 U6813 ( .A(n5654), .ZN(n5656) );
  OAI22_X1 U6814 ( .A1(n5656), .A2(n5697), .B1(n5655), .B2(n5696), .ZN(U2828)
         );
  AOI22_X1 U6815 ( .A1(n3114), .A2(n4499), .B1(n5684), .B2(EBX_REG_29__SCAN_IN), .ZN(n5657) );
  OAI21_X1 U6816 ( .B1(n5703), .B2(n5694), .A(n5657), .ZN(U2830) );
  INV_X1 U6817 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5658) );
  INV_X1 U6818 ( .A(n5775), .ZN(n5706) );
  OAI222_X1 U6819 ( .A1(n5932), .A2(n5697), .B1(n5658), .B2(n5696), .C1(n5706), 
        .C2(n5694), .ZN(U2832) );
  AOI22_X1 U6820 ( .A1(n5939), .A2(n4499), .B1(n5684), .B2(EBX_REG_26__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U6821 ( .B1(n5786), .B2(n5694), .A(n5659), .ZN(U2833) );
  AOI22_X1 U6822 ( .A1(n5953), .A2(n4499), .B1(n5684), .B2(EBX_REG_25__SCAN_IN), .ZN(n5660) );
  OAI21_X1 U6823 ( .B1(n5794), .B2(n5694), .A(n5660), .ZN(U2834) );
  INV_X1 U6824 ( .A(EBX_REG_24__SCAN_IN), .ZN(n7094) );
  OAI222_X1 U6825 ( .A1(n5956), .A2(n5697), .B1(n7094), .B2(n5696), .C1(n5799), 
        .C2(n5694), .ZN(U2835) );
  AOI22_X1 U6826 ( .A1(n5970), .A2(n4499), .B1(n5684), .B2(EBX_REG_23__SCAN_IN), .ZN(n5661) );
  OAI21_X1 U6827 ( .B1(n5715), .B2(n5694), .A(n5661), .ZN(U2836) );
  OAI222_X1 U6828 ( .A1(n5981), .A2(n5697), .B1(n5662), .B2(n5696), .C1(n5718), 
        .C2(n5694), .ZN(U2837) );
  AOI22_X1 U6829 ( .A1(n5987), .A2(n4499), .B1(n5684), .B2(EBX_REG_21__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U6830 ( .B1(n5721), .B2(n5694), .A(n5663), .ZN(U2838) );
  AOI22_X1 U6831 ( .A1(n6002), .A2(n4499), .B1(EBX_REG_20__SCAN_IN), .B2(n5684), .ZN(n5664) );
  OAI21_X1 U6832 ( .B1(n5824), .B2(n5694), .A(n5664), .ZN(U2839) );
  INV_X1 U6833 ( .A(n5838), .ZN(n5726) );
  OAI222_X1 U6834 ( .A1(n5726), .A2(n5694), .B1(n5697), .B2(n6007), .C1(n5696), 
        .C2(n5665), .ZN(U2840) );
  AOI22_X1 U6835 ( .A1(n6019), .A2(n4499), .B1(n5684), .B2(EBX_REG_18__SCAN_IN), .ZN(n5666) );
  OAI21_X1 U6836 ( .B1(n5846), .B2(n5694), .A(n5666), .ZN(U2841) );
  AOI22_X1 U6837 ( .A1(n6027), .A2(n4499), .B1(n5684), .B2(EBX_REG_17__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6838 ( .B1(n5731), .B2(n5694), .A(n5667), .ZN(U2842) );
  INV_X1 U6839 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5668) );
  OAI222_X1 U6840 ( .A1(n5669), .A2(n5697), .B1(n5668), .B2(n5696), .C1(n5866), 
        .C2(n5694), .ZN(U2843) );
  INV_X1 U6841 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5671) );
  INV_X1 U6842 ( .A(n5670), .ZN(n5875) );
  OAI222_X1 U6843 ( .A1(n6053), .A2(n5697), .B1(n5671), .B2(n5696), .C1(n5875), 
        .C2(n5694), .ZN(U2844) );
  OAI222_X1 U6844 ( .A1(n6066), .A2(n5697), .B1(n5672), .B2(n5696), .C1(n5739), 
        .C2(n5694), .ZN(U2845) );
  NAND2_X1 U6845 ( .A1(n5674), .A2(n5675), .ZN(n5676) );
  INV_X1 U6846 ( .A(n5574), .ZN(n5678) );
  AOI21_X1 U6847 ( .B1(n5679), .B2(n5682), .A(n5678), .ZN(n6185) );
  AOI22_X1 U6848 ( .A1(n6185), .A2(n4499), .B1(EBX_REG_13__SCAN_IN), .B2(n5684), .ZN(n5680) );
  OAI21_X1 U6849 ( .B1(n5889), .B2(n5694), .A(n5680), .ZN(U2846) );
  XOR2_X1 U6850 ( .A(n5681), .B(n3110), .Z(n5896) );
  OAI21_X1 U6851 ( .B1(n5688), .B2(n5683), .A(n5682), .ZN(n6194) );
  INV_X1 U6852 ( .A(n6194), .ZN(n6087) );
  AOI22_X1 U6853 ( .A1(n6087), .A2(n4499), .B1(n5684), .B2(EBX_REG_12__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6854 ( .B1(n6195), .B2(n5694), .A(n5685), .ZN(U2847) );
  AND2_X1 U6855 ( .A1(n5583), .A2(n5686), .ZN(n5687) );
  OR2_X1 U6856 ( .A1(n3110), .A2(n5687), .ZN(n6335) );
  INV_X1 U6857 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5693) );
  INV_X1 U6858 ( .A(n5688), .ZN(n5692) );
  NAND2_X1 U6859 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  NAND2_X1 U6860 ( .A1(n5692), .A2(n5691), .ZN(n6206) );
  OAI222_X1 U6861 ( .A1(n6335), .A2(n5694), .B1(n5696), .B2(n5693), .C1(n6206), 
        .C2(n5697), .ZN(U2848) );
  INV_X1 U6862 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5695) );
  OAI222_X1 U6863 ( .A1(n6379), .A2(n5697), .B1(n5696), .B2(n5695), .C1(n5694), 
        .C2(n5751), .ZN(U2849) );
  NAND2_X1 U6864 ( .A1(n5746), .A2(n5698), .ZN(n5700) );
  AOI22_X1 U6865 ( .A1(n5732), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5748), .ZN(n5699) );
  OAI21_X1 U6866 ( .B1(n5758), .B2(n5700), .A(n5699), .ZN(U2860) );
  AOI22_X1 U6867 ( .A1(n5732), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5748), .ZN(n5702) );
  NAND2_X1 U6868 ( .A1(n5733), .A2(DATAI_13_), .ZN(n5701) );
  OAI211_X1 U6869 ( .C1(n5703), .C2(n5747), .A(n5702), .B(n5701), .ZN(U2862)
         );
  AOI22_X1 U6870 ( .A1(n5732), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5748), .ZN(n5705) );
  NAND2_X1 U6871 ( .A1(n5733), .A2(DATAI_11_), .ZN(n5704) );
  OAI211_X1 U6872 ( .C1(n5706), .C2(n5747), .A(n5705), .B(n5704), .ZN(U2864)
         );
  AOI22_X1 U6873 ( .A1(n5732), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5748), .ZN(n5708) );
  NAND2_X1 U6874 ( .A1(n5733), .A2(DATAI_10_), .ZN(n5707) );
  OAI211_X1 U6875 ( .C1(n5786), .C2(n5747), .A(n5708), .B(n5707), .ZN(U2865)
         );
  AOI22_X1 U6876 ( .A1(n5732), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5748), .ZN(n5710) );
  NAND2_X1 U6877 ( .A1(n5733), .A2(DATAI_9_), .ZN(n5709) );
  OAI211_X1 U6878 ( .C1(n5794), .C2(n5747), .A(n5710), .B(n5709), .ZN(U2866)
         );
  AOI22_X1 U6879 ( .A1(n5732), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5748), .ZN(n5712) );
  NAND2_X1 U6880 ( .A1(n5733), .A2(DATAI_8_), .ZN(n5711) );
  OAI211_X1 U6881 ( .C1(n5799), .C2(n5747), .A(n5712), .B(n5711), .ZN(U2867)
         );
  AOI22_X1 U6882 ( .A1(n5732), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5748), .ZN(n5714) );
  NAND2_X1 U6883 ( .A1(n5733), .A2(DATAI_7_), .ZN(n5713) );
  OAI211_X1 U6884 ( .C1(n5715), .C2(n5747), .A(n5714), .B(n5713), .ZN(U2868)
         );
  AOI22_X1 U6885 ( .A1(n5732), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5748), .ZN(n5717) );
  NAND2_X1 U6886 ( .A1(n5733), .A2(DATAI_6_), .ZN(n5716) );
  OAI211_X1 U6887 ( .C1(n5718), .C2(n5747), .A(n5717), .B(n5716), .ZN(U2869)
         );
  AOI22_X1 U6888 ( .A1(n5732), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5748), .ZN(n5720) );
  NAND2_X1 U6889 ( .A1(n5733), .A2(DATAI_5_), .ZN(n5719) );
  OAI211_X1 U6890 ( .C1(n5721), .C2(n5747), .A(n5720), .B(n5719), .ZN(U2870)
         );
  AOI22_X1 U6891 ( .A1(n5732), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5748), .ZN(n5723) );
  NAND2_X1 U6892 ( .A1(n5733), .A2(DATAI_4_), .ZN(n5722) );
  OAI211_X1 U6893 ( .C1(n5824), .C2(n5747), .A(n5723), .B(n5722), .ZN(U2871)
         );
  AOI22_X1 U6894 ( .A1(n5732), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5748), .ZN(n5725) );
  NAND2_X1 U6895 ( .A1(n5733), .A2(DATAI_3_), .ZN(n5724) );
  OAI211_X1 U6896 ( .C1(n5726), .C2(n5747), .A(n5725), .B(n5724), .ZN(U2872)
         );
  AOI22_X1 U6897 ( .A1(n5732), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5748), .ZN(n5728) );
  NAND2_X1 U6898 ( .A1(n5733), .A2(DATAI_2_), .ZN(n5727) );
  OAI211_X1 U6899 ( .C1(n5846), .C2(n5747), .A(n5728), .B(n5727), .ZN(U2873)
         );
  AOI22_X1 U6900 ( .A1(n5732), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5748), .ZN(n5730) );
  NAND2_X1 U6901 ( .A1(n5733), .A2(DATAI_1_), .ZN(n5729) );
  OAI211_X1 U6902 ( .C1(n5731), .C2(n5747), .A(n5730), .B(n5729), .ZN(U2874)
         );
  AOI22_X1 U6903 ( .A1(n5732), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5748), .ZN(n5735) );
  NAND2_X1 U6904 ( .A1(n5733), .A2(DATAI_0_), .ZN(n5734) );
  OAI211_X1 U6905 ( .C1(n5866), .C2(n5747), .A(n5735), .B(n5734), .ZN(U2875)
         );
  AOI22_X1 U6906 ( .A1(n5749), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5748), .ZN(n5736) );
  OAI21_X1 U6907 ( .B1(n5875), .B2(n5747), .A(n5736), .ZN(U2876) );
  INV_X1 U6908 ( .A(DATAI_14_), .ZN(n5737) );
  OAI222_X1 U6909 ( .A1(n5739), .A2(n5747), .B1(n5746), .B2(n5738), .C1(n5737), 
        .C2(n5744), .ZN(U2877) );
  INV_X1 U6910 ( .A(DATAI_13_), .ZN(n5740) );
  OAI222_X1 U6911 ( .A1(n5889), .A2(n5747), .B1(n5746), .B2(n5741), .C1(n5740), 
        .C2(n5744), .ZN(U2878) );
  OAI222_X1 U6912 ( .A1(n5744), .A2(n5743), .B1(n5747), .B2(n6195), .C1(n5742), 
        .C2(n5746), .ZN(U2879) );
  INV_X1 U6913 ( .A(DATAI_11_), .ZN(n6823) );
  OAI222_X1 U6914 ( .A1(n6335), .A2(n5747), .B1(n5746), .B2(n5745), .C1(n5744), 
        .C2(n6823), .ZN(U2880) );
  AOI22_X1 U6915 ( .A1(n5749), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5748), .ZN(n5750) );
  OAI21_X1 U6916 ( .B1(n5751), .B2(n5747), .A(n5750), .ZN(U2881) );
  NAND2_X1 U6917 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5752)
         );
  OAI211_X1 U6918 ( .C1(n5754), .C2(n6370), .A(n5753), .B(n5752), .ZN(n5755)
         );
  AOI21_X1 U6919 ( .B1(n5756), .B2(n6366), .A(n5755), .ZN(n5757) );
  OAI21_X1 U6920 ( .B1(n5758), .B2(n6334), .A(n5757), .ZN(U2955) );
  OAI21_X1 U6921 ( .B1(n5761), .B2(n5760), .A(n5759), .ZN(n5762) );
  XNOR2_X1 U6922 ( .A(n5762), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5919)
         );
  NAND2_X1 U6923 ( .A1(n5763), .A2(n6350), .ZN(n5764) );
  NAND2_X1 U6924 ( .A1(n6377), .A2(REIP_REG_29__SCAN_IN), .ZN(n5914) );
  OAI211_X1 U6925 ( .C1(n6356), .C2(n5765), .A(n5764), .B(n5914), .ZN(n5766)
         );
  AOI21_X1 U6926 ( .B1(n5767), .B2(n6365), .A(n5766), .ZN(n5768) );
  OAI21_X1 U6927 ( .B1(n5919), .B2(n6339), .A(n5768), .ZN(U2957) );
  NAND2_X1 U6928 ( .A1(n3122), .A2(n5769), .ZN(n5770) );
  XNOR2_X1 U6929 ( .A(n5770), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5938)
         );
  NAND2_X1 U6930 ( .A1(n5771), .A2(n6350), .ZN(n5772) );
  NAND2_X1 U6931 ( .A1(n6377), .A2(REIP_REG_27__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U6932 ( .C1(n6356), .C2(n5773), .A(n5772), .B(n5930), .ZN(n5774)
         );
  AOI21_X1 U6933 ( .B1(n5775), .B2(n6365), .A(n5774), .ZN(n5776) );
  OAI21_X1 U6934 ( .B1(n5938), .B2(n6339), .A(n5776), .ZN(U2959) );
  NOR2_X1 U6935 ( .A1(n6396), .A2(n7062), .ZN(n5943) );
  NOR2_X1 U6936 ( .A1(n5777), .A2(n6370), .ZN(n5778) );
  AOI211_X1 U6937 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5943), 
        .B(n5778), .ZN(n5785) );
  INV_X1 U6938 ( .A(n5779), .ZN(n5781) );
  NAND2_X1 U6939 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  XNOR2_X1 U6940 ( .A(n5783), .B(n5782), .ZN(n5940) );
  NAND2_X1 U6941 ( .A1(n5940), .A2(n6366), .ZN(n5784) );
  OAI211_X1 U6942 ( .C1(n5786), .C2(n6334), .A(n5785), .B(n5784), .ZN(U2960)
         );
  OAI21_X1 U6943 ( .B1(n5789), .B2(n5788), .A(n5787), .ZN(n5947) );
  NAND2_X1 U6944 ( .A1(n5790), .A2(n6350), .ZN(n5791) );
  NAND2_X1 U6945 ( .A1(n6377), .A2(REIP_REG_25__SCAN_IN), .ZN(n5949) );
  OAI211_X1 U6946 ( .C1(n6356), .C2(n3193), .A(n5791), .B(n5949), .ZN(n5792)
         );
  AOI21_X1 U6947 ( .B1(n5947), .B2(n6366), .A(n5792), .ZN(n5793) );
  OAI21_X1 U6948 ( .B1(n5794), .B2(n6334), .A(n5793), .ZN(U2961) );
  NAND3_X1 U6949 ( .A1(n4407), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U6950 ( .A(n5798), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5963)
         );
  NAND2_X1 U6951 ( .A1(n6377), .A2(REIP_REG_24__SCAN_IN), .ZN(n5957) );
  OAI21_X1 U6952 ( .B1(n6356), .B2(n7044), .A(n5957), .ZN(n5801) );
  NOR2_X1 U6953 ( .A1(n5799), .A2(n6334), .ZN(n5800) );
  OAI21_X1 U6954 ( .B1(n5963), .B2(n6339), .A(n5803), .ZN(U2962) );
  NAND4_X1 U6955 ( .A1(n5820), .A2(n5976), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n4407), .ZN(n5804) );
  NAND2_X1 U6956 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  XNOR2_X1 U6957 ( .A(n5806), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5972)
         );
  NAND2_X1 U6958 ( .A1(n6377), .A2(REIP_REG_23__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U6959 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5807)
         );
  OAI211_X1 U6960 ( .C1(n5808), .C2(n6370), .A(n5965), .B(n5807), .ZN(n5809)
         );
  AOI21_X1 U6961 ( .B1(n5810), .B2(n6365), .A(n5809), .ZN(n5811) );
  OAI21_X1 U6962 ( .B1(n5972), .B2(n6339), .A(n5811), .ZN(U2963) );
  AOI21_X1 U6963 ( .B1(n5814), .B2(n5813), .A(n5812), .ZN(n5989) );
  NOR2_X1 U6964 ( .A1(n6396), .A2(n6756), .ZN(n5982) );
  AOI21_X1 U6965 ( .B1(n6358), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5982), 
        .ZN(n5815) );
  OAI21_X1 U6966 ( .B1(n5816), .B2(n6370), .A(n5815), .ZN(n5817) );
  AOI21_X1 U6967 ( .B1(n5818), .B2(n6365), .A(n5817), .ZN(n5819) );
  OAI21_X1 U6968 ( .B1(n5989), .B2(n6339), .A(n5819), .ZN(U2965) );
  OR2_X1 U6969 ( .A1(n5820), .A2(n5830), .ZN(n5822) );
  AOI21_X1 U6970 ( .B1(n5823), .B2(n5822), .A(n5821), .ZN(n6004) );
  INV_X1 U6971 ( .A(n5824), .ZN(n5828) );
  NAND2_X1 U6972 ( .A1(n6377), .A2(REIP_REG_20__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U6973 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5825)
         );
  OAI211_X1 U6974 ( .C1(n5826), .C2(n6370), .A(n5998), .B(n5825), .ZN(n5827)
         );
  AOI21_X1 U6975 ( .B1(n5828), .B2(n6365), .A(n5827), .ZN(n5829) );
  OAI21_X1 U6976 ( .B1(n6004), .B2(n6339), .A(n5829), .ZN(U2966) );
  INV_X1 U6977 ( .A(n5830), .ZN(n5832) );
  NAND2_X1 U6978 ( .A1(n5832), .A2(n5831), .ZN(n5834) );
  XOR2_X1 U6979 ( .A(n5834), .B(n5833), .Z(n6013) );
  NAND2_X1 U6980 ( .A1(n6377), .A2(REIP_REG_19__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U6981 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5835)
         );
  OAI211_X1 U6982 ( .C1(n6370), .C2(n5836), .A(n6005), .B(n5835), .ZN(n5837)
         );
  AOI21_X1 U6983 ( .B1(n5838), .B2(n6365), .A(n5837), .ZN(n5839) );
  OAI21_X1 U6984 ( .B1(n6013), .B2(n6339), .A(n5839), .ZN(U2967) );
  INV_X1 U6985 ( .A(n5840), .ZN(n5872) );
  NAND2_X1 U6986 ( .A1(n4407), .A2(n6031), .ZN(n5869) );
  INV_X1 U6987 ( .A(n5870), .ZN(n5841) );
  AOI21_X2 U6988 ( .B1(n5872), .B2(n5869), .A(n5841), .ZN(n5861) );
  NOR3_X1 U6989 ( .A1(n5861), .A2(n5853), .A3(n7026), .ZN(n5844) );
  NOR2_X1 U6990 ( .A1(n5852), .A2(n5842), .ZN(n5843) );
  MUX2_X1 U6991 ( .A(n5844), .B(n5843), .S(n4524), .Z(n5845) );
  XNOR2_X1 U6992 ( .A(n5845), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6021)
         );
  INV_X1 U6993 ( .A(n5846), .ZN(n5850) );
  NAND2_X1 U6994 ( .A1(n6377), .A2(REIP_REG_18__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U6995 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5847)
         );
  OAI211_X1 U6996 ( .C1(n6370), .C2(n5848), .A(n6014), .B(n5847), .ZN(n5849)
         );
  AOI21_X1 U6997 ( .B1(n5850), .B2(n6365), .A(n5849), .ZN(n5851) );
  OAI21_X1 U6998 ( .B1(n6021), .B2(n6339), .A(n5851), .ZN(U2968) );
  NAND2_X1 U6999 ( .A1(n5861), .A2(n5853), .ZN(n5854) );
  NAND2_X1 U7000 ( .A1(n6350), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U7001 ( .A1(n6377), .A2(REIP_REG_17__SCAN_IN), .ZN(n6023) );
  OAI211_X1 U7002 ( .C1(n6356), .C2(n3201), .A(n5856), .B(n6023), .ZN(n5857)
         );
  AOI21_X1 U7003 ( .B1(n5858), .B2(n6365), .A(n5857), .ZN(n5859) );
  OAI21_X1 U7004 ( .B1(n6029), .B2(n6339), .A(n5859), .ZN(U2969) );
  XNOR2_X1 U7005 ( .A(n4407), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5860)
         );
  XNOR2_X1 U7006 ( .A(n5861), .B(n5860), .ZN(n6030) );
  NAND2_X1 U7007 ( .A1(n6030), .A2(n6366), .ZN(n5865) );
  NOR2_X1 U7008 ( .A1(n6396), .A2(n6750), .ZN(n6033) );
  NOR2_X1 U7009 ( .A1(n6370), .A2(n5862), .ZN(n5863) );
  AOI211_X1 U7010 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6033), 
        .B(n5863), .ZN(n5864) );
  OAI211_X1 U7011 ( .C1(n6334), .C2(n5866), .A(n5865), .B(n5864), .ZN(U2970)
         );
  INV_X1 U7012 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U7013 ( .A1(n6396), .A2(n6985), .ZN(n6049) );
  NOR2_X1 U7014 ( .A1(n6370), .A2(n5867), .ZN(n5868) );
  AOI211_X1 U7015 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6049), 
        .B(n5868), .ZN(n5874) );
  NAND2_X1 U7016 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  XNOR2_X1 U7017 ( .A(n5872), .B(n5871), .ZN(n6047) );
  NAND2_X1 U7018 ( .A1(n6047), .A2(n6366), .ZN(n5873) );
  OAI211_X1 U7019 ( .C1(n5875), .C2(n6334), .A(n5874), .B(n5873), .ZN(U2971)
         );
  XNOR2_X1 U7020 ( .A(n4407), .B(n6062), .ZN(n5876) );
  XNOR2_X1 U7021 ( .A(n5877), .B(n5876), .ZN(n6070) );
  NAND2_X1 U7022 ( .A1(n6377), .A2(REIP_REG_14__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7023 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5878)
         );
  OAI211_X1 U7024 ( .C1(n6370), .C2(n5879), .A(n6065), .B(n5878), .ZN(n5880)
         );
  AOI21_X1 U7025 ( .B1(n5881), .B2(n6365), .A(n5880), .ZN(n5882) );
  OAI21_X1 U7026 ( .B1(n6339), .B2(n6070), .A(n5882), .ZN(U2972) );
  AND2_X1 U7027 ( .A1(n6377), .A2(REIP_REG_13__SCAN_IN), .ZN(n6075) );
  NOR2_X1 U7028 ( .A1(n6370), .A2(n6187), .ZN(n5883) );
  AOI211_X1 U7029 ( .C1(n6358), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6075), 
        .B(n5883), .ZN(n5888) );
  OAI21_X1 U7030 ( .B1(n5886), .B2(n5885), .A(n5884), .ZN(n6071) );
  NAND2_X1 U7031 ( .A1(n6071), .A2(n6366), .ZN(n5887) );
  OAI211_X1 U7032 ( .C1(n5889), .C2(n6334), .A(n5888), .B(n5887), .ZN(U2973)
         );
  NAND2_X1 U7033 ( .A1(n3123), .A2(n5898), .ZN(n6094) );
  NOR2_X1 U7034 ( .A1(n4407), .A2(n6099), .ZN(n6092) );
  AOI21_X1 U7035 ( .B1(n6094), .B2(n6090), .A(n6092), .ZN(n5892) );
  OAI21_X1 U7036 ( .B1(n4407), .B2(n6082), .A(n5890), .ZN(n5891) );
  XNOR2_X1 U7037 ( .A(n5892), .B(n5891), .ZN(n6089) );
  INV_X1 U7038 ( .A(n6198), .ZN(n5894) );
  NAND2_X1 U7039 ( .A1(n6377), .A2(REIP_REG_12__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7040 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5893)
         );
  OAI211_X1 U7041 ( .C1(n6370), .C2(n5894), .A(n6081), .B(n5893), .ZN(n5895)
         );
  AOI21_X1 U7042 ( .B1(n5896), .B2(n6365), .A(n5895), .ZN(n5897) );
  OAI21_X1 U7043 ( .B1(n6089), .B2(n6339), .A(n5897), .ZN(U2974) );
  INV_X1 U7044 ( .A(n5898), .ZN(n5900) );
  NOR2_X1 U7045 ( .A1(n5900), .A2(n5899), .ZN(n5902) );
  XOR2_X1 U7046 ( .A(n5902), .B(n5901), .Z(n6372) );
  AOI22_X1 U7047 ( .A1(n6358), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6377), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U7048 ( .B1(n5904), .B2(n6370), .A(n5903), .ZN(n5905) );
  AOI21_X1 U7049 ( .B1(n5906), .B2(n6365), .A(n5905), .ZN(n5907) );
  OAI21_X1 U7050 ( .B1(n6372), .B2(n6339), .A(n5907), .ZN(U2976) );
  XNOR2_X1 U7051 ( .A(n4407), .B(n7064), .ZN(n5908) );
  XNOR2_X1 U7052 ( .A(n5909), .B(n5908), .ZN(n6385) );
  NAND2_X1 U7053 ( .A1(n6385), .A2(n6366), .ZN(n5912) );
  OAI22_X1 U7054 ( .A1(n6356), .A2(n6981), .B1(n6396), .B2(n6737), .ZN(n5910)
         );
  AOI21_X1 U7055 ( .B1(n6350), .B2(n6212), .A(n5910), .ZN(n5911) );
  OAI211_X1 U7056 ( .C1(n6334), .C2(n6215), .A(n5912), .B(n5911), .ZN(U2977)
         );
  NAND2_X1 U7057 ( .A1(n5913), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5915) );
  OAI211_X1 U7058 ( .C1(n5916), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5915), .B(n5914), .ZN(n5917) );
  AOI21_X1 U7059 ( .B1(n3114), .B2(n6410), .A(n5917), .ZN(n5918) );
  OAI21_X1 U7060 ( .B1(n5919), .B2(n6101), .A(n5918), .ZN(U2989) );
  INV_X1 U7061 ( .A(n5920), .ZN(n5922) );
  NAND3_X1 U7062 ( .A1(n5936), .A2(n5922), .A3(n5921), .ZN(n5924) );
  OAI211_X1 U7063 ( .C1(n5931), .C2(n5925), .A(n5924), .B(n5923), .ZN(n5926)
         );
  AOI21_X1 U7064 ( .B1(n5927), .B2(n6410), .A(n5926), .ZN(n5928) );
  OAI21_X1 U7065 ( .B1(n5929), .B2(n6101), .A(n5928), .ZN(U2990) );
  INV_X1 U7066 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5935) );
  OAI21_X1 U7067 ( .B1(n5931), .B2(n5935), .A(n5930), .ZN(n5934) );
  NOR2_X1 U7068 ( .A1(n5932), .A2(n6398), .ZN(n5933) );
  AOI211_X1 U7069 ( .C1(n5936), .C2(n5935), .A(n5934), .B(n5933), .ZN(n5937)
         );
  OAI21_X1 U7070 ( .B1(n5938), .B2(n6101), .A(n5937), .ZN(U2991) );
  INV_X1 U7071 ( .A(n5939), .ZN(n5946) );
  NAND2_X1 U7072 ( .A1(n5940), .A2(n6412), .ZN(n5945) );
  INV_X1 U7073 ( .A(n5958), .ZN(n5948) );
  XNOR2_X1 U7074 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5941) );
  NOR2_X1 U7075 ( .A1(n5951), .A2(n5941), .ZN(n5942) );
  AOI211_X1 U7076 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5948), .A(n5943), .B(n5942), .ZN(n5944) );
  OAI211_X1 U7077 ( .C1(n6398), .C2(n5946), .A(n5945), .B(n5944), .ZN(U2992)
         );
  INV_X1 U7078 ( .A(n5947), .ZN(n5955) );
  NAND2_X1 U7079 ( .A1(n5948), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5950) );
  OAI211_X1 U7080 ( .C1(n5951), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5950), .B(n5949), .ZN(n5952) );
  AOI21_X1 U7081 ( .B1(n5953), .B2(n6410), .A(n5952), .ZN(n5954) );
  OAI21_X1 U7082 ( .B1(n5955), .B2(n6101), .A(n5954), .ZN(U2993) );
  INV_X1 U7083 ( .A(n5956), .ZN(n5961) );
  AOI21_X1 U7084 ( .B1(n5964), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5959) );
  OAI21_X1 U7085 ( .B1(n5959), .B2(n5958), .A(n5957), .ZN(n5960) );
  AOI21_X1 U7086 ( .B1(n5961), .B2(n6410), .A(n5960), .ZN(n5962) );
  OAI21_X1 U7087 ( .B1(n5963), .B2(n6101), .A(n5962), .ZN(U2994) );
  NAND2_X1 U7088 ( .A1(n5964), .A2(n5967), .ZN(n5966) );
  OAI211_X1 U7089 ( .C1(n5968), .C2(n5967), .A(n5966), .B(n5965), .ZN(n5969)
         );
  AOI21_X1 U7090 ( .B1(n5970), .B2(n6410), .A(n5969), .ZN(n5971) );
  OAI21_X1 U7091 ( .B1(n5972), .B2(n6101), .A(n5971), .ZN(U2995) );
  INV_X1 U7092 ( .A(n5974), .ZN(n5983) );
  NOR3_X1 U7093 ( .A1(n5985), .A2(n5976), .A3(n5975), .ZN(n5977) );
  AOI211_X1 U7094 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5983), .A(n5978), .B(n5977), .ZN(n5979) );
  OAI211_X1 U7095 ( .C1(n6398), .C2(n5981), .A(n5980), .B(n5979), .ZN(U2996)
         );
  AOI21_X1 U7096 ( .B1(n5983), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5982), 
        .ZN(n5984) );
  OAI21_X1 U7097 ( .B1(n5985), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5984), 
        .ZN(n5986) );
  AOI21_X1 U7098 ( .B1(n5987), .B2(n6410), .A(n5986), .ZN(n5988) );
  OAI21_X1 U7099 ( .B1(n5989), .B2(n6101), .A(n5988), .ZN(U2997) );
  INV_X1 U7100 ( .A(n6011), .ZN(n5992) );
  NOR3_X1 U7101 ( .A1(n5992), .A2(n5991), .A3(n5990), .ZN(n6001) );
  INV_X1 U7102 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7103 ( .B1(n5993), .B2(n7026), .A(n6039), .ZN(n5994) );
  AND2_X1 U7104 ( .A1(n5995), .A2(n5994), .ZN(n6025) );
  NAND2_X1 U7105 ( .A1(n6392), .A2(n7026), .ZN(n5996) );
  AND2_X1 U7106 ( .A1(n6025), .A2(n5996), .ZN(n6017) );
  INV_X1 U7107 ( .A(n6017), .ZN(n5997) );
  AOI21_X1 U7108 ( .B1(n6016), .B2(n6415), .A(n5997), .ZN(n6006) );
  OAI21_X1 U7109 ( .B1(n6006), .B2(n5999), .A(n5998), .ZN(n6000) );
  AOI211_X1 U7110 ( .C1(n6002), .C2(n6410), .A(n6001), .B(n6000), .ZN(n6003)
         );
  OAI21_X1 U7111 ( .B1(n6004), .B2(n6101), .A(n6003), .ZN(U2998) );
  OAI21_X1 U7112 ( .B1(n6006), .B2(n6010), .A(n6005), .ZN(n6009) );
  NOR2_X1 U7113 ( .A1(n6007), .A2(n6398), .ZN(n6008) );
  AOI211_X1 U7114 ( .C1(n6011), .C2(n6010), .A(n6009), .B(n6008), .ZN(n6012)
         );
  OAI21_X1 U7115 ( .B1(n6013), .B2(n6101), .A(n6012), .ZN(U2999) );
  NAND3_X1 U7116 ( .A1(n6022), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6016), .ZN(n6015) );
  OAI211_X1 U7117 ( .C1(n6017), .C2(n6016), .A(n6015), .B(n6014), .ZN(n6018)
         );
  AOI21_X1 U7118 ( .B1(n6019), .B2(n6410), .A(n6018), .ZN(n6020) );
  OAI21_X1 U7119 ( .B1(n6021), .B2(n6101), .A(n6020), .ZN(U3000) );
  NAND2_X1 U7120 ( .A1(n6022), .A2(n7026), .ZN(n6024) );
  OAI211_X1 U7121 ( .C1(n6025), .C2(n7026), .A(n6024), .B(n6023), .ZN(n6026)
         );
  AOI21_X1 U7122 ( .B1(n6027), .B2(n6410), .A(n6026), .ZN(n6028) );
  OAI21_X1 U7123 ( .B1(n6029), .B2(n6101), .A(n6028), .ZN(U3001) );
  INV_X1 U7124 ( .A(n6030), .ZN(n6046) );
  INV_X1 U7125 ( .A(n6042), .ZN(n6035) );
  NOR4_X1 U7126 ( .A1(n6084), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6031), 
        .A4(n6035), .ZN(n6032) );
  AOI211_X1 U7127 ( .C1(n6034), .C2(n6410), .A(n6033), .B(n6032), .ZN(n6045)
         );
  NOR3_X1 U7128 ( .A1(n6084), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6035), 
        .ZN(n6048) );
  INV_X1 U7129 ( .A(n6415), .ZN(n6043) );
  NAND2_X1 U7130 ( .A1(n6037), .A2(n6036), .ZN(n6041) );
  NAND2_X1 U7131 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U7132 ( .A1(n6041), .A2(n6040), .ZN(n6079) );
  INV_X1 U7133 ( .A(n6079), .ZN(n6095) );
  OAI21_X1 U7134 ( .B1(n6043), .B2(n6042), .A(n6095), .ZN(n6050) );
  OAI21_X1 U7135 ( .B1(n6048), .B2(n6050), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n6044) );
  OAI211_X1 U7136 ( .C1(n6046), .C2(n6101), .A(n6045), .B(n6044), .ZN(U3002)
         );
  NAND2_X1 U7137 ( .A1(n6047), .A2(n6412), .ZN(n6052) );
  AOI211_X1 U7138 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6050), .A(n6049), .B(n6048), .ZN(n6051) );
  OAI211_X1 U7139 ( .C1(n6398), .C2(n6053), .A(n6052), .B(n6051), .ZN(U3003)
         );
  NOR2_X1 U7140 ( .A1(n6055), .A2(n6054), .ZN(n6061) );
  INV_X1 U7141 ( .A(n6060), .ZN(n6056) );
  NAND2_X1 U7142 ( .A1(n6056), .A2(n6072), .ZN(n6078) );
  INV_X1 U7143 ( .A(n6416), .ZN(n6057) );
  NOR2_X1 U7144 ( .A1(n6057), .A2(n6063), .ZN(n6058) );
  AOI211_X1 U7145 ( .C1(n6060), .C2(n6059), .A(n6058), .B(n6079), .ZN(n6073)
         );
  OAI21_X1 U7146 ( .B1(n6061), .B2(n6078), .A(n6073), .ZN(n6068) );
  NAND3_X1 U7147 ( .A1(n6098), .A2(n6063), .A3(n6062), .ZN(n6064) );
  OAI211_X1 U7148 ( .C1(n6066), .C2(n6398), .A(n6065), .B(n6064), .ZN(n6067)
         );
  AOI21_X1 U7149 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6068), .A(n6067), 
        .ZN(n6069) );
  OAI21_X1 U7150 ( .B1(n6070), .B2(n6101), .A(n6069), .ZN(U3004) );
  NAND2_X1 U7151 ( .A1(n6071), .A2(n6412), .ZN(n6077) );
  NOR2_X1 U7152 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  AOI211_X1 U7153 ( .C1(n6410), .C2(n6185), .A(n6075), .B(n6074), .ZN(n6076)
         );
  OAI211_X1 U7154 ( .C1(n6084), .C2(n6078), .A(n6077), .B(n6076), .ZN(U3005)
         );
  AOI221_X1 U7155 ( .B1(n6395), .B2(n6099), .C1(n6080), .C2(n6099), .A(n6079), 
        .ZN(n6083) );
  OAI21_X1 U7156 ( .B1(n6083), .B2(n6082), .A(n6081), .ZN(n6086) );
  NOR3_X1 U7157 ( .A1(n6084), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n6099), 
        .ZN(n6085) );
  AOI211_X1 U7158 ( .C1(n6410), .C2(n6087), .A(n6086), .B(n6085), .ZN(n6088)
         );
  OAI21_X1 U7159 ( .B1(n6089), .B2(n6101), .A(n6088), .ZN(U3006) );
  INV_X1 U7160 ( .A(n6090), .ZN(n6091) );
  NOR2_X1 U7161 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  XNOR2_X1 U7162 ( .A(n6094), .B(n6093), .ZN(n6340) );
  NOR2_X1 U7163 ( .A1(n6095), .A2(n6099), .ZN(n6097) );
  OAI22_X1 U7164 ( .A1(n6206), .A2(n6398), .B1(n6396), .B2(n6741), .ZN(n6096)
         );
  AOI211_X1 U7165 ( .C1(n6099), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6100)
         );
  OAI21_X1 U7166 ( .B1(n6340), .B2(n6101), .A(n6100), .ZN(U3007) );
  NAND2_X1 U7167 ( .A1(n6102), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6110)
         );
  NAND2_X1 U7168 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6103) );
  OAI211_X1 U7169 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6104), .B(n6103), .ZN(n6109) );
  NOR2_X1 U7170 ( .A1(n6398), .A2(n6276), .ZN(n6105) );
  AOI211_X1 U7171 ( .C1(n6107), .C2(n6412), .A(n6106), .B(n6105), .ZN(n6108)
         );
  NAND3_X1 U7172 ( .A1(n6110), .A2(n6109), .A3(n6108), .ZN(U3014) );
  INV_X1 U7173 ( .A(n6111), .ZN(n6112) );
  OAI22_X1 U7174 ( .A1(n6114), .A2(n6113), .B1(n6112), .B2(n6145), .ZN(n6116)
         );
  MUX2_X1 U7175 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6116), .S(n6115), 
        .Z(U3456) );
  AOI21_X1 U7176 ( .B1(n6117), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n7028), 
        .ZN(n6118) );
  AND2_X1 U7177 ( .A1(n6119), .A2(n6118), .ZN(n6122) );
  INV_X1 U7178 ( .A(n6122), .ZN(n6124) );
  AOI211_X1 U7179 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6122), .A(n6121), .B(n6120), .ZN(n6123) );
  AOI21_X1 U7180 ( .B1(n6461), .B2(n6124), .A(n6123), .ZN(n6125) );
  OAI21_X1 U7181 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6126), .A(n6125), 
        .ZN(n6127) );
  OAI21_X1 U7182 ( .B1(n6128), .B2(n6827), .A(n6127), .ZN(n6129) );
  OAI21_X1 U7183 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6130), .A(n6129), 
        .ZN(n6139) );
  AOI21_X1 U7184 ( .B1(n6130), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7185 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6131), 
        .ZN(n6132) );
  NAND4_X1 U7186 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n6136)
         );
  AOI211_X1 U7187 ( .C1(n6139), .C2(n6138), .A(n6137), .B(n6136), .ZN(n6153)
         );
  INV_X1 U7188 ( .A(n6140), .ZN(n6142) );
  AOI22_X1 U7189 ( .A1(n6153), .A2(n6154), .B1(n6300), .B2(READY_N), .ZN(n6141) );
  AOI21_X1 U7190 ( .B1(n6143), .B2(n6142), .A(n6141), .ZN(n6780) );
  INV_X1 U7191 ( .A(n6780), .ZN(n6144) );
  OAI21_X1 U7192 ( .B1(n6145), .B2(n6713), .A(n6144), .ZN(n6146) );
  AOI21_X1 U7193 ( .B1(READY_N), .B2(n6592), .A(n6780), .ZN(n6161) );
  MUX2_X1 U7194 ( .A(n6146), .B(n6161), .S(STATE2_REG_0__SCAN_IN), .Z(n6151)
         );
  INV_X1 U7195 ( .A(n6147), .ZN(n6148) );
  AOI21_X1 U7196 ( .B1(n6149), .B2(n6779), .A(n6148), .ZN(n6150) );
  OAI211_X1 U7197 ( .C1(n6153), .C2(n6152), .A(n6151), .B(n6150), .ZN(U3148)
         );
  NAND2_X1 U7198 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n6160) );
  NOR2_X1 U7199 ( .A1(READY_N), .A2(n7027), .ZN(n6715) );
  AOI21_X1 U7200 ( .B1(n6155), .B2(n6715), .A(n6154), .ZN(n6157) );
  MUX2_X1 U7201 ( .A(n6157), .B(n6156), .S(n6780), .Z(n6158) );
  OAI211_X1 U7202 ( .C1(n6161), .C2(n6160), .A(n6159), .B(n6158), .ZN(U3149)
         );
  AND2_X1 U7203 ( .A1(n6303), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U7204 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6163) );
  OAI21_X1 U7205 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6163), .A(n6800), .ZN(n6162)
         );
  OAI21_X1 U7206 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6800), .A(n6162), .ZN(
        U2791) );
  OAI21_X1 U7207 ( .B1(n6163), .B2(BS16_N), .A(n6778), .ZN(n6776) );
  OAI21_X1 U7208 ( .B1(n6778), .B2(n6467), .A(n6776), .ZN(U2792) );
  OAI21_X1 U7209 ( .B1(n6165), .B2(n6164), .A(n6339), .ZN(U2793) );
  INV_X1 U7210 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6777) );
  INV_X1 U7211 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6166) );
  NOR2_X1 U7212 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6818) );
  NOR4_X1 U7213 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_30__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6801) );
  OAI211_X1 U7214 ( .C1(n6777), .C2(n6166), .A(n6818), .B(n6801), .ZN(n6174)
         );
  OR4_X1 U7215 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n6173) );
  INV_X1 U7216 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n7045) );
  INV_X1 U7217 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7033) );
  INV_X1 U7218 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6878) );
  INV_X1 U7219 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6897) );
  NAND4_X1 U7220 ( .A1(n7045), .A2(n7033), .A3(n6878), .A4(n6897), .ZN(n6172)
         );
  NOR4_X1 U7221 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U7222 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(
        n6169) );
  NOR4_X1 U7223 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6168) );
  NOR4_X1 U7224 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6167) );
  NAND4_X1 U7225 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n6171)
         );
  INV_X1 U7226 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6923) );
  NOR3_X1 U7227 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6176) );
  OAI21_X1 U7228 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6176), .A(n6785), .ZN(n6175)
         );
  OAI21_X1 U7229 ( .B1(n6785), .B2(n6923), .A(n6175), .ZN(U2794) );
  AOI21_X1 U7230 ( .B1(n6782), .B2(n6777), .A(n6176), .ZN(n6178) );
  INV_X1 U7231 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6177) );
  INV_X1 U7232 ( .A(n6785), .ZN(n6787) );
  AOI22_X1 U7233 ( .A1(n6785), .A2(n6178), .B1(n6177), .B2(n6787), .ZN(U2795)
         );
  NOR3_X1 U7234 ( .A1(n6232), .A2(REIP_REG_13__SCAN_IN), .A3(n6179), .ZN(n6180) );
  AOI211_X1 U7235 ( .C1(n6250), .C2(EBX_REG_13__SCAN_IN), .A(n6249), .B(n6180), 
        .ZN(n6191) );
  INV_X1 U7236 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6743) );
  NAND3_X1 U7237 ( .A1(n6263), .A2(n6181), .A3(n6743), .ZN(n6193) );
  INV_X1 U7238 ( .A(n6181), .ZN(n6182) );
  NAND2_X1 U7239 ( .A1(n6263), .A2(n6182), .ZN(n6203) );
  NAND2_X1 U7240 ( .A1(n6183), .A2(n6203), .ZN(n6202) );
  INV_X1 U7241 ( .A(n6202), .ZN(n6201) );
  AOI21_X1 U7242 ( .B1(n6193), .B2(n6201), .A(n6746), .ZN(n6184) );
  AOI21_X1 U7243 ( .B1(n6185), .B2(n6252), .A(n6184), .ZN(n6186) );
  OAI21_X1 U7244 ( .B1(n6247), .B2(n6187), .A(n6186), .ZN(n6188) );
  AOI21_X1 U7245 ( .B1(n6189), .B2(n6241), .A(n6188), .ZN(n6190) );
  OAI211_X1 U7246 ( .C1(n6192), .C2(n6266), .A(n6191), .B(n6190), .ZN(U2814)
         );
  OAI211_X1 U7247 ( .C1(n6266), .C2(n3736), .A(n6264), .B(n6193), .ZN(n6197)
         );
  OAI22_X1 U7248 ( .A1(n6195), .A2(n6207), .B1(n6277), .B2(n6194), .ZN(n6196)
         );
  AOI211_X1 U7249 ( .C1(EBX_REG_12__SCAN_IN), .C2(n6250), .A(n6197), .B(n6196), 
        .ZN(n6200) );
  NAND2_X1 U7250 ( .A1(n6198), .A2(n6259), .ZN(n6199) );
  OAI211_X1 U7251 ( .C1(n6201), .C2(n6743), .A(n6200), .B(n6199), .ZN(U2815)
         );
  AOI22_X1 U7252 ( .A1(n6332), .A2(n6259), .B1(REIP_REG_11__SCAN_IN), .B2(
        n6202), .ZN(n6211) );
  OAI22_X1 U7253 ( .A1(n6951), .A2(n6266), .B1(n6204), .B2(n6203), .ZN(n6205)
         );
  AOI211_X1 U7254 ( .C1(n6250), .C2(EBX_REG_11__SCAN_IN), .A(n6249), .B(n6205), 
        .ZN(n6210) );
  OAI22_X1 U7255 ( .A1(n6335), .A2(n6207), .B1(n6277), .B2(n6206), .ZN(n6208)
         );
  INV_X1 U7256 ( .A(n6208), .ZN(n6209) );
  NAND3_X1 U7257 ( .A1(n6211), .A2(n6210), .A3(n6209), .ZN(U2816) );
  AOI22_X1 U7258 ( .A1(n6212), .A2(n6259), .B1(n6252), .B2(n6384), .ZN(n6219)
         );
  OAI21_X1 U7259 ( .B1(n6266), .B2(n6981), .A(n6264), .ZN(n6213) );
  AOI211_X1 U7260 ( .C1(n6250), .C2(EBX_REG_9__SCAN_IN), .A(n6214), .B(n6213), 
        .ZN(n6218) );
  INV_X1 U7261 ( .A(n6215), .ZN(n6216) );
  AOI22_X1 U7262 ( .A1(n6241), .A2(n6216), .B1(REIP_REG_9__SCAN_IN), .B2(n6225), .ZN(n6217) );
  NAND3_X1 U7263 ( .A1(n6219), .A2(n6218), .A3(n6217), .ZN(U2818) );
  AOI22_X1 U7264 ( .A1(n6221), .A2(n6259), .B1(n6252), .B2(n6220), .ZN(n6230)
         );
  AOI22_X1 U7265 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6234), .B1(n6223), 
        .B2(n6222), .ZN(n6229) );
  AOI21_X1 U7266 ( .B1(n6250), .B2(EBX_REG_8__SCAN_IN), .A(n6249), .ZN(n6228)
         );
  INV_X1 U7267 ( .A(n6224), .ZN(n6226) );
  AOI22_X1 U7268 ( .A1(n6241), .A2(n6226), .B1(REIP_REG_8__SCAN_IN), .B2(n6225), .ZN(n6227) );
  NAND4_X1 U7269 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(U2819)
         );
  INV_X1 U7270 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6244) );
  NOR3_X1 U7271 ( .A1(n6232), .A2(REIP_REG_7__SCAN_IN), .A3(n6231), .ZN(n6233)
         );
  AOI211_X1 U7272 ( .C1(n6234), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6249), 
        .B(n6233), .ZN(n6243) );
  INV_X1 U7273 ( .A(n6235), .ZN(n6342) );
  INV_X1 U7274 ( .A(n6255), .ZN(n6236) );
  AOI21_X1 U7275 ( .B1(n6263), .B2(n6732), .A(n6236), .ZN(n6238) );
  OAI22_X1 U7276 ( .A1(n6238), .A2(n6969), .B1(n6277), .B2(n6237), .ZN(n6240)
         );
  NOR2_X1 U7277 ( .A1(n6247), .A2(n6341), .ZN(n6239) );
  AOI211_X1 U7278 ( .C1(n6342), .C2(n6241), .A(n6240), .B(n6239), .ZN(n6242)
         );
  OAI211_X1 U7279 ( .C1(n6244), .C2(n6269), .A(n6243), .B(n6242), .ZN(U2820)
         );
  INV_X1 U7280 ( .A(n6245), .ZN(n6246) );
  AOI21_X1 U7281 ( .B1(n6263), .B2(n6246), .A(REIP_REG_5__SCAN_IN), .ZN(n6256)
         );
  OAI22_X1 U7282 ( .A1(n6357), .A2(n6266), .B1(n6349), .B2(n6247), .ZN(n6248)
         );
  AOI211_X1 U7283 ( .C1(n6250), .C2(EBX_REG_5__SCAN_IN), .A(n6249), .B(n6248), 
        .ZN(n6254) );
  AOI22_X1 U7284 ( .A1(n6273), .A2(n6352), .B1(n6252), .B2(n6251), .ZN(n6253)
         );
  OAI211_X1 U7285 ( .C1(n6256), .C2(n6255), .A(n6254), .B(n6253), .ZN(U2822)
         );
  INV_X1 U7286 ( .A(n6257), .ZN(n6260) );
  AOI22_X1 U7287 ( .A1(n6260), .A2(n6259), .B1(REIP_REG_4__SCAN_IN), .B2(n6258), .ZN(n6275) );
  INV_X1 U7288 ( .A(n6261), .ZN(n6272) );
  NAND3_X1 U7289 ( .A1(n6263), .A2(n6262), .A3(n6727), .ZN(n6265) );
  OAI211_X1 U7290 ( .C1(n6266), .C2(n6864), .A(n6265), .B(n6264), .ZN(n6271)
         );
  OAI22_X1 U7291 ( .A1(n6269), .A2(n6925), .B1(n6268), .B2(n6267), .ZN(n6270)
         );
  AOI211_X1 U7292 ( .C1(n6273), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6274)
         );
  OAI211_X1 U7293 ( .C1(n6277), .C2(n6276), .A(n6275), .B(n6274), .ZN(U2823)
         );
  INV_X1 U7294 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6928) );
  AOI22_X1 U7295 ( .A1(n6282), .A2(EAX_REG_29__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U7296 ( .B1(n6306), .B2(n6928), .A(n6278), .ZN(U2894) );
  INV_X1 U7297 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6929) );
  AOI22_X1 U7298 ( .A1(n6282), .A2(EAX_REG_27__SCAN_IN), .B1(n6300), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U7299 ( .B1(n6929), .B2(n6299), .A(n6279), .ZN(U2896) );
  INV_X1 U7300 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n7095) );
  AOI22_X1 U7301 ( .A1(n6282), .A2(EAX_REG_26__SCAN_IN), .B1(n6300), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6280) );
  OAI21_X1 U7302 ( .B1(n7095), .B2(n6299), .A(n6280), .ZN(U2897) );
  INV_X1 U7303 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n7057) );
  AOI22_X1 U7304 ( .A1(n6282), .A2(EAX_REG_23__SCAN_IN), .B1(n6300), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n6281) );
  OAI21_X1 U7305 ( .B1(n7057), .B2(n6299), .A(n6281), .ZN(U2900) );
  AOI22_X1 U7306 ( .A1(n6282), .A2(EAX_REG_19__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6283) );
  OAI21_X1 U7307 ( .B1(n6306), .B2(n7000), .A(n6283), .ZN(U2904) );
  INV_X1 U7308 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6331) );
  AOI22_X1 U7309 ( .A1(n6300), .A2(LWORD_REG_15__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7310 ( .B1(n6331), .B2(n6302), .A(n6284), .ZN(U2908) );
  INV_X1 U7311 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n7011) );
  INV_X1 U7312 ( .A(n6302), .ZN(n6304) );
  AOI22_X1 U7313 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6304), .B1(n6300), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6285) );
  OAI21_X1 U7314 ( .B1(n7011), .B2(n6299), .A(n6285), .ZN(U2909) );
  INV_X1 U7315 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7316 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6304), .B1(n6303), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7317 ( .B1(n6306), .B2(n6931), .A(n6286), .ZN(U2910) );
  AOI22_X1 U7318 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6304), .B1(n6303), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7319 ( .B1(n6306), .B2(n7015), .A(n6287), .ZN(U2911) );
  INV_X1 U7320 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U7321 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6304), .B1(n6303), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6288) );
  OAI21_X1 U7322 ( .B1(n6306), .B2(n6903), .A(n6288), .ZN(U2912) );
  INV_X1 U7323 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U7324 ( .A1(n6300), .A2(LWORD_REG_10__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6289) );
  OAI21_X1 U7325 ( .B1(n6290), .B2(n6302), .A(n6289), .ZN(U2913) );
  AOI22_X1 U7326 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6304), .B1(n6303), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6291) );
  OAI21_X1 U7327 ( .B1(n6306), .B2(n7092), .A(n6291), .ZN(U2914) );
  AOI222_X1 U7328 ( .A1(n6300), .A2(LWORD_REG_8__SCAN_IN), .B1(n6304), .B2(
        EAX_REG_8__SCAN_IN), .C1(DATAO_REG_8__SCAN_IN), .C2(n6303), .ZN(n6292)
         );
  INV_X1 U7329 ( .A(n6292), .ZN(U2915) );
  AOI22_X1 U7330 ( .A1(n6300), .A2(LWORD_REG_7__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7331 ( .B1(n3672), .B2(n6302), .A(n6293), .ZN(U2916) );
  AOI22_X1 U7332 ( .A1(n6300), .A2(LWORD_REG_6__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6294) );
  OAI21_X1 U7333 ( .B1(n4650), .B2(n6302), .A(n6294), .ZN(U2917) );
  INV_X1 U7334 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6988) );
  INV_X1 U7335 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6888) );
  OAI222_X1 U7336 ( .A1(n6299), .A2(n6988), .B1(n6302), .B2(n6295), .C1(n6306), 
        .C2(n6888), .ZN(U2918) );
  AOI22_X1 U7337 ( .A1(n6300), .A2(LWORD_REG_4__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7338 ( .B1(n6297), .B2(n6302), .A(n6296), .ZN(U2919) );
  AOI222_X1 U7339 ( .A1(n6303), .A2(DATAO_REG_3__SCAN_IN), .B1(n6304), .B2(
        EAX_REG_3__SCAN_IN), .C1(n6300), .C2(LWORD_REG_3__SCAN_IN), .ZN(n6298)
         );
  INV_X1 U7340 ( .A(n6298), .ZN(U2920) );
  INV_X1 U7341 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n7080) );
  INV_X1 U7342 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6879) );
  OAI222_X1 U7343 ( .A1(n6306), .A2(n7080), .B1(n6302), .B2(n6952), .C1(n6879), 
        .C2(n6299), .ZN(U2921) );
  AOI22_X1 U7344 ( .A1(n6300), .A2(LWORD_REG_1__SCAN_IN), .B1(n6303), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U7345 ( .B1(n4648), .B2(n6302), .A(n6301), .ZN(U2922) );
  AOI22_X1 U7346 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6304), .B1(n6303), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6305) );
  OAI21_X1 U7347 ( .B1(n6306), .B2(n4651), .A(n6305), .ZN(U2923) );
  INV_X1 U7348 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U7349 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_1_), .ZN(n6307) );
  OAI21_X1 U7350 ( .B1(n6308), .B2(n6330), .A(n6307), .ZN(U2925) );
  AOI22_X1 U7351 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_2_), .ZN(n6309) );
  OAI21_X1 U7352 ( .B1(n6906), .B2(n6330), .A(n6309), .ZN(U2926) );
  INV_X1 U7353 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6311) );
  AOI22_X1 U7354 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_4_), .ZN(n6310) );
  OAI21_X1 U7355 ( .B1(n6311), .B2(n6330), .A(n6310), .ZN(U2928) );
  INV_X1 U7356 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7024) );
  AOI22_X1 U7357 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_5_), .ZN(n6312) );
  OAI21_X1 U7358 ( .B1(n7024), .B2(n6330), .A(n6312), .ZN(U2929) );
  AOI22_X1 U7359 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_6_), .ZN(n6313) );
  OAI21_X1 U7360 ( .B1(n7014), .B2(n6330), .A(n6313), .ZN(U2930) );
  AOI21_X1 U7361 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6328), .A(n6314), .ZN(n6315) );
  OAI21_X1 U7362 ( .B1(n3998), .B2(n6330), .A(n6315), .ZN(U2933) );
  AOI22_X1 U7363 ( .A1(n6328), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6324), .ZN(n6316) );
  NAND2_X1 U7364 ( .A1(n6327), .A2(DATAI_10_), .ZN(n6322) );
  NAND2_X1 U7365 ( .A1(n6316), .A2(n6322), .ZN(U2934) );
  INV_X1 U7366 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6319) );
  AOI21_X1 U7367 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6328), .A(n6317), .ZN(
        n6318) );
  OAI21_X1 U7368 ( .B1(n6319), .B2(n6330), .A(n6318), .ZN(U2936) );
  INV_X1 U7369 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U7370 ( .A1(n6327), .A2(DATAI_14_), .ZN(n6325) );
  INV_X1 U7371 ( .A(n6325), .ZN(n6320) );
  AOI21_X1 U7372 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6328), .A(n6320), .ZN(
        n6321) );
  OAI21_X1 U7373 ( .B1(n6821), .B2(n6330), .A(n6321), .ZN(U2938) );
  AOI22_X1 U7374 ( .A1(n6328), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6324), .ZN(n6323) );
  NAND2_X1 U7375 ( .A1(n6323), .A2(n6322), .ZN(U2949) );
  AOI22_X1 U7376 ( .A1(n6328), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6324), .ZN(n6326) );
  NAND2_X1 U7377 ( .A1(n6326), .A2(n6325), .ZN(U2953) );
  AOI22_X1 U7378 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6328), .B1(n6327), .B2(
        DATAI_15_), .ZN(n6329) );
  OAI21_X1 U7379 ( .B1(n6331), .B2(n6330), .A(n6329), .ZN(U2954) );
  AOI22_X1 U7380 ( .A1(n6377), .A2(REIP_REG_11__SCAN_IN), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6338) );
  INV_X1 U7381 ( .A(n6332), .ZN(n6333) );
  OAI22_X1 U7382 ( .A1(n6335), .A2(n6334), .B1(n6333), .B2(n6370), .ZN(n6336)
         );
  INV_X1 U7383 ( .A(n6336), .ZN(n6337) );
  OAI211_X1 U7384 ( .C1(n6340), .C2(n6339), .A(n6338), .B(n6337), .ZN(U2975)
         );
  INV_X1 U7385 ( .A(n6341), .ZN(n6343) );
  AOI222_X1 U7386 ( .A1(n6344), .A2(n6366), .B1(n6343), .B2(n6350), .C1(n6342), 
        .C2(n6365), .ZN(n6346) );
  OAI211_X1 U7387 ( .C1(n6347), .C2(n6356), .A(n6346), .B(n6345), .ZN(U2979)
         );
  INV_X1 U7388 ( .A(n6348), .ZN(n6353) );
  INV_X1 U7389 ( .A(n6349), .ZN(n6351) );
  AOI222_X1 U7390 ( .A1(n6353), .A2(n6366), .B1(n6352), .B2(n6365), .C1(n6351), 
        .C2(n6350), .ZN(n6355) );
  OAI211_X1 U7391 ( .C1(n6357), .C2(n6356), .A(n6355), .B(n6354), .ZN(U2981)
         );
  AOI22_X1 U7392 ( .A1(n6377), .A2(REIP_REG_2__SCAN_IN), .B1(n6358), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U7393 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  XOR2_X1 U7394 ( .A(n6362), .B(n6361), .Z(n6401) );
  INV_X1 U7395 ( .A(n6363), .ZN(n6364) );
  AOI22_X1 U7396 ( .A1(n6401), .A2(n6366), .B1(n6365), .B2(n6364), .ZN(n6367)
         );
  OAI211_X1 U7397 ( .C1(n6370), .C2(n6369), .A(n6368), .B(n6367), .ZN(U2984)
         );
  AOI21_X1 U7398 ( .B1(n6373), .B2(n6415), .A(n6371), .ZN(n6391) );
  INV_X1 U7399 ( .A(n6372), .ZN(n6381) );
  INV_X1 U7400 ( .A(n6373), .ZN(n6375) );
  NAND2_X1 U7401 ( .A1(n6375), .A2(n6374), .ZN(n6388) );
  AOI221_X1 U7402 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n7064), .C2(n6383), .A(n6388), 
        .ZN(n6376) );
  AOI21_X1 U7403 ( .B1(n6377), .B2(REIP_REG_10__SCAN_IN), .A(n6376), .ZN(n6378) );
  OAI21_X1 U7404 ( .B1(n6379), .B2(n6398), .A(n6378), .ZN(n6380) );
  AOI21_X1 U7405 ( .B1(n6381), .B2(n6412), .A(n6380), .ZN(n6382) );
  OAI21_X1 U7406 ( .B1(n6391), .B2(n6383), .A(n6382), .ZN(U3008) );
  AOI22_X1 U7407 ( .A1(n6384), .A2(n6410), .B1(n6377), .B2(REIP_REG_9__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U7408 ( .A1(n6385), .A2(n6412), .ZN(n6386) );
  OAI211_X1 U7409 ( .C1(n6388), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6387), 
        .B(n6386), .ZN(n6389) );
  INV_X1 U7410 ( .A(n6389), .ZN(n6390) );
  OAI21_X1 U7411 ( .B1(n6391), .B2(n7064), .A(n6390), .ZN(U3009) );
  NAND2_X1 U7412 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6392), .ZN(n6405)
         );
  OAI21_X1 U7413 ( .B1(n6805), .B2(n6404), .A(n6393), .ZN(n6394) );
  AND2_X1 U7414 ( .A1(n6395), .A2(n6394), .ZN(n6400) );
  OAI22_X1 U7415 ( .A1(n6398), .A2(n6397), .B1(n6869), .B2(n6396), .ZN(n6399)
         );
  AOI211_X1 U7416 ( .C1(n6401), .C2(n6412), .A(n6400), .B(n6399), .ZN(n6402)
         );
  OAI221_X1 U7417 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6405), .C1(n6404), .C2(n6403), .A(n6402), .ZN(U3016) );
  OAI21_X1 U7418 ( .B1(n6407), .B2(n4189), .A(n6406), .ZN(n6408) );
  AOI21_X1 U7419 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6414) );
  NAND2_X1 U7420 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  AND2_X1 U7421 ( .A1(n6414), .A2(n6413), .ZN(n6418) );
  OAI211_X1 U7422 ( .C1(n6416), .C2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4189), 
        .B(n6415), .ZN(n6417) );
  NAND2_X1 U7423 ( .A1(n6418), .A2(n6417), .ZN(U3017) );
  NOR2_X1 U7424 ( .A1(n6420), .A2(n6419), .ZN(U3019) );
  AND2_X1 U7425 ( .A1(n6431), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6423)
         );
  AOI21_X1 U7426 ( .B1(n6421), .B2(n6583), .A(n6423), .ZN(n6428) );
  NOR2_X1 U7427 ( .A1(n6428), .A2(n6651), .ZN(n6422) );
  AOI21_X1 U7428 ( .B1(n6431), .B2(STATE2_REG_2__SCAN_IN), .A(n6422), .ZN(
        n6460) );
  INV_X1 U7429 ( .A(n6423), .ZN(n6453) );
  OAI22_X1 U7430 ( .A1(n6454), .A2(n6665), .B1(n6544), .B2(n6453), .ZN(n6424)
         );
  INV_X1 U7431 ( .A(n6424), .ZN(n6434) );
  NAND3_X1 U7432 ( .A1(n6427), .A2(n6426), .A3(n6425), .ZN(n6429) );
  NAND3_X1 U7433 ( .A1(n6429), .A2(n6586), .A3(n6428), .ZN(n6430) );
  OAI211_X1 U7434 ( .C1(n6586), .C2(n6431), .A(n6430), .B(n6585), .ZN(n6457)
         );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6457), .B1(n6662), 
        .B2(n6456), .ZN(n6433) );
  OAI211_X1 U7436 ( .C1(n6460), .C2(n6553), .A(n6434), .B(n6433), .ZN(U3044)
         );
  OAI22_X1 U7437 ( .A1(n6454), .A2(n6671), .B1(n6507), .B2(n6453), .ZN(n6435)
         );
  INV_X1 U7438 ( .A(n6435), .ZN(n6437) );
  AOI22_X1 U7439 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6457), .B1(n6668), 
        .B2(n6456), .ZN(n6436) );
  OAI211_X1 U7440 ( .C1(n6460), .C2(n6556), .A(n6437), .B(n6436), .ZN(U3045)
         );
  OAI22_X1 U7441 ( .A1(n6454), .A2(n6677), .B1(n7112), .B2(n6453), .ZN(n6438)
         );
  INV_X1 U7442 ( .A(n6438), .ZN(n6440) );
  AOI22_X1 U7443 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6457), .B1(n6674), 
        .B2(n6456), .ZN(n6439) );
  OAI211_X1 U7444 ( .C1(n6460), .C2(n7113), .A(n6440), .B(n6439), .ZN(U3046)
         );
  OAI22_X1 U7445 ( .A1(n6454), .A2(n6683), .B1(n6606), .B2(n6453), .ZN(n6441)
         );
  INV_X1 U7446 ( .A(n6441), .ZN(n6443) );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6457), .B1(n6680), 
        .B2(n6456), .ZN(n6442) );
  OAI211_X1 U7448 ( .C1(n6460), .C2(n6562), .A(n6443), .B(n6442), .ZN(U3047)
         );
  OAI22_X1 U7449 ( .A1(n6454), .A2(n6689), .B1(n6613), .B2(n6453), .ZN(n6444)
         );
  INV_X1 U7450 ( .A(n6444), .ZN(n6446) );
  AOI22_X1 U7451 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6457), .B1(n6686), 
        .B2(n6456), .ZN(n6445) );
  OAI211_X1 U7452 ( .C1(n6460), .C2(n6565), .A(n6446), .B(n6445), .ZN(U3048)
         );
  OAI22_X1 U7453 ( .A1(n6454), .A2(n6695), .B1(n6523), .B2(n6453), .ZN(n6447)
         );
  INV_X1 U7454 ( .A(n6447), .ZN(n6449) );
  AOI22_X1 U7455 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6457), .B1(n6692), 
        .B2(n6456), .ZN(n6448) );
  OAI211_X1 U7456 ( .C1(n6460), .C2(n6568), .A(n6449), .B(n6448), .ZN(U3049)
         );
  OAI22_X1 U7457 ( .A1(n6454), .A2(n6701), .B1(n6625), .B2(n6453), .ZN(n6450)
         );
  INV_X1 U7458 ( .A(n6450), .ZN(n6452) );
  AOI22_X1 U7459 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6457), .B1(n6698), 
        .B2(n6456), .ZN(n6451) );
  OAI211_X1 U7460 ( .C1(n6460), .C2(n6574), .A(n6452), .B(n6451), .ZN(U3050)
         );
  OAI22_X1 U7461 ( .A1(n6454), .A2(n6712), .B1(n6633), .B2(n6453), .ZN(n6455)
         );
  INV_X1 U7462 ( .A(n6455), .ZN(n6459) );
  AOI22_X1 U7463 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6457), .B1(n6707), 
        .B2(n6456), .ZN(n6458) );
  OAI211_X1 U7464 ( .C1(n6460), .C2(n6580), .A(n6459), .B(n6458), .ZN(U3051)
         );
  AND3_X1 U7465 ( .A1(n6462), .A2(n6461), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6501) );
  NAND2_X1 U7466 ( .A1(n6501), .A2(n7028), .ZN(n6470) );
  INV_X1 U7467 ( .A(n6470), .ZN(n6490) );
  INV_X1 U7468 ( .A(n6463), .ZN(n6645) );
  INV_X1 U7469 ( .A(n6464), .ZN(n6465) );
  OAI22_X1 U7470 ( .A1(n6466), .A2(n6653), .B1(n6645), .B2(n6465), .ZN(n6489)
         );
  AOI22_X1 U7471 ( .A1(n6648), .A2(n6490), .B1(n6489), .B2(n6649), .ZN(n6476)
         );
  INV_X1 U7472 ( .A(n6474), .ZN(n6468) );
  OAI22_X1 U7473 ( .A1(n6494), .A2(n6655), .B1(n6495), .B2(n6653), .ZN(n6472)
         );
  AOI211_X1 U7474 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6470), .A(n6658), .B(
        n6469), .ZN(n6471) );
  AOI22_X1 U7475 ( .A1(n6491), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6662), 
        .B2(n6534), .ZN(n6475) );
  OAI211_X1 U7476 ( .C1(n6665), .C2(n6494), .A(n6476), .B(n6475), .ZN(U3052)
         );
  AOI22_X1 U7477 ( .A1(n6666), .A2(n6490), .B1(n6489), .B2(n6667), .ZN(n6478)
         );
  AOI22_X1 U7478 ( .A1(n6491), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6668), 
        .B2(n6534), .ZN(n6477) );
  OAI211_X1 U7479 ( .C1(n6671), .C2(n6494), .A(n6478), .B(n6477), .ZN(U3053)
         );
  AOI22_X1 U7480 ( .A1(n6672), .A2(n6490), .B1(n6489), .B2(n6673), .ZN(n6480)
         );
  AOI22_X1 U7481 ( .A1(n6491), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6674), 
        .B2(n6534), .ZN(n6479) );
  OAI211_X1 U7482 ( .C1(n6677), .C2(n6494), .A(n6480), .B(n6479), .ZN(U3054)
         );
  AOI22_X1 U7483 ( .A1(n6678), .A2(n6490), .B1(n6489), .B2(n6679), .ZN(n6482)
         );
  AOI22_X1 U7484 ( .A1(n6491), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6680), 
        .B2(n6534), .ZN(n6481) );
  OAI211_X1 U7485 ( .C1(n6683), .C2(n6494), .A(n6482), .B(n6481), .ZN(U3055)
         );
  AOI22_X1 U7486 ( .A1(n6684), .A2(n6490), .B1(n6489), .B2(n6685), .ZN(n6484)
         );
  AOI22_X1 U7487 ( .A1(n6491), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6686), 
        .B2(n6534), .ZN(n6483) );
  OAI211_X1 U7488 ( .C1(n6689), .C2(n6494), .A(n6484), .B(n6483), .ZN(U3056)
         );
  AOI22_X1 U7489 ( .A1(n6690), .A2(n6490), .B1(n6489), .B2(n6691), .ZN(n6486)
         );
  AOI22_X1 U7490 ( .A1(n6491), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6692), 
        .B2(n6534), .ZN(n6485) );
  OAI211_X1 U7491 ( .C1(n6695), .C2(n6494), .A(n6486), .B(n6485), .ZN(U3057)
         );
  AOI22_X1 U7492 ( .A1(n6696), .A2(n6490), .B1(n6489), .B2(n6697), .ZN(n6488)
         );
  AOI22_X1 U7493 ( .A1(n6491), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6698), 
        .B2(n6534), .ZN(n6487) );
  OAI211_X1 U7494 ( .C1(n6701), .C2(n6494), .A(n6488), .B(n6487), .ZN(U3058)
         );
  AOI22_X1 U7495 ( .A1(n6703), .A2(n6490), .B1(n6489), .B2(n6704), .ZN(n6493)
         );
  AOI22_X1 U7496 ( .A1(n6491), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6707), 
        .B2(n6534), .ZN(n6492) );
  OAI211_X1 U7497 ( .C1(n6712), .C2(n6494), .A(n6493), .B(n6492), .ZN(U3059)
         );
  INV_X1 U7498 ( .A(n6504), .ZN(n6499) );
  OR2_X1 U7499 ( .A1(n6496), .A2(n6495), .ZN(n6540) );
  OR2_X1 U7500 ( .A1(n6653), .A2(n6540), .ZN(n6497) );
  NAND2_X1 U7501 ( .A1(n6501), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6531) );
  AND2_X1 U7502 ( .A1(n6497), .A2(n6531), .ZN(n6503) );
  OAI21_X1 U7503 ( .B1(n6586), .B2(n6501), .A(n6585), .ZN(n6498) );
  NOR2_X1 U7504 ( .A1(n6544), .A2(n6531), .ZN(n6500) );
  AOI21_X1 U7505 ( .B1(n6533), .B2(n6662), .A(n6500), .ZN(n6506) );
  INV_X1 U7506 ( .A(n6501), .ZN(n6502) );
  OAI22_X1 U7507 ( .A1(n6504), .A2(n6503), .B1(n6592), .B2(n6502), .ZN(n6535)
         );
  AOI22_X1 U7508 ( .A1(n6535), .A2(n6649), .B1(n6589), .B2(n6534), .ZN(n6505)
         );
  OAI211_X1 U7509 ( .C1(n6539), .C2(n6968), .A(n6506), .B(n6505), .ZN(U3060)
         );
  INV_X1 U7510 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6511) );
  NOR2_X1 U7511 ( .A1(n6507), .A2(n6531), .ZN(n6508) );
  AOI21_X1 U7512 ( .B1(n6533), .B2(n6668), .A(n6508), .ZN(n6510) );
  AOI22_X1 U7513 ( .A1(n6535), .A2(n6667), .B1(n6599), .B2(n6534), .ZN(n6509)
         );
  OAI211_X1 U7514 ( .C1(n6539), .C2(n6511), .A(n6510), .B(n6509), .ZN(U3061)
         );
  INV_X1 U7515 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6515) );
  NOR2_X1 U7516 ( .A1(n7112), .A2(n6531), .ZN(n6512) );
  AOI21_X1 U7517 ( .B1(n6533), .B2(n6674), .A(n6512), .ZN(n6514) );
  AOI22_X1 U7518 ( .A1(n6535), .A2(n6673), .B1(n7117), .B2(n6534), .ZN(n6513)
         );
  OAI211_X1 U7519 ( .C1(n6539), .C2(n6515), .A(n6514), .B(n6513), .ZN(U3062)
         );
  INV_X1 U7520 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n7089) );
  NOR2_X1 U7521 ( .A1(n6606), .A2(n6531), .ZN(n6516) );
  AOI21_X1 U7522 ( .B1(n6533), .B2(n6680), .A(n6516), .ZN(n6518) );
  AOI22_X1 U7523 ( .A1(n6535), .A2(n6679), .B1(n6609), .B2(n6534), .ZN(n6517)
         );
  OAI211_X1 U7524 ( .C1(n6539), .C2(n7089), .A(n6518), .B(n6517), .ZN(U3063)
         );
  INV_X1 U7525 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6522) );
  NOR2_X1 U7526 ( .A1(n6613), .A2(n6531), .ZN(n6519) );
  AOI21_X1 U7527 ( .B1(n6533), .B2(n6686), .A(n6519), .ZN(n6521) );
  AOI22_X1 U7528 ( .A1(n6535), .A2(n6685), .B1(n6616), .B2(n6534), .ZN(n6520)
         );
  OAI211_X1 U7529 ( .C1(n6539), .C2(n6522), .A(n6521), .B(n6520), .ZN(U3064)
         );
  NOR2_X1 U7530 ( .A1(n6523), .A2(n6531), .ZN(n6524) );
  AOI21_X1 U7531 ( .B1(n6533), .B2(n6692), .A(n6524), .ZN(n6526) );
  AOI22_X1 U7532 ( .A1(n6535), .A2(n6691), .B1(n6621), .B2(n6534), .ZN(n6525)
         );
  OAI211_X1 U7533 ( .C1(n6539), .C2(n3912), .A(n6526), .B(n6525), .ZN(U3065)
         );
  INV_X1 U7534 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6530) );
  NOR2_X1 U7535 ( .A1(n6625), .A2(n6531), .ZN(n6527) );
  AOI21_X1 U7536 ( .B1(n6533), .B2(n6698), .A(n6527), .ZN(n6529) );
  AOI22_X1 U7537 ( .A1(n6535), .A2(n6697), .B1(n6628), .B2(n6534), .ZN(n6528)
         );
  OAI211_X1 U7538 ( .C1(n6539), .C2(n6530), .A(n6529), .B(n6528), .ZN(U3066)
         );
  INV_X1 U7539 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6538) );
  NOR2_X1 U7540 ( .A1(n6633), .A2(n6531), .ZN(n6532) );
  AOI21_X1 U7541 ( .B1(n6533), .B2(n6707), .A(n6532), .ZN(n6537) );
  AOI22_X1 U7542 ( .A1(n6535), .A2(n6704), .B1(n6636), .B2(n6534), .ZN(n6536)
         );
  OAI211_X1 U7543 ( .C1(n6539), .C2(n6538), .A(n6537), .B(n6536), .ZN(U3067)
         );
  INV_X1 U7544 ( .A(n6540), .ZN(n6541) );
  INV_X1 U7545 ( .A(n6569), .ZN(n6575) );
  AOI21_X1 U7546 ( .B1(n6542), .B2(n6541), .A(n6575), .ZN(n6547) );
  NOR2_X1 U7547 ( .A1(n6547), .A2(n6651), .ZN(n6543) );
  AOI21_X1 U7548 ( .B1(n6550), .B2(STATE2_REG_2__SCAN_IN), .A(n6543), .ZN(
        n6581) );
  OAI22_X1 U7549 ( .A1(n6570), .A2(n6545), .B1(n6569), .B2(n6544), .ZN(n6546)
         );
  INV_X1 U7550 ( .A(n6546), .ZN(n6552) );
  NAND3_X1 U7551 ( .A1(n6548), .A2(n6586), .A3(n6547), .ZN(n6549) );
  OAI211_X1 U7552 ( .C1(n6550), .C2(n6586), .A(n6549), .B(n6585), .ZN(n6577)
         );
  AOI22_X1 U7553 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6577), .B1(n6589), 
        .B2(n6576), .ZN(n6551) );
  OAI211_X1 U7554 ( .C1(n6581), .C2(n6553), .A(n6552), .B(n6551), .ZN(U3076)
         );
  AOI22_X1 U7555 ( .A1(n6576), .A2(n6599), .B1(n6575), .B2(n6666), .ZN(n6555)
         );
  AOI22_X1 U7556 ( .A1(n6577), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6668), 
        .B2(n7116), .ZN(n6554) );
  OAI211_X1 U7557 ( .C1(n6581), .C2(n6556), .A(n6555), .B(n6554), .ZN(U3077)
         );
  AOI22_X1 U7558 ( .A1(n6576), .A2(n7117), .B1(n6575), .B2(n6672), .ZN(n6558)
         );
  AOI22_X1 U7559 ( .A1(n6577), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6674), 
        .B2(n7116), .ZN(n6557) );
  OAI211_X1 U7560 ( .C1(n6581), .C2(n7113), .A(n6558), .B(n6557), .ZN(U3078)
         );
  OAI22_X1 U7561 ( .A1(n6570), .A2(n6607), .B1(n6569), .B2(n6606), .ZN(n6559)
         );
  INV_X1 U7562 ( .A(n6559), .ZN(n6561) );
  AOI22_X1 U7563 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6577), .B1(n6609), 
        .B2(n6576), .ZN(n6560) );
  OAI211_X1 U7564 ( .C1(n6581), .C2(n6562), .A(n6561), .B(n6560), .ZN(U3079)
         );
  AOI22_X1 U7565 ( .A1(n6576), .A2(n6616), .B1(n6575), .B2(n6684), .ZN(n6564)
         );
  AOI22_X1 U7566 ( .A1(n6577), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6686), 
        .B2(n7116), .ZN(n6563) );
  OAI211_X1 U7567 ( .C1(n6581), .C2(n6565), .A(n6564), .B(n6563), .ZN(U3080)
         );
  AOI22_X1 U7568 ( .A1(n6576), .A2(n6621), .B1(n6575), .B2(n6690), .ZN(n6567)
         );
  AOI22_X1 U7569 ( .A1(n6577), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6692), 
        .B2(n7116), .ZN(n6566) );
  OAI211_X1 U7570 ( .C1(n6581), .C2(n6568), .A(n6567), .B(n6566), .ZN(U3081)
         );
  OAI22_X1 U7571 ( .A1(n6570), .A2(n6626), .B1(n6569), .B2(n6625), .ZN(n6571)
         );
  INV_X1 U7572 ( .A(n6571), .ZN(n6573) );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6577), .B1(n6628), 
        .B2(n6576), .ZN(n6572) );
  OAI211_X1 U7574 ( .C1(n6581), .C2(n6574), .A(n6573), .B(n6572), .ZN(U3082)
         );
  AOI22_X1 U7575 ( .A1(n6576), .A2(n6636), .B1(n6575), .B2(n6703), .ZN(n6579)
         );
  AOI22_X1 U7576 ( .A1(n6577), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6707), 
        .B2(n7116), .ZN(n6578) );
  OAI211_X1 U7577 ( .C1(n6581), .C2(n6580), .A(n6579), .B(n6578), .ZN(U3083)
         );
  OAI21_X1 U7578 ( .B1(n6596), .B2(n6582), .A(n6586), .ZN(n6594) );
  INV_X1 U7579 ( .A(n6594), .ZN(n6588) );
  AND2_X1 U7580 ( .A1(n6590), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6620)
         );
  AOI21_X1 U7581 ( .B1(n6584), .B2(n6583), .A(n6620), .ZN(n6593) );
  OAI21_X1 U7582 ( .B1(n6586), .B2(n6590), .A(n6585), .ZN(n6587) );
  INV_X1 U7583 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U7584 ( .A1(n6637), .A2(n6589), .B1(n6648), .B2(n6620), .ZN(n6598)
         );
  INV_X1 U7585 ( .A(n6590), .ZN(n6591) );
  OAI22_X1 U7586 ( .A1(n6594), .A2(n6593), .B1(n6592), .B2(n6591), .ZN(n6638)
         );
  AOI22_X1 U7587 ( .A1(n6638), .A2(n6649), .B1(n6662), .B2(n6652), .ZN(n6597)
         );
  OAI211_X1 U7588 ( .C1(n6641), .C2(n6991), .A(n6598), .B(n6597), .ZN(U3108)
         );
  INV_X1 U7589 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7590 ( .A1(n6637), .A2(n6599), .B1(n6666), .B2(n6620), .ZN(n6601)
         );
  AOI22_X1 U7591 ( .A1(n6638), .A2(n6667), .B1(n6668), .B2(n6652), .ZN(n6600)
         );
  OAI211_X1 U7592 ( .C1(n6641), .C2(n6602), .A(n6601), .B(n6600), .ZN(U3109)
         );
  INV_X1 U7593 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7594 ( .A1(n6637), .A2(n7117), .B1(n6672), .B2(n6620), .ZN(n6604)
         );
  AOI22_X1 U7595 ( .A1(n6638), .A2(n6673), .B1(n6674), .B2(n6652), .ZN(n6603)
         );
  OAI211_X1 U7596 ( .C1(n6641), .C2(n6605), .A(n6604), .B(n6603), .ZN(U3110)
         );
  INV_X1 U7597 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6612) );
  INV_X1 U7598 ( .A(n6620), .ZN(n6632) );
  OAI22_X1 U7599 ( .A1(n6711), .A2(n6607), .B1(n6606), .B2(n6632), .ZN(n6608)
         );
  INV_X1 U7600 ( .A(n6608), .ZN(n6611) );
  AOI22_X1 U7601 ( .A1(n6638), .A2(n6679), .B1(n6637), .B2(n6609), .ZN(n6610)
         );
  OAI211_X1 U7602 ( .C1(n6641), .C2(n6612), .A(n6611), .B(n6610), .ZN(U3111)
         );
  INV_X1 U7603 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6619) );
  OAI22_X1 U7604 ( .A1(n6711), .A2(n6614), .B1(n6613), .B2(n6632), .ZN(n6615)
         );
  INV_X1 U7605 ( .A(n6615), .ZN(n6618) );
  AOI22_X1 U7606 ( .A1(n6638), .A2(n6685), .B1(n6637), .B2(n6616), .ZN(n6617)
         );
  OAI211_X1 U7607 ( .C1(n6641), .C2(n6619), .A(n6618), .B(n6617), .ZN(U3112)
         );
  INV_X1 U7608 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6624) );
  AOI22_X1 U7609 ( .A1(n6637), .A2(n6621), .B1(n6690), .B2(n6620), .ZN(n6623)
         );
  AOI22_X1 U7610 ( .A1(n6638), .A2(n6691), .B1(n6692), .B2(n6652), .ZN(n6622)
         );
  OAI211_X1 U7611 ( .C1(n6641), .C2(n6624), .A(n6623), .B(n6622), .ZN(U3113)
         );
  INV_X1 U7612 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6631) );
  OAI22_X1 U7613 ( .A1(n6711), .A2(n6626), .B1(n6625), .B2(n6632), .ZN(n6627)
         );
  INV_X1 U7614 ( .A(n6627), .ZN(n6630) );
  AOI22_X1 U7615 ( .A1(n6638), .A2(n6697), .B1(n6637), .B2(n6628), .ZN(n6629)
         );
  OAI211_X1 U7616 ( .C1(n6641), .C2(n6631), .A(n6630), .B(n6629), .ZN(U3114)
         );
  INV_X1 U7617 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n7049) );
  OAI22_X1 U7618 ( .A1(n6711), .A2(n6634), .B1(n6633), .B2(n6632), .ZN(n6635)
         );
  INV_X1 U7619 ( .A(n6635), .ZN(n6640) );
  AOI22_X1 U7620 ( .A1(n6638), .A2(n6704), .B1(n6637), .B2(n6636), .ZN(n6639)
         );
  OAI211_X1 U7621 ( .C1(n6641), .C2(n7049), .A(n6640), .B(n6639), .ZN(U3115)
         );
  INV_X1 U7622 ( .A(n6642), .ZN(n6646) );
  INV_X1 U7623 ( .A(n6643), .ZN(n6644) );
  OAI22_X1 U7624 ( .A1(n6646), .A2(n6653), .B1(n6645), .B2(n6644), .ZN(n6705)
         );
  NAND2_X1 U7625 ( .A1(n6647), .A2(n7028), .ZN(n6659) );
  INV_X1 U7626 ( .A(n6659), .ZN(n6702) );
  AOI22_X1 U7627 ( .A1(n6705), .A2(n6649), .B1(n6648), .B2(n6702), .ZN(n6664)
         );
  NOR3_X1 U7628 ( .A1(n6652), .A2(n6706), .A3(n6651), .ZN(n6656) );
  OAI22_X1 U7629 ( .A1(n6656), .A2(n6655), .B1(n6654), .B2(n6653), .ZN(n6661)
         );
  AOI211_X1 U7630 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6659), .A(n6658), .B(
        n6657), .ZN(n6660) );
  NAND2_X1 U7631 ( .A1(n6661), .A2(n6660), .ZN(n6708) );
  AOI22_X1 U7632 ( .A1(n6708), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6662), 
        .B2(n6706), .ZN(n6663) );
  OAI211_X1 U7633 ( .C1(n6665), .C2(n6711), .A(n6664), .B(n6663), .ZN(U3116)
         );
  AOI22_X1 U7634 ( .A1(n6705), .A2(n6667), .B1(n6666), .B2(n6702), .ZN(n6670)
         );
  AOI22_X1 U7635 ( .A1(n6708), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6668), 
        .B2(n6706), .ZN(n6669) );
  OAI211_X1 U7636 ( .C1(n6671), .C2(n6711), .A(n6670), .B(n6669), .ZN(U3117)
         );
  AOI22_X1 U7637 ( .A1(n6705), .A2(n6673), .B1(n6672), .B2(n6702), .ZN(n6676)
         );
  AOI22_X1 U7638 ( .A1(n6708), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6674), 
        .B2(n6706), .ZN(n6675) );
  OAI211_X1 U7639 ( .C1(n6677), .C2(n6711), .A(n6676), .B(n6675), .ZN(U3118)
         );
  AOI22_X1 U7640 ( .A1(n6705), .A2(n6679), .B1(n6678), .B2(n6702), .ZN(n6682)
         );
  AOI22_X1 U7641 ( .A1(n6708), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6680), 
        .B2(n6706), .ZN(n6681) );
  OAI211_X1 U7642 ( .C1(n6683), .C2(n6711), .A(n6682), .B(n6681), .ZN(U3119)
         );
  AOI22_X1 U7643 ( .A1(n6705), .A2(n6685), .B1(n6684), .B2(n6702), .ZN(n6688)
         );
  AOI22_X1 U7644 ( .A1(n6708), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6686), 
        .B2(n6706), .ZN(n6687) );
  OAI211_X1 U7645 ( .C1(n6689), .C2(n6711), .A(n6688), .B(n6687), .ZN(U3120)
         );
  AOI22_X1 U7646 ( .A1(n6705), .A2(n6691), .B1(n6690), .B2(n6702), .ZN(n6694)
         );
  AOI22_X1 U7647 ( .A1(n6708), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6692), 
        .B2(n6706), .ZN(n6693) );
  OAI211_X1 U7648 ( .C1(n6695), .C2(n6711), .A(n6694), .B(n6693), .ZN(U3121)
         );
  AOI22_X1 U7649 ( .A1(n6705), .A2(n6697), .B1(n6696), .B2(n6702), .ZN(n6700)
         );
  AOI22_X1 U7650 ( .A1(n6708), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6698), 
        .B2(n6706), .ZN(n6699) );
  OAI211_X1 U7651 ( .C1(n6701), .C2(n6711), .A(n6700), .B(n6699), .ZN(U3122)
         );
  AOI22_X1 U7652 ( .A1(n6705), .A2(n6704), .B1(n6703), .B2(n6702), .ZN(n6710)
         );
  AOI22_X1 U7653 ( .A1(n6708), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6707), 
        .B2(n6706), .ZN(n6709) );
  OAI211_X1 U7654 ( .C1(n6712), .C2(n6711), .A(n6710), .B(n6709), .ZN(U3123)
         );
  OAI211_X1 U7655 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6715), .A(n6714), .B(
        n6713), .ZN(n6716) );
  NAND2_X1 U7656 ( .A1(n6717), .A2(n6716), .ZN(U3150) );
  AND2_X1 U7657 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6718), .ZN(U3151) );
  INV_X1 U7658 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U7659 ( .A1(n6778), .A2(n7012), .ZN(U3152) );
  AND2_X1 U7660 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6718), .ZN(U3153) );
  INV_X1 U7661 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6990) );
  NOR2_X1 U7662 ( .A1(n6778), .A2(n6990), .ZN(U3154) );
  INV_X1 U7663 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6957) );
  NOR2_X1 U7664 ( .A1(n6778), .A2(n6957), .ZN(U3155) );
  AND2_X1 U7665 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6718), .ZN(U3156) );
  NOR2_X1 U7666 ( .A1(n6778), .A2(n7045), .ZN(U3157) );
  NOR2_X1 U7667 ( .A1(n6778), .A2(n6897), .ZN(U3158) );
  NOR2_X1 U7668 ( .A1(n6778), .A2(n6878), .ZN(U3159) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6718), .ZN(U3160) );
  AND2_X1 U7670 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6718), .ZN(U3161) );
  AND2_X1 U7671 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6718), .ZN(U3162) );
  AND2_X1 U7672 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6718), .ZN(U3163) );
  AND2_X1 U7673 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6718), .ZN(U3164) );
  INV_X1 U7674 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U7675 ( .A1(n6778), .A2(n6963), .ZN(U3165) );
  AND2_X1 U7676 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6718), .ZN(U3166) );
  AND2_X1 U7677 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6718), .ZN(U3167) );
  AND2_X1 U7678 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6718), .ZN(U3168) );
  INV_X1 U7679 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6904) );
  NOR2_X1 U7680 ( .A1(n6778), .A2(n6904), .ZN(U3169) );
  AND2_X1 U7681 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6718), .ZN(U3170) );
  NOR2_X1 U7682 ( .A1(n6778), .A2(n7033), .ZN(U3171) );
  AND2_X1 U7683 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6718), .ZN(U3172) );
  AND2_X1 U7684 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6718), .ZN(U3173) );
  INV_X1 U7685 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7003) );
  NOR2_X1 U7686 ( .A1(n6778), .A2(n7003), .ZN(U3174) );
  AND2_X1 U7687 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6718), .ZN(U3175) );
  AND2_X1 U7688 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6718), .ZN(U3176) );
  INV_X1 U7689 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U7690 ( .A1(n6778), .A2(n6911), .ZN(U3177) );
  AND2_X1 U7691 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6718), .ZN(U3178) );
  AND2_X1 U7692 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6718), .ZN(U3179) );
  AND2_X1 U7693 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6718), .ZN(U3180) );
  AOI22_X1 U7694 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .B1(
        n6719), .B2(n6965), .ZN(n6723) );
  AOI221_X1 U7695 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4601), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6720) );
  AOI221_X1 U7696 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6720), .C2(HOLD), .A(n6943), .ZN(n6722) );
  OAI22_X1 U7697 ( .A1(n6724), .A2(n6723), .B1(n6722), .B2(n6721), .ZN(U3183)
         );
  NAND2_X1 U7698 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6789), .ZN(n6767) );
  INV_X1 U7699 ( .A(n6767), .ZN(n6771) );
  AOI22_X1 U7700 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6800), .ZN(n6725) );
  OAI21_X1 U7701 ( .B1(n6869), .B2(n6773), .A(n6725), .ZN(U3184) );
  AOI22_X1 U7702 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6800), .ZN(n6726) );
  OAI21_X1 U7703 ( .B1(n6728), .B2(n6773), .A(n6726), .ZN(U3185) );
  INV_X1 U7704 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6894) );
  OAI222_X1 U7705 ( .A1(n6767), .A2(n6728), .B1(n6894), .B2(n6789), .C1(n6727), 
        .C2(n6773), .ZN(U3186) );
  AOI22_X1 U7706 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6800), .ZN(n6729) );
  OAI21_X1 U7707 ( .B1(n6730), .B2(n6773), .A(n6729), .ZN(U3187) );
  AOI22_X1 U7708 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6800), .ZN(n6731) );
  OAI21_X1 U7709 ( .B1(n6732), .B2(n6773), .A(n6731), .ZN(U3188) );
  AOI22_X1 U7710 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6800), .ZN(n6733) );
  OAI21_X1 U7711 ( .B1(n6969), .B2(n6773), .A(n6733), .ZN(U3189) );
  AOI22_X1 U7712 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6800), .ZN(n6734) );
  OAI21_X1 U7713 ( .B1(n6735), .B2(n6773), .A(n6734), .ZN(U3190) );
  AOI22_X1 U7714 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6800), .ZN(n6736) );
  OAI21_X1 U7715 ( .B1(n6737), .B2(n6773), .A(n6736), .ZN(U3191) );
  AOI22_X1 U7716 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6800), .ZN(n6738) );
  OAI21_X1 U7717 ( .B1(n6739), .B2(n6773), .A(n6738), .ZN(U3192) );
  AOI22_X1 U7718 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6800), .ZN(n6740) );
  OAI21_X1 U7719 ( .B1(n6741), .B2(n6773), .A(n6740), .ZN(U3193) );
  AOI22_X1 U7720 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6800), .ZN(n6742) );
  OAI21_X1 U7721 ( .B1(n6743), .B2(n6773), .A(n6742), .ZN(U3194) );
  AOI22_X1 U7722 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6800), .ZN(n6744) );
  OAI21_X1 U7723 ( .B1(n6746), .B2(n6773), .A(n6744), .ZN(U3195) );
  AOI22_X1 U7724 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6800), .ZN(n6745) );
  OAI21_X1 U7725 ( .B1(n6746), .B2(n6767), .A(n6745), .ZN(U3196) );
  AOI22_X1 U7726 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6800), .ZN(n6747) );
  OAI21_X1 U7727 ( .B1(n6985), .B2(n6773), .A(n6747), .ZN(U3197) );
  AOI22_X1 U7728 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6800), .ZN(n6748) );
  OAI21_X1 U7729 ( .B1(n6985), .B2(n6767), .A(n6748), .ZN(U3198) );
  AOI22_X1 U7730 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6800), .ZN(n6749) );
  OAI21_X1 U7731 ( .B1(n6750), .B2(n6767), .A(n6749), .ZN(U3199) );
  AOI22_X1 U7732 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6800), .ZN(n6751) );
  OAI21_X1 U7733 ( .B1(n6753), .B2(n6773), .A(n6751), .ZN(U3200) );
  INV_X1 U7734 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7065) );
  OAI222_X1 U7735 ( .A1(n6767), .A2(n6753), .B1(n7065), .B2(n6789), .C1(n6752), 
        .C2(n6773), .ZN(U3201) );
  AOI22_X1 U7736 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6800), .ZN(n6754) );
  OAI21_X1 U7737 ( .B1(n6987), .B2(n6773), .A(n6754), .ZN(U3202) );
  AOI22_X1 U7738 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6800), .ZN(n6755) );
  OAI21_X1 U7739 ( .B1(n6756), .B2(n6773), .A(n6755), .ZN(U3203) );
  INV_X1 U7740 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6997) );
  OAI222_X1 U7741 ( .A1(n6767), .A2(n6756), .B1(n6997), .B2(n6789), .C1(n6758), 
        .C2(n6773), .ZN(U3204) );
  AOI22_X1 U7742 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6800), .ZN(n6757) );
  OAI21_X1 U7743 ( .B1(n6758), .B2(n6767), .A(n6757), .ZN(U3205) );
  AOI22_X1 U7744 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6800), .ZN(n6759) );
  OAI21_X1 U7745 ( .B1(n6761), .B2(n6773), .A(n6759), .ZN(U3206) );
  AOI22_X1 U7746 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6800), .ZN(n6760) );
  OAI21_X1 U7747 ( .B1(n6761), .B2(n6767), .A(n6760), .ZN(U3207) );
  AOI22_X1 U7748 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6800), .ZN(n6762) );
  OAI21_X1 U7749 ( .B1(n7062), .B2(n6773), .A(n6762), .ZN(U3208) );
  AOI22_X1 U7750 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6800), .ZN(n6763) );
  OAI21_X1 U7751 ( .B1(n6764), .B2(n6773), .A(n6763), .ZN(U3209) );
  INV_X1 U7752 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6982) );
  OAI222_X1 U7753 ( .A1(n6767), .A2(n6764), .B1(n6982), .B2(n6789), .C1(n6768), 
        .C2(n6773), .ZN(U3210) );
  AOI22_X1 U7754 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6765), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6800), .ZN(n6766) );
  OAI21_X1 U7755 ( .B1(n6768), .B2(n6767), .A(n6766), .ZN(U3211) );
  AOI22_X1 U7756 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6800), .ZN(n6769) );
  OAI21_X1 U7757 ( .B1(n6770), .B2(n6773), .A(n6769), .ZN(U3212) );
  INV_X1 U7758 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7759 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6771), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6800), .ZN(n6772) );
  OAI21_X1 U7760 ( .B1(n6774), .B2(n6773), .A(n6772), .ZN(U3213) );
  MUX2_X1 U7761 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6800), .Z(U3445) );
  MUX2_X1 U7762 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6800), .Z(U3446) );
  MUX2_X1 U7763 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6800), .Z(U3447) );
  MUX2_X1 U7764 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6800), .Z(U3448) );
  OAI21_X1 U7765 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6778), .A(n6776), .ZN(
        n6775) );
  INV_X1 U7766 ( .A(n6775), .ZN(U3451) );
  OAI21_X1 U7767 ( .B1(n6778), .B2(n6777), .A(n6776), .ZN(U3452) );
  AOI221_X1 U7768 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7027), .C1(
        STATE2_REG_3__SCAN_IN), .C2(n6780), .A(n6779), .ZN(n6781) );
  INV_X1 U7769 ( .A(n6781), .ZN(U3453) );
  AOI21_X1 U7770 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6783) );
  AOI22_X1 U7771 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6783), .B2(n6782), .ZN(n6784) );
  INV_X1 U7772 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7773 ( .A1(n6785), .A2(n6784), .B1(n6955), .B2(n6787), .ZN(U3468)
         );
  INV_X1 U7774 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U7775 ( .A1(n6787), .A2(REIP_REG_1__SCAN_IN), .ZN(n6786) );
  AOI22_X1 U7776 ( .A1(n6788), .A2(n6787), .B1(n7077), .B2(n6786), .ZN(U3469)
         );
  INV_X1 U7777 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7035) );
  AOI22_X1 U7778 ( .A1(n6789), .A2(READREQUEST_REG_SCAN_IN), .B1(n7035), .B2(
        n6800), .ZN(U3470) );
  AND2_X1 U7779 ( .A1(n6300), .A2(n4601), .ZN(n6791) );
  NOR3_X1 U7780 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6799) );
  OAI211_X1 U7781 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6794), .A(n6793), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6796) );
  AOI21_X1 U7782 ( .B1(n6796), .B2(STATE2_REG_0__SCAN_IN), .A(n6795), .ZN(
        n6798) );
  NAND2_X1 U7783 ( .A1(n6799), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6797) );
  OAI21_X1 U7784 ( .B1(n6799), .B2(n6798), .A(n6797), .ZN(U3472) );
  MUX2_X1 U7785 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6800), .Z(U3473) );
  INV_X1 U7786 ( .A(n6801), .ZN(n6820) );
  INV_X1 U7787 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6803) );
  NAND4_X1 U7788 ( .A1(n6803), .A2(n6802), .A3(INSTQUEUE_REG_12__7__SCAN_IN), 
        .A4(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U7789 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), 
        .ZN(n6804) );
  NOR3_X1 U7790 ( .A1(n6806), .A2(n6805), .A3(n6804), .ZN(n6817) );
  INV_X1 U7791 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6862) );
  AND4_X1 U7792 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__0__SCAN_IN), .A3(n6862), .A4(n6991), .ZN(n6816) );
  OR4_X1 U7793 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(
        INSTQUEUE_REG_8__1__SCAN_IN), .A3(INSTQUEUE_REG_15__1__SCAN_IN), .A4(
        n3324), .ZN(n6808) );
  NOR2_X1 U7794 ( .A1(n6808), .A2(n6807), .ZN(n6809) );
  NAND4_X1 U7795 ( .A1(n7027), .A2(n6810), .A3(n7028), .A4(n6809), .ZN(n6814)
         );
  INV_X1 U7796 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6812) );
  INV_X1 U7797 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6811) );
  NAND4_X1 U7798 ( .A1(n6812), .A2(n6811), .A3(n3288), .A4(
        INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U7799 ( .A1(n6814), .A2(n6813), .ZN(n6815) );
  NAND4_X1 U7800 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6819)
         );
  NOR2_X1 U7801 ( .A1(n6820), .A2(n6819), .ZN(n6860) );
  NAND4_X1 U7802 ( .A1(DATAI_13_), .A2(DATAWIDTH_REG_25__SCAN_IN), .A3(n7044), 
        .A4(n6821), .ZN(n6822) );
  NOR3_X1 U7803 ( .A1(REIP_REG_29__SCAN_IN), .A2(LWORD_REG_9__SCAN_IN), .A3(
        n6822), .ZN(n6836) );
  INV_X1 U7804 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6984) );
  NOR4_X1 U7805 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(
        INSTQUEUE_REG_4__5__SCAN_IN), .A3(INSTQUEUE_REG_14__2__SCAN_IN), .A4(
        n6984), .ZN(n6834) );
  INV_X1 U7806 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6824) );
  OR4_X1 U7807 ( .A1(n6824), .A2(n6823), .A3(INSTQUEUE_REG_12__3__SCAN_IN), 
        .A4(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6831) );
  NAND4_X1 U7808 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        REIP_REG_26__SCAN_IN), .A3(DATAI_31_), .A4(ADDRESS_REG_17__SCAN_IN), 
        .ZN(n6830) );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6825) );
  NOR4_X1 U7810 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(
        INSTQUEUE_REG_4__2__SCAN_IN), .A3(INSTQUEUE_REG_10__2__SCAN_IN), .A4(
        n6825), .ZN(n6826) );
  INV_X1 U7811 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6940) );
  NAND4_X1 U7812 ( .A1(n6827), .A2(n6826), .A3(n7089), .A4(
        INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6829) );
  INV_X1 U7813 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6828) );
  NOR4_X1 U7814 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6833)
         );
  INV_X1 U7815 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6945) );
  NOR4_X1 U7816 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(
        INSTQUEUE_REG_8__6__SCAN_IN), .A3(n6922), .A4(n6945), .ZN(n6832) );
  AND3_X1 U7817 ( .A1(n6834), .A2(n6833), .A3(n6832), .ZN(n6835) );
  NAND4_X1 U7818 ( .A1(DATAO_REG_26__SCAN_IN), .A2(n6836), .A3(n6835), .A4(
        n7094), .ZN(n6858) );
  NOR4_X1 U7819 ( .A1(W_R_N_REG_SCAN_IN), .A2(EAX_REG_22__SCAN_IN), .A3(
        LWORD_REG_12__SCAN_IN), .A4(n4645), .ZN(n6840) );
  NOR4_X1 U7820 ( .A1(n6869), .A2(n7033), .A3(n7011), .A4(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6839) );
  INV_X1 U7821 ( .A(DATAI_8_), .ZN(n6875) );
  NOR4_X1 U7822 ( .A1(n4195), .A2(n6875), .A3(n6879), .A4(n6878), .ZN(n6838)
         );
  NOR4_X1 U7823 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .A3(PHYADDRPOINTER_REG_4__SCAN_IN), 
        .A4(n4506), .ZN(n6837) );
  NAND4_X1 U7824 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6857)
         );
  NOR4_X1 U7825 ( .A1(HOLD), .A2(UWORD_REG_3__SCAN_IN), .A3(
        ADDRESS_REG_20__SCAN_IN), .A4(n6998), .ZN(n6844) );
  INV_X1 U7826 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n7071) );
  NOR4_X1 U7827 ( .A1(DATAI_7_), .A2(LWORD_REG_2__SCAN_IN), .A3(n7071), .A4(
        n7077), .ZN(n6843) );
  NOR4_X1 U7828 ( .A1(EAX_REG_21__SCAN_IN), .A2(DATAO_REG_5__SCAN_IN), .A3(
        n6981), .A4(n6987), .ZN(n6842) );
  NOR4_X1 U7829 ( .A1(EBX_REG_30__SCAN_IN), .A2(CODEFETCH_REG_SCAN_IN), .A3(
        ADDRESS_REG_26__SCAN_IN), .A4(n6985), .ZN(n6841) );
  NAND4_X1 U7830 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6856)
         );
  NAND4_X1 U7831 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_24__SCAN_IN), 
        .A3(LWORD_REG_11__SCAN_IN), .A4(n6891), .ZN(n6845) );
  NOR3_X1 U7832 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4651), .A3(n6845), .ZN(n6854) );
  NOR4_X1 U7833 ( .A1(EAX_REG_25__SCAN_IN), .A2(BYTEENABLE_REG_2__SCAN_IN), 
        .A3(n6967), .A4(n5655), .ZN(n6846) );
  NAND3_X1 U7834 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(NA_N), .A3(n6846), .ZN(
        n6852) );
  NOR4_X1 U7835 ( .A1(DATAI_16_), .A2(DATAO_REG_27__SCAN_IN), .A3(
        LWORD_REG_13__SCAN_IN), .A4(n6928), .ZN(n6850) );
  NOR4_X1 U7836 ( .A1(EBX_REG_4__SCAN_IN), .A2(BYTEENABLE_REG_1__SCAN_IN), 
        .A3(DATAO_REG_3__SCAN_IN), .A4(n6912), .ZN(n6849) );
  NOR4_X1 U7837 ( .A1(EBX_REG_27__SCAN_IN), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .A3(EAX_REG_2__SCAN_IN), .A4(DATAO_REG_8__SCAN_IN), .ZN(n6848) );
  NOR4_X1 U7838 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        LWORD_REG_8__SCAN_IN), .A3(n6937), .A4(n6943), .ZN(n6847) );
  NAND4_X1 U7839 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6851)
         );
  NOR4_X1 U7840 ( .A1(n4601), .A2(n4644), .A3(n6852), .A4(n6851), .ZN(n6853)
         );
  NAND4_X1 U7841 ( .A1(n6854), .A2(n6853), .A3(n6909), .A4(n6906), .ZN(n6855)
         );
  NOR4_X1 U7842 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6859)
         );
  AOI21_X1 U7843 ( .B1(n6860), .B2(n6859), .A(DATAO_REG_23__SCAN_IN), .ZN(
        n7109) );
  AOI22_X1 U7844 ( .A1(n6862), .A2(keyinput71), .B1(keyinput9), .B2(n4020), 
        .ZN(n6861) );
  OAI221_X1 U7845 ( .B1(n6862), .B2(keyinput71), .C1(n4020), .C2(keyinput9), 
        .A(n6861), .ZN(n6873) );
  INV_X1 U7846 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7847 ( .A1(n6865), .A2(keyinput50), .B1(keyinput57), .B2(n6864), 
        .ZN(n6863) );
  OAI221_X1 U7848 ( .B1(n6865), .B2(keyinput50), .C1(n6864), .C2(keyinput57), 
        .A(n6863), .ZN(n6872) );
  XOR2_X1 U7849 ( .A(n4385), .B(keyinput2), .Z(n6868) );
  XNOR2_X1 U7850 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput43), .ZN(
        n6867) );
  XNOR2_X1 U7851 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .B(keyinput113), .ZN(
        n6866) );
  NAND3_X1 U7852 ( .A1(n6868), .A2(n6867), .A3(n6866), .ZN(n6871) );
  XNOR2_X1 U7853 ( .A(n6869), .B(keyinput24), .ZN(n6870) );
  NOR4_X1 U7854 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6920)
         );
  AOI22_X1 U7855 ( .A1(n6876), .A2(keyinput41), .B1(keyinput22), .B2(n6875), 
        .ZN(n6874) );
  OAI221_X1 U7856 ( .B1(n6876), .B2(keyinput41), .C1(n6875), .C2(keyinput22), 
        .A(n6874), .ZN(n6886) );
  AOI22_X1 U7857 ( .A1(n6879), .A2(keyinput17), .B1(keyinput86), .B2(n6878), 
        .ZN(n6877) );
  OAI221_X1 U7858 ( .B1(n6879), .B2(keyinput17), .C1(n6878), .C2(keyinput86), 
        .A(n6877), .ZN(n6885) );
  AOI22_X1 U7859 ( .A1(n5517), .A2(keyinput76), .B1(n4195), .B2(keyinput16), 
        .ZN(n6880) );
  OAI221_X1 U7860 ( .B1(n5517), .B2(keyinput76), .C1(n4195), .C2(keyinput16), 
        .A(n6880), .ZN(n6884) );
  XNOR2_X1 U7861 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(keyinput62), .ZN(
        n6882) );
  XNOR2_X1 U7862 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .B(keyinput28), .ZN(n6881)
         );
  NAND2_X1 U7863 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  NOR4_X1 U7864 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6919)
         );
  INV_X1 U7865 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6889) );
  AOI22_X1 U7866 ( .A1(n6889), .A2(keyinput122), .B1(keyinput54), .B2(n6888), 
        .ZN(n6887) );
  OAI221_X1 U7867 ( .B1(n6889), .B2(keyinput122), .C1(n6888), .C2(keyinput54), 
        .A(n6887), .ZN(n6901) );
  AOI22_X1 U7868 ( .A1(n4651), .A2(keyinput35), .B1(n6891), .B2(keyinput91), 
        .ZN(n6890) );
  OAI221_X1 U7869 ( .B1(n4651), .B2(keyinput35), .C1(n6891), .C2(keyinput91), 
        .A(n6890), .ZN(n6900) );
  INV_X1 U7870 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7871 ( .A1(n6894), .A2(keyinput21), .B1(n6893), .B2(keyinput42), 
        .ZN(n6892) );
  OAI221_X1 U7872 ( .B1(n6894), .B2(keyinput21), .C1(n6893), .C2(keyinput42), 
        .A(n6892), .ZN(n6899) );
  INV_X1 U7873 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7874 ( .A1(n6897), .A2(keyinput60), .B1(n6896), .B2(keyinput100), 
        .ZN(n6895) );
  OAI221_X1 U7875 ( .B1(n6897), .B2(keyinput60), .C1(n6896), .C2(keyinput100), 
        .A(n6895), .ZN(n6898) );
  NOR4_X1 U7876 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6918)
         );
  AOI22_X1 U7877 ( .A1(n6904), .A2(keyinput79), .B1(keyinput101), .B2(n6903), 
        .ZN(n6902) );
  OAI221_X1 U7878 ( .B1(n6904), .B2(keyinput79), .C1(n6903), .C2(keyinput101), 
        .A(n6902), .ZN(n6916) );
  INV_X1 U7879 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6907) );
  AOI22_X1 U7880 ( .A1(n6907), .A2(keyinput67), .B1(keyinput11), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U7881 ( .B1(n6907), .B2(keyinput67), .C1(n6906), .C2(keyinput11), 
        .A(n6905), .ZN(n6915) );
  AOI22_X1 U7882 ( .A1(n4378), .A2(keyinput48), .B1(n6909), .B2(keyinput4), 
        .ZN(n6908) );
  OAI221_X1 U7883 ( .B1(n4378), .B2(keyinput48), .C1(n6909), .C2(keyinput4), 
        .A(n6908), .ZN(n6914) );
  AOI22_X1 U7884 ( .A1(n6912), .A2(keyinput94), .B1(keyinput83), .B2(n6911), 
        .ZN(n6910) );
  OAI221_X1 U7885 ( .B1(n6912), .B2(keyinput94), .C1(n6911), .C2(keyinput83), 
        .A(n6910), .ZN(n6913) );
  NOR4_X1 U7886 ( .A1(n6916), .A2(n6915), .A3(n6914), .A4(n6913), .ZN(n6917)
         );
  NAND4_X1 U7887 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(n7107)
         );
  AOI22_X1 U7888 ( .A1(n6923), .A2(keyinput69), .B1(n6922), .B2(keyinput3), 
        .ZN(n6921) );
  OAI221_X1 U7889 ( .B1(n6923), .B2(keyinput69), .C1(n6922), .C2(keyinput3), 
        .A(n6921), .ZN(n6935) );
  INV_X1 U7890 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U7891 ( .A1(n6926), .A2(keyinput108), .B1(n6925), .B2(keyinput126), 
        .ZN(n6924) );
  OAI221_X1 U7892 ( .B1(n6926), .B2(keyinput108), .C1(n6925), .C2(keyinput126), 
        .A(n6924), .ZN(n6934) );
  AOI22_X1 U7893 ( .A1(n6929), .A2(keyinput39), .B1(keyinput45), .B2(n6928), 
        .ZN(n6927) );
  OAI221_X1 U7894 ( .B1(n6929), .B2(keyinput39), .C1(n6928), .C2(keyinput45), 
        .A(n6927), .ZN(n6933) );
  AOI22_X1 U7895 ( .A1(n4746), .A2(keyinput47), .B1(keyinput87), .B2(n6931), 
        .ZN(n6930) );
  OAI221_X1 U7896 ( .B1(n4746), .B2(keyinput47), .C1(n6931), .C2(keyinput87), 
        .A(n6930), .ZN(n6932) );
  NOR4_X1 U7897 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(n6979)
         );
  AOI22_X1 U7898 ( .A1(n6937), .A2(keyinput115), .B1(keyinput18), .B2(n5462), 
        .ZN(n6936) );
  OAI221_X1 U7899 ( .B1(n6937), .B2(keyinput115), .C1(n5462), .C2(keyinput18), 
        .A(n6936), .ZN(n6949) );
  INV_X1 U7900 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6939) );
  AOI22_X1 U7901 ( .A1(n6940), .A2(keyinput44), .B1(keyinput119), .B2(n6939), 
        .ZN(n6938) );
  OAI221_X1 U7902 ( .B1(n6940), .B2(keyinput44), .C1(n6939), .C2(keyinput119), 
        .A(n6938), .ZN(n6948) );
  INV_X1 U7903 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7904 ( .A1(n6943), .A2(keyinput65), .B1(keyinput49), .B2(n6942), 
        .ZN(n6941) );
  OAI221_X1 U7905 ( .B1(n6943), .B2(keyinput65), .C1(n6942), .C2(keyinput49), 
        .A(n6941), .ZN(n6947) );
  AOI22_X1 U7906 ( .A1(n5658), .A2(keyinput34), .B1(n6945), .B2(keyinput14), 
        .ZN(n6944) );
  OAI221_X1 U7907 ( .B1(n5658), .B2(keyinput34), .C1(n6945), .C2(keyinput14), 
        .A(n6944), .ZN(n6946) );
  NOR4_X1 U7908 ( .A1(n6949), .A2(n6948), .A3(n6947), .A4(n6946), .ZN(n6978)
         );
  AOI22_X1 U7909 ( .A1(n6952), .A2(keyinput114), .B1(n6951), .B2(keyinput31), 
        .ZN(n6950) );
  OAI221_X1 U7910 ( .B1(n6952), .B2(keyinput114), .C1(n6951), .C2(keyinput31), 
        .A(n6950), .ZN(n6961) );
  AOI22_X1 U7911 ( .A1(n5655), .A2(keyinput75), .B1(n6812), .B2(keyinput8), 
        .ZN(n6953) );
  OAI221_X1 U7912 ( .B1(n5655), .B2(keyinput75), .C1(n6812), .C2(keyinput8), 
        .A(n6953), .ZN(n6960) );
  AOI22_X1 U7913 ( .A1(n6955), .A2(keyinput55), .B1(n4601), .B2(keyinput70), 
        .ZN(n6954) );
  OAI221_X1 U7914 ( .B1(n6955), .B2(keyinput55), .C1(n4601), .C2(keyinput70), 
        .A(n6954), .ZN(n6959) );
  AOI22_X1 U7915 ( .A1(n4644), .A2(keyinput78), .B1(keyinput58), .B2(n6957), 
        .ZN(n6956) );
  OAI221_X1 U7916 ( .B1(n4644), .B2(keyinput78), .C1(n6957), .C2(keyinput58), 
        .A(n6956), .ZN(n6958) );
  NOR4_X1 U7917 ( .A1(n6961), .A2(n6960), .A3(n6959), .A4(n6958), .ZN(n6977)
         );
  AOI22_X1 U7918 ( .A1(n6963), .A2(keyinput84), .B1(n3998), .B2(keyinput33), 
        .ZN(n6962) );
  OAI221_X1 U7919 ( .B1(n6963), .B2(keyinput84), .C1(n3998), .C2(keyinput33), 
        .A(n6962), .ZN(n6975) );
  AOI22_X1 U7920 ( .A1(n6803), .A2(keyinput102), .B1(keyinput125), .B2(n6965), 
        .ZN(n6964) );
  OAI221_X1 U7921 ( .B1(n6803), .B2(keyinput102), .C1(n6965), .C2(keyinput125), 
        .A(n6964), .ZN(n6974) );
  AOI22_X1 U7922 ( .A1(n6968), .A2(keyinput93), .B1(keyinput95), .B2(n6967), 
        .ZN(n6966) );
  OAI221_X1 U7923 ( .B1(n6968), .B2(keyinput93), .C1(n6967), .C2(keyinput95), 
        .A(n6966), .ZN(n6973) );
  XOR2_X1 U7924 ( .A(n6969), .B(keyinput23), .Z(n6971) );
  XNOR2_X1 U7925 ( .A(STATE2_REG_1__SCAN_IN), .B(keyinput81), .ZN(n6970) );
  NAND2_X1 U7926 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  NOR4_X1 U7927 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n6976)
         );
  NAND4_X1 U7928 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n7106)
         );
  AOI22_X1 U7929 ( .A1(n6982), .A2(keyinput124), .B1(n6981), .B2(keyinput38), 
        .ZN(n6980) );
  OAI221_X1 U7930 ( .B1(n6982), .B2(keyinput124), .C1(n6981), .C2(keyinput38), 
        .A(n6980), .ZN(n6995) );
  AOI22_X1 U7931 ( .A1(n6985), .A2(keyinput25), .B1(n6984), .B2(keyinput127), 
        .ZN(n6983) );
  OAI221_X1 U7932 ( .B1(n6985), .B2(keyinput25), .C1(n6984), .C2(keyinput127), 
        .A(n6983), .ZN(n6994) );
  AOI22_X1 U7933 ( .A1(n6988), .A2(keyinput106), .B1(n6987), .B2(keyinput104), 
        .ZN(n6986) );
  OAI221_X1 U7934 ( .B1(n6988), .B2(keyinput106), .C1(n6987), .C2(keyinput104), 
        .A(n6986), .ZN(n6993) );
  AOI22_X1 U7935 ( .A1(n6991), .A2(keyinput19), .B1(keyinput20), .B2(n6990), 
        .ZN(n6989) );
  OAI221_X1 U7936 ( .B1(n6991), .B2(keyinput19), .C1(n6990), .C2(keyinput20), 
        .A(n6989), .ZN(n6992) );
  NOR4_X1 U7937 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n7042)
         );
  AOI22_X1 U7938 ( .A1(n6998), .A2(keyinput37), .B1(keyinput12), .B2(n6997), 
        .ZN(n6996) );
  OAI221_X1 U7939 ( .B1(n6998), .B2(keyinput37), .C1(n6997), .C2(keyinput12), 
        .A(n6996), .ZN(n7009) );
  AOI22_X1 U7940 ( .A1(n7001), .A2(keyinput74), .B1(keyinput64), .B2(n7000), 
        .ZN(n6999) );
  OAI221_X1 U7941 ( .B1(n7001), .B2(keyinput74), .C1(n7000), .C2(keyinput64), 
        .A(n6999), .ZN(n7008) );
  AOI22_X1 U7942 ( .A1(n4497), .A2(keyinput61), .B1(keyinput27), .B2(n7003), 
        .ZN(n7002) );
  OAI221_X1 U7943 ( .B1(n4497), .B2(keyinput61), .C1(n7003), .C2(keyinput27), 
        .A(n7002), .ZN(n7007) );
  INV_X1 U7944 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n7005) );
  AOI22_X1 U7945 ( .A1(n3904), .A2(keyinput103), .B1(keyinput80), .B2(n7005), 
        .ZN(n7004) );
  OAI221_X1 U7946 ( .B1(n3904), .B2(keyinput103), .C1(n7005), .C2(keyinput80), 
        .A(n7004), .ZN(n7006) );
  NOR4_X1 U7947 ( .A1(n7009), .A2(n7008), .A3(n7007), .A4(n7006), .ZN(n7041)
         );
  AOI22_X1 U7948 ( .A1(n7012), .A2(keyinput73), .B1(keyinput99), .B2(n7011), 
        .ZN(n7010) );
  OAI221_X1 U7949 ( .B1(n7012), .B2(keyinput73), .C1(n7011), .C2(keyinput99), 
        .A(n7010), .ZN(n7022) );
  AOI22_X1 U7950 ( .A1(n7015), .A2(keyinput88), .B1(n7014), .B2(keyinput0), 
        .ZN(n7013) );
  OAI221_X1 U7951 ( .B1(n7015), .B2(keyinput88), .C1(n7014), .C2(keyinput0), 
        .A(n7013), .ZN(n7021) );
  XNOR2_X1 U7952 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput66), .ZN(n7019)
         );
  XNOR2_X1 U7953 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput77), .ZN(n7018)
         );
  XNOR2_X1 U7954 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(keyinput89), .ZN(
        n7017) );
  XNOR2_X1 U7955 ( .A(keyinput72), .B(EAX_REG_16__SCAN_IN), .ZN(n7016) );
  NAND4_X1 U7956 ( .A1(n7019), .A2(n7018), .A3(n7017), .A4(n7016), .ZN(n7020)
         );
  NOR3_X1 U7957 ( .A1(n7022), .A2(n7021), .A3(n7020), .ZN(n7040) );
  AOI22_X1 U7958 ( .A1(n4189), .A2(keyinput6), .B1(keyinput90), .B2(n7024), 
        .ZN(n7023) );
  OAI221_X1 U7959 ( .B1(n4189), .B2(keyinput6), .C1(n7024), .C2(keyinput90), 
        .A(n7023), .ZN(n7031) );
  AOI22_X1 U7960 ( .A1(n7027), .A2(keyinput118), .B1(keyinput85), .B2(n7026), 
        .ZN(n7025) );
  OAI221_X1 U7961 ( .B1(n7027), .B2(keyinput118), .C1(n7026), .C2(keyinput85), 
        .A(n7025), .ZN(n7030) );
  XNOR2_X1 U7962 ( .A(n7028), .B(keyinput32), .ZN(n7029) );
  OR3_X1 U7963 ( .A1(n7031), .A2(n7030), .A3(n7029), .ZN(n7038) );
  INV_X1 U7964 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n7034) );
  AOI22_X1 U7965 ( .A1(n7034), .A2(keyinput121), .B1(keyinput52), .B2(n7033), 
        .ZN(n7032) );
  OAI221_X1 U7966 ( .B1(n7034), .B2(keyinput121), .C1(n7033), .C2(keyinput52), 
        .A(n7032), .ZN(n7037) );
  XNOR2_X1 U7967 ( .A(n7035), .B(keyinput36), .ZN(n7036) );
  NOR3_X1 U7968 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(n7039) );
  NAND4_X1 U7969 ( .A1(n7042), .A2(n7041), .A3(n7040), .A4(n7039), .ZN(n7105)
         );
  AOI22_X1 U7970 ( .A1(n7045), .A2(keyinput46), .B1(n7044), .B2(keyinput56), 
        .ZN(n7043) );
  OAI221_X1 U7971 ( .B1(n7045), .B2(keyinput46), .C1(n7044), .C2(keyinput56), 
        .A(n7043), .ZN(n7056) );
  INV_X1 U7972 ( .A(DATAI_31_), .ZN(n7048) );
  AOI22_X1 U7973 ( .A1(n7048), .A2(keyinput63), .B1(n7047), .B2(keyinput120), 
        .ZN(n7046) );
  OAI221_X1 U7974 ( .B1(n7048), .B2(keyinput63), .C1(n7047), .C2(keyinput120), 
        .A(n7046), .ZN(n7055) );
  XOR2_X1 U7975 ( .A(n7049), .B(keyinput96), .Z(n7053) );
  XNOR2_X1 U7976 ( .A(keyinput111), .B(EAX_REG_30__SCAN_IN), .ZN(n7052) );
  XNOR2_X1 U7977 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .B(keyinput68), .ZN(n7051) );
  XNOR2_X1 U7978 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput92), .ZN(n7050)
         );
  NAND4_X1 U7979 ( .A1(n7053), .A2(n7052), .A3(n7051), .A4(n7050), .ZN(n7054)
         );
  NOR3_X1 U7980 ( .A1(n7056), .A2(n7055), .A3(n7054), .ZN(n7103) );
  AOI22_X1 U7981 ( .A1(keyinput53), .A2(n6828), .B1(keyinput117), .B2(n7057), 
        .ZN(n7058) );
  OAI21_X1 U7982 ( .B1(n6828), .B2(keyinput53), .A(n7058), .ZN(n7069) );
  AOI22_X1 U7983 ( .A1(n6811), .A2(keyinput10), .B1(keyinput123), .B2(n6823), 
        .ZN(n7059) );
  OAI221_X1 U7984 ( .B1(n6811), .B2(keyinput10), .C1(n6823), .C2(keyinput123), 
        .A(n7059), .ZN(n7068) );
  INV_X1 U7985 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U7986 ( .A1(n7062), .A2(keyinput109), .B1(n7061), .B2(keyinput82), 
        .ZN(n7060) );
  OAI221_X1 U7987 ( .B1(n7062), .B2(keyinput109), .C1(n7061), .C2(keyinput82), 
        .A(n7060), .ZN(n7067) );
  AOI22_X1 U7988 ( .A1(n7065), .A2(keyinput51), .B1(n7064), .B2(keyinput98), 
        .ZN(n7063) );
  OAI221_X1 U7989 ( .B1(n7065), .B2(keyinput51), .C1(n7064), .C2(keyinput98), 
        .A(n7063), .ZN(n7066) );
  NOR4_X1 U7990 ( .A1(n7069), .A2(n7068), .A3(n7067), .A4(n7066), .ZN(n7102)
         );
  INV_X1 U7991 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n7072) );
  AOI22_X1 U7992 ( .A1(n7072), .A2(keyinput112), .B1(keyinput105), .B2(n7071), 
        .ZN(n7070) );
  OAI221_X1 U7993 ( .B1(n7072), .B2(keyinput112), .C1(n7071), .C2(keyinput105), 
        .A(n7070), .ZN(n7084) );
  INV_X1 U7994 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n7074) );
  AOI22_X1 U7995 ( .A1(n7075), .A2(keyinput110), .B1(n7074), .B2(keyinput7), 
        .ZN(n7073) );
  OAI221_X1 U7996 ( .B1(n7075), .B2(keyinput110), .C1(n7074), .C2(keyinput7), 
        .A(n7073), .ZN(n7083) );
  AOI22_X1 U7997 ( .A1(n7077), .A2(keyinput107), .B1(n3324), .B2(keyinput5), 
        .ZN(n7076) );
  OAI221_X1 U7998 ( .B1(n7077), .B2(keyinput107), .C1(n3324), .C2(keyinput5), 
        .A(n7076), .ZN(n7082) );
  AOI22_X1 U7999 ( .A1(n7080), .A2(keyinput26), .B1(n7079), .B2(keyinput116), 
        .ZN(n7078) );
  OAI221_X1 U8000 ( .B1(n7080), .B2(keyinput26), .C1(n7079), .C2(keyinput116), 
        .A(n7078), .ZN(n7081) );
  NOR4_X1 U8001 ( .A1(n7084), .A2(n7083), .A3(n7082), .A4(n7081), .ZN(n7101)
         );
  INV_X1 U8002 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n7086) );
  AOI22_X1 U8003 ( .A1(n7086), .A2(keyinput59), .B1(keyinput29), .B2(n5740), 
        .ZN(n7085) );
  OAI221_X1 U8004 ( .B1(n7086), .B2(keyinput59), .C1(n5740), .C2(keyinput29), 
        .A(n7085), .ZN(n7099) );
  INV_X1 U8005 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n7088) );
  AOI22_X1 U8006 ( .A1(n7089), .A2(keyinput30), .B1(n7088), .B2(keyinput13), 
        .ZN(n7087) );
  OAI221_X1 U8007 ( .B1(n7089), .B2(keyinput30), .C1(n7088), .C2(keyinput13), 
        .A(n7087), .ZN(n7098) );
  AOI22_X1 U8008 ( .A1(n7092), .A2(keyinput15), .B1(n7091), .B2(keyinput1), 
        .ZN(n7090) );
  OAI221_X1 U8009 ( .B1(n7092), .B2(keyinput15), .C1(n7091), .C2(keyinput1), 
        .A(n7090), .ZN(n7097) );
  AOI22_X1 U8010 ( .A1(n7095), .A2(keyinput97), .B1(n7094), .B2(keyinput40), 
        .ZN(n7093) );
  OAI221_X1 U8011 ( .B1(n7095), .B2(keyinput97), .C1(n7094), .C2(keyinput40), 
        .A(n7093), .ZN(n7096) );
  NOR4_X1 U8012 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7100)
         );
  NAND4_X1 U8013 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7104)
         );
  NOR4_X1 U8014 ( .A1(n7107), .A2(n7106), .A3(n7105), .A4(n7104), .ZN(n7108)
         );
  OAI21_X1 U8015 ( .B1(keyinput117), .B2(n7109), .A(n7108), .ZN(n7123) );
  NAND2_X1 U8016 ( .A1(n7110), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n7119) );
  OAI22_X1 U8017 ( .A1(n7114), .A2(n7113), .B1(n7112), .B2(n7111), .ZN(n7115)
         );
  AOI21_X1 U8018 ( .B1(n7117), .B2(n7116), .A(n7115), .ZN(n7118) );
  OAI211_X1 U8019 ( .C1(n7121), .C2(n7120), .A(n7119), .B(n7118), .ZN(n7122)
         );
  XNOR2_X1 U8020 ( .A(n7123), .B(n7122), .ZN(U3086) );
  BUF_X1 U3542 ( .A(n4285), .Z(n5388) );
  OR2_X1 U4186 ( .A1(n5365), .A2(n6207), .ZN(n3170) );
  CLKBUF_X1 U3565 ( .A(n3513), .Z(n3535) );
  CLKBUF_X1 U3568 ( .A(n3426), .Z(n4763) );
  CLKBUF_X1 U3978 ( .A(n3419), .Z(n4602) );
  CLKBUF_X1 U4560 ( .A(n4712), .Z(n5612) );
endmodule

