

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656;

  CLKBUF_X2 U3651 ( .A(n4519), .Z(n4724) );
  CLKBUF_X2 U3652 ( .A(n3846), .Z(n3937) );
  CLKBUF_X1 U3654 ( .A(n3860), .Z(n4229) );
  NAND2_X1 U3655 ( .A1(n3919), .A2(n3860), .ZN(n3904) );
  AND2_X2 U3656 ( .A1(n3667), .A2(n4939), .ZN(n3876) );
  CLKBUF_X1 U3657 ( .A(n7489), .Z(n3617) );
  NOR2_X1 U3658 ( .A1(n5744), .A2(n5743), .ZN(n7489) );
  AND2_X1 U3659 ( .A1(n3749), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3763)
         );
  AND2_X2 U3660 ( .A1(n4222), .A2(n5000), .ZN(n3951) );
  NAND2_X1 U3661 ( .A1(n3661), .A2(n5000), .ZN(n3924) );
  INV_X1 U3662 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U3663 ( .A1(n3856), .A2(n3652), .ZN(n3926) );
  BUF_X1 U3664 ( .A(n4777), .Z(n3644) );
  NOR2_X2 U3665 ( .A1(n5196), .A2(n3645), .ZN(n3925) );
  INV_X1 U3666 ( .A(n6443), .ZN(n3618) );
  CLKBUF_X3 U3667 ( .A(n4778), .Z(n4789) );
  OR2_X1 U3668 ( .A1(n4257), .A2(n4256), .ZN(n6115) );
  INV_X1 U3670 ( .A(n7483), .ZN(n7491) );
  NAND2_X2 U3671 ( .A1(n6384), .A2(n4195), .ZN(n6374) );
  AND2_X4 U3672 ( .A1(n3751), .A2(n5282), .ZN(n3851) );
  AND2_X4 U3673 ( .A1(n5268), .A2(n3743), .ZN(n4519) );
  AND2_X4 U3674 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4939) );
  AOI211_X2 U3675 ( .C1(n6600), .C2(n6599), .A(n6598), .B(n6597), .ZN(n6601)
         );
  NAND2_X1 U3676 ( .A1(n6463), .A2(n6462), .ZN(n6461) );
  NAND2_X1 U3677 ( .A1(n6048), .A2(n4174), .ZN(n6482) );
  NOR2_X2 U3678 ( .A1(n6131), .A2(n6070), .ZN(n6069) );
  OR2_X1 U3679 ( .A1(n6146), .A2(n6129), .ZN(n6131) );
  OR2_X1 U3680 ( .A1(n6184), .A2(n6172), .ZN(n6170) );
  CLKBUF_X2 U3681 ( .A(n5894), .Z(n5933) );
  NAND2_X1 U3682 ( .A1(n3969), .A2(n3970), .ZN(n4020) );
  OR2_X1 U3683 ( .A1(n4934), .A2(n3934), .ZN(n3970) );
  OAI21_X1 U3684 ( .B1(n3895), .B2(n3921), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3897) );
  NAND2_X1 U3685 ( .A1(n4985), .A2(n4229), .ZN(n4437) );
  NAND2_X4 U3686 ( .A1(n4969), .A2(n4789), .ZN(n4865) );
  NAND2_X4 U3687 ( .A1(n4792), .A2(n4789), .ZN(n4977) );
  NAND2_X2 U3688 ( .A1(n5069), .A2(n3645), .ZN(n4792) );
  NAND2_X1 U3689 ( .A1(n4967), .A2(n3900), .ZN(n3908) );
  NAND4_X1 U3690 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3857)
         );
  AOI21_X1 U3691 ( .B1(n4547), .B2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n3629), 
        .ZN(n3844) );
  CLKBUF_X2 U3692 ( .A(n4547), .Z(n4702) );
  BUF_X2 U3693 ( .A(n3974), .Z(n4677) );
  BUF_X2 U3694 ( .A(n4318), .Z(n4722) );
  BUF_X2 U3695 ( .A(n3867), .Z(n4708) );
  BUF_X2 U3696 ( .A(n4109), .Z(n4723) );
  AND2_X2 U3697 ( .A1(n3763), .A2(n3667), .ZN(n4109) );
  AND2_X2 U3698 ( .A1(n3763), .A2(n5279), .ZN(n4318) );
  CLKBUF_X2 U3699 ( .A(n4524), .Z(n4725) );
  CLKBUF_X2 U3700 ( .A(n3876), .Z(n4709) );
  CLKBUF_X2 U3701 ( .A(n4518), .Z(n4593) );
  AND2_X1 U3702 ( .A1(n3752), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3757)
         );
  NOR2_X4 U3703 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3667) );
  AOI21_X1 U3704 ( .B1(n6128), .B2(n6142), .A(n6066), .ZN(n6372) );
  AOI21_X1 U3705 ( .B1(n6143), .B2(n6141), .A(n6127), .ZN(n6382) );
  NAND2_X1 U3706 ( .A1(n6461), .A2(n3656), .ZN(n6446) );
  NAND2_X1 U3707 ( .A1(n6482), .A2(n3694), .ZN(n3690) );
  NAND2_X1 U3708 ( .A1(n3622), .A2(n4173), .ZN(n6048) );
  NAND2_X1 U3709 ( .A1(n6033), .A2(n6034), .ZN(n3622) );
  NAND2_X1 U3710 ( .A1(n3623), .A2(n4171), .ZN(n6033) );
  NAND2_X1 U3711 ( .A1(n5988), .A2(n5989), .ZN(n3623) );
  NOR2_X1 U3712 ( .A1(n3640), .A2(n6471), .ZN(n3639) );
  NAND2_X1 U3713 ( .A1(n3634), .A2(n7163), .ZN(n7162) );
  NAND2_X1 U3714 ( .A1(n7158), .A2(n4104), .ZN(n3634) );
  NOR2_X1 U3715 ( .A1(n3702), .A2(n3701), .ZN(n3700) );
  NAND2_X1 U3716 ( .A1(n4873), .A2(n4872), .ZN(n4875) );
  NAND2_X1 U3717 ( .A1(n4102), .A2(n4101), .ZN(n7158) );
  INV_X2 U3718 ( .A(n4172), .ZN(n6443) );
  OAI21_X1 U3719 ( .B1(n4317), .B2(n4418), .A(n4316), .ZN(n5701) );
  NAND2_X1 U3720 ( .A1(n3625), .A2(n3624), .ZN(n7157) );
  OAI21_X1 U3721 ( .B1(n5033), .B2(n5039), .A(n5034), .ZN(n3625) );
  NAND2_X1 U3722 ( .A1(n6164), .A2(n6144), .ZN(n6146) );
  AND2_X1 U3723 ( .A1(n4122), .A2(n4146), .ZN(n4301) );
  NAND2_X1 U3724 ( .A1(n3627), .A2(n3626), .ZN(n5033) );
  NOR2_X2 U3725 ( .A1(n6170), .A2(n6165), .ZN(n6164) );
  NAND2_X2 U3726 ( .A1(n4086), .A2(n4052), .ZN(n5050) );
  NOR2_X1 U3727 ( .A1(n4965), .A2(n5234), .ZN(n4276) );
  NOR2_X1 U3728 ( .A1(n5051), .A2(n3655), .ZN(n3709) );
  NOR3_X1 U3729 ( .A1(n6313), .A2(n6302), .A3(n3675), .ZN(n6221) );
  NAND2_X1 U3730 ( .A1(n4001), .A2(n4000), .ZN(n3635) );
  CLKBUF_X1 U3731 ( .A(n5045), .Z(n6703) );
  OR2_X2 U3732 ( .A1(n7183), .A2(n7146), .ZN(n7190) );
  NOR2_X1 U3733 ( .A1(n6647), .A2(n4826), .ZN(n6640) );
  OR2_X1 U3734 ( .A1(n6021), .A2(n6022), .ZN(n6647) );
  NAND2_X1 U3735 ( .A1(n4030), .A2(n4031), .ZN(n5286) );
  NAND2_X1 U3736 ( .A1(n3989), .A2(n4003), .ZN(n4006) );
  OR2_X1 U3737 ( .A1(n5977), .A2(n6003), .ZN(n6021) );
  NOR2_X1 U3738 ( .A1(n5782), .A2(n3658), .ZN(n5979) );
  NAND2_X1 U3739 ( .A1(n7138), .A2(n4798), .ZN(n5782) );
  NOR2_X2 U3740 ( .A1(n7136), .A2(n7135), .ZN(n7138) );
  OR2_X1 U3741 ( .A1(n6088), .A2(n5025), .ZN(n7136) );
  NAND2_X1 U3742 ( .A1(n3918), .A2(n3917), .ZN(n3969) );
  AOI21_X1 U3743 ( .B1(n3668), .B2(n4969), .A(n3669), .ZN(n6087) );
  NAND2_X1 U3744 ( .A1(n3897), .A2(n3896), .ZN(n4024) );
  OAI211_X1 U3745 ( .C1(n4764), .C2(n3909), .A(n4903), .B(n3646), .ZN(n3910)
         );
  OR2_X1 U3746 ( .A1(n4004), .A2(n4003), .ZN(n4005) );
  NOR2_X2 U3747 ( .A1(n4260), .A2(n3906), .ZN(n4772) );
  INV_X1 U3748 ( .A(n3924), .ZN(n4985) );
  AND2_X2 U3749 ( .A1(n3929), .A2(n3903), .ZN(n4907) );
  BUF_X2 U3750 ( .A(n4780), .Z(n4975) );
  AND2_X1 U3751 ( .A1(n5230), .A2(n3902), .ZN(n3929) );
  OR2_X1 U3752 ( .A1(n3904), .A2(n4778), .ZN(n4936) );
  AND2_X2 U3753 ( .A1(n4229), .A2(n5196), .ZN(n4984) );
  OR2_X1 U3754 ( .A1(n3961), .A2(n3960), .ZN(n4166) );
  AND2_X1 U3755 ( .A1(n3901), .A2(n3900), .ZN(n5230) );
  NAND4_X1 U3756 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n4777)
         );
  INV_X1 U3757 ( .A(n3919), .ZN(n5000) );
  CLKBUF_X1 U3758 ( .A(n3919), .Z(n3920) );
  BUF_X2 U3759 ( .A(n3857), .Z(n5196) );
  AND4_X2 U3760 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n5073)
         );
  AND4_X1 U3761 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3882)
         );
  AND4_X1 U3762 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  AND4_X1 U3763 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  AND4_X1 U3764 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3883)
         );
  AND4_X1 U3765 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3769)
         );
  AND3_X1 U3766 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n3792) );
  AND4_X1 U3767 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3884)
         );
  AND4_X1 U3768 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3791)
         );
  AND4_X1 U3769 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3801)
         );
  AND4_X1 U3770 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AND4_X1 U3771 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3802)
         );
  AND4_X1 U3772 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  AND4_X1 U3773 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3843)
         );
  AND4_X1 U3774 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AND4_X1 U3775 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  AND4_X1 U3776 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3887)
         );
  AND4_X1 U3777 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3771)
         );
  AND4_X1 U3778 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3770)
         );
  AND4_X1 U3779 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3889)
         );
  AND4_X1 U3780 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3888)
         );
  BUF_X2 U3781 ( .A(n3866), .Z(n4730) );
  BUF_X2 U3782 ( .A(n3942), .Z(n4700) );
  BUF_X2 U3783 ( .A(n4065), .Z(n3936) );
  BUF_X2 U3784 ( .A(n3845), .Z(n4707) );
  BUF_X2 U3785 ( .A(n3851), .Z(n4731) );
  AND2_X1 U3786 ( .A1(n3773), .A2(n3772), .ZN(n3774) );
  NAND2_X1 U3787 ( .A1(n4065), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3632) );
  NAND2_X1 U3788 ( .A1(n3866), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3631)
         );
  NAND2_X1 U3789 ( .A1(n3867), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3630)
         );
  CLKBUF_X2 U3790 ( .A(n3861), .Z(n4547) );
  INV_X2 U3791 ( .A(n7553), .ZN(n7556) );
  AND2_X1 U3792 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5268) );
  NOR2_X1 U3793 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3743) );
  INV_X1 U3794 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3628) );
  INV_X1 U3795 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3750) );
  NOR2_X2 U3796 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4286) );
  NAND2_X2 U3797 ( .A1(n3620), .A2(n3619), .ZN(n4086) );
  INV_X1 U3798 ( .A(n3621), .ZN(n3619) );
  INV_X1 U3799 ( .A(n4051), .ZN(n3620) );
  NAND2_X1 U3800 ( .A1(n4051), .A2(n3621), .ZN(n4052) );
  OAI21_X2 U3801 ( .B1(n4018), .B2(n4017), .A(n3638), .ZN(n3621) );
  AOI21_X2 U3802 ( .B1(n7162), .B2(n3706), .A(n3705), .ZN(n5952) );
  NAND2_X1 U3803 ( .A1(n5033), .A2(n5039), .ZN(n3624) );
  NAND2_X1 U3804 ( .A1(n3633), .A2(n7259), .ZN(n3626) );
  OAI21_X1 U3805 ( .B1(n3633), .B2(n7259), .A(n7150), .ZN(n3627) );
  NOR2_X2 U3806 ( .A1(n3628), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3762)
         );
  XNOR2_X2 U3807 ( .A(n6422), .B(n6421), .ZN(n6596) );
  AND2_X2 U3808 ( .A1(n3636), .A2(n6401), .ZN(n6422) );
  OR2_X2 U3809 ( .A1(n6427), .A2(n6426), .ZN(n3636) );
  NAND3_X1 U3810 ( .A1(n3632), .A2(n3631), .A3(n3630), .ZN(n3629) );
  AND2_X2 U3811 ( .A1(n3757), .A2(n5279), .ZN(n3867) );
  AND2_X2 U3812 ( .A1(n3762), .A2(n3757), .ZN(n3866) );
  AND2_X2 U3813 ( .A1(n3762), .A2(n3763), .ZN(n4065) );
  XNOR2_X1 U3814 ( .A(n7151), .B(n3633), .ZN(n7257) );
  NAND2_X1 U3815 ( .A1(n4015), .A2(n5134), .ZN(n3633) );
  AOI21_X2 U3816 ( .B1(n3690), .B2(n3641), .A(n3639), .ZN(n6463) );
  NAND2_X1 U3817 ( .A1(n4163), .A2(n4162), .ZN(n5988) );
  OAI21_X1 U3818 ( .B1(n7163), .B2(n3634), .A(n7162), .ZN(n7241) );
  INV_X1 U3819 ( .A(n3635), .ZN(n4014) );
  NAND2_X1 U3820 ( .A1(n3635), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5133)
         );
  NAND3_X1 U3821 ( .A1(n6602), .A2(n7186), .A3(n3636), .ZN(n6431) );
  NAND3_X1 U3822 ( .A1(n6602), .A2(n7314), .A3(n3636), .ZN(n6608) );
  NAND2_X1 U3823 ( .A1(n3860), .A2(n4262), .ZN(n3637) );
  NAND2_X1 U3824 ( .A1(n3860), .A2(n4262), .ZN(n3901) );
  AND4_X2 U3825 ( .A1(n3889), .A2(n3887), .A3(n3888), .A4(n3886), .ZN(n4262)
         );
  OR2_X1 U3826 ( .A1(n6295), .A2(n6202), .ZN(n6287) );
  AND4_X1 U3827 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3886)
         );
  BUF_X4 U3828 ( .A(n4261), .Z(n5052) );
  XNOR2_X2 U3829 ( .A(n4018), .B(n4017), .ZN(n4261) );
  NOR2_X2 U3830 ( .A1(n6227), .A2(n6230), .ZN(n6229) );
  NAND2_X1 U3831 ( .A1(n3965), .A2(n3964), .ZN(n3638) );
  INV_X1 U3832 ( .A(n4175), .ZN(n3640) );
  AND2_X1 U3833 ( .A1(n3691), .A2(n4175), .ZN(n3641) );
  CLKBUF_X1 U3834 ( .A(n5988), .Z(n3642) );
  OAI21_X1 U3835 ( .B1(n5046), .B2(STATE2_REG_0__SCAN_IN), .A(n3950), .ZN(
        n3643) );
  NAND2_X1 U3836 ( .A1(n3965), .A2(n3964), .ZN(n4016) );
  OAI21_X1 U3837 ( .B1(n5046), .B2(STATE2_REG_0__SCAN_IN), .A(n3950), .ZN(
        n3967) );
  NAND2_X2 U3838 ( .A1(n4907), .A2(n3645), .ZN(n4764) );
  AOI21_X2 U3839 ( .B1(n3859), .B2(n3992), .A(n3858), .ZN(n3931) );
  NOR2_X1 U3840 ( .A1(n4928), .A2(n3860), .ZN(n4970) );
  BUF_X4 U3841 ( .A(n4777), .Z(n3645) );
  OAI21_X1 U3842 ( .B1(n5050), .B2(n4418), .A(n4605), .ZN(n5233) );
  AND2_X4 U3843 ( .A1(n3644), .A2(n3907), .ZN(n3992) );
  INV_X2 U3844 ( .A(n3644), .ZN(n3905) );
  AND2_X1 U3845 ( .A1(n3645), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4222) );
  AOI211_X1 U3846 ( .C1(n3992), .C2(n7535), .A(READY_N), .B(n7200), .ZN(n7201)
         );
  XNOR2_X1 U3847 ( .A(n4086), .B(n4085), .ZN(n5242) );
  NAND2_X2 U3848 ( .A1(n4016), .A2(n3968), .ZN(n4018) );
  INV_X2 U3849 ( .A(n3857), .ZN(n3907) );
  NAND2_X4 U3850 ( .A1(n3738), .A2(n3828), .ZN(n3900) );
  NAND4_X4 U3851 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3860)
         );
  NOR2_X2 U3852 ( .A1(n6278), .A2(n3726), .ZN(n6168) );
  NAND2_X2 U3853 ( .A1(n6446), .A2(n4178), .ZN(n6442) );
  NAND2_X1 U3854 ( .A1(n4154), .A2(n4165), .ZN(n4172) );
  INV_X2 U3855 ( .A(n6443), .ZN(n6483) );
  NAND2_X1 U3856 ( .A1(n3904), .A2(n3819), .ZN(n3902) );
  NAND2_X1 U3857 ( .A1(n4262), .A2(n3919), .ZN(n3819) );
  AND2_X1 U3858 ( .A1(n4117), .A2(n4116), .ZN(n4119) );
  NAND2_X1 U3859 ( .A1(n3710), .A2(n3709), .ZN(n4118) );
  INV_X1 U3860 ( .A(n4058), .ZN(n4059) );
  NAND2_X1 U3861 ( .A1(n3730), .A2(n4559), .ZN(n3729) );
  INV_X1 U3862 ( .A(n6273), .ZN(n3730) );
  INV_X1 U3863 ( .A(n6477), .ZN(n3695) );
  INV_X1 U3864 ( .A(n3700), .ZN(n3692) );
  INV_X1 U3865 ( .A(n4146), .ZN(n4144) );
  OR2_X1 U3866 ( .A1(n3904), .A2(n3908), .ZN(n4260) );
  NAND2_X1 U3867 ( .A1(n6215), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5744) );
  NOR2_X1 U3868 ( .A1(n3718), .A2(n3716), .ZN(n3715) );
  INV_X1 U3869 ( .A(n6348), .ZN(n3716) );
  NAND2_X1 U3870 ( .A1(n6215), .A2(n4776), .ZN(n7467) );
  NAND2_X1 U3871 ( .A1(n3949), .A2(n3948), .ZN(n3993) );
  NOR3_X1 U3872 ( .A1(n3947), .A2(n3946), .A3(n3945), .ZN(n3948) );
  INV_X1 U3873 ( .A(n3935), .ZN(n3947) );
  NAND2_X1 U3874 ( .A1(n4121), .A2(n4120), .ZN(n4146) );
  INV_X1 U3875 ( .A(n4119), .ZN(n4120) );
  AND2_X1 U3876 ( .A1(n4142), .A2(n4141), .ZN(n4145) );
  AND2_X1 U3877 ( .A1(n3860), .A2(n5073), .ZN(n3996) );
  NAND2_X1 U3878 ( .A1(n3905), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U3879 ( .A1(n4696), .A2(n3734), .ZN(n3733) );
  INV_X1 U3880 ( .A(n6128), .ZN(n4696) );
  INV_X1 U3881 ( .A(n6143), .ZN(n3734) );
  NAND2_X1 U3882 ( .A1(n3725), .A2(n3735), .ZN(n3724) );
  INV_X1 U3883 ( .A(n6293), .ZN(n3725) );
  NAND2_X1 U3884 ( .A1(n4438), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4747) );
  NOR2_X1 U3885 ( .A1(n3649), .A2(n3713), .ZN(n3712) );
  INV_X1 U3886 ( .A(n5975), .ZN(n3713) );
  INV_X1 U3887 ( .A(n4286), .ZN(n4743) );
  NOR2_X1 U3888 ( .A1(n3689), .A2(n6288), .ZN(n3687) );
  INV_X1 U3889 ( .A(n6281), .ZN(n3689) );
  NOR2_X1 U3890 ( .A1(n4789), .A2(n4975), .ZN(n4870) );
  NAND2_X1 U3891 ( .A1(n3740), .A2(n3684), .ZN(n3683) );
  INV_X1 U3892 ( .A(n5995), .ZN(n3684) );
  INV_X1 U3893 ( .A(n4870), .ZN(n4860) );
  AND2_X1 U3894 ( .A1(n4999), .A2(n4998), .ZN(n5007) );
  NAND2_X1 U3895 ( .A1(n3920), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4036) );
  OR2_X1 U3896 ( .A1(n3984), .A2(n3983), .ZN(n4009) );
  OR2_X1 U3897 ( .A1(n4046), .A2(n4045), .ZN(n4078) );
  AND2_X1 U3898 ( .A1(n5048), .A2(n4060), .ZN(n5830) );
  INV_X1 U3899 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6706) );
  AND2_X2 U3900 ( .A1(n3802), .A2(n3801), .ZN(n3919) );
  NAND2_X1 U3901 ( .A1(n4036), .A2(n4035), .ZN(n4253) );
  AND2_X1 U3902 ( .A1(n5266), .A2(n5265), .ZN(n6969) );
  AND2_X2 U3903 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5279) );
  AND2_X1 U3904 ( .A1(n5276), .A2(n5275), .ZN(n6957) );
  INV_X1 U3905 ( .A(n5744), .ZN(n5733) );
  NAND2_X1 U3906 ( .A1(n6069), .A2(n6058), .ZN(n4872) );
  INV_X1 U3907 ( .A(n4780), .ZN(n4969) );
  NAND2_X1 U3908 ( .A1(n4906), .A2(n4905), .ZN(n5228) );
  OR3_X1 U3909 ( .A1(n4904), .A2(READY_N), .A3(n6110), .ZN(n4905) );
  NOR2_X1 U3910 ( .A1(n5195), .A2(READY_N), .ZN(n5199) );
  NAND2_X1 U3911 ( .A1(n6180), .A2(n3727), .ZN(n3726) );
  INV_X1 U3912 ( .A(n3729), .ZN(n3727) );
  CLKBUF_X1 U3913 ( .A(n6227), .Z(n6228) );
  NOR2_X1 U3914 ( .A1(n3720), .A2(n3719), .ZN(n3718) );
  INV_X1 U3915 ( .A(n4403), .ZN(n3719) );
  INV_X1 U3916 ( .A(n6352), .ZN(n3720) );
  NAND2_X1 U3917 ( .A1(n6016), .A2(n3665), .ZN(n3717) );
  AND2_X1 U3918 ( .A1(n6115), .A2(n7522), .ZN(n5197) );
  OAI21_X2 U3919 ( .B1(n6442), .B2(n4181), .A(n4180), .ZN(n6617) );
  NAND2_X1 U3920 ( .A1(n4838), .A2(n3676), .ZN(n3675) );
  INV_X1 U3921 ( .A(n6231), .ZN(n3676) );
  NOR2_X1 U3922 ( .A1(n6443), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3702)
         );
  INV_X1 U3923 ( .A(n6485), .ZN(n3701) );
  INV_X1 U3924 ( .A(n6482), .ZN(n3697) );
  NOR2_X1 U3925 ( .A1(n3618), .A2(n3699), .ZN(n3698) );
  NAND2_X1 U3926 ( .A1(n6485), .A2(n3666), .ZN(n3699) );
  AND2_X1 U3927 ( .A1(n5037), .A2(n5036), .ZN(n7256) );
  INV_X1 U3928 ( .A(n5007), .ZN(n5014) );
  NAND2_X1 U3929 ( .A1(n5286), .A2(n4034), .ZN(n4925) );
  XNOR2_X1 U3930 ( .A(n5286), .B(n5284), .ZN(n5045) );
  INV_X1 U3931 ( .A(n6679), .ZN(n5748) );
  AND2_X1 U3932 ( .A1(n6667), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U3933 ( .A1(n4907), .A2(n3992), .ZN(n6988) );
  AND2_X1 U3934 ( .A1(n6125), .A2(REIP_REG_30__SCAN_IN), .ZN(n3679) );
  AND2_X1 U3935 ( .A1(n4882), .A2(n4876), .ZN(n7412) );
  XNOR2_X1 U3936 ( .A(n3680), .B(n6058), .ZN(n6527) );
  INV_X1 U3937 ( .A(n6057), .ZN(n3680) );
  NOR2_X1 U3938 ( .A1(n4759), .A2(n6120), .ZN(n4760) );
  XNOR2_X1 U3939 ( .A(n4753), .B(n4752), .ZN(n6062) );
  NOR2_X1 U3940 ( .A1(n6140), .A2(n3663), .ZN(n4753) );
  INV_X1 U3941 ( .A(n6053), .ZN(n6054) );
  XNOR2_X1 U3942 ( .A(n4201), .B(n6512), .ZN(n6522) );
  OR2_X1 U3943 ( .A1(n6101), .A2(n6100), .ZN(n6103) );
  INV_X1 U3944 ( .A(n7301), .ZN(n7313) );
  INV_X1 U3945 ( .A(n7521), .ZN(n7512) );
  OAI21_X1 U3946 ( .B1(n3996), .B2(n3908), .A(n3924), .ZN(n3890) );
  INV_X1 U3947 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3749) );
  AND2_X1 U3948 ( .A1(n4253), .A2(n4767), .ZN(n4241) );
  OR2_X1 U3949 ( .A1(n4220), .A2(n3925), .ZN(n4242) );
  OR2_X1 U3950 ( .A1(n4115), .A2(n4114), .ZN(n4148) );
  OR2_X1 U3951 ( .A1(n4036), .A2(n3994), .ZN(n3950) );
  AOI22_X1 U3952 ( .A1(n4065), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3793) );
  NAND2_X1 U3953 ( .A1(n4208), .A2(n4207), .ZN(n4212) );
  NAND2_X1 U3954 ( .A1(n7520), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U3955 ( .A1(n3673), .A2(EBX_REG_1__SCAN_IN), .ZN(n3672) );
  AND2_X1 U3956 ( .A1(n6407), .A2(n4286), .ZN(n4606) );
  NAND2_X1 U3957 ( .A1(n4436), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4452)
         );
  NOR2_X1 U3958 ( .A1(n4361), .A2(n6254), .ZN(n4385) );
  INV_X1 U3959 ( .A(n6001), .ZN(n4374) );
  AND2_X1 U3960 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4295), .ZN(n4304)
         );
  INV_X1 U3961 ( .A(n4296), .ZN(n4295) );
  NAND2_X1 U3962 ( .A1(n3687), .A2(n6275), .ZN(n3686) );
  OR2_X1 U3963 ( .A1(n4075), .A2(n4074), .ZN(n4082) );
  NAND2_X1 U3964 ( .A1(n4984), .A2(n3920), .ZN(n5003) );
  NAND2_X1 U3965 ( .A1(n4006), .A2(n3991), .ZN(n4017) );
  OR2_X1 U3966 ( .A1(n4036), .A2(n3990), .ZN(n3991) );
  AND2_X1 U3967 ( .A1(n4902), .A2(n4911), .ZN(n5010) );
  OR2_X1 U3968 ( .A1(n6090), .A2(n6665), .ZN(n5829) );
  AND2_X1 U3969 ( .A1(n4059), .A2(n4026), .ZN(n5151) );
  AND2_X1 U3970 ( .A1(n7592), .A2(n5824), .ZN(n6707) );
  NAND2_X1 U3971 ( .A1(n3846), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3811)
         );
  OAI21_X1 U3972 ( .B1(n5044), .B2(n7526), .A(n7505), .ZN(n5055) );
  AND2_X1 U3973 ( .A1(n4025), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4058)
         );
  AND2_X1 U3974 ( .A1(n4210), .A2(n4211), .ZN(n4254) );
  OR2_X1 U3975 ( .A1(n4212), .A2(n4209), .ZN(n4210) );
  AND2_X1 U3976 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n7016), .ZN(n4209)
         );
  INV_X1 U3977 ( .A(n4254), .ZN(n4771) );
  OR2_X1 U3978 ( .A1(n4212), .A2(n4211), .ZN(n4251) );
  AND2_X1 U3979 ( .A1(n4985), .A2(n4918), .ZN(n6111) );
  INV_X1 U3980 ( .A(n4534), .ZN(n4535) );
  NAND2_X1 U3981 ( .A1(n3674), .A2(n3670), .ZN(n3669) );
  OR2_X1 U3982 ( .A1(n4977), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3674)
         );
  INV_X1 U3983 ( .A(n3671), .ZN(n3670) );
  OAI21_X1 U3984 ( .B1(n4865), .B2(EBX_REG_1__SCAN_IN), .A(n3672), .ZN(n3671)
         );
  OR2_X1 U3985 ( .A1(n7492), .A2(n4743), .ZN(n4591) );
  AND2_X1 U3986 ( .A1(n4796), .A2(n4795), .ZN(n5778) );
  AND2_X1 U3987 ( .A1(n5197), .A2(n4949), .ZN(n7019) );
  OR2_X1 U3988 ( .A1(n4698), .A2(n6073), .ZN(n4759) );
  NAND2_X1 U3989 ( .A1(n6068), .A2(n3732), .ZN(n3731) );
  INV_X1 U3990 ( .A(n3733), .ZN(n3732) );
  AND2_X1 U3991 ( .A1(n4671), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4672)
         );
  OR2_X1 U3992 ( .A1(n4676), .A2(n4675), .ZN(n6143) );
  NOR2_X1 U3993 ( .A1(n4586), .A2(n7479), .ZN(n4587) );
  INV_X1 U3994 ( .A(n6278), .ZN(n3728) );
  NAND2_X1 U3995 ( .A1(n3722), .A2(n6197), .ZN(n3721) );
  INV_X1 U3996 ( .A(n3724), .ZN(n3722) );
  NOR2_X1 U3997 ( .A1(n4486), .A2(n6220), .ZN(n4487) );
  NAND2_X1 U3998 ( .A1(n4487), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4534)
         );
  NOR2_X1 U3999 ( .A1(n4452), .A2(n6234), .ZN(n4453) );
  AND2_X1 U4000 ( .A1(n4414), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4419)
         );
  NOR2_X1 U4001 ( .A1(n4401), .A2(n4386), .ZN(n4414) );
  OR2_X1 U4002 ( .A1(n4399), .A2(n4398), .ZN(n4400) );
  NAND2_X1 U4003 ( .A1(n4385), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4401)
         );
  CLKBUF_X1 U4004 ( .A(n5999), .Z(n6000) );
  NAND2_X1 U4005 ( .A1(n4357), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4361)
         );
  INV_X1 U4006 ( .A(n5960), .ZN(n4333) );
  INV_X1 U4007 ( .A(n4315), .ZN(n4316) );
  AND2_X1 U4008 ( .A1(n4304), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4312)
         );
  AOI21_X1 U4009 ( .B1(n4311), .B2(n4429), .A(n4310), .ZN(n5784) );
  AOI21_X1 U4010 ( .B1(n4301), .B2(n4429), .A(n4300), .ZN(n5030) );
  CLKBUF_X1 U4011 ( .A(n5027), .Z(n5028) );
  NAND2_X1 U4012 ( .A1(n4285), .A2(n4429), .ZN(n4294) );
  AND3_X1 U4013 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4287) );
  AOI21_X1 U4014 ( .B1(n5242), .B2(n4429), .A(n4283), .ZN(n5023) );
  CLKBUF_X1 U4015 ( .A(n5021), .Z(n5022) );
  AND2_X1 U4016 ( .A1(n6365), .A2(n4197), .ZN(n6357) );
  NAND2_X1 U4017 ( .A1(n6384), .A2(n3703), .ZN(n6366) );
  NOR2_X1 U4018 ( .A1(n3651), .A2(n3704), .ZN(n3703) );
  INV_X1 U4019 ( .A(n4195), .ZN(n3704) );
  AND2_X1 U4020 ( .A1(n4857), .A2(n4856), .ZN(n6172) );
  XNOR2_X1 U4021 ( .A(n3618), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6393)
         );
  NAND2_X1 U4022 ( .A1(n6443), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6401) );
  AND2_X1 U4023 ( .A1(n4851), .A2(n4850), .ZN(n6281) );
  NOR2_X1 U4024 ( .A1(n6287), .A2(n3685), .ZN(n6283) );
  INV_X1 U4025 ( .A(n3687), .ZN(n3685) );
  AND2_X1 U4026 ( .A1(n4849), .A2(n4848), .ZN(n6288) );
  NOR2_X1 U4027 ( .A1(n6287), .A2(n6288), .ZN(n6286) );
  AND3_X1 U4028 ( .A1(n4835), .A2(n4840), .A3(n4834), .ZN(n6302) );
  AOI21_X1 U4029 ( .B1(n3694), .B2(n3692), .A(n3647), .ZN(n3691) );
  AND2_X1 U4030 ( .A1(n4814), .A2(n4813), .ZN(n6003) );
  INV_X1 U4031 ( .A(n5948), .ZN(n3681) );
  AND2_X1 U4032 ( .A1(n7256), .A2(n7252), .ZN(n6628) );
  NOR2_X1 U4033 ( .A1(n5782), .A2(n3683), .ZN(n5993) );
  NAND2_X1 U4034 ( .A1(n3682), .A2(n3740), .ZN(n5994) );
  AOI21_X1 U4035 ( .B1(n7167), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3707), 
        .ZN(n3706) );
  NOR2_X1 U4036 ( .A1(n7167), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3705)
         );
  INV_X1 U4037 ( .A(n4130), .ZN(n3707) );
  XNOR2_X1 U4038 ( .A(n4161), .B(n5990), .ZN(n5953) );
  OR2_X1 U4039 ( .A1(n5038), .A2(n7256), .ZN(n6509) );
  OR2_X1 U4040 ( .A1(n5057), .A2(n4007), .ZN(n4013) );
  NAND2_X1 U4041 ( .A1(n5015), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5136)
         );
  INV_X1 U4042 ( .A(n4047), .ZN(n4048) );
  NAND3_X1 U4043 ( .A1(n3905), .A2(n4986), .A3(n5069), .ZN(n3906) );
  INV_X1 U4044 ( .A(n4033), .ZN(n4030) );
  NAND2_X1 U4045 ( .A1(n4064), .A2(n4063), .ZN(n5284) );
  NOR2_X1 U4046 ( .A1(n5242), .A2(n5098), .ZN(n5105) );
  OAI21_X1 U4047 ( .B1(n5750), .B2(n6853), .A(n5749), .ZN(n5791) );
  OR2_X1 U4048 ( .A1(n6703), .A2(n7587), .ZN(n6797) );
  AND2_X1 U4049 ( .A1(n5146), .A2(n5206), .ZN(n5670) );
  INV_X1 U4050 ( .A(n5670), .ZN(n5678) );
  NAND3_X1 U4051 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4049), .A3(n5055), .ZN(
        n6678) );
  NAND2_X1 U4052 ( .A1(n4049), .A2(n5055), .ZN(n6679) );
  AOI21_X1 U4053 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6784), .A(n6679), .ZN(
        n7602) );
  INV_X1 U4054 ( .A(n7599), .ZN(n7587) );
  NOR2_X1 U4055 ( .A1(n4255), .A2(n4771), .ZN(n4256) );
  AOI21_X1 U4056 ( .B1(n4253), .B2(n4254), .A(n4252), .ZN(n4257) );
  OAI21_X1 U4057 ( .B1(n4255), .B2(n4251), .A(n4250), .ZN(n4252) );
  AND2_X1 U4058 ( .A1(n5281), .A2(n5280), .ZN(n6984) );
  OR2_X1 U4059 ( .A1(n4892), .A2(n6986), .ZN(n4896) );
  AND2_X1 U4060 ( .A1(n7599), .A2(n6667), .ZN(n6009) );
  NAND2_X1 U4061 ( .A1(n5733), .A2(n4878), .ZN(n7473) );
  AND2_X1 U4062 ( .A1(n6215), .A2(n5735), .ZN(n7483) );
  INV_X1 U4063 ( .A(n7467), .ZN(n7496) );
  AND2_X1 U4064 ( .A1(n6215), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7490) );
  INV_X1 U4065 ( .A(n7473), .ZN(n7333) );
  INV_X1 U4066 ( .A(n7490), .ZN(n7478) );
  INV_X1 U4067 ( .A(n3969), .ZN(n3972) );
  OR2_X1 U4068 ( .A1(n6069), .A2(n3673), .ZN(n4873) );
  INV_X1 U4069 ( .A(n6304), .ZN(n7139) );
  AND2_X2 U4070 ( .A1(n4973), .A2(n7522), .ZN(n7143) );
  NAND2_X1 U4071 ( .A1(n7143), .A2(n6060), .ZN(n6304) );
  INV_X1 U4072 ( .A(n7567), .ZN(n7582) );
  AND2_X1 U4073 ( .A1(n7564), .A2(n6063), .ZN(n7578) );
  AND2_X1 U4074 ( .A1(n7564), .A2(n5231), .ZN(n7579) );
  NAND2_X1 U4075 ( .A1(n5935), .A2(n5229), .ZN(n7564) );
  INV_X1 U4076 ( .A(n7184), .ZN(n7563) );
  INV_X1 U4077 ( .A(n3718), .ZN(n3714) );
  XNOR2_X1 U4078 ( .A(n6378), .B(n6554), .ZN(n6559) );
  NAND2_X1 U4079 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  NAND2_X1 U4080 ( .A1(n6374), .A2(n6444), .ZN(n6376) );
  NAND2_X1 U4081 ( .A1(n6375), .A2(n6443), .ZN(n6377) );
  AND2_X1 U4082 ( .A1(n6585), .A2(n4187), .ZN(n6571) );
  AND2_X1 U4083 ( .A1(n6603), .A2(n6514), .ZN(n6585) );
  INV_X1 U4084 ( .A(n3698), .ZN(n3693) );
  NAND2_X1 U4085 ( .A1(n3697), .A2(n3700), .ZN(n3696) );
  INV_X1 U4086 ( .A(n7310), .ZN(n7275) );
  NAND2_X1 U4087 ( .A1(n7162), .A2(n4130), .ZN(n7169) );
  INV_X1 U4088 ( .A(n7252), .ZN(n7298) );
  INV_X1 U4089 ( .A(n6509), .ZN(n7260) );
  NAND2_X1 U4090 ( .A1(n5014), .A2(n5001), .ZN(n7301) );
  INV_X1 U4091 ( .A(n7280), .ZN(n7248) );
  INV_X1 U4092 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6784) );
  CLKBUF_X1 U4093 ( .A(n5046), .Z(n5047) );
  CLKBUF_X1 U4094 ( .A(n4925), .Z(n6090) );
  INV_X1 U4095 ( .A(n7015), .ZN(n6082) );
  AND2_X1 U4096 ( .A1(n4772), .A2(n5196), .ZN(n6958) );
  INV_X1 U4097 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6667) );
  INV_X1 U4098 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7520) );
  CLKBUF_X1 U4099 ( .A(n4903), .Z(n4904) );
  OR2_X1 U4100 ( .A1(n7518), .A2(n4924), .ZN(n7521) );
  INV_X1 U4101 ( .A(n6952), .ZN(n6684) );
  INV_X1 U4102 ( .A(n6839), .ZN(n7649) );
  OR2_X1 U4103 ( .A1(n6786), .A2(n5057), .ZN(n6839) );
  NOR2_X2 U4104 ( .A1(n5182), .A2(n5057), .ZN(n6895) );
  INV_X1 U4105 ( .A(n6929), .ZN(n6917) );
  AND2_X1 U4106 ( .A1(n7185), .A2(DATAI_16_), .ZN(n7606) );
  AND2_X1 U4107 ( .A1(n7185), .A2(DATAI_17_), .ZN(n7611) );
  AND2_X1 U4108 ( .A1(n7185), .A2(DATAI_18_), .ZN(n7617) );
  AND2_X1 U4109 ( .A1(n7185), .A2(DATAI_19_), .ZN(n7624) );
  AND2_X1 U4110 ( .A1(n7185), .A2(DATAI_20_), .ZN(n7629) );
  AND2_X1 U4111 ( .A1(n7185), .A2(DATAI_21_), .ZN(n7635) );
  AND2_X1 U4112 ( .A1(n7185), .A2(DATAI_22_), .ZN(n7641) );
  NOR2_X1 U4113 ( .A1(n5058), .A2(n5057), .ZN(n6952) );
  AND2_X1 U4114 ( .A1(n5059), .A2(n5057), .ZN(n6951) );
  AND2_X1 U4115 ( .A1(n7185), .A2(DATAI_23_), .ZN(n7648) );
  NOR2_X1 U4116 ( .A1(n7200), .A2(n6667), .ZN(n7526) );
  AND2_X1 U4117 ( .A1(n4258), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7522) );
  INV_X1 U4118 ( .A(READY_N), .ZN(n7546) );
  INV_X1 U4119 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U4120 ( .A1(n7547), .A2(STATE_REG_1__SCAN_IN), .ZN(n7553) );
  OAI21_X1 U4121 ( .B1(n6527), .B2(n7493), .A(n3677), .ZN(U2797) );
  INV_X1 U4122 ( .A(n3678), .ZN(n3677) );
  OAI21_X1 U4123 ( .B1(n6522), .B2(n7501), .A(n4763), .ZN(U2955) );
  AOI21_X1 U4124 ( .B1(n6319), .B2(n7185), .A(n6107), .ZN(n6108) );
  NAND2_X1 U4125 ( .A1(n3723), .A2(n3735), .ZN(n6211) );
  OR2_X1 U4126 ( .A1(n4935), .A2(n3908), .ZN(n3646) );
  NAND2_X1 U4127 ( .A1(n3728), .A2(n4559), .ZN(n6272) );
  AND2_X1 U4128 ( .A1(n6483), .A2(n4821), .ZN(n3647) );
  OR3_X1 U4129 ( .A1(n6313), .A2(n6302), .A3(n6231), .ZN(n3648) );
  NAND2_X1 U4130 ( .A1(n4333), .A2(n5947), .ZN(n3649) );
  OR2_X1 U4131 ( .A1(n6287), .A2(n3686), .ZN(n3650) );
  AND2_X1 U4132 ( .A1(n6483), .A2(n6554), .ZN(n3651) );
  AND4_X1 U4133 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3652)
         );
  XOR2_X1 U4134 ( .A(n6359), .B(n6358), .Z(n3653) );
  NOR2_X1 U4135 ( .A1(n6210), .A2(n3724), .ZN(n6196) );
  NOR2_X1 U4136 ( .A1(n6210), .A2(n3721), .ZN(n6195) );
  NOR2_X1 U4137 ( .A1(n6278), .A2(n3729), .ZN(n6181) );
  NAND2_X1 U4138 ( .A1(n6444), .A2(n4177), .ZN(n3654) );
  NAND2_X1 U4139 ( .A1(n4144), .A2(n4143), .ZN(n4154) );
  NAND2_X1 U4140 ( .A1(n4194), .A2(n4193), .ZN(n6384) );
  AND2_X1 U4141 ( .A1(n4098), .A2(n4097), .ZN(n3655) );
  AND2_X1 U4142 ( .A1(n3654), .A2(n4176), .ZN(n3656) );
  OAI21_X1 U4143 ( .B1(n4284), .B2(n4007), .A(n4100), .ZN(n4103) );
  NOR2_X1 U4144 ( .A1(n6124), .A2(n3679), .ZN(n3657) );
  OR2_X1 U4145 ( .A1(n3683), .A2(n3681), .ZN(n3658) );
  NAND2_X1 U4146 ( .A1(n6461), .A2(n4176), .ZN(n6454) );
  NOR2_X1 U4147 ( .A1(n3698), .A2(n3695), .ZN(n3694) );
  NAND2_X2 U4148 ( .A1(n4006), .A2(n4005), .ZN(n5057) );
  OR2_X1 U4149 ( .A1(n3900), .A2(n5906), .ZN(n3659) );
  AND2_X2 U4150 ( .A1(n7501), .A2(n4756), .ZN(n7183) );
  NOR2_X1 U4151 ( .A1(n5699), .A2(n3649), .ZN(n5945) );
  XNOR2_X1 U4152 ( .A(n6016), .B(n4403), .ZN(n6351) );
  AND2_X1 U4153 ( .A1(n3717), .A2(n3714), .ZN(n3660) );
  AND2_X1 U4154 ( .A1(n3696), .A2(n3693), .ZN(n6476) );
  NOR3_X1 U4155 ( .A1(n6287), .A2(n3686), .A3(n6185), .ZN(n3688) );
  AND2_X1 U4156 ( .A1(n3900), .A2(n4262), .ZN(n3661) );
  INV_X1 U4157 ( .A(n6210), .ZN(n3723) );
  AND2_X1 U4158 ( .A1(n3711), .A2(n4333), .ZN(n3662) );
  OR2_X1 U4159 ( .A1(n3731), .A2(n6053), .ZN(n3663) );
  NAND2_X1 U4160 ( .A1(n4262), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4418) );
  INV_X1 U4161 ( .A(n4418), .ZN(n4429) );
  NOR2_X1 U4162 ( .A1(n6313), .A2(n6231), .ZN(n3664) );
  OR2_X1 U4163 ( .A1(n6352), .A2(n4403), .ZN(n3665) );
  NAND2_X1 U4164 ( .A1(n4266), .A2(n4265), .ZN(n4964) );
  NAND2_X1 U4165 ( .A1(n5197), .A2(n6975), .ZN(n7501) );
  INV_X1 U4166 ( .A(n7501), .ZN(n7186) );
  INV_X1 U4167 ( .A(n7185), .ZN(n7174) );
  AND2_X2 U4168 ( .A1(n7599), .A2(n4754), .ZN(n7185) );
  XNOR2_X1 U4169 ( .A(n3669), .B(n4978), .ZN(n4974) );
  INV_X1 U4170 ( .A(n4789), .ZN(n3673) );
  INV_X1 U4171 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6254) );
  INV_X1 U4172 ( .A(n5782), .ZN(n3682) );
  NAND3_X1 U4173 ( .A1(n6486), .A2(n6046), .A3(n6484), .ZN(n3666) );
  INV_X1 U4174 ( .A(n3617), .ZN(n7476) );
  AND2_X4 U4175 ( .A1(n5282), .A2(n3667), .ZN(n4518) );
  AND2_X2 U4176 ( .A1(n3757), .A2(n3667), .ZN(n3845) );
  INV_X1 U4177 ( .A(n4978), .ZN(n3668) );
  OAI21_X2 U4178 ( .B1(n6126), .B2(n7467), .A(n3657), .ZN(n3678) );
  INV_X1 U4179 ( .A(n3688), .ZN(n6184) );
  NAND2_X1 U4180 ( .A1(n3690), .A2(n3691), .ZN(n6469) );
  NAND2_X1 U4181 ( .A1(n5952), .A2(n5953), .ZN(n4163) );
  NAND2_X1 U4182 ( .A1(n4118), .A2(n3708), .ZN(n4284) );
  OAI21_X1 U4183 ( .B1(n4086), .B2(n5051), .A(n3655), .ZN(n3708) );
  INV_X1 U4184 ( .A(n4086), .ZN(n3710) );
  INV_X1 U4185 ( .A(n5699), .ZN(n3711) );
  NAND2_X1 U4186 ( .A1(n3711), .A2(n3712), .ZN(n5973) );
  NAND2_X1 U4187 ( .A1(n3717), .A2(n3715), .ZN(n6308) );
  INV_X1 U4188 ( .A(n6308), .ZN(n4435) );
  NOR2_X1 U4189 ( .A1(n6140), .A2(n3733), .ZN(n6066) );
  NOR2_X1 U4190 ( .A1(n6140), .A2(n6143), .ZN(n6127) );
  OR2_X2 U4191 ( .A1(n6140), .A2(n3731), .ZN(n6067) );
  INV_X1 U4192 ( .A(n4118), .ZN(n4121) );
  NAND2_X1 U4193 ( .A1(n4964), .A2(n4966), .ZN(n4965) );
  NAND2_X1 U4194 ( .A1(n4420), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3776) );
  AND2_X1 U4195 ( .A1(n4485), .A2(n4484), .ZN(n3735) );
  INV_X1 U4196 ( .A(n3937), .ZN(n7507) );
  AND2_X1 U4197 ( .A1(n4056), .A2(n5004), .ZN(n3736) );
  OR2_X1 U4198 ( .A1(n3739), .A2(n4867), .ZN(n3737) );
  AND4_X1 U4199 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3738)
         );
  AND2_X1 U4200 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3739) );
  NAND3_X1 U4201 ( .A1(n4800), .A2(n4840), .A3(n4799), .ZN(n3740) );
  INV_X1 U4202 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6220) );
  OR2_X1 U4203 ( .A1(n7200), .A2(n4950), .ZN(n6985) );
  INV_X1 U4204 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7016) );
  AND2_X1 U4205 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5753), .ZN(n3741) );
  OR2_X1 U4206 ( .A1(n3914), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3742)
         );
  NAND2_X1 U4207 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  OR2_X1 U4208 ( .A1(n4096), .A2(n4095), .ZN(n4123) );
  INV_X1 U4209 ( .A(n3993), .ZN(n3994) );
  AND2_X1 U4210 ( .A1(n4205), .A2(n4204), .ZN(n4217) );
  INV_X1 U4211 ( .A(n4145), .ZN(n4143) );
  INV_X1 U4212 ( .A(n4166), .ZN(n3990) );
  AND2_X1 U4213 ( .A1(n3899), .A2(n3898), .ZN(n3913) );
  AND2_X1 U4214 ( .A1(n6784), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4231)
         );
  INV_X1 U4215 ( .A(n6280), .ZN(n4559) );
  INV_X1 U4216 ( .A(n6156), .ZN(n4652) );
  OAI21_X1 U4217 ( .B1(n3659), .B2(n4314), .A(n4313), .ZN(n4315) );
  OR2_X1 U4218 ( .A1(n4140), .A2(n4139), .ZN(n4156) );
  OAI21_X1 U4219 ( .B1(n3637), .B2(n5000), .A(n3900), .ZN(n4929) );
  NAND2_X1 U4220 ( .A1(n5045), .A2(n4049), .ZN(n4077) );
  OR2_X1 U4221 ( .A1(n4697), .A2(n6132), .ZN(n4698) );
  OR2_X1 U4222 ( .A1(n4619), .A2(n4618), .ZN(n4644) );
  INV_X1 U4223 ( .A(n5030), .ZN(n4302) );
  INV_X1 U4224 ( .A(n4747), .ZN(n4690) );
  INV_X1 U4225 ( .A(n4437), .ZN(n4438) );
  NOR2_X1 U4226 ( .A1(n5003), .A2(n4164), .ZN(n4165) );
  NAND2_X1 U4227 ( .A1(n3972), .A2(n3971), .ZN(n3973) );
  NAND2_X1 U4228 ( .A1(n4077), .A2(n4076), .ZN(n4085) );
  AND4_X1 U4229 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3856)
         );
  INV_X1 U4230 ( .A(n4085), .ZN(n5051) );
  NAND2_X1 U4231 ( .A1(n3951), .A2(n4984), .ZN(n4255) );
  AND2_X1 U4232 ( .A1(n4626), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4627)
         );
  NAND2_X1 U4233 ( .A1(n4672), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4697)
         );
  NAND2_X1 U4234 ( .A1(n4587), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4625)
         );
  INV_X1 U4235 ( .A(n4605), .ZN(n4751) );
  NAND2_X1 U4236 ( .A1(n6443), .A2(n4867), .ZN(n6100) );
  NAND2_X1 U4237 ( .A1(n4029), .A2(n4028), .ZN(n4031) );
  INV_X1 U4238 ( .A(n6783), .ZN(n6769) );
  INV_X1 U4239 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U4240 ( .A1(n4627), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4670)
         );
  AND2_X1 U4241 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4535), .ZN(n4536)
         );
  INV_X1 U4242 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6234) );
  OR3_X1 U4243 ( .A1(n7280), .A2(n7524), .A3(n6993), .ZN(n4775) );
  AND2_X1 U4244 ( .A1(n4759), .A2(n4699), .ZN(n6072) );
  INV_X1 U4245 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7479) );
  AND2_X1 U4246 ( .A1(n4517), .A2(n4516), .ZN(n6197) );
  AND2_X1 U4247 ( .A1(n4419), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4436)
         );
  NOR2_X1 U4248 ( .A1(n4334), .A2(n4329), .ZN(n4357) );
  AND2_X1 U4249 ( .A1(n4332), .A2(n4331), .ZN(n5960) );
  NAND2_X1 U4250 ( .A1(n6101), .A2(n6483), .ZN(n6102) );
  NAND2_X1 U4251 ( .A1(n5014), .A2(n6111), .ZN(n7252) );
  INV_X1 U4252 ( .A(n5047), .ZN(n6665) );
  NAND2_X1 U4253 ( .A1(n5105), .A2(n5057), .ZN(n6697) );
  INV_X1 U4254 ( .A(n6710), .ZN(n6750) );
  NAND2_X1 U4255 ( .A1(n5672), .A2(n5243), .ZN(n5251) );
  INV_X1 U4256 ( .A(n5052), .ZN(n5206) );
  AND2_X1 U4257 ( .A1(n7594), .A2(n7593), .ZN(n7600) );
  NOR2_X2 U4258 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7599) );
  NAND2_X1 U4259 ( .A1(n5909), .A2(n5206), .ZN(n5182) );
  NAND2_X1 U4260 ( .A1(n5909), .A2(n5908), .ZN(n6905) );
  INV_X1 U4261 ( .A(n5829), .ZN(n5679) );
  OR2_X1 U4262 ( .A1(n6090), .A2(n5047), .ZN(n7590) );
  INV_X1 U4263 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5906) );
  INV_X1 U4264 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7200) );
  INV_X1 U4265 ( .A(n4764), .ZN(n4765) );
  NAND2_X1 U4266 ( .A1(n5195), .A2(n4896), .ZN(n7205) );
  OAI21_X1 U4267 ( .B1(n6496), .B2(n7493), .A(n4888), .ZN(n4889) );
  NAND2_X1 U4268 ( .A1(n4536), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4586)
         );
  NOR3_X1 U4269 ( .A1(n7473), .A2(n7064), .A3(n6018), .ZN(n7410) );
  OR2_X1 U4270 ( .A1(n7205), .A2(n4775), .ZN(n6215) );
  NAND2_X1 U4271 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4334)
         );
  INV_X1 U4272 ( .A(n7423), .ZN(n7449) );
  INV_X1 U4273 ( .A(n7143), .ZN(n6314) );
  AND2_X1 U4274 ( .A1(n7564), .A2(n6060), .ZN(n6061) );
  INV_X1 U4275 ( .A(n7564), .ZN(n7581) );
  OAI21_X1 U4276 ( .B1(n5228), .B2(n5227), .A(n7522), .ZN(n5229) );
  NOR2_X1 U4277 ( .A1(n5198), .A2(n6988), .ZN(n5894) );
  NOR2_X1 U4278 ( .A1(n5199), .A2(n5933), .ZN(n5860) );
  INV_X1 U4279 ( .A(n5935), .ZN(n5893) );
  INV_X1 U4280 ( .A(n6417), .ZN(n7580) );
  NAND2_X1 U4281 ( .A1(n4453), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4486)
         );
  NAND2_X1 U4282 ( .A1(n4287), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4296)
         );
  NOR2_X1 U4283 ( .A1(n4260), .A2(n4259), .ZN(n6975) );
  NAND2_X1 U4284 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  INV_X1 U4285 ( .A(n6628), .ZN(n7226) );
  INV_X1 U4286 ( .A(n7240), .ZN(n7314) );
  AND2_X1 U4287 ( .A1(n5242), .A2(n5050), .ZN(n5909) );
  NOR2_X1 U4288 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7517) );
  INV_X1 U4289 ( .A(n6697), .ZN(n6686) );
  NOR2_X1 U4290 ( .A1(n5104), .A2(n5057), .ZN(n6710) );
  NOR2_X2 U4291 ( .A1(n5251), .A2(n6785), .ZN(n6760) );
  OR4_X1 U4292 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n6774) );
  INV_X1 U4293 ( .A(n5057), .ZN(n6785) );
  NOR2_X2 U4294 ( .A1(n5213), .A2(n5057), .ZN(n6827) );
  INV_X1 U4295 ( .A(n6852), .ZN(n6841) );
  AND2_X1 U4296 ( .A1(n5909), .A2(n5145), .ZN(n6919) );
  AND2_X1 U4297 ( .A1(n5670), .A2(n5057), .ZN(n6929) );
  INV_X1 U4298 ( .A(n6932), .ZN(n6939) );
  NAND2_X1 U4299 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6115), .ZN(n7505) );
  INV_X1 U4300 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U4301 ( .A1(n5197), .A2(n4765), .ZN(n5195) );
  INV_X1 U4302 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7535) );
  INV_X1 U4303 ( .A(n4889), .ZN(n4890) );
  INV_X1 U4304 ( .A(n7412), .ZN(n7493) );
  AND2_X1 U4305 ( .A1(n5731), .A2(n7467), .ZN(n7319) );
  NAND2_X1 U4306 ( .A1(n7564), .A2(n6318), .ZN(n7567) );
  INV_X1 U4307 ( .A(n7579), .ZN(n6354) );
  INV_X1 U4308 ( .A(n7019), .ZN(n7050) );
  NAND2_X1 U4309 ( .A1(n5199), .A2(n5196), .ZN(n5935) );
  AOI21_X1 U4310 ( .B1(n6612), .B2(n7298), .A(n7275), .ZN(n7307) );
  NAND2_X1 U4311 ( .A1(n5014), .A2(n5013), .ZN(n7240) );
  INV_X1 U4312 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6967) );
  INV_X1 U4313 ( .A(n5103), .ZN(n6701) );
  NAND2_X1 U4314 ( .A1(n5244), .A2(n6785), .ZN(n6772) );
  OR2_X1 U4315 ( .A1(n5213), .A2(n6785), .ZN(n6783) );
  INV_X1 U4316 ( .A(n6794), .ZN(n6831) );
  NAND2_X1 U4317 ( .A1(n5176), .A2(n5057), .ZN(n6852) );
  AOI22_X1 U4318 ( .A1(n6862), .A2(n6858), .B1(n6856), .B2(n6855), .ZN(n6897)
         );
  INV_X1 U4319 ( .A(n5907), .ZN(n6909) );
  OR2_X1 U4320 ( .A1(n5678), .A2(n5057), .ZN(n6932) );
  AND2_X1 U4321 ( .A1(n5711), .A2(n5710), .ZN(n6943) );
  AND2_X1 U4322 ( .A1(n7602), .A2(n5054), .ZN(n6956) );
  INV_X1 U4323 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7533) );
  OR2_X1 U4324 ( .A1(n7553), .A2(n6998), .ZN(n7095) );
  AND2_X2 U4325 ( .A1(n5279), .A2(n4939), .ZN(n3846) );
  NAND2_X1 U4326 ( .A1(n3846), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3748)
         );
  NAND2_X1 U4327 ( .A1(n4519), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3747) );
  INV_X1 U4328 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3744) );
  AND2_X2 U4329 ( .A1(n3744), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3751)
         );
  NAND2_X1 U4331 ( .A1(n4420), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3746) );
  NOR2_X4 U4332 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U4333 ( .A1(n3851), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3745) );
  NAND2_X1 U4334 ( .A1(n4065), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3756) );
  AND2_X2 U4335 ( .A1(n3763), .A2(n3751), .ZN(n3974) );
  NAND2_X1 U4336 ( .A1(n3974), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3755) );
  INV_X1 U4337 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3752) );
  NAND2_X1 U4338 ( .A1(n3866), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3754)
         );
  NAND2_X1 U4339 ( .A1(n3867), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4340 ( .A1(n4318), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3761)
         );
  AND2_X2 U4341 ( .A1(n3762), .A2(n5282), .ZN(n3861) );
  NAND2_X1 U4342 ( .A1(n3861), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4343 ( .A1(n3845), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4344 ( .A1(n4518), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3758) );
  AND2_X2 U4345 ( .A1(n3762), .A2(n4939), .ZN(n3942) );
  NAND2_X1 U4346 ( .A1(n3942), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3767)
         );
  NAND2_X1 U4347 ( .A1(n4109), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4348 ( .A1(n3876), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3765) );
  AND2_X4 U4349 ( .A1(n5282), .A2(n5279), .ZN(n4524) );
  NAND2_X1 U4350 ( .A1(n4524), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3764)
         );
  AND4_X1 U4351 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  XNOR2_X1 U4352 ( .A(n6998), .B(STATE_REG_1__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U4353 ( .A1(n5196), .A2(n4877), .ZN(n3909) );
  NAND2_X1 U4354 ( .A1(n3851), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4355 ( .A1(n3846), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3773)
         );
  NAND2_X1 U4356 ( .A1(n4519), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4357 ( .A1(n4065), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3780) );
  NAND2_X1 U4358 ( .A1(n3974), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4359 ( .A1(n3866), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3778)
         );
  NAND2_X1 U4360 ( .A1(n3867), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3777)
         );
  NAND2_X1 U4361 ( .A1(n3861), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4362 ( .A1(n4318), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3783)
         );
  NAND2_X1 U4363 ( .A1(n3845), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4364 ( .A1(n4518), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3781) );
  NAND2_X1 U4365 ( .A1(n3876), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4366 ( .A1(n4524), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3787)
         );
  NAND2_X1 U4367 ( .A1(n4109), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4368 ( .A1(n3942), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3785)
         );
  AOI22_X1 U4369 ( .A1(n3861), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4370 ( .A1(n4318), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3845), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4371 ( .A1(n3974), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4372 ( .A1(n4109), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4373 ( .A1(n4420), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3851), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4374 ( .A1(n3942), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4375 ( .A1(n3846), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4376 ( .A1(n3861), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3806) );
  NAND2_X1 U4377 ( .A1(n3974), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4378 ( .A1(n4065), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4379 ( .A1(n4109), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4380 ( .A1(n4518), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3810) );
  NAND2_X1 U4381 ( .A1(n4524), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3809)
         );
  NAND2_X1 U4382 ( .A1(n3866), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3808)
         );
  NAND2_X1 U4383 ( .A1(n4318), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3807)
         );
  NAND2_X1 U4384 ( .A1(n4420), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U4385 ( .A1(n3942), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3813)
         );
  NAND2_X1 U4386 ( .A1(n3867), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3812)
         );
  NAND2_X1 U4387 ( .A1(n3845), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4388 ( .A1(n3851), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4389 ( .A1(n3876), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4390 ( .A1(n4519), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4391 ( .A1(n3861), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4392 ( .A1(n3851), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3845), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4393 ( .A1(n3974), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4394 ( .A1(n3876), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4395 ( .A1(n4109), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4396 ( .A1(n4065), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4397 ( .A1(n4420), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4398 ( .A1(n3866), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4399 ( .A1(n3902), .A2(n3900), .ZN(n3859) );
  NAND2_X1 U4400 ( .A1(n3974), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4401 ( .A1(n4420), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3831) );
  NAND2_X1 U4402 ( .A1(n3851), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4403 ( .A1(n3846), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3829)
         );
  NAND2_X1 U4404 ( .A1(n3942), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3836)
         );
  NAND2_X1 U4405 ( .A1(n4109), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U4406 ( .A1(n3876), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4407 ( .A1(n4524), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3833)
         );
  NAND2_X1 U4408 ( .A1(n4318), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3840)
         );
  NAND2_X1 U4409 ( .A1(n3845), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4410 ( .A1(n4518), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3838) );
  NAND2_X1 U4411 ( .A1(n4519), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4412 ( .A1(n3861), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4413 ( .A1(n4109), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3845), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4414 ( .A1(n3866), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4415 ( .A1(n4420), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3846), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4416 ( .A1(n4065), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4417 ( .A1(n3942), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4418 ( .A1(n4318), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4419 ( .A1(n3851), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U4420 ( .A1(n3926), .A2(n3857), .ZN(n4778) );
  INV_X1 U4421 ( .A(n4936), .ZN(n3858) );
  NAND2_X1 U4422 ( .A1(n4318), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3865)
         );
  NAND2_X1 U4423 ( .A1(n3861), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4424 ( .A1(n3845), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4425 ( .A1(n4518), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4426 ( .A1(n4065), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4427 ( .A1(n3866), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3870)
         );
  NAND2_X1 U4428 ( .A1(n3974), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4429 ( .A1(n3867), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3868)
         );
  NAND2_X1 U4430 ( .A1(n3851), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4431 ( .A1(n4420), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4432 ( .A1(n4519), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4433 ( .A1(n3846), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3872)
         );
  NAND2_X1 U4434 ( .A1(n3942), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3880)
         );
  NAND2_X1 U4435 ( .A1(n4109), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4436 ( .A1(n3876), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3878) );
  NAND2_X1 U4437 ( .A1(n4524), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3877)
         );
  NAND2_X1 U4438 ( .A1(n5073), .A2(n3926), .ZN(n4926) );
  NOR2_X2 U4439 ( .A1(n4929), .A2(n4926), .ZN(n4911) );
  OAI211_X1 U4440 ( .C1(n3909), .C2(n4229), .A(n3931), .B(n4911), .ZN(n3895)
         );
  OAI21_X1 U4441 ( .B1(n3902), .B2(n5073), .A(n3907), .ZN(n3885) );
  INV_X1 U4442 ( .A(n3885), .ZN(n3891) );
  NAND4_X1 U4443 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n4967)
         );
  NAND2_X1 U4444 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  NAND2_X1 U4445 ( .A1(n3892), .A2(n3905), .ZN(n3894) );
  AND2_X1 U4446 ( .A1(n3926), .A2(n3905), .ZN(n4008) );
  NAND2_X1 U4447 ( .A1(n4008), .A2(n3637), .ZN(n3893) );
  NAND2_X1 U4448 ( .A1(n3894), .A2(n3893), .ZN(n3921) );
  NAND2_X1 U4449 ( .A1(n3951), .A2(n3637), .ZN(n3896) );
  NAND2_X1 U4450 ( .A1(n4024), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4451 ( .A1(n7517), .A2(n4049), .ZN(n4755) );
  INV_X1 U4452 ( .A(n4755), .ZN(n4062) );
  NAND2_X1 U4453 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U4454 ( .A1(n6967), .A2(n6784), .ZN(n5824) );
  NAND2_X1 U4455 ( .A1(n4062), .A2(n6707), .ZN(n3899) );
  INV_X1 U4456 ( .A(n4258), .ZN(n4027) );
  NAND2_X1 U4457 ( .A1(n4027), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3898) );
  NOR2_X1 U4458 ( .A1(n4926), .A2(n4967), .ZN(n3903) );
  INV_X1 U4459 ( .A(n5073), .ZN(n4986) );
  NAND2_X1 U4461 ( .A1(n4772), .A2(n3907), .ZN(n4903) );
  NAND2_X1 U4462 ( .A1(n5069), .A2(n5073), .ZN(n4928) );
  NAND2_X1 U4463 ( .A1(n4970), .A2(n3925), .ZN(n4935) );
  NAND2_X1 U4464 ( .A1(n3910), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3912) );
  NAND3_X1 U4465 ( .A1(n3911), .A2(n3913), .A3(n3912), .ZN(n4022) );
  INV_X1 U4466 ( .A(n3912), .ZN(n3915) );
  INV_X1 U4467 ( .A(n3913), .ZN(n3914) );
  NAND2_X1 U4468 ( .A1(n3915), .A2(n3742), .ZN(n3916) );
  NAND2_X1 U4469 ( .A1(n4022), .A2(n3916), .ZN(n4019) );
  NAND2_X1 U4470 ( .A1(n4024), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3918) );
  MUX2_X1 U4471 ( .A(n4258), .B(n4755), .S(n6784), .Z(n3917) );
  NAND2_X1 U4472 ( .A1(n3921), .A2(n5003), .ZN(n3923) );
  OR2_X1 U4473 ( .A1(n3905), .A2(n5073), .ZN(n3922) );
  NAND2_X1 U4474 ( .A1(n3923), .A2(n3922), .ZN(n4934) );
  AOI21_X1 U4475 ( .B1(n3924), .B2(n3925), .A(n3926), .ZN(n3928) );
  INV_X1 U4476 ( .A(n3992), .ZN(n4010) );
  AND2_X1 U4477 ( .A1(n7517), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U4478 ( .B1(n4010), .B2(n3637), .A(n7523), .ZN(n3927) );
  NOR2_X1 U4479 ( .A1(n3928), .A2(n3927), .ZN(n3933) );
  INV_X1 U4480 ( .A(n3929), .ZN(n3930) );
  NAND3_X1 U4481 ( .A1(n4437), .A2(n5196), .A3(n3930), .ZN(n3932) );
  NAND3_X1 U4482 ( .A1(n3933), .A2(n3932), .A3(n3931), .ZN(n3934) );
  XNOR2_X1 U4483 ( .A(n4019), .B(n4020), .ZN(n5046) );
  AOI22_X1 U4484 ( .A1(n4731), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4485 ( .A1(n4707), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4486 ( .A1(n4677), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4487 ( .A1(n3936), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4488 ( .A1(n4593), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4489 ( .A1(n4701), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4490 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3946)
         );
  AOI22_X1 U4491 ( .A1(n4722), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4492 ( .A1(n4700), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3943) );
  INV_X1 U4493 ( .A(n3967), .ZN(n3965) );
  NAND2_X1 U4494 ( .A1(n3951), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4495 ( .A1(n4722), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4496 ( .A1(n4677), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4497 ( .A1(n3936), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4498 ( .A1(n4547), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4499 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3961)
         );
  AOI22_X1 U4500 ( .A1(n4701), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4501 ( .A1(n4700), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4502 ( .A1(n4723), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4503 ( .A1(n3937), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4504 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  OR2_X1 U4505 ( .A1(n4036), .A2(n4166), .ZN(n3962) );
  OAI211_X1 U4506 ( .C1(n3994), .C2(n4035), .A(n3963), .B(n3962), .ZN(n3966)
         );
  INV_X1 U4507 ( .A(n3966), .ZN(n3964) );
  NAND2_X1 U4508 ( .A1(n3643), .A2(n3966), .ZN(n3968) );
  INV_X1 U4509 ( .A(n3970), .ZN(n3971) );
  NAND2_X1 U4510 ( .A1(n4020), .A2(n3973), .ZN(n4267) );
  INV_X1 U4511 ( .A(n4036), .ZN(n3986) );
  AOI22_X1 U4512 ( .A1(n4547), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4513 ( .A1(n3974), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4514 ( .A1(n3936), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4515 ( .A1(n3937), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4516 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3984)
         );
  AOI22_X1 U4517 ( .A1(n4701), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4518 ( .A1(n4700), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4519 ( .A1(n4722), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4520 ( .A1(n4723), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4521 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3983)
         );
  XNOR2_X1 U4522 ( .A(n3990), .B(n4009), .ZN(n3985) );
  NAND2_X1 U4523 ( .A1(n3986), .A2(n3985), .ZN(n4002) );
  OAI21_X1 U4524 ( .B1(n4267), .B2(STATE2_REG_0__SCAN_IN), .A(n4002), .ZN(
        n3989) );
  INV_X1 U4525 ( .A(n4009), .ZN(n3995) );
  NAND2_X1 U4526 ( .A1(n3951), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3988) );
  AOI21_X1 U4527 ( .B1(n3920), .B2(n4166), .A(n4049), .ZN(n3987) );
  OAI211_X1 U4528 ( .C1(n3995), .C2(n3645), .A(n3988), .B(n3987), .ZN(n4003)
         );
  NAND2_X1 U4529 ( .A1(n4261), .A2(n4984), .ZN(n4001) );
  NAND2_X1 U4530 ( .A1(n4009), .A2(n3993), .ZN(n4080) );
  NAND2_X1 U4531 ( .A1(n3992), .A2(n4080), .ZN(n4055) );
  INV_X1 U4532 ( .A(n4055), .ZN(n3999) );
  NAND2_X1 U4533 ( .A1(n3995), .A2(n3994), .ZN(n3998) );
  INV_X1 U4534 ( .A(n3996), .ZN(n3997) );
  AOI21_X1 U4535 ( .B1(n3999), .B2(n3998), .A(n3997), .ZN(n4000) );
  INV_X1 U4536 ( .A(n4002), .ZN(n4004) );
  INV_X1 U4537 ( .A(n4984), .ZN(n4007) );
  INV_X1 U4538 ( .A(n4008), .ZN(n5004) );
  OAI21_X1 U4539 ( .B1(n4010), .B2(n4009), .A(n5004), .ZN(n4011) );
  INV_X1 U4540 ( .A(n4011), .ZN(n4012) );
  NAND2_X1 U4541 ( .A1(n4013), .A2(n4012), .ZN(n5015) );
  NAND2_X1 U4542 ( .A1(n5133), .A2(n5136), .ZN(n4015) );
  INV_X1 U4543 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U4544 ( .A1(n4014), .A2(n5138), .ZN(n5134) );
  INV_X1 U4545 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7259) );
  INV_X1 U4546 ( .A(n4019), .ZN(n4021) );
  NAND2_X1 U4547 ( .A1(n4021), .A2(n4020), .ZN(n4023) );
  NAND2_X1 U4548 ( .A1(n4023), .A2(n4022), .ZN(n4033) );
  NAND2_X1 U4549 ( .A1(n4024), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4029) );
  INV_X1 U4550 ( .A(n7592), .ZN(n4025) );
  NAND2_X1 U4551 ( .A1(n7592), .A2(n5904), .ZN(n4026) );
  AOI22_X1 U4552 ( .A1(n5151), .A2(n4062), .B1(n4027), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4028) );
  INV_X1 U4553 ( .A(n4031), .ZN(n4032) );
  NAND2_X1 U4554 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  INV_X1 U4555 ( .A(n4925), .ZN(n4050) );
  INV_X1 U4556 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4557 ( .A1(n4701), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4558 ( .A1(n4318), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4559 ( .A1(n4730), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4560 ( .A1(n4709), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U4561 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4046)
         );
  AOI22_X1 U4562 ( .A1(n3936), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4563 ( .A1(n4700), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4564 ( .A1(n4707), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4565 ( .A1(n3937), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U4566 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4045)
         );
  AOI22_X1 U4567 ( .A1(n4253), .A2(n4078), .B1(n3951), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4047) );
  AOI21_X1 U4568 ( .B1(n4050), .B2(n4049), .A(n4048), .ZN(n4051) );
  INV_X1 U4569 ( .A(n4080), .ZN(n4053) );
  NAND2_X1 U4570 ( .A1(n3992), .A2(n4053), .ZN(n4054) );
  MUX2_X1 U4571 ( .A(n4055), .B(n4054), .S(n4078), .Z(n4056) );
  OAI21_X1 U4572 ( .B1(n5050), .B2(n4007), .A(n3736), .ZN(n4057) );
  INV_X1 U4573 ( .A(n4057), .ZN(n7150) );
  INV_X1 U4574 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U4575 ( .A1(n4024), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4064) );
  NAND2_X1 U4576 ( .A1(n4058), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U4577 ( .A1(n4059), .A2(n6706), .ZN(n4060) );
  NOR2_X1 U4578 ( .A1(n4258), .A2(n6706), .ZN(n4061) );
  AOI21_X1 U4579 ( .B1(n5830), .B2(n4062), .A(n4061), .ZN(n4063) );
  AOI22_X1 U4580 ( .A1(n4722), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4581 ( .A1(n4677), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4582 ( .A1(n3936), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4583 ( .A1(n4547), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U4584 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4075)
         );
  AOI22_X1 U4585 ( .A1(n4701), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4586 ( .A1(n4700), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4587 ( .A1(n4723), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4588 ( .A1(n3937), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U4589 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4074)
         );
  AOI22_X1 U4590 ( .A1(n4253), .A2(n4082), .B1(n3951), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4076) );
  INV_X1 U4591 ( .A(n4078), .ZN(n4079) );
  NAND2_X1 U4592 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  NAND2_X1 U4593 ( .A1(n4081), .A2(n4082), .ZN(n4125) );
  OAI211_X1 U4594 ( .C1(n4082), .C2(n4081), .A(n4125), .B(n3992), .ZN(n4083)
         );
  INV_X1 U4595 ( .A(n4083), .ZN(n4084) );
  AOI21_X1 U4596 ( .B1(n5242), .B2(n4984), .A(n4084), .ZN(n5034) );
  INV_X1 U4597 ( .A(n7157), .ZN(n4102) );
  AOI22_X1 U4598 ( .A1(n3936), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U4599 ( .A1(n4722), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4600 ( .A1(n4708), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4601 ( .A1(n3937), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4087) );
  NAND4_X1 U4602 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4096)
         );
  AOI22_X1 U4603 ( .A1(n4701), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4604 ( .A1(n4730), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U4605 ( .A1(n4700), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4606 ( .A1(n4109), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4091) );
  NAND4_X1 U4607 ( .A1(n4094), .A2(n4093), .A3(n4092), .A4(n4091), .ZN(n4095)
         );
  NAND2_X1 U4608 ( .A1(n4253), .A2(n4123), .ZN(n4098) );
  NAND2_X1 U4609 ( .A1(n3951), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4097) );
  XNOR2_X1 U4610 ( .A(n4125), .B(n4123), .ZN(n4099) );
  NAND2_X1 U4611 ( .A1(n4099), .A2(n3992), .ZN(n4100) );
  XNOR2_X1 U4612 ( .A(n4103), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n7156)
         );
  INV_X1 U4613 ( .A(n7156), .ZN(n4101) );
  NAND2_X1 U4614 ( .A1(n4103), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4104)
         );
  AOI22_X1 U4615 ( .A1(n4722), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4616 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n4677), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4617 ( .A1(n3936), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U4618 ( .A1(n4547), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U4619 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4115)
         );
  AOI22_X1 U4620 ( .A1(n4701), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4621 ( .A1(n4700), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4622 ( .A1(n4109), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U4623 ( .A1(n3937), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U4624 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4114)
         );
  NAND2_X1 U4625 ( .A1(n4253), .A2(n4148), .ZN(n4117) );
  NAND2_X1 U4626 ( .A1(n3951), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4116) );
  NAND2_X1 U4627 ( .A1(n4118), .A2(n4119), .ZN(n4122) );
  NAND2_X1 U4628 ( .A1(n4301), .A2(n4984), .ZN(n4128) );
  INV_X1 U4629 ( .A(n4123), .ZN(n4124) );
  OR2_X1 U4630 ( .A1(n4125), .A2(n4124), .ZN(n4147) );
  XNOR2_X1 U4631 ( .A(n4147), .B(n4148), .ZN(n4126) );
  NAND2_X1 U4632 ( .A1(n4126), .A2(n3992), .ZN(n4127) );
  NAND2_X1 U4633 ( .A1(n4128), .A2(n4127), .ZN(n4129) );
  INV_X1 U4634 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7229) );
  XNOR2_X1 U4635 ( .A(n4129), .B(n7229), .ZN(n7163) );
  NAND2_X1 U4636 ( .A1(n4129), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4130)
         );
  AOI22_X1 U4637 ( .A1(n4700), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4638 ( .A1(n4677), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4639 ( .A1(n4702), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4640 ( .A1(n4701), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4131) );
  NAND4_X1 U4641 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4140)
         );
  AOI22_X1 U4642 ( .A1(n4722), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4643 ( .A1(n3936), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U4644 ( .A1(n4709), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U4645 ( .A1(n4731), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U4646 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4139)
         );
  NAND2_X1 U4647 ( .A1(n4253), .A2(n4156), .ZN(n4142) );
  NAND2_X1 U4648 ( .A1(n3951), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4141) );
  NAND2_X1 U4649 ( .A1(n4146), .A2(n4145), .ZN(n4311) );
  NAND3_X1 U4650 ( .A1(n4154), .A2(n4984), .A3(n4311), .ZN(n4152) );
  INV_X1 U4651 ( .A(n4147), .ZN(n4149) );
  NAND2_X1 U4652 ( .A1(n4149), .A2(n4148), .ZN(n4155) );
  XNOR2_X1 U4653 ( .A(n4155), .B(n4156), .ZN(n4150) );
  NAND2_X1 U4654 ( .A1(n4150), .A2(n3992), .ZN(n4151) );
  NAND2_X1 U4655 ( .A1(n4152), .A2(n4151), .ZN(n7167) );
  AOI22_X1 U4656 ( .A1(n4253), .A2(n4166), .B1(n3951), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4153) );
  XNOR2_X1 U4657 ( .A(n4154), .B(n4153), .ZN(n4317) );
  OR2_X1 U4658 ( .A1(n4317), .A2(n4007), .ZN(n4160) );
  INV_X1 U4659 ( .A(n4155), .ZN(n4157) );
  NAND2_X1 U4660 ( .A1(n4157), .A2(n4156), .ZN(n4168) );
  XNOR2_X1 U4661 ( .A(n4168), .B(n4166), .ZN(n4158) );
  NAND2_X1 U4662 ( .A1(n4158), .A2(n3992), .ZN(n4159) );
  NAND2_X1 U4663 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  INV_X1 U4664 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U4665 ( .A1(n4161), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4162)
         );
  NAND2_X1 U4666 ( .A1(n4166), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U4667 ( .A1(n3992), .A2(n4166), .ZN(n4167) );
  OR2_X1 U4668 ( .A1(n4168), .A2(n4167), .ZN(n4169) );
  NAND2_X1 U4669 ( .A1(n4172), .A2(n4169), .ZN(n4170) );
  INV_X1 U4670 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5991) );
  XNOR2_X1 U4671 ( .A(n4170), .B(n5991), .ZN(n5989) );
  NAND2_X1 U4672 ( .A1(n4170), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4171)
         );
  XNOR2_X1 U4673 ( .A(n4172), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6034)
         );
  INV_X1 U4674 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7265) );
  OR2_X1 U4675 ( .A1(n3618), .A2(n7265), .ZN(n4173) );
  INV_X1 U4676 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U4677 ( .A1(n6444), .A2(n6046), .ZN(n4174) );
  INV_X1 U4678 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6486) );
  INV_X1 U4679 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U4680 ( .A1(n4172), .A2(n6486), .ZN(n6485) );
  XNOR2_X1 U4681 ( .A(n4172), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6477)
         );
  INV_X1 U4682 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4821) );
  XNOR2_X1 U4683 ( .A(n6444), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6471)
         );
  NAND2_X1 U4684 ( .A1(n6469), .A2(n6471), .ZN(n6470) );
  INV_X1 U4685 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U4686 ( .A1(n6444), .A2(n6499), .ZN(n4175) );
  XNOR2_X1 U4687 ( .A(n6444), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6462)
         );
  INV_X1 U4688 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U4689 ( .A1(n6483), .A2(n7285), .ZN(n4176) );
  INV_X1 U4690 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4177) );
  OR2_X1 U4691 ( .A1(n6483), .A2(n4177), .ZN(n4178) );
  NOR2_X1 U4692 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4179) );
  NOR2_X1 U4693 ( .A1(n6444), .A2(n4179), .ZN(n4181) );
  NAND2_X1 U4694 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U4695 ( .A1(n6483), .A2(n6500), .ZN(n4180) );
  NOR2_X1 U4696 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6412) );
  INV_X1 U4697 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6402) );
  INV_X1 U4698 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4182) );
  NAND3_X1 U4699 ( .A1(n6412), .A2(n6402), .A3(n4182), .ZN(n4184) );
  INV_X1 U4700 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6433) );
  INV_X1 U4701 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4183) );
  NAND2_X1 U4702 ( .A1(n6433), .A2(n4183), .ZN(n7209) );
  NOR2_X1 U4703 ( .A1(n4184), .A2(n7209), .ZN(n4185) );
  NAND2_X1 U4704 ( .A1(n6617), .A2(n4185), .ZN(n4186) );
  NAND2_X1 U4705 ( .A1(n4186), .A2(n6443), .ZN(n4192) );
  INV_X1 U4706 ( .A(n6617), .ZN(n4190) );
  AND2_X1 U4707 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7217) );
  AND2_X1 U4708 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U4709 ( .A1(n7217), .A2(n6514), .ZN(n6413) );
  INV_X1 U4710 ( .A(n6413), .ZN(n4188) );
  NAND2_X1 U4711 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6515) );
  INV_X1 U4712 ( .A(n6515), .ZN(n4187) );
  AND2_X1 U4713 ( .A1(n4188), .A2(n4187), .ZN(n4189) );
  NAND2_X1 U4714 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  NAND2_X1 U4715 ( .A1(n4192), .A2(n4191), .ZN(n6392) );
  NAND2_X1 U4716 ( .A1(n6392), .A2(n6393), .ZN(n4194) );
  INV_X1 U4717 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6573) );
  OR2_X1 U4718 ( .A1(n6483), .A2(n6573), .ZN(n4193) );
  INV_X1 U4719 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U4720 ( .A1(n6483), .A2(n6562), .ZN(n4195) );
  INV_X1 U4721 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6554) );
  INV_X1 U4722 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4867) );
  XNOR2_X1 U4723 ( .A(n6483), .B(n4867), .ZN(n6359) );
  AOI21_X1 U4724 ( .B1(n6366), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6359), 
        .ZN(n4200) );
  AND2_X1 U4725 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U4726 ( .A1(n6533), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6523) );
  AND2_X1 U4727 ( .A1(n6483), .A2(n6523), .ZN(n4198) );
  NOR2_X1 U4728 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4196) );
  OR2_X1 U4729 ( .A1(n6444), .A2(n4196), .ZN(n6365) );
  INV_X1 U4730 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6545) );
  OR2_X1 U4731 ( .A1(n6444), .A2(n6545), .ZN(n4197) );
  OAI21_X2 U4732 ( .B1(n6374), .B2(n4198), .A(n6357), .ZN(n6101) );
  NAND2_X1 U4733 ( .A1(n6101), .A2(n4867), .ZN(n4199) );
  NAND3_X1 U4734 ( .A1(n4200), .A2(n4199), .A3(n3737), .ZN(n4201) );
  INV_X1 U4735 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6512) );
  XNOR2_X1 U4736 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U4737 ( .A1(n4231), .A2(n4230), .ZN(n4203) );
  NAND2_X1 U4738 ( .A1(n6967), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4202) );
  NAND2_X1 U4739 ( .A1(n4203), .A2(n4202), .ZN(n4218) );
  NAND2_X1 U4740 ( .A1(n5904), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U4741 ( .A1(n3750), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U4742 ( .A1(n4218), .A2(n4217), .ZN(n4206) );
  NAND2_X1 U4743 ( .A1(n4206), .A2(n4205), .ZN(n4215) );
  XNOR2_X1 U4744 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U4745 ( .A1(n4215), .A2(n4213), .ZN(n4208) );
  NAND2_X1 U4746 ( .A1(n6706), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4207) );
  INV_X1 U4747 ( .A(n4251), .ZN(n4769) );
  INV_X1 U4748 ( .A(n4213), .ZN(n4214) );
  XNOR2_X1 U4749 ( .A(n4215), .B(n4214), .ZN(n4768) );
  INV_X1 U4750 ( .A(n4768), .ZN(n4216) );
  INV_X1 U4751 ( .A(n3951), .ZN(n4233) );
  OAI21_X1 U4752 ( .B1(n4769), .B2(n4216), .A(n4233), .ZN(n4249) );
  INV_X1 U4753 ( .A(n4217), .ZN(n4219) );
  XNOR2_X1 U4754 ( .A(n4219), .B(n4218), .ZN(n4767) );
  INV_X1 U4755 ( .A(n4241), .ZN(n4247) );
  AND2_X1 U4756 ( .A1(n3907), .A2(n4229), .ZN(n4220) );
  INV_X1 U4757 ( .A(n4242), .ZN(n4246) );
  INV_X1 U4758 ( .A(n4231), .ZN(n4221) );
  OAI21_X1 U4759 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6784), .A(n4221), 
        .ZN(n4225) );
  INV_X1 U4760 ( .A(n4225), .ZN(n4224) );
  INV_X1 U4761 ( .A(n4222), .ZN(n4223) );
  AOI21_X1 U4762 ( .B1(n4224), .B2(n3904), .A(n4223), .ZN(n4228) );
  INV_X1 U4763 ( .A(n4253), .ZN(n4226) );
  OAI21_X1 U4764 ( .B1(n4226), .B2(n4225), .A(n4255), .ZN(n4227) );
  OAI21_X1 U4765 ( .B1(n4228), .B2(n4242), .A(n4227), .ZN(n4236) );
  INV_X1 U4766 ( .A(n4236), .ZN(n4240) );
  INV_X1 U4767 ( .A(n4229), .ZN(n6317) );
  INV_X1 U4768 ( .A(n4230), .ZN(n4232) );
  XNOR2_X1 U4769 ( .A(n4232), .B(n4231), .ZN(n4766) );
  NOR2_X1 U4770 ( .A1(n4233), .A2(n4766), .ZN(n4234) );
  AOI211_X1 U4771 ( .C1(n5196), .C2(n4253), .A(n6317), .B(n4234), .ZN(n4237)
         );
  INV_X1 U4772 ( .A(n4237), .ZN(n4239) );
  NAND2_X1 U4773 ( .A1(n4766), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4774 ( .A1(n4237), .A2(n4236), .B1(n4255), .B2(n4235), .ZN(n4238)
         );
  AOI21_X1 U4775 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4245) );
  INV_X1 U4776 ( .A(n4767), .ZN(n4243) );
  AOI211_X1 U4777 ( .C1(n4243), .C2(n3951), .A(n4242), .B(n4241), .ZN(n4244)
         );
  OAI222_X1 U4778 ( .A1(n4247), .A2(n4246), .B1(n4007), .B2(n4768), .C1(n4245), 
        .C2(n4244), .ZN(n4248) );
  AOI22_X1 U4779 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4049), .B1(n4249), .B2(n4248), .ZN(n4250) );
  OR2_X1 U4780 ( .A1(n4926), .A2(n3905), .ZN(n4259) );
  NAND2_X1 U4781 ( .A1(n5052), .A2(n4429), .ZN(n4266) );
  AOI22_X1 U4782 ( .A1(n4745), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5906), .ZN(n4264) );
  NOR2_X1 U4783 ( .A1(n3908), .A2(n5906), .ZN(n4277) );
  NAND2_X1 U4784 ( .A1(n4277), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4263) );
  AND2_X1 U4785 ( .A1(n4264), .A2(n4263), .ZN(n4265) );
  AOI21_X1 U4786 ( .B1(n5057), .B2(n3661), .A(n5906), .ZN(n4981) );
  INV_X2 U4787 ( .A(n3659), .ZN(n4745) );
  AOI22_X1 U4788 ( .A1(n4277), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n4745), .B2(EAX_REG_0__SCAN_IN), .ZN(n4268) );
  OAI21_X1 U4789 ( .B1(n4267), .B2(n4418), .A(n4268), .ZN(n4980) );
  INV_X1 U4790 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n7325) );
  NOR2_X1 U4791 ( .A1(n7325), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4269) );
  OR2_X1 U4792 ( .A1(n4980), .A2(n4269), .ZN(n4983) );
  MUX2_X1 U4793 ( .A(n4286), .B(n4981), .S(n4983), .Z(n4966) );
  NAND2_X1 U4794 ( .A1(n4277), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4274) );
  INV_X1 U4795 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4271) );
  NAND2_X1 U4796 ( .A1(n7200), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4605) );
  NAND2_X1 U4797 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4278) );
  OAI21_X1 U4798 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4278), .ZN(n7155) );
  NAND2_X1 U4799 ( .A1(n4286), .A2(n7155), .ZN(n4270) );
  OAI21_X1 U4800 ( .B1(n4271), .B2(n4605), .A(n4270), .ZN(n4272) );
  AOI21_X1 U4801 ( .B1(n4745), .B2(EAX_REG_2__SCAN_IN), .A(n4272), .ZN(n4273)
         );
  AND2_X1 U4802 ( .A1(n4274), .A2(n4273), .ZN(n5234) );
  NAND2_X1 U4803 ( .A1(n4965), .A2(n5234), .ZN(n4275) );
  OAI21_X1 U4804 ( .B1(n4276), .B2(n5233), .A(n4275), .ZN(n5020) );
  INV_X1 U4805 ( .A(n4277), .ZN(n4291) );
  INV_X1 U4806 ( .A(n4278), .ZN(n4280) );
  INV_X1 U4807 ( .A(n4287), .ZN(n4279) );
  OAI21_X1 U4808 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4280), .A(n4279), 
        .ZN(n5964) );
  AOI22_X1 U4809 ( .A1(n4286), .A2(n5964), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U4810 ( .A1(n4745), .A2(EAX_REG_3__SCAN_IN), .ZN(n4281) );
  OAI211_X1 U4811 ( .C1(n4291), .C2(n3744), .A(n4282), .B(n4281), .ZN(n4283)
         );
  NOR2_X2 U4812 ( .A1(n5020), .A2(n5023), .ZN(n5021) );
  INV_X1 U4813 ( .A(n4284), .ZN(n4285) );
  OAI21_X1 U4814 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4287), .A(n4296), 
        .ZN(n7340) );
  INV_X1 U4815 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4288) );
  AOI21_X1 U4816 ( .B1(n4288), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4289) );
  AOI21_X1 U4817 ( .B1(n4745), .B2(EAX_REG_4__SCAN_IN), .A(n4289), .ZN(n4290)
         );
  OAI21_X1 U4818 ( .B1(n4291), .B2(n7520), .A(n4290), .ZN(n4292) );
  OAI21_X1 U4819 ( .B1(n4743), .B2(n7340), .A(n4292), .ZN(n4293) );
  NAND2_X1 U4820 ( .A1(n4294), .A2(n4293), .ZN(n5239) );
  NAND2_X1 U4821 ( .A1(n5021), .A2(n5239), .ZN(n5029) );
  INV_X1 U4822 ( .A(n5029), .ZN(n4303) );
  INV_X1 U4823 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4299) );
  INV_X1 U4824 ( .A(n4304), .ZN(n4305) );
  INV_X1 U4825 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7344) );
  NAND2_X1 U4826 ( .A1(n7344), .A2(n4296), .ZN(n4297) );
  NAND2_X1 U4827 ( .A1(n4305), .A2(n4297), .ZN(n7353) );
  AOI22_X1 U4828 ( .A1(n7353), .A2(n4286), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4298) );
  OAI21_X1 U4829 ( .B1(n3659), .B2(n4299), .A(n4298), .ZN(n4300) );
  NAND2_X1 U4830 ( .A1(n4303), .A2(n4302), .ZN(n5027) );
  INV_X1 U4831 ( .A(n4312), .ZN(n4307) );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U4833 ( .A1(n4305), .A2(n7355), .ZN(n4306) );
  NAND2_X1 U4834 ( .A1(n4307), .A2(n4306), .ZN(n7363) );
  INV_X1 U4835 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4308) );
  OAI22_X1 U4836 ( .A1(n3659), .A2(n4308), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7355), .ZN(n4309) );
  MUX2_X1 U4837 ( .A(n7363), .B(n4309), .S(n4743), .Z(n4310) );
  NOR2_X2 U4838 ( .A1(n5027), .A2(n5784), .ZN(n5700) );
  INV_X1 U4839 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4314) );
  OAI21_X1 U4840 ( .B1(n4312), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4334), 
        .ZN(n7374) );
  AOI22_X1 U4841 ( .A1(n7374), .A2(n4286), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U4842 ( .A1(n5700), .A2(n5701), .ZN(n5699) );
  AOI22_X1 U4843 ( .A1(n4745), .A2(EAX_REG_8__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U4844 ( .A1(n4731), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4845 ( .A1(n3936), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4846 ( .A1(n4318), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U4847 ( .A1(n4708), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4319) );
  NAND4_X1 U4848 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4328)
         );
  AOI22_X1 U4849 ( .A1(n4730), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4850 ( .A1(n4701), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4851 ( .A1(n4700), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U4852 ( .A1(n3937), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U4853 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4327)
         );
  OR2_X1 U4854 ( .A1(n4328), .A2(n4327), .ZN(n4330) );
  INV_X1 U4855 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4329) );
  XNOR2_X1 U4856 ( .A(n4334), .B(n4329), .ZN(n7381) );
  AOI22_X1 U4857 ( .A1(n4429), .A2(n4330), .B1(n4286), .B2(n7381), .ZN(n4331)
         );
  XOR2_X1 U4858 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4357), .Z(n7392) );
  AOI22_X1 U4859 ( .A1(n4745), .A2(EAX_REG_9__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4860 ( .A1(n4730), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4861 ( .A1(n4708), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U4862 ( .A1(n4731), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4863 ( .A1(n4722), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4335) );
  NAND4_X1 U4864 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4344)
         );
  AOI22_X1 U4865 ( .A1(n3936), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4701), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U4866 ( .A1(n4723), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U4867 ( .A1(n4677), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4868 ( .A1(n4700), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4339) );
  NAND4_X1 U4869 ( .A1(n4342), .A2(n4341), .A3(n4340), .A4(n4339), .ZN(n4343)
         );
  OAI21_X1 U4870 ( .B1(n4344), .B2(n4343), .A(n4429), .ZN(n4345) );
  OAI211_X1 U4871 ( .C1(n7392), .C2(n4743), .A(n4346), .B(n4345), .ZN(n5947)
         );
  AOI22_X1 U4872 ( .A1(n4723), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4873 ( .A1(n3936), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4874 ( .A1(n4702), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4875 ( .A1(n4700), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U4876 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4356)
         );
  AOI22_X1 U4877 ( .A1(n4701), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4878 ( .A1(n4730), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4879 ( .A1(n4707), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U4880 ( .A1(n3937), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4351) );
  NAND4_X1 U4881 ( .A1(n4354), .A2(n4353), .A3(n4352), .A4(n4351), .ZN(n4355)
         );
  NOR2_X1 U4882 ( .A1(n4356), .A2(n4355), .ZN(n4360) );
  XNOR2_X1 U4883 ( .A(n4361), .B(n6254), .ZN(n6247) );
  NAND2_X1 U4884 ( .A1(n6247), .A2(n4286), .ZN(n4359) );
  AOI22_X1 U4885 ( .A1(n4745), .A2(EAX_REG_10__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4358) );
  OAI211_X1 U4886 ( .C1(n4360), .C2(n4418), .A(n4359), .B(n4358), .ZN(n5975)
         );
  XOR2_X1 U4887 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4385), .Z(n7172) );
  AOI22_X1 U4888 ( .A1(n4745), .A2(EAX_REG_11__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4889 ( .A1(n4677), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4890 ( .A1(n4702), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4891 ( .A1(n4701), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U4892 ( .A1(n4731), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U4893 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4371)
         );
  AOI22_X1 U4894 ( .A1(n4722), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4895 ( .A1(n3936), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4896 ( .A1(n4723), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U4897 ( .A1(n4700), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4366) );
  NAND4_X1 U4898 ( .A1(n4369), .A2(n4368), .A3(n4367), .A4(n4366), .ZN(n4370)
         );
  OAI21_X1 U4899 ( .B1(n4371), .B2(n4370), .A(n4429), .ZN(n4372) );
  OAI211_X1 U4900 ( .C1(n7172), .C2(n4743), .A(n4373), .B(n4372), .ZN(n6001)
         );
  NOR2_X2 U4901 ( .A1(n5973), .A2(n4374), .ZN(n5999) );
  AOI22_X1 U4902 ( .A1(n4700), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4903 ( .A1(n4677), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4904 ( .A1(n4709), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4905 ( .A1(n4701), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4906 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4384)
         );
  AOI22_X1 U4907 ( .A1(n3936), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4908 ( .A1(n4731), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U4909 ( .A1(n4708), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4380) );
  AOI22_X1 U4910 ( .A1(n4702), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4379) );
  NAND4_X1 U4911 ( .A1(n4382), .A2(n4381), .A3(n4380), .A4(n4379), .ZN(n4383)
         );
  NOR2_X1 U4912 ( .A1(n4384), .A2(n4383), .ZN(n4389) );
  INV_X1 U4913 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4386) );
  XNOR2_X1 U4914 ( .A(n4401), .B(n4386), .ZN(n6491) );
  NAND2_X1 U4915 ( .A1(n6491), .A2(n4286), .ZN(n4388) );
  AOI22_X1 U4916 ( .A1(n4745), .A2(EAX_REG_12__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4387) );
  OAI211_X1 U4917 ( .C1(n4389), .C2(n4418), .A(n4388), .B(n4387), .ZN(n6017)
         );
  NAND2_X1 U4918 ( .A1(n5999), .A2(n6017), .ZN(n6016) );
  AOI22_X1 U4919 ( .A1(n4701), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U4920 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n3936), .B1(n4730), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4921 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n4707), .B1(n4708), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4922 ( .A1(n3937), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4390) );
  NAND4_X1 U4923 ( .A1(n4393), .A2(n4392), .A3(n4391), .A4(n4390), .ZN(n4399)
         );
  AOI22_X1 U4924 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n4722), .B1(n4702), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4925 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n4731), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4926 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n4677), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U4927 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4723), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4394) );
  NAND4_X1 U4928 ( .A1(n4397), .A2(n4396), .A3(n4395), .A4(n4394), .ZN(n4398)
         );
  NAND2_X1 U4929 ( .A1(n4429), .A2(n4400), .ZN(n4403) );
  XNOR2_X1 U4930 ( .A(n4414), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n7400)
         );
  INV_X1 U4931 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7045) );
  INV_X1 U4932 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n7397) );
  OAI22_X1 U4933 ( .A1(n3659), .A2(n7045), .B1(n4605), .B2(n7397), .ZN(n4402)
         );
  AOI21_X1 U4934 ( .B1(n7400), .B2(n4286), .A(n4402), .ZN(n6352) );
  AOI22_X1 U4935 ( .A1(n3936), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4701), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U4936 ( .A1(n4722), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4937 ( .A1(n4677), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4938 ( .A1(n4723), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4404) );
  NAND4_X1 U4939 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4413)
         );
  AOI22_X1 U4940 ( .A1(n4730), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4941 ( .A1(n4593), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4942 ( .A1(n4731), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4943 ( .A1(n4700), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4944 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4412)
         );
  NOR2_X1 U4945 ( .A1(n4413), .A2(n4412), .ZN(n4417) );
  NAND2_X1 U4946 ( .A1(n4745), .A2(EAX_REG_14__SCAN_IN), .ZN(n4416) );
  XNOR2_X1 U4947 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4419), .ZN(n7417)
         );
  AOI22_X1 U4948 ( .A1(n4286), .A2(n7417), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4415) );
  OAI211_X1 U4949 ( .C1(n4418), .C2(n4417), .A(n4416), .B(n4415), .ZN(n6348)
         );
  XOR2_X1 U4950 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4436), .Z(n7432) );
  AOI22_X1 U4951 ( .A1(n4745), .A2(EAX_REG_15__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U4952 ( .A1(n4701), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U4953 ( .A1(n3936), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4423) );
  AOI22_X1 U4954 ( .A1(n4702), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4422) );
  AOI22_X1 U4955 ( .A1(n3937), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4421) );
  NAND4_X1 U4956 ( .A1(n4424), .A2(n4423), .A3(n4422), .A4(n4421), .ZN(n4431)
         );
  AOI22_X1 U4957 ( .A1(n4700), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4958 ( .A1(n4722), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U4959 ( .A1(n4730), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U4960 ( .A1(n4723), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4425) );
  NAND4_X1 U4961 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), .ZN(n4430)
         );
  OAI21_X1 U4962 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4432) );
  OAI211_X1 U4963 ( .C1(n7432), .C2(n4743), .A(n4433), .B(n4432), .ZN(n4434)
         );
  INV_X1 U4964 ( .A(n4434), .ZN(n6309) );
  NAND2_X1 U4965 ( .A1(n4435), .A2(n4434), .ZN(n6227) );
  XNOR2_X1 U4966 ( .A(n4452), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6232)
         );
  INV_X1 U4967 ( .A(n6232), .ZN(n6456) );
  AOI22_X1 U4968 ( .A1(n3936), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U4969 ( .A1(n4730), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U4970 ( .A1(n4709), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U4971 ( .A1(n4707), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4439) );
  NAND4_X1 U4972 ( .A1(n4442), .A2(n4441), .A3(n4440), .A4(n4439), .ZN(n4448)
         );
  AOI22_X1 U4973 ( .A1(n4677), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U4974 ( .A1(n4723), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4975 ( .A1(n4708), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U4976 ( .A1(n4701), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4443) );
  NAND4_X1 U4977 ( .A1(n4446), .A2(n4445), .A3(n4444), .A4(n4443), .ZN(n4447)
         );
  NOR2_X1 U4978 ( .A1(n4448), .A2(n4447), .ZN(n4450) );
  AOI22_X1 U4979 ( .A1(n4745), .A2(EAX_REG_16__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U4980 ( .B1(n4747), .B2(n4450), .A(n4449), .ZN(n4451) );
  AOI21_X1 U4981 ( .B1(n6456), .B2(n4286), .A(n4451), .ZN(n6230) );
  OR2_X1 U4982 ( .A1(n4453), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4454)
         );
  NAND2_X1 U4983 ( .A1(n4454), .A2(n4486), .ZN(n7435) );
  INV_X1 U4984 ( .A(n7435), .ZN(n4469) );
  AOI22_X1 U4985 ( .A1(n4677), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4986 ( .A1(n4701), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U4987 ( .A1(n4702), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U4988 ( .A1(n4700), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4455) );
  NAND4_X1 U4989 ( .A1(n4458), .A2(n4457), .A3(n4456), .A4(n4455), .ZN(n4464)
         );
  AOI22_X1 U4990 ( .A1(n4730), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U4991 ( .A1(n4723), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U4992 ( .A1(n4731), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U4993 ( .A1(n3936), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4459) );
  NAND4_X1 U4994 ( .A1(n4462), .A2(n4461), .A3(n4460), .A4(n4459), .ZN(n4463)
         );
  OR2_X1 U4995 ( .A1(n4464), .A2(n4463), .ZN(n4467) );
  INV_X1 U4996 ( .A(EAX_REG_17__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U4997 ( .A1(n5906), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4465)
         );
  OAI211_X1 U4998 ( .C1(n3659), .C2(n7558), .A(n4743), .B(n4465), .ZN(n4466)
         );
  AOI21_X1 U4999 ( .B1(n4690), .B2(n4467), .A(n4466), .ZN(n4468) );
  AOI21_X1 U5000 ( .B1(n4469), .B2(n4286), .A(n4468), .ZN(n6300) );
  NAND2_X1 U5001 ( .A1(n6229), .A2(n6300), .ZN(n6210) );
  AOI22_X1 U5002 ( .A1(n4701), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5003 ( .A1(n4677), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5004 ( .A1(n4731), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5005 ( .A1(n4709), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4470) );
  NAND4_X1 U5006 ( .A1(n4473), .A2(n4472), .A3(n4471), .A4(n4470), .ZN(n4479)
         );
  AOI22_X1 U5007 ( .A1(n3936), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5008 ( .A1(n4730), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5009 ( .A1(n4722), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4475) );
  AOI22_X1 U5010 ( .A1(n4707), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4474) );
  NAND4_X1 U5011 ( .A1(n4477), .A2(n4476), .A3(n4475), .A4(n4474), .ZN(n4478)
         );
  NOR2_X1 U5012 ( .A1(n4479), .A2(n4478), .ZN(n4483) );
  NAND2_X1 U5013 ( .A1(n7200), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4480)
         );
  NAND2_X1 U5014 ( .A1(n4743), .A2(n4480), .ZN(n4481) );
  AOI21_X1 U5015 ( .B1(n4745), .B2(EAX_REG_18__SCAN_IN), .A(n4481), .ZN(n4482)
         );
  OAI21_X1 U5016 ( .B1(n4747), .B2(n4483), .A(n4482), .ZN(n4485) );
  XNOR2_X1 U5017 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4486), .ZN(n6450)
         );
  NAND2_X1 U5018 ( .A1(n4286), .A2(n6450), .ZN(n4484) );
  OR2_X1 U5019 ( .A1(n4487), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4488)
         );
  NAND2_X1 U5020 ( .A1(n4488), .A2(n4534), .ZN(n7448) );
  AOI22_X1 U5021 ( .A1(n4701), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U5022 ( .A1(n3936), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5023 ( .A1(n4723), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U5024 ( .A1(n4708), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4489) );
  NAND4_X1 U5025 ( .A1(n4492), .A2(n4491), .A3(n4490), .A4(n4489), .ZN(n4498)
         );
  AOI22_X1 U5026 ( .A1(n4677), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4496) );
  AOI22_X1 U5027 ( .A1(n4731), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5028 ( .A1(n4707), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5029 ( .A1(n3937), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4493) );
  NAND4_X1 U5030 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), .ZN(n4497)
         );
  NOR2_X1 U5031 ( .A1(n4498), .A2(n4497), .ZN(n4501) );
  OAI21_X1 U5032 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n7535), .A(n7200), 
        .ZN(n4500) );
  NAND2_X1 U5033 ( .A1(n4745), .A2(EAX_REG_19__SCAN_IN), .ZN(n4499) );
  OAI211_X1 U5034 ( .C1(n4747), .C2(n4501), .A(n4500), .B(n4499), .ZN(n4502)
         );
  OAI21_X1 U5035 ( .B1(n7448), .B2(n4743), .A(n4502), .ZN(n6293) );
  AOI22_X1 U5036 ( .A1(n3936), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5037 ( .A1(n4722), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5038 ( .A1(n3937), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5039 ( .A1(n4723), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4503) );
  NAND4_X1 U5040 ( .A1(n4506), .A2(n4505), .A3(n4504), .A4(n4503), .ZN(n4512)
         );
  AOI22_X1 U5041 ( .A1(n4701), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5042 ( .A1(n4730), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5043 ( .A1(n4707), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4518), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4508) );
  AOI22_X1 U5044 ( .A1(n4700), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4524), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4507) );
  NAND4_X1 U5045 ( .A1(n4510), .A2(n4509), .A3(n4508), .A4(n4507), .ZN(n4511)
         );
  NOR2_X1 U5046 ( .A1(n4512), .A2(n4511), .ZN(n4515) );
  INV_X1 U5047 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6436) );
  AOI21_X1 U5048 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6436), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4513) );
  AOI21_X1 U5049 ( .B1(n4745), .B2(EAX_REG_20__SCAN_IN), .A(n4513), .ZN(n4514)
         );
  OAI21_X1 U5050 ( .B1(n4747), .B2(n4515), .A(n4514), .ZN(n4517) );
  XNOR2_X1 U5051 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4534), .ZN(n6438)
         );
  NAND2_X1 U5052 ( .A1(n4286), .A2(n6438), .ZN(n4516) );
  AOI22_X1 U5053 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n4731), .B1(n4702), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5054 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4708), .B1(n4707), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5055 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4730), .B1(n4518), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5056 ( .A1(n4700), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4519), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4520) );
  NAND4_X1 U5057 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4530)
         );
  AOI22_X1 U5058 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3936), .B1(n4722), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5059 ( .A1(n4701), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5060 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n4723), .B1(n4524), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5061 ( .A1(n4677), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4525) );
  NAND4_X1 U5062 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4529)
         );
  NOR2_X1 U5063 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  OR2_X1 U5064 ( .A1(n4747), .A2(n4531), .ZN(n4542) );
  NAND2_X1 U5065 ( .A1(n5906), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4532)
         );
  NAND2_X1 U5066 ( .A1(n4743), .A2(n4532), .ZN(n4533) );
  AOI21_X1 U5067 ( .B1(n4745), .B2(EAX_REG_21__SCAN_IN), .A(n4533), .ZN(n4541)
         );
  INV_X1 U5068 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4538) );
  INV_X1 U5069 ( .A(n4536), .ZN(n4537) );
  NAND2_X1 U5070 ( .A1(n4538), .A2(n4537), .ZN(n4539) );
  NAND2_X1 U5071 ( .A1(n4586), .A2(n4539), .ZN(n7471) );
  NOR2_X1 U5072 ( .A1(n7471), .A2(n4743), .ZN(n4540) );
  AOI21_X1 U5073 ( .B1(n4542), .B2(n4541), .A(n4540), .ZN(n6285) );
  NAND2_X1 U5074 ( .A1(n6195), .A2(n6285), .ZN(n6278) );
  AOI22_X1 U5075 ( .A1(n4700), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4723), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4546) );
  AOI22_X1 U5076 ( .A1(n3936), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4677), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5077 ( .A1(n4722), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5078 ( .A1(n3937), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4543) );
  NAND4_X1 U5079 ( .A1(n4546), .A2(n4545), .A3(n4544), .A4(n4543), .ZN(n4553)
         );
  AOI22_X1 U5080 ( .A1(n4701), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4551) );
  AOI22_X1 U5081 ( .A1(n4730), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5082 ( .A1(n4547), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5083 ( .A1(n4709), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4548) );
  NAND4_X1 U5084 ( .A1(n4551), .A2(n4550), .A3(n4549), .A4(n4548), .ZN(n4552)
         );
  NOR2_X1 U5085 ( .A1(n4553), .A2(n4552), .ZN(n4556) );
  OAI21_X1 U5086 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7479), .A(n4743), .ZN(
        n4554) );
  AOI21_X1 U5087 ( .B1(n4745), .B2(EAX_REG_22__SCAN_IN), .A(n4554), .ZN(n4555)
         );
  OAI21_X1 U5088 ( .B1(n4747), .B2(n4556), .A(n4555), .ZN(n4558) );
  XNOR2_X1 U5089 ( .A(n4586), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n7484)
         );
  NAND2_X1 U5090 ( .A1(n7484), .A2(n4286), .ZN(n4557) );
  NAND2_X1 U5091 ( .A1(n4558), .A2(n4557), .ZN(n6280) );
  AOI22_X1 U5092 ( .A1(n4722), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5093 ( .A1(n4677), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5094 ( .A1(n3936), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5095 ( .A1(n4702), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4560) );
  NAND4_X1 U5096 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4569)
         );
  AOI22_X1 U5097 ( .A1(n4701), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5098 ( .A1(n4700), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5099 ( .A1(n4723), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5100 ( .A1(n3937), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4564) );
  NAND4_X1 U5101 ( .A1(n4567), .A2(n4566), .A3(n4565), .A4(n4564), .ZN(n4568)
         );
  OR2_X1 U5102 ( .A1(n4569), .A2(n4568), .ZN(n4581) );
  AOI22_X1 U5103 ( .A1(n4722), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5104 ( .A1(n4677), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5105 ( .A1(n3936), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5106 ( .A1(n4702), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4570) );
  NAND4_X1 U5107 ( .A1(n4573), .A2(n4572), .A3(n4571), .A4(n4570), .ZN(n4579)
         );
  AOI22_X1 U5108 ( .A1(n4701), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4577) );
  AOI22_X1 U5109 ( .A1(n4700), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5110 ( .A1(n4723), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5111 ( .A1(n3937), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4574) );
  NAND4_X1 U5112 ( .A1(n4577), .A2(n4576), .A3(n4575), .A4(n4574), .ZN(n4578)
         );
  OR2_X1 U5113 ( .A1(n4579), .A2(n4578), .ZN(n4580) );
  NAND2_X1 U5114 ( .A1(n4580), .A2(n4581), .ZN(n4620) );
  OAI21_X1 U5115 ( .B1(n4581), .B2(n4580), .A(n4620), .ZN(n4585) );
  NAND2_X1 U5116 ( .A1(n5906), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4582)
         );
  NAND2_X1 U5117 ( .A1(n4743), .A2(n4582), .ZN(n4583) );
  AOI21_X1 U5118 ( .B1(n4745), .B2(EAX_REG_23__SCAN_IN), .A(n4583), .ZN(n4584)
         );
  OAI21_X1 U5119 ( .B1(n4747), .B2(n4585), .A(n4584), .ZN(n4592) );
  INV_X1 U5120 ( .A(n4587), .ZN(n4589) );
  INV_X1 U5121 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5122 ( .A1(n4589), .A2(n4588), .ZN(n4590) );
  NAND2_X1 U5123 ( .A1(n4625), .A2(n4590), .ZN(n7492) );
  NAND2_X1 U5124 ( .A1(n4592), .A2(n4591), .ZN(n6273) );
  AOI22_X1 U5125 ( .A1(n4701), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5126 ( .A1(n3936), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U5127 ( .A1(n4723), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5128 ( .A1(n4708), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4594) );
  NAND4_X1 U5129 ( .A1(n4597), .A2(n4596), .A3(n4595), .A4(n4594), .ZN(n4603)
         );
  AOI22_X1 U5130 ( .A1(n4677), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5131 ( .A1(n4731), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5132 ( .A1(n4722), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5133 ( .A1(n3937), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4598) );
  NAND4_X1 U5134 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4602)
         );
  NOR2_X1 U5135 ( .A1(n4603), .A2(n4602), .ZN(n4621) );
  XNOR2_X1 U5136 ( .A(n4620), .B(n4621), .ZN(n4604) );
  OR2_X1 U5137 ( .A1(n4747), .A2(n4604), .ZN(n4609) );
  INV_X1 U5138 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6187) );
  NOR2_X1 U5139 ( .A1(n4605), .A2(n6187), .ZN(n4607) );
  XNOR2_X1 U5140 ( .A(n4625), .B(n6187), .ZN(n6407) );
  AOI211_X1 U5141 ( .C1(n4745), .C2(EAX_REG_24__SCAN_IN), .A(n4607), .B(n4606), 
        .ZN(n4608) );
  NAND2_X1 U5142 ( .A1(n4609), .A2(n4608), .ZN(n6180) );
  AOI22_X1 U5143 ( .A1(n4722), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5144 ( .A1(n4677), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5145 ( .A1(n3936), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4611) );
  AOI22_X1 U5146 ( .A1(n4702), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4610) );
  NAND4_X1 U5147 ( .A1(n4613), .A2(n4612), .A3(n4611), .A4(n4610), .ZN(n4619)
         );
  AOI22_X1 U5148 ( .A1(n4701), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4617) );
  AOI22_X1 U5149 ( .A1(n4700), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5150 ( .A1(n4723), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4615) );
  AOI22_X1 U5151 ( .A1(n3937), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4614) );
  NAND4_X1 U5152 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4618)
         );
  NOR2_X1 U5153 ( .A1(n4621), .A2(n4620), .ZN(n4645) );
  XNOR2_X1 U5154 ( .A(n4644), .B(n4645), .ZN(n4622) );
  OR2_X1 U5155 ( .A1(n4747), .A2(n4622), .ZN(n4633) );
  NAND2_X1 U5156 ( .A1(n7200), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4623)
         );
  NAND2_X1 U5157 ( .A1(n4743), .A2(n4623), .ZN(n4624) );
  AOI21_X1 U5158 ( .B1(n4745), .B2(EAX_REG_25__SCAN_IN), .A(n4624), .ZN(n4632)
         );
  INV_X1 U5159 ( .A(n4625), .ZN(n4626) );
  INV_X1 U5160 ( .A(n4627), .ZN(n4629) );
  INV_X1 U5161 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5162 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  NAND2_X1 U5163 ( .A1(n4670), .A2(n4630), .ZN(n6396) );
  NOR2_X1 U5164 ( .A1(n6396), .A2(n4743), .ZN(n4631) );
  AOI21_X1 U5165 ( .B1(n4633), .B2(n4632), .A(n4631), .ZN(n6169) );
  NAND2_X1 U5166 ( .A1(n6168), .A2(n6169), .ZN(n6154) );
  INV_X1 U5167 ( .A(n6154), .ZN(n4653) );
  AOI22_X1 U5168 ( .A1(n4677), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4637) );
  AOI22_X1 U5169 ( .A1(n4700), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5170 ( .A1(n4723), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5171 ( .A1(n4701), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4634) );
  NAND4_X1 U5172 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4643)
         );
  AOI22_X1 U5173 ( .A1(n4722), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5174 ( .A1(n3936), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5175 ( .A1(n4702), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5176 ( .A1(n4731), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4638) );
  NAND4_X1 U5177 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4642)
         );
  NOR2_X1 U5178 ( .A1(n4643), .A2(n4642), .ZN(n4655) );
  NAND2_X1 U5179 ( .A1(n4645), .A2(n4644), .ZN(n4654) );
  XOR2_X1 U5180 ( .A(n4655), .B(n4654), .Z(n4646) );
  NAND2_X1 U5181 ( .A1(n4646), .A2(n4690), .ZN(n4649) );
  INV_X1 U5182 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U5183 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6158), .A(n4743), .ZN(
        n4647) );
  AOI21_X1 U5184 ( .B1(n4745), .B2(EAX_REG_26__SCAN_IN), .A(n4647), .ZN(n4648)
         );
  NAND2_X1 U5185 ( .A1(n4649), .A2(n4648), .ZN(n4651) );
  XNOR2_X1 U5186 ( .A(n4670), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6386)
         );
  NAND2_X1 U5187 ( .A1(n6386), .A2(n4286), .ZN(n4650) );
  NAND2_X1 U5188 ( .A1(n4651), .A2(n4650), .ZN(n6156) );
  NAND2_X1 U5189 ( .A1(n4653), .A2(n4652), .ZN(n6140) );
  NOR2_X1 U5190 ( .A1(n4655), .A2(n4654), .ZN(n4689) );
  AOI22_X1 U5191 ( .A1(n4722), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5192 ( .A1(n4677), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5193 ( .A1(n3936), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5194 ( .A1(n4702), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4656) );
  NAND4_X1 U5195 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4665)
         );
  AOI22_X1 U5196 ( .A1(n4701), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5197 ( .A1(n4700), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5198 ( .A1(n4723), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5199 ( .A1(n3937), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4660) );
  NAND4_X1 U5200 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4664)
         );
  OR2_X1 U5201 ( .A1(n4665), .A2(n4664), .ZN(n4688) );
  INV_X1 U5202 ( .A(n4688), .ZN(n4666) );
  XNOR2_X1 U5203 ( .A(n4689), .B(n4666), .ZN(n4669) );
  NAND2_X1 U5204 ( .A1(n7200), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4667)
         );
  OAI211_X1 U5205 ( .C1(n3659), .C2(n5093), .A(n4743), .B(n4667), .ZN(n4668)
         );
  AOI21_X1 U5206 ( .B1(n4669), .B2(n4690), .A(n4668), .ZN(n4676) );
  INV_X1 U5207 ( .A(n4670), .ZN(n4671) );
  INV_X1 U5208 ( .A(n4672), .ZN(n4673) );
  INV_X1 U5209 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U5210 ( .A1(n4673), .A2(n6147), .ZN(n4674) );
  NAND2_X1 U5211 ( .A1(n4697), .A2(n4674), .ZN(n6380) );
  NOR2_X1 U5212 ( .A1(n6380), .A2(n4743), .ZN(n4675) );
  INV_X1 U5213 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6132) );
  XNOR2_X1 U5214 ( .A(n4697), .B(n6132), .ZN(n6370) );
  INV_X1 U5215 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5216 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n3936), .B1(n4677), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5217 ( .A1(n4723), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5218 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n4700), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5219 ( .A1(n4731), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4678) );
  NAND4_X1 U5220 ( .A1(n4681), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4687)
         );
  AOI22_X1 U5221 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4722), .B1(n4702), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5222 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n4730), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5223 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n4707), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5224 ( .A1(n4701), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4682) );
  NAND4_X1 U5225 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4686)
         );
  NOR2_X1 U5226 ( .A1(n4687), .A2(n4686), .ZN(n4717) );
  NAND2_X1 U5227 ( .A1(n4689), .A2(n4688), .ZN(n4716) );
  XOR2_X1 U5228 ( .A(n4717), .B(n4716), .Z(n4691) );
  NAND2_X1 U5229 ( .A1(n4691), .A2(n4690), .ZN(n4693) );
  AOI21_X1 U5230 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5906), .A(n4286), 
        .ZN(n4692) );
  OAI211_X1 U5231 ( .C1(n3659), .C2(n4694), .A(n4693), .B(n4692), .ZN(n4695)
         );
  OAI21_X1 U5232 ( .B1(n4743), .B2(n6370), .A(n4695), .ZN(n6128) );
  INV_X1 U5233 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U5234 ( .A1(n4698), .A2(n6073), .ZN(n4699) );
  OAI21_X1 U5235 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6073), .A(n4743), .ZN(
        n4720) );
  AOI22_X1 U5236 ( .A1(n4701), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5237 ( .A1(n3936), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5238 ( .A1(n4731), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5239 ( .A1(n4722), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4725), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4703) );
  NAND4_X1 U5240 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4715)
         );
  AOI22_X1 U5241 ( .A1(n4677), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5242 ( .A1(n4723), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5243 ( .A1(n4708), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5244 ( .A1(n4709), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4710) );
  NAND4_X1 U5245 ( .A1(n4713), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4714)
         );
  NOR2_X1 U5246 ( .A1(n4715), .A2(n4714), .ZN(n4739) );
  OR2_X1 U5247 ( .A1(n4717), .A2(n4716), .ZN(n4738) );
  XNOR2_X1 U5248 ( .A(n4739), .B(n4738), .ZN(n4718) );
  NOR2_X1 U5249 ( .A1(n4718), .A2(n4747), .ZN(n4719) );
  AOI211_X1 U5250 ( .C1(n4745), .C2(EAX_REG_29__SCAN_IN), .A(n4720), .B(n4719), 
        .ZN(n4721) );
  AOI21_X1 U5251 ( .B1(n4286), .B2(n6072), .A(n4721), .ZN(n6068) );
  AOI22_X1 U5252 ( .A1(n4723), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5253 ( .A1(n4677), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4708), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5254 ( .A1(n4702), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4593), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U5255 ( .A1(n4725), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4724), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4726) );
  NAND4_X1 U5256 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4737)
         );
  AOI22_X1 U5257 ( .A1(n3936), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5258 ( .A1(n4700), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5259 ( .A1(n4701), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5260 ( .A1(n4731), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4732) );
  NAND4_X1 U5261 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4736)
         );
  NOR2_X1 U5262 ( .A1(n4737), .A2(n4736), .ZN(n4741) );
  NOR2_X1 U5263 ( .A1(n4739), .A2(n4738), .ZN(n4740) );
  XOR2_X1 U5264 ( .A(n4741), .B(n4740), .Z(n4748) );
  NAND2_X1 U5265 ( .A1(n7200), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4742)
         );
  NAND2_X1 U5266 ( .A1(n4743), .A2(n4742), .ZN(n4744) );
  AOI21_X1 U5267 ( .B1(n4745), .B2(EAX_REG_30__SCAN_IN), .A(n4744), .ZN(n4746)
         );
  OAI21_X1 U5268 ( .B1(n4748), .B2(n4747), .A(n4746), .ZN(n4750) );
  XNOR2_X1 U5269 ( .A(n4759), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6105)
         );
  NAND2_X1 U5270 ( .A1(n6105), .A2(n4286), .ZN(n4749) );
  NAND2_X1 U5271 ( .A1(n4750), .A2(n4749), .ZN(n6053) );
  AOI22_X1 U5272 ( .A1(n4745), .A2(EAX_REG_31__SCAN_IN), .B1(n4751), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5273 ( .A1(n4049), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4950) );
  INV_X1 U5274 ( .A(n4950), .ZN(n4774) );
  NAND2_X1 U5275 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4774), .ZN(n7197) );
  INV_X1 U5276 ( .A(n7197), .ZN(n4754) );
  NAND2_X1 U5277 ( .A1(n7587), .A2(n4755), .ZN(n7206) );
  NAND2_X1 U5278 ( .A1(n7206), .A2(n4049), .ZN(n4756) );
  NAND2_X1 U5279 ( .A1(n4049), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4758) );
  NAND2_X1 U5280 ( .A1(n7535), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4757) );
  AND2_X1 U5281 ( .A1(n4758), .A2(n4757), .ZN(n7146) );
  INV_X1 U5282 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6120) );
  XNOR2_X1 U5283 ( .A(n4760), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5734)
         );
  AND2_X2 U5284 ( .A1(n6009), .A2(n4049), .ZN(n7280) );
  AND2_X1 U5285 ( .A1(n7280), .A2(REIP_REG_31__SCAN_IN), .ZN(n6518) );
  AOI21_X1 U5286 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6518), 
        .ZN(n4761) );
  OAI21_X1 U5287 ( .B1(n7190), .B2(n5734), .A(n4761), .ZN(n4762) );
  AOI21_X1 U5288 ( .B1(n6062), .B2(n7185), .A(n4762), .ZN(n4763) );
  NAND3_X1 U5289 ( .A1(n4768), .A2(n4767), .A3(n4766), .ZN(n4770) );
  AOI21_X1 U5290 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n6110) );
  INV_X1 U5291 ( .A(n6110), .ZN(n4773) );
  NAND2_X1 U5292 ( .A1(n4773), .A2(n4772), .ZN(n4892) );
  INV_X1 U5293 ( .A(n7522), .ZN(n6986) );
  AND2_X1 U5294 ( .A1(n4286), .A2(n4774), .ZN(n7524) );
  NAND2_X1 U5295 ( .A1(n7200), .A2(n6667), .ZN(n7203) );
  NOR3_X1 U5296 ( .A1(n4049), .A2(n7533), .A3(n7203), .ZN(n6993) );
  NOR2_X1 U5297 ( .A1(n5734), .A2(n6667), .ZN(n4776) );
  NAND2_X1 U5298 ( .A1(n6062), .A2(n7496), .ZN(n4891) );
  NAND2_X1 U5299 ( .A1(n5196), .A2(n3645), .ZN(n4780) );
  INV_X1 U5300 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5301 ( .A1(n4792), .A2(n4779), .B1(n4789), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4978) );
  INV_X1 U5302 ( .A(n4865), .ZN(n4817) );
  INV_X1 U5303 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U5304 ( .A1(n4817), .A2(n7129), .ZN(n4783) );
  NAND2_X1 U5305 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4781)
         );
  OAI211_X1 U5306 ( .C1(n4975), .C2(EBX_REG_2__SCAN_IN), .A(n4792), .B(n4781), 
        .ZN(n4782) );
  AND2_X1 U5307 ( .A1(n4783), .A2(n4782), .ZN(n6086) );
  NAND2_X1 U5308 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  INV_X1 U5309 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5310 ( .A1(n4870), .A2(n4784), .ZN(n4788) );
  NAND2_X1 U5311 ( .A1(n4792), .A2(n5039), .ZN(n4786) );
  NAND2_X1 U5312 ( .A1(n4969), .A2(n4784), .ZN(n4785) );
  NAND3_X1 U5313 ( .A1(n4786), .A2(n4789), .A3(n4785), .ZN(n4787) );
  AND2_X1 U5314 ( .A1(n4788), .A2(n4787), .ZN(n5025) );
  NAND2_X1 U5315 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4790)
         );
  OAI211_X1 U5316 ( .C1(n4975), .C2(EBX_REG_4__SCAN_IN), .A(n4792), .B(n4790), 
        .ZN(n4791) );
  OAI21_X1 U5317 ( .B1(n4865), .B2(EBX_REG_4__SCAN_IN), .A(n4791), .ZN(n7135)
         );
  MUX2_X1 U5318 ( .A(n4860), .B(n4792), .S(EBX_REG_5__SCAN_IN), .Z(n4796) );
  INV_X1 U5319 ( .A(n4792), .ZN(n4793) );
  NAND2_X1 U5320 ( .A1(n4793), .A2(n4975), .ZN(n4840) );
  NAND2_X1 U5321 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4975), .ZN(n4794)
         );
  AND2_X1 U5322 ( .A1(n4840), .A2(n4794), .ZN(n4795) );
  MUX2_X1 U5323 ( .A(n4865), .B(n4789), .S(EBX_REG_6__SCAN_IN), .Z(n4797) );
  OAI21_X1 U5324 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4977), .A(n4797), 
        .ZN(n5780) );
  NOR2_X1 U5325 ( .A1(n5778), .A2(n5780), .ZN(n4798) );
  MUX2_X1 U5326 ( .A(n4860), .B(n4792), .S(EBX_REG_7__SCAN_IN), .Z(n4800) );
  NAND2_X1 U5327 ( .A1(n4975), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4799)
         );
  NAND2_X1 U5328 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4801)
         );
  OAI211_X1 U5329 ( .C1(n4975), .C2(EBX_REG_8__SCAN_IN), .A(n4792), .B(n4801), 
        .ZN(n4802) );
  OAI21_X1 U5330 ( .B1(n4865), .B2(EBX_REG_8__SCAN_IN), .A(n4802), .ZN(n5995)
         );
  OR2_X1 U5331 ( .A1(n4860), .A2(EBX_REG_9__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U5332 ( .A1(n4792), .A2(n7265), .ZN(n4805) );
  INV_X1 U5333 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U5334 ( .A1(n4969), .A2(n4803), .ZN(n4804) );
  NAND3_X1 U5335 ( .A1(n4805), .A2(n4789), .A3(n4804), .ZN(n4806) );
  NAND2_X1 U5336 ( .A1(n4807), .A2(n4806), .ZN(n5948) );
  INV_X1 U5337 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U5338 ( .A1(n4817), .A2(n6249), .ZN(n4810) );
  NAND2_X1 U5339 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4808) );
  OAI211_X1 U5340 ( .C1(n4975), .C2(EBX_REG_10__SCAN_IN), .A(n4792), .B(n4808), 
        .ZN(n4809) );
  AND2_X1 U5341 ( .A1(n4810), .A2(n4809), .ZN(n5978) );
  NAND2_X1 U5342 ( .A1(n5979), .A2(n5978), .ZN(n5977) );
  INV_X1 U5343 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U5344 ( .A1(n4870), .A2(n6008), .ZN(n4814) );
  NAND2_X1 U5345 ( .A1(n4792), .A2(n6484), .ZN(n4812) );
  NAND2_X1 U5346 ( .A1(n4969), .A2(n6008), .ZN(n4811) );
  NAND3_X1 U5347 ( .A1(n4812), .A2(n4789), .A3(n4811), .ZN(n4813) );
  NAND2_X1 U5348 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4815) );
  OAI211_X1 U5349 ( .C1(n4975), .C2(EBX_REG_12__SCAN_IN), .A(n4792), .B(n4815), 
        .ZN(n4816) );
  OAI21_X1 U5350 ( .B1(n4865), .B2(EBX_REG_12__SCAN_IN), .A(n4816), .ZN(n6022)
         );
  INV_X1 U5351 ( .A(EBX_REG_14__SCAN_IN), .ZN(n7413) );
  NAND2_X1 U5352 ( .A1(n4817), .A2(n7413), .ZN(n4820) );
  NAND2_X1 U5353 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4818) );
  OAI211_X1 U5354 ( .C1(n4975), .C2(EBX_REG_14__SCAN_IN), .A(n4792), .B(n4818), 
        .ZN(n4819) );
  AND2_X1 U5355 ( .A1(n4820), .A2(n4819), .ZN(n6638) );
  OR2_X1 U5356 ( .A1(n4860), .A2(EBX_REG_13__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U5357 ( .A1(n4792), .A2(n4821), .ZN(n4823) );
  INV_X1 U5358 ( .A(EBX_REG_13__SCAN_IN), .ZN(n7396) );
  NAND2_X1 U5359 ( .A1(n4969), .A2(n7396), .ZN(n4822) );
  NAND3_X1 U5360 ( .A1(n4823), .A2(n4789), .A3(n4822), .ZN(n4824) );
  NAND2_X1 U5361 ( .A1(n4825), .A2(n4824), .ZN(n6646) );
  NAND2_X1 U5362 ( .A1(n6638), .A2(n6646), .ZN(n4826) );
  OR2_X1 U5363 ( .A1(n4860), .A2(EBX_REG_15__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U5364 ( .A1(n4792), .A2(n7285), .ZN(n4829) );
  INV_X1 U5365 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4827) );
  NAND2_X1 U5366 ( .A1(n4969), .A2(n4827), .ZN(n4828) );
  NAND3_X1 U5367 ( .A1(n4829), .A2(n4789), .A3(n4828), .ZN(n4830) );
  NAND2_X1 U5368 ( .A1(n4831), .A2(n4830), .ZN(n6311) );
  NAND2_X1 U5369 ( .A1(n6640), .A2(n6311), .ZN(n6313) );
  NAND2_X1 U5370 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4832) );
  OAI211_X1 U5371 ( .C1(n4975), .C2(EBX_REG_16__SCAN_IN), .A(n4792), .B(n4832), 
        .ZN(n4833) );
  OAI21_X1 U5372 ( .B1(n4865), .B2(EBX_REG_16__SCAN_IN), .A(n4833), .ZN(n6231)
         );
  MUX2_X1 U5373 ( .A(n4860), .B(n4792), .S(EBX_REG_17__SCAN_IN), .Z(n4835) );
  NAND2_X1 U5374 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n4975), .ZN(n4834) );
  MUX2_X1 U5375 ( .A(n4865), .B(n4789), .S(EBX_REG_18__SCAN_IN), .Z(n4837) );
  OR2_X1 U5376 ( .A1(n4977), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4836)
         );
  NAND2_X1 U5377 ( .A1(n4837), .A2(n4836), .ZN(n6222) );
  INV_X1 U5378 ( .A(n6222), .ZN(n4838) );
  MUX2_X1 U5379 ( .A(n4860), .B(n4792), .S(EBX_REG_19__SCAN_IN), .Z(n4842) );
  NAND2_X1 U5380 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n4975), .ZN(n4839) );
  AND2_X1 U5381 ( .A1(n4840), .A2(n4839), .ZN(n4841) );
  NAND2_X1 U5382 ( .A1(n4842), .A2(n4841), .ZN(n6296) );
  NAND2_X1 U5383 ( .A1(n6221), .A2(n6296), .ZN(n6295) );
  NAND2_X1 U5384 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4843) );
  OAI211_X1 U5385 ( .C1(n4975), .C2(EBX_REG_20__SCAN_IN), .A(n4792), .B(n4843), 
        .ZN(n4844) );
  OAI21_X1 U5386 ( .B1(n4865), .B2(EBX_REG_20__SCAN_IN), .A(n4844), .ZN(n6202)
         );
  INV_X1 U5387 ( .A(EBX_REG_21__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U5388 ( .A1(n4870), .A2(n4845), .ZN(n4849) );
  INV_X1 U5389 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U5390 ( .A1(n4792), .A2(n6609), .ZN(n4847) );
  NAND2_X1 U5391 ( .A1(n4969), .A2(n4845), .ZN(n4846) );
  NAND3_X1 U5392 ( .A1(n4847), .A2(n4789), .A3(n4846), .ZN(n4848) );
  MUX2_X1 U5393 ( .A(n4865), .B(n4789), .S(EBX_REG_22__SCAN_IN), .Z(n4851) );
  INV_X1 U5394 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6594) );
  INV_X1 U5395 ( .A(n4977), .ZN(n4868) );
  NAND2_X1 U5396 ( .A1(n6594), .A2(n4868), .ZN(n4850) );
  MUX2_X1 U5397 ( .A(n4860), .B(n4792), .S(EBX_REG_23__SCAN_IN), .Z(n4853) );
  NAND2_X1 U5398 ( .A1(n4975), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5399 ( .A1(n4853), .A2(n4852), .ZN(n6275) );
  MUX2_X1 U5400 ( .A(n4865), .B(n4789), .S(EBX_REG_24__SCAN_IN), .Z(n4854) );
  OAI21_X1 U5401 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n4977), .A(n4854), 
        .ZN(n6185) );
  OR2_X1 U5402 ( .A1(n4860), .A2(EBX_REG_25__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5403 ( .A1(n4792), .A2(n6573), .ZN(n4855) );
  OAI211_X1 U5404 ( .C1(EBX_REG_25__SCAN_IN), .C2(n4975), .A(n4855), .B(n4789), 
        .ZN(n4856) );
  NAND2_X1 U5405 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4858) );
  OAI211_X1 U5406 ( .C1(n4975), .C2(EBX_REG_26__SCAN_IN), .A(n4792), .B(n4858), 
        .ZN(n4859) );
  OAI21_X1 U5407 ( .B1(n4865), .B2(EBX_REG_26__SCAN_IN), .A(n4859), .ZN(n6165)
         );
  MUX2_X1 U5408 ( .A(n4860), .B(n4792), .S(EBX_REG_27__SCAN_IN), .Z(n4862) );
  NAND2_X1 U5409 ( .A1(n4975), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5410 ( .A1(n4862), .A2(n4861), .ZN(n6144) );
  NAND2_X1 U5411 ( .A1(n4789), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4863) );
  OAI211_X1 U5412 ( .C1(n4975), .C2(EBX_REG_28__SCAN_IN), .A(n4792), .B(n4863), 
        .ZN(n4864) );
  OAI21_X1 U5413 ( .B1(n4865), .B2(EBX_REG_28__SCAN_IN), .A(n4864), .ZN(n6129)
         );
  NOR2_X1 U5414 ( .A1(n4975), .A2(EBX_REG_29__SCAN_IN), .ZN(n4866) );
  AOI21_X1 U5415 ( .B1(n4868), .B2(n4867), .A(n4866), .ZN(n6055) );
  INV_X1 U5416 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4869) );
  AOI22_X1 U5417 ( .A1(n6055), .A2(n4789), .B1(n4870), .B2(n4869), .ZN(n6070)
         );
  AND2_X1 U5418 ( .A1(n4975), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4871)
         );
  AOI21_X1 U5419 ( .B1(n4977), .B2(EBX_REG_30__SCAN_IN), .A(n4871), .ZN(n6058)
         );
  AOI22_X1 U5420 ( .A1(n4977), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4975), .ZN(n4874) );
  XNOR2_X2 U5421 ( .A(n4875), .B(n4874), .ZN(n6496) );
  INV_X1 U5422 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6260) );
  NOR2_X1 U5423 ( .A1(n5744), .A2(n6260), .ZN(n4882) );
  NOR2_X1 U5424 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4883) );
  NOR2_X1 U5425 ( .A1(n4975), .A2(n4883), .ZN(n4876) );
  INV_X1 U5426 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7096) );
  INV_X1 U5427 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7094) );
  NOR2_X1 U5428 ( .A1(n7096), .A2(n7094), .ZN(n4881) );
  NAND2_X1 U5429 ( .A1(n4877), .A2(n7547), .ZN(n7194) );
  NAND2_X1 U5430 ( .A1(n3907), .A2(n7194), .ZN(n4993) );
  AND3_X1 U5431 ( .A1(n4993), .A2(n4883), .A3(n3645), .ZN(n4878) );
  NAND2_X1 U5432 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4880) );
  INV_X1 U5433 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7086) );
  INV_X1 U5434 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7482) );
  INV_X1 U5435 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7082) );
  INV_X1 U5436 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7078) );
  NAND3_X1 U5437 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n7331) );
  INV_X1 U5438 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7328) );
  NOR2_X1 U5439 ( .A1(n7331), .A2(n7328), .ZN(n6241) );
  NAND2_X1 U5440 ( .A1(n6241), .A2(REIP_REG_5__SCAN_IN), .ZN(n6244) );
  NAND3_X1 U5441 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .ZN(n6243) );
  INV_X1 U5442 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7061) );
  NOR3_X1 U5443 ( .A1(n6244), .A2(n6243), .A3(n7061), .ZN(n6252) );
  NAND2_X1 U5444 ( .A1(n6252), .A2(REIP_REG_10__SCAN_IN), .ZN(n6018) );
  INV_X1 U5445 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7064) );
  NOR2_X1 U5446 ( .A1(n6018), .A2(n7064), .ZN(n6007) );
  NAND4_X1 U5447 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .A4(n6007), .ZN(n6213) );
  NAND3_X1 U5448 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n6212) );
  INV_X1 U5449 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7074) );
  NOR2_X1 U5450 ( .A1(n6212), .A2(n7074), .ZN(n7447) );
  NAND2_X1 U5451 ( .A1(n7447), .A2(REIP_REG_19__SCAN_IN), .ZN(n6199) );
  NOR3_X1 U5452 ( .A1(n7078), .A2(n6213), .A3(n6199), .ZN(n7461) );
  NAND2_X1 U5453 ( .A1(REIP_REG_21__SCAN_IN), .A2(n7461), .ZN(n7472) );
  NOR3_X1 U5454 ( .A1(n7482), .A2(n7082), .A3(n7472), .ZN(n6186) );
  NAND2_X1 U5455 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6186), .ZN(n6174) );
  NOR2_X1 U5456 ( .A1(n7086), .A2(n6174), .ZN(n6173) );
  AND2_X1 U5457 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6173), .ZN(n4879) );
  NAND2_X1 U5458 ( .A1(n6215), .A2(n4879), .ZN(n6160) );
  NAND2_X1 U5459 ( .A1(n7473), .A2(n6215), .ZN(n6217) );
  OAI21_X1 U5460 ( .B1(n4880), .B2(n6160), .A(n6217), .ZN(n6137) );
  OAI21_X1 U5461 ( .B1(n4881), .B2(n7473), .A(n6137), .ZN(n6125) );
  INV_X1 U5462 ( .A(n4882), .ZN(n4885) );
  INV_X1 U5463 ( .A(n4883), .ZN(n5740) );
  OR2_X1 U5464 ( .A1(n7194), .A2(n5740), .ZN(n6987) );
  NAND2_X1 U5465 ( .A1(n3992), .A2(n6987), .ZN(n5742) );
  INV_X1 U5466 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4884) );
  OAI22_X1 U5467 ( .A1(n4885), .A2(n5742), .B1(n4884), .B2(n7478), .ZN(n4887)
         );
  NAND2_X1 U5468 ( .A1(n7333), .A2(n6173), .ZN(n6159) );
  INV_X1 U5469 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7090) );
  INV_X1 U5470 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7088) );
  NOR3_X1 U5471 ( .A1(n6159), .A2(n7090), .A3(n7088), .ZN(n6135) );
  NAND3_X1 U5472 ( .A1(n6135), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n6123) );
  NOR3_X1 U5473 ( .A1(n6123), .A2(REIP_REG_31__SCAN_IN), .A3(n7096), .ZN(n4886) );
  AOI211_X1 U5474 ( .C1(REIP_REG_31__SCAN_IN), .C2(n6125), .A(n4887), .B(n4886), .ZN(n4888) );
  NAND2_X1 U5475 ( .A1(n4891), .A2(n4890), .ZN(U2796) );
  INV_X1 U5476 ( .A(n7523), .ZN(n4895) );
  NAND2_X1 U5477 ( .A1(n4764), .A2(n4892), .ZN(n4893) );
  OAI21_X1 U5478 ( .B1(n6115), .B2(n3925), .A(n4893), .ZN(n6118) );
  OAI21_X1 U5479 ( .B1(n6118), .B2(n6986), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4894) );
  OAI21_X1 U5480 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4895), .A(n4894), .ZN(
        U2790) );
  INV_X1 U5481 ( .A(n4896), .ZN(n4898) );
  INV_X1 U5482 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7555) );
  INV_X1 U5483 ( .A(n6009), .ZN(n4897) );
  OAI211_X1 U5484 ( .C1(n4898), .C2(n7555), .A(n5195), .B(n4897), .ZN(U2788)
         );
  INV_X1 U5485 ( .A(n7205), .ZN(n4900) );
  NAND2_X1 U5486 ( .A1(n3905), .A2(n5196), .ZN(n4914) );
  INV_X1 U5487 ( .A(n4914), .ZN(n5732) );
  OR2_X1 U5488 ( .A1(n3992), .A2(n5732), .ZN(n6116) );
  OAI21_X1 U5489 ( .B1(n6009), .B2(READREQUEST_REG_SCAN_IN), .A(n4900), .ZN(
        n4899) );
  OAI21_X1 U5490 ( .B1(n4900), .B2(n6116), .A(n4899), .ZN(U3474) );
  INV_X1 U5491 ( .A(n3925), .ZN(n4901) );
  NOR2_X1 U5492 ( .A1(n4437), .A2(n4901), .ZN(n4902) );
  NAND2_X1 U5493 ( .A1(n6115), .A2(n5010), .ZN(n4906) );
  INV_X1 U5494 ( .A(n5228), .ZN(n4921) );
  OR2_X1 U5495 ( .A1(n4764), .A2(n3907), .ZN(n5012) );
  OAI21_X1 U5496 ( .B1(n6958), .B2(n4907), .A(n7546), .ZN(n4908) );
  AOI21_X1 U5497 ( .B1(n7194), .B2(n5012), .A(n4908), .ZN(n4916) );
  AOI21_X1 U5498 ( .B1(n3645), .B2(n3637), .A(n3992), .ZN(n4909) );
  OR2_X1 U5499 ( .A1(n3929), .A2(n4909), .ZN(n4932) );
  NAND2_X1 U5500 ( .A1(n4437), .A2(n3905), .ZN(n4910) );
  NAND3_X1 U5501 ( .A1(n4932), .A2(n4911), .A3(n4910), .ZN(n4913) );
  INV_X1 U5502 ( .A(n4772), .ZN(n4912) );
  NAND2_X1 U5503 ( .A1(n4913), .A2(n4912), .ZN(n4990) );
  OAI21_X1 U5504 ( .B1(n4986), .B2(n4914), .A(n4990), .ZN(n4915) );
  AOI21_X1 U5505 ( .B1(n6115), .B2(n4916), .A(n4915), .ZN(n4920) );
  INV_X1 U5506 ( .A(n6115), .ZN(n4919) );
  NAND2_X1 U5507 ( .A1(n4984), .A2(n3645), .ZN(n4917) );
  NOR2_X1 U5508 ( .A1(n4917), .A2(n4926), .ZN(n4918) );
  NAND2_X1 U5509 ( .A1(n4919), .A2(n6111), .ZN(n4972) );
  NAND3_X1 U5510 ( .A1(n4921), .A2(n4920), .A3(n4972), .ZN(n6962) );
  NAND2_X1 U5511 ( .A1(n6962), .A2(n7522), .ZN(n4923) );
  NAND2_X1 U5512 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7526), .ZN(n7531) );
  INV_X1 U5513 ( .A(n7531), .ZN(n7199) );
  NAND2_X1 U5514 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7199), .ZN(n4922) );
  NAND2_X1 U5515 ( .A1(n4923), .A2(n4922), .ZN(n7518) );
  AND2_X1 U5516 ( .A1(n4049), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U5517 ( .A1(n4926), .A2(n3908), .ZN(n4927) );
  OAI211_X1 U5518 ( .C1(n4928), .C2(n3907), .A(n4927), .B(n4792), .ZN(n4930)
         );
  NOR2_X1 U5519 ( .A1(n4930), .A2(n4929), .ZN(n4931) );
  NAND2_X1 U5520 ( .A1(n4932), .A2(n4931), .ZN(n4933) );
  NOR2_X1 U5521 ( .A1(n4934), .A2(n4933), .ZN(n5002) );
  NAND3_X1 U5522 ( .A1(n4904), .A2(n4935), .A3(n4936), .ZN(n4937) );
  NOR2_X1 U5523 ( .A1(n4937), .A2(n4907), .ZN(n4938) );
  AND2_X1 U5524 ( .A1(n5002), .A2(n4938), .ZN(n5267) );
  OR2_X1 U5525 ( .A1(n6090), .A2(n5267), .ZN(n4943) );
  OR2_X1 U5526 ( .A1(n5010), .A2(n6111), .ZN(n5271) );
  INV_X1 U5527 ( .A(n4939), .ZN(n4944) );
  NAND2_X1 U5528 ( .A1(n4944), .A2(n3750), .ZN(n5269) );
  NAND2_X1 U5529 ( .A1(n4939), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U5530 ( .A1(n5269), .A2(n7504), .ZN(n4941) );
  XNOR2_X1 U5531 ( .A(n3750), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4940)
         );
  AOI22_X1 U5532 ( .A1(n5271), .A2(n4941), .B1(n6958), .B2(n4940), .ZN(n4942)
         );
  NAND2_X1 U5533 ( .A1(n4943), .A2(n4942), .ZN(n5264) );
  INV_X1 U5534 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U5535 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6512), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5138), .ZN(n6669) );
  NOR3_X1 U5536 ( .A1(n6667), .A2(n6666), .A3(n6669), .ZN(n4946) );
  NOR3_X1 U5537 ( .A1(n4944), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7505), 
        .ZN(n4945) );
  AOI211_X1 U5538 ( .C1(n5264), .C2(n7517), .A(n4946), .B(n4945), .ZN(n4948)
         );
  NOR2_X1 U5539 ( .A1(n4939), .A2(n7505), .ZN(n6671) );
  OAI21_X1 U5540 ( .B1(n7512), .B2(n6671), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4947) );
  OAI21_X1 U5541 ( .B1(n7512), .B2(n4948), .A(n4947), .ZN(U3459) );
  INV_X1 U5542 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4952) );
  INV_X1 U5543 ( .A(n6958), .ZN(n6661) );
  AOI21_X1 U5544 ( .B1(n6661), .B2(n6988), .A(n7194), .ZN(n4949) );
  NAND2_X1 U5545 ( .A1(n7019), .A2(n3645), .ZN(n5096) );
  INV_X2 U5546 ( .A(n6985), .ZN(n7048) );
  NOR2_X4 U5547 ( .A1(n7048), .A2(n7019), .ZN(n7031) );
  AOI22_X1 U5548 ( .A1(n7048), .A2(UWORD_REG_6__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4951) );
  OAI21_X1 U5549 ( .B1(n4952), .B2(n5096), .A(n4951), .ZN(U2901) );
  INV_X1 U5550 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5551 ( .A1(n7048), .A2(UWORD_REG_7__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4953) );
  OAI21_X1 U5552 ( .B1(n4954), .B2(n5096), .A(n4953), .ZN(U2900) );
  INV_X1 U5553 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U5554 ( .A1(n7048), .A2(UWORD_REG_5__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4955) );
  OAI21_X1 U5555 ( .B1(n4956), .B2(n5096), .A(n4955), .ZN(U2902) );
  INV_X1 U5556 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U5557 ( .A1(n7048), .A2(UWORD_REG_8__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U5558 ( .B1(n4958), .B2(n5096), .A(n4957), .ZN(U2899) );
  INV_X1 U5559 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U5560 ( .A1(n7048), .A2(UWORD_REG_9__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4959) );
  OAI21_X1 U5561 ( .B1(n4960), .B2(n5096), .A(n4959), .ZN(U2898) );
  AOI21_X1 U5562 ( .B1(n6958), .B2(n7517), .A(n7512), .ZN(n4963) );
  OAI22_X1 U5563 ( .A1(n4267), .A2(n5267), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4437), .ZN(n6961) );
  OAI22_X1 U5564 ( .A1(n6667), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7505), .ZN(n4961) );
  AOI21_X1 U5565 ( .B1(n6961), .B2(n7517), .A(n4961), .ZN(n4962) );
  OAI22_X1 U5566 ( .A1(n4963), .A2(n3752), .B1(n7512), .B2(n4962), .ZN(U3461)
         );
  OAI21_X1 U5567 ( .B1(n4964), .B2(n4966), .A(n4965), .ZN(n5987) );
  INV_X1 U5568 ( .A(n3900), .ZN(n6060) );
  NAND3_X1 U5569 ( .A1(n3920), .A2(n6060), .A3(n4967), .ZN(n5226) );
  INV_X1 U5570 ( .A(n5226), .ZN(n4968) );
  NAND3_X1 U5571 ( .A1(n4970), .A2(n4969), .A3(n4968), .ZN(n4971) );
  NAND2_X1 U5572 ( .A1(n4972), .A2(n4971), .ZN(n4973) );
  NAND2_X2 U5573 ( .A1(n7143), .A2(n3900), .ZN(n7127) );
  INV_X1 U5574 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4976) );
  XNOR2_X1 U5575 ( .A(n4974), .B(n4975), .ZN(n5142) );
  OAI222_X1 U5576 ( .A1(n5987), .A2(n7127), .B1(n4976), .B2(n7143), .C1(n5142), 
        .C2(n6304), .ZN(U2858) );
  NOR2_X1 U5577 ( .A1(n4977), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4979)
         );
  OR2_X1 U5578 ( .A1(n4979), .A2(n4978), .ZN(n7320) );
  INV_X1 U5579 ( .A(n4980), .ZN(n4982) );
  MUX2_X1 U5580 ( .A(n4983), .B(n4982), .S(n4981), .Z(n7323) );
  INV_X1 U5581 ( .A(n7323), .ZN(n5232) );
  OAI222_X1 U5582 ( .A1(n6304), .A2(n7320), .B1(n4779), .B2(n7143), .C1(n7127), 
        .C2(n5232), .ZN(U2859) );
  NAND2_X1 U5583 ( .A1(n4985), .A2(n4984), .ZN(n4991) );
  INV_X1 U5584 ( .A(n7194), .ZN(n4987) );
  OAI211_X1 U5585 ( .C1(n3907), .C2(n4987), .A(n4986), .B(n7546), .ZN(n4988)
         );
  OR2_X1 U5586 ( .A1(n6110), .A2(n4988), .ZN(n4989) );
  OAI211_X1 U5587 ( .C1(n6115), .C2(n4991), .A(n4990), .B(n4989), .ZN(n4992)
         );
  NAND2_X1 U5588 ( .A1(n4992), .A2(n7522), .ZN(n4999) );
  NAND3_X1 U5589 ( .A1(n4907), .A2(n4993), .A3(n7546), .ZN(n4996) );
  NAND2_X1 U5590 ( .A1(n3908), .A2(n3645), .ZN(n4994) );
  NAND2_X1 U5591 ( .A1(n4994), .A2(n5073), .ZN(n4995) );
  NAND2_X1 U5592 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  NAND2_X1 U5593 ( .A1(n5197), .A2(n4997), .ZN(n4998) );
  OAI21_X1 U5594 ( .B1(n3646), .B2(n5000), .A(n6988), .ZN(n5001) );
  OAI21_X1 U5595 ( .B1(n5004), .B2(n5003), .A(n5002), .ZN(n5005) );
  NAND2_X1 U5596 ( .A1(n5014), .A2(n5005), .ZN(n5037) );
  NOR2_X1 U5597 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5037), .ZN(n5006)
         );
  AOI21_X1 U5598 ( .B1(n5007), .B2(n7248), .A(n5006), .ZN(n7300) );
  OAI21_X1 U5599 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n7252), .A(n7300), 
        .ZN(n5137) );
  NAND2_X1 U5600 ( .A1(n5014), .A2(n6958), .ZN(n5036) );
  INV_X1 U5601 ( .A(n5036), .ZN(n5009) );
  NAND3_X1 U5602 ( .A1(n6666), .A2(n7252), .A3(n5037), .ZN(n5008) );
  OAI21_X1 U5603 ( .B1(n5137), .B2(n5009), .A(n5008), .ZN(n5019) );
  NOR2_X1 U5604 ( .A1(n5010), .A2(n6975), .ZN(n6109) );
  OR2_X1 U5605 ( .A1(n3646), .A2(n3920), .ZN(n5011) );
  NAND4_X1 U5606 ( .A1(n6109), .A2(n5012), .A3(n4904), .A4(n5011), .ZN(n5013)
         );
  OAI21_X1 U5607 ( .B1(n5015), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5136), 
        .ZN(n7144) );
  INV_X1 U5608 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5016) );
  OAI22_X1 U5609 ( .A1(n7240), .A2(n7144), .B1(n7248), .B2(n5016), .ZN(n5017)
         );
  INV_X1 U5610 ( .A(n5017), .ZN(n5018) );
  OAI211_X1 U5611 ( .C1(n7301), .C2(n7320), .A(n5019), .B(n5018), .ZN(U3018)
         );
  AOI21_X1 U5612 ( .B1(n5023), .B2(n5020), .A(n5022), .ZN(n5966) );
  INV_X1 U5613 ( .A(n5966), .ZN(n5944) );
  INV_X1 U5614 ( .A(n7136), .ZN(n5024) );
  AOI21_X1 U5615 ( .B1(n5025), .B2(n6088), .A(n5024), .ZN(n5941) );
  AOI22_X1 U5616 ( .A1(n7139), .A2(n5941), .B1(EBX_REG_3__SCAN_IN), .B2(n6314), 
        .ZN(n5026) );
  OAI21_X1 U5617 ( .B1(n5944), .B2(n7127), .A(n5026), .ZN(U2856) );
  NAND2_X1 U5618 ( .A1(n5029), .A2(n5030), .ZN(n5031) );
  NAND2_X1 U5619 ( .A1(n5028), .A2(n5031), .ZN(n7341) );
  INV_X1 U5620 ( .A(EBX_REG_5__SCAN_IN), .ZN(n5032) );
  XNOR2_X1 U5621 ( .A(n7138), .B(n5778), .ZN(n7342) );
  INV_X1 U5622 ( .A(n7342), .ZN(n7239) );
  OAI222_X1 U5623 ( .A1(n7341), .A2(n7127), .B1(n5032), .B2(n7143), .C1(n6304), 
        .C2(n7239), .ZN(U2854) );
  XNOR2_X1 U5624 ( .A(n5034), .B(n5039), .ZN(n5035) );
  XNOR2_X1 U5625 ( .A(n5033), .B(n5035), .ZN(n5968) );
  AOI21_X1 U5626 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5954) );
  NAND2_X1 U5627 ( .A1(n5036), .A2(n6666), .ZN(n5139) );
  INV_X1 U5628 ( .A(n5139), .ZN(n5038) );
  NAND2_X1 U5629 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5955) );
  INV_X1 U5630 ( .A(n5955), .ZN(n7255) );
  AOI21_X1 U5631 ( .B1(n7260), .B2(n7255), .A(n7298), .ZN(n7230) );
  NOR2_X1 U5632 ( .A1(n5954), .A2(n7230), .ZN(n7219) );
  NAND2_X1 U5633 ( .A1(n7219), .A2(n5039), .ZN(n5043) );
  NAND2_X1 U5634 ( .A1(n7298), .A2(n5954), .ZN(n7262) );
  OAI211_X1 U5635 ( .C1(n7256), .C2(n7255), .A(n7300), .B(n7262), .ZN(n7224)
         );
  INV_X1 U5636 ( .A(n5941), .ZN(n5040) );
  INV_X1 U5637 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7054) );
  OAI22_X1 U5638 ( .A1(n7301), .A2(n5040), .B1(n7054), .B2(n7248), .ZN(n5041)
         );
  AOI21_X1 U5639 ( .B1(n7224), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5041), 
        .ZN(n5042) );
  OAI211_X1 U5640 ( .C1(n5968), .C2(n7240), .A(n5043), .B(n5042), .ZN(U3015)
         );
  INV_X1 U5641 ( .A(n7203), .ZN(n5044) );
  INV_X1 U5642 ( .A(n4267), .ZN(n5905) );
  AND2_X1 U5643 ( .A1(n6703), .A2(n5905), .ZN(n5680) );
  INV_X1 U5644 ( .A(n7590), .ZN(n5049) );
  INV_X1 U5645 ( .A(n5048), .ZN(n6950) );
  AOI21_X1 U5646 ( .B1(n5680), .B2(n5049), .A(n6950), .ZN(n5056) );
  NOR2_X1 U5647 ( .A1(n5050), .A2(n5051), .ZN(n5146) );
  NAND2_X1 U5648 ( .A1(n5146), .A2(n5052), .ZN(n5058) );
  INV_X1 U5649 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U5650 ( .A1(n7599), .A2(n7535), .ZN(n6853) );
  OAI21_X1 U5651 ( .B1(n5059), .B2(n7174), .A(n6853), .ZN(n5053) );
  NAND3_X1 U5652 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5708) );
  AOI22_X1 U5653 ( .A1(n5056), .A2(n5053), .B1(n7587), .B2(n5708), .ZN(n5054)
         );
  INV_X1 U5654 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5062) );
  NOR2_X2 U5655 ( .A1(n6678), .A2(n4262), .ZN(n7640) );
  INV_X1 U5656 ( .A(DATAI_6_), .ZN(n5787) );
  NOR2_X2 U5657 ( .A1(n5787), .A2(n6679), .ZN(n6820) );
  OAI22_X1 U5658 ( .A1(n5056), .A2(n7587), .B1(n5708), .B2(n5906), .ZN(n6948)
         );
  AOI22_X1 U5659 ( .A1(n7640), .A2(n6950), .B1(n6820), .B2(n6948), .ZN(n5061)
         );
  NAND2_X1 U5660 ( .A1(n7185), .A2(DATAI_30_), .ZN(n6742) );
  INV_X1 U5661 ( .A(n6742), .ZN(n7642) );
  AOI22_X1 U5662 ( .A1(n7641), .A2(n6952), .B1(n6951), .B2(n7642), .ZN(n5060)
         );
  OAI211_X1 U5663 ( .C1(n6956), .C2(n5062), .A(n5061), .B(n5060), .ZN(U3146)
         );
  INV_X1 U5664 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5065) );
  NOR2_X2 U5665 ( .A1(n6678), .A2(n6317), .ZN(n7634) );
  INV_X1 U5666 ( .A(DATAI_5_), .ZN(n5238) );
  NOR2_X2 U5667 ( .A1(n5238), .A2(n6679), .ZN(n6816) );
  AOI22_X1 U5668 ( .A1(n7634), .A2(n6950), .B1(n6816), .B2(n6948), .ZN(n5064)
         );
  NAND2_X1 U5669 ( .A1(n7185), .A2(DATAI_29_), .ZN(n6737) );
  INV_X1 U5670 ( .A(n6737), .ZN(n7636) );
  AOI22_X1 U5671 ( .A1(n7635), .A2(n6952), .B1(n6951), .B2(n7636), .ZN(n5063)
         );
  OAI211_X1 U5672 ( .C1(n6956), .C2(n5065), .A(n5064), .B(n5063), .ZN(U3145)
         );
  INV_X1 U5673 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5068) );
  NOR2_X2 U5674 ( .A1(n6678), .A2(n6060), .ZN(n7647) );
  INV_X1 U5675 ( .A(DATAI_7_), .ZN(n5704) );
  NOR2_X2 U5676 ( .A1(n5704), .A2(n6679), .ZN(n6825) );
  AOI22_X1 U5677 ( .A1(n7647), .A2(n6950), .B1(n6825), .B2(n6948), .ZN(n5067)
         );
  NAND2_X1 U5678 ( .A1(n7185), .A2(DATAI_31_), .ZN(n6749) );
  INV_X1 U5679 ( .A(n6749), .ZN(n7651) );
  AOI22_X1 U5680 ( .A1(n7648), .A2(n6952), .B1(n6951), .B2(n7651), .ZN(n5066)
         );
  OAI211_X1 U5681 ( .C1(n6956), .C2(n5068), .A(n5067), .B(n5066), .ZN(U3147)
         );
  INV_X1 U5682 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5072) );
  NOR2_X2 U5683 ( .A1(n6678), .A2(n5069), .ZN(n7622) );
  INV_X1 U5684 ( .A(DATAI_3_), .ZN(n7566) );
  NOR2_X2 U5685 ( .A1(n7566), .A2(n6679), .ZN(n6809) );
  AOI22_X1 U5686 ( .A1(n7622), .A2(n6950), .B1(n6809), .B2(n6948), .ZN(n5071)
         );
  NAND2_X1 U5687 ( .A1(n7185), .A2(DATAI_27_), .ZN(n6728) );
  INV_X1 U5688 ( .A(n6728), .ZN(n7623) );
  AOI22_X1 U5689 ( .A1(n7624), .A2(n6952), .B1(n6951), .B2(n7623), .ZN(n5070)
         );
  OAI211_X1 U5690 ( .C1(n6956), .C2(n5072), .A(n5071), .B(n5070), .ZN(U3143)
         );
  INV_X1 U5691 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5076) );
  NOR2_X2 U5692 ( .A1(n6678), .A2(n5073), .ZN(n7616) );
  INV_X1 U5693 ( .A(DATAI_2_), .ZN(n5237) );
  NOR2_X2 U5694 ( .A1(n5237), .A2(n6679), .ZN(n6805) );
  AOI22_X1 U5695 ( .A1(n7616), .A2(n6950), .B1(n6805), .B2(n6948), .ZN(n5075)
         );
  NAND2_X1 U5696 ( .A1(n7185), .A2(DATAI_26_), .ZN(n6723) );
  INV_X1 U5697 ( .A(n6723), .ZN(n7618) );
  AOI22_X1 U5698 ( .A1(n7617), .A2(n6952), .B1(n6951), .B2(n7618), .ZN(n5074)
         );
  OAI211_X1 U5699 ( .C1(n6956), .C2(n5076), .A(n5075), .B(n5074), .ZN(U3142)
         );
  INV_X1 U5700 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5079) );
  NOR2_X2 U5701 ( .A1(n6678), .A2(n3905), .ZN(n7596) );
  INV_X1 U5702 ( .A(DATAI_0_), .ZN(n6346) );
  NOR2_X2 U5703 ( .A1(n6346), .A2(n6679), .ZN(n6798) );
  AOI22_X1 U5704 ( .A1(n7596), .A2(n6950), .B1(n6798), .B2(n6948), .ZN(n5078)
         );
  NAND2_X1 U5705 ( .A1(n7185), .A2(DATAI_24_), .ZN(n6714) );
  INV_X1 U5706 ( .A(n6714), .ZN(n7597) );
  AOI22_X1 U5707 ( .A1(n7606), .A2(n6952), .B1(n6951), .B2(n7597), .ZN(n5077)
         );
  OAI211_X1 U5708 ( .C1(n6956), .C2(n5079), .A(n5078), .B(n5077), .ZN(U3140)
         );
  INV_X1 U5709 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U5710 ( .A1(n7048), .A2(UWORD_REG_14__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5080) );
  OAI21_X1 U5711 ( .B1(n5081), .B2(n5096), .A(n5080), .ZN(U2893) );
  INV_X1 U5712 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5083) );
  AOI22_X1 U5713 ( .A1(n7048), .A2(UWORD_REG_0__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5082) );
  OAI21_X1 U5714 ( .B1(n5083), .B2(n5096), .A(n5082), .ZN(U2907) );
  AOI22_X1 U5715 ( .A1(n7048), .A2(UWORD_REG_1__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5084) );
  OAI21_X1 U5716 ( .B1(n7558), .B2(n5096), .A(n5084), .ZN(U2906) );
  INV_X1 U5717 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5086) );
  AOI22_X1 U5718 ( .A1(n7048), .A2(UWORD_REG_2__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5085) );
  OAI21_X1 U5719 ( .B1(n5086), .B2(n5096), .A(n5085), .ZN(U2905) );
  INV_X1 U5720 ( .A(EAX_REG_19__SCAN_IN), .ZN(n7565) );
  AOI22_X1 U5721 ( .A1(n7048), .A2(UWORD_REG_3__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5087) );
  OAI21_X1 U5722 ( .B1(n7565), .B2(n5096), .A(n5087), .ZN(U2904) );
  INV_X1 U5723 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5089) );
  AOI22_X1 U5724 ( .A1(n7048), .A2(UWORD_REG_4__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5088) );
  OAI21_X1 U5725 ( .B1(n5089), .B2(n5096), .A(n5088), .ZN(U2903) );
  INV_X1 U5726 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U5727 ( .A1(n7048), .A2(UWORD_REG_10__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5090) );
  OAI21_X1 U5728 ( .B1(n5091), .B2(n5096), .A(n5090), .ZN(U2897) );
  INV_X1 U5729 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5093) );
  AOI22_X1 U5730 ( .A1(n7048), .A2(UWORD_REG_11__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5092) );
  OAI21_X1 U5731 ( .B1(n5093), .B2(n5096), .A(n5092), .ZN(U2896) );
  AOI22_X1 U5732 ( .A1(n7048), .A2(UWORD_REG_12__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5094) );
  OAI21_X1 U5733 ( .B1(n4694), .B2(n5096), .A(n5094), .ZN(U2895) );
  INV_X1 U5734 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5097) );
  AOI22_X1 U5735 ( .A1(n7048), .A2(UWORD_REG_13__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5095) );
  OAI21_X1 U5736 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(U2894) );
  NAND2_X1 U5737 ( .A1(n6706), .A2(n5904), .ZN(n5789) );
  NOR2_X1 U5738 ( .A1(n5789), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5102)
         );
  NAND2_X1 U5739 ( .A1(n5050), .A2(n5206), .ZN(n5098) );
  OR2_X1 U5740 ( .A1(n6703), .A2(n4267), .ZN(n7589) );
  NAND2_X1 U5741 ( .A1(n6090), .A2(n5047), .ZN(n5795) );
  NOR2_X1 U5742 ( .A1(n7589), .A2(n5795), .ZN(n5106) );
  AOI211_X1 U5743 ( .C1(n5105), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n5106), .ZN(n5100) );
  INV_X1 U5744 ( .A(n5102), .ZN(n5108) );
  NOR2_X1 U5745 ( .A1(n6784), .A2(n5108), .ZN(n6695) );
  INV_X1 U5746 ( .A(n6695), .ZN(n5099) );
  OAI21_X1 U5747 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5100), .A(n5099), .ZN(
        n5101) );
  OAI211_X1 U5748 ( .C1(n5102), .C2(n7200), .A(n5748), .B(n5101), .ZN(n5103)
         );
  INV_X1 U5749 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5112) );
  INV_X1 U5750 ( .A(n5105), .ZN(n5104) );
  OAI21_X1 U5751 ( .B1(n5106), .B2(n6695), .A(n7599), .ZN(n5107) );
  OAI21_X1 U5752 ( .B1(n5108), .B2(n5906), .A(n5107), .ZN(n6694) );
  AOI22_X1 U5753 ( .A1(n7616), .A2(n6695), .B1(n6805), .B2(n6694), .ZN(n5109)
         );
  OAI21_X1 U5754 ( .B1(n6723), .B2(n6697), .A(n5109), .ZN(n5110) );
  AOI21_X1 U5755 ( .B1(n7617), .B2(n6710), .A(n5110), .ZN(n5111) );
  OAI21_X1 U5756 ( .B1(n6701), .B2(n5112), .A(n5111), .ZN(U3030) );
  INV_X1 U5757 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U5758 ( .A1(n7634), .A2(n6695), .B1(n6816), .B2(n6694), .ZN(n5113)
         );
  OAI21_X1 U5759 ( .B1(n6737), .B2(n6697), .A(n5113), .ZN(n5114) );
  AOI21_X1 U5760 ( .B1(n7635), .B2(n6710), .A(n5114), .ZN(n5115) );
  OAI21_X1 U5761 ( .B1(n6701), .B2(n5116), .A(n5115), .ZN(U3033) );
  INV_X1 U5762 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U5763 ( .A1(n7640), .A2(n6695), .B1(n6820), .B2(n6694), .ZN(n5117)
         );
  OAI21_X1 U5764 ( .B1(n6742), .B2(n6697), .A(n5117), .ZN(n5118) );
  AOI21_X1 U5765 ( .B1(n7641), .B2(n6710), .A(n5118), .ZN(n5119) );
  OAI21_X1 U5766 ( .B1(n6701), .B2(n5120), .A(n5119), .ZN(U3034) );
  INV_X1 U5767 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5124) );
  AOI22_X1 U5768 ( .A1(n7622), .A2(n6695), .B1(n6809), .B2(n6694), .ZN(n5121)
         );
  OAI21_X1 U5769 ( .B1(n6728), .B2(n6697), .A(n5121), .ZN(n5122) );
  AOI21_X1 U5770 ( .B1(n7624), .B2(n6710), .A(n5122), .ZN(n5123) );
  OAI21_X1 U5771 ( .B1(n6701), .B2(n5124), .A(n5123), .ZN(U3031) );
  INV_X1 U5772 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U5773 ( .A1(n7596), .A2(n6695), .B1(n6798), .B2(n6694), .ZN(n5125)
         );
  OAI21_X1 U5774 ( .B1(n6714), .B2(n6697), .A(n5125), .ZN(n5126) );
  AOI21_X1 U5775 ( .B1(n7606), .B2(n6710), .A(n5126), .ZN(n5127) );
  OAI21_X1 U5776 ( .B1(n6701), .B2(n5128), .A(n5127), .ZN(U3028) );
  INV_X1 U5777 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U5778 ( .A1(n7647), .A2(n6695), .B1(n6825), .B2(n6694), .ZN(n5129)
         );
  OAI21_X1 U5779 ( .B1(n6749), .B2(n6697), .A(n5129), .ZN(n5130) );
  AOI21_X1 U5780 ( .B1(n7648), .B2(n6710), .A(n5130), .ZN(n5131) );
  OAI21_X1 U5781 ( .B1(n6701), .B2(n5132), .A(n5131), .ZN(U3035) );
  NAND2_X1 U5782 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  XOR2_X1 U5783 ( .A(n5136), .B(n5135), .Z(n5984) );
  OAI222_X1 U5784 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5139), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n7226), .C1(n5138), .C2(n5137), 
        .ZN(n5141) );
  AND2_X1 U5785 ( .A1(n7280), .A2(REIP_REG_1__SCAN_IN), .ZN(n5983) );
  INV_X1 U5786 ( .A(n5983), .ZN(n5140) );
  OAI211_X1 U5787 ( .C1(n7301), .C2(n5142), .A(n5141), .B(n5140), .ZN(n5143)
         );
  AOI21_X1 U5788 ( .B1(n7314), .B2(n5984), .A(n5143), .ZN(n5144) );
  INV_X1 U5789 ( .A(n5144), .ZN(U3017) );
  NAND2_X1 U5790 ( .A1(n5829), .A2(n7599), .ZN(n5823) );
  AND2_X1 U5791 ( .A1(n5052), .A2(n6785), .ZN(n5145) );
  AOI211_X1 U5792 ( .C1(n6797), .C2(n5823), .A(n6919), .B(n6929), .ZN(n5150)
         );
  NAND3_X1 U5793 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6967), .ZN(n5684) );
  NOR2_X1 U5794 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5684), .ZN(n6915)
         );
  NOR2_X1 U5795 ( .A1(n6915), .A2(n7533), .ZN(n5149) );
  INV_X1 U5796 ( .A(n5151), .ZN(n5147) );
  NAND2_X1 U5797 ( .A1(n5147), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U5798 ( .A1(n5748), .A2(n6711), .ZN(n6789) );
  INV_X1 U5799 ( .A(n6789), .ZN(n5148) );
  OAI21_X1 U5800 ( .B1(n5679), .B2(n6853), .A(n5148), .ZN(n5825) );
  INV_X1 U5801 ( .A(n6707), .ZN(n5831) );
  NAND2_X1 U5802 ( .A1(n5830), .A2(n5831), .ZN(n5753) );
  NOR4_X2 U5803 ( .A1(n5150), .A2(n5149), .A3(n5825), .A4(n3741), .ZN(n6922)
         );
  INV_X1 U5804 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5155) );
  INV_X1 U5805 ( .A(n7606), .ZN(n6865) );
  NAND2_X1 U5806 ( .A1(n6703), .A2(n7599), .ZN(n6788) );
  NAND2_X1 U5807 ( .A1(n5151), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6796) );
  OAI22_X1 U5808 ( .A1(n6788), .A2(n5829), .B1(n6796), .B2(n5753), .ZN(n6914)
         );
  AOI22_X1 U5809 ( .A1(n7596), .A2(n6915), .B1(n6798), .B2(n6914), .ZN(n5152)
         );
  OAI21_X1 U5810 ( .B1(n6917), .B2(n6865), .A(n5152), .ZN(n5153) );
  AOI21_X1 U5811 ( .B1(n7597), .B2(n6919), .A(n5153), .ZN(n5154) );
  OAI21_X1 U5812 ( .B1(n6922), .B2(n5155), .A(n5154), .ZN(U3116) );
  INV_X1 U5813 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5159) );
  INV_X1 U5814 ( .A(n7617), .ZN(n6872) );
  AOI22_X1 U5815 ( .A1(n7616), .A2(n6915), .B1(n6805), .B2(n6914), .ZN(n5156)
         );
  OAI21_X1 U5816 ( .B1(n6917), .B2(n6872), .A(n5156), .ZN(n5157) );
  AOI21_X1 U5817 ( .B1(n7618), .B2(n6919), .A(n5157), .ZN(n5158) );
  OAI21_X1 U5818 ( .B1(n6922), .B2(n5159), .A(n5158), .ZN(U3118) );
  INV_X1 U5819 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5163) );
  INV_X1 U5820 ( .A(n7624), .ZN(n6876) );
  AOI22_X1 U5821 ( .A1(n7622), .A2(n6915), .B1(n6809), .B2(n6914), .ZN(n5160)
         );
  OAI21_X1 U5822 ( .B1(n6917), .B2(n6876), .A(n5160), .ZN(n5161) );
  AOI21_X1 U5823 ( .B1(n7623), .B2(n6919), .A(n5161), .ZN(n5162) );
  OAI21_X1 U5824 ( .B1(n6922), .B2(n5163), .A(n5162), .ZN(U3119) );
  INV_X1 U5825 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5167) );
  INV_X1 U5826 ( .A(n7648), .ZN(n6893) );
  AOI22_X1 U5827 ( .A1(n7647), .A2(n6915), .B1(n6825), .B2(n6914), .ZN(n5164)
         );
  OAI21_X1 U5828 ( .B1(n6917), .B2(n6893), .A(n5164), .ZN(n5165) );
  AOI21_X1 U5829 ( .B1(n7651), .B2(n6919), .A(n5165), .ZN(n5166) );
  OAI21_X1 U5830 ( .B1(n6922), .B2(n5167), .A(n5166), .ZN(U3123) );
  INV_X1 U5831 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5171) );
  INV_X1 U5832 ( .A(n7641), .ZN(n6887) );
  AOI22_X1 U5833 ( .A1(n7640), .A2(n6915), .B1(n6820), .B2(n6914), .ZN(n5168)
         );
  OAI21_X1 U5834 ( .B1(n6917), .B2(n6887), .A(n5168), .ZN(n5169) );
  AOI21_X1 U5835 ( .B1(n7642), .B2(n6919), .A(n5169), .ZN(n5170) );
  OAI21_X1 U5836 ( .B1(n6922), .B2(n5171), .A(n5170), .ZN(U3122) );
  INV_X1 U5837 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5175) );
  INV_X1 U5838 ( .A(n7635), .ZN(n6883) );
  AOI22_X1 U5839 ( .A1(n7634), .A2(n6915), .B1(n6816), .B2(n6914), .ZN(n5172)
         );
  OAI21_X1 U5840 ( .B1(n6917), .B2(n6883), .A(n5172), .ZN(n5173) );
  AOI21_X1 U5841 ( .B1(n7636), .B2(n6919), .A(n5173), .ZN(n5174) );
  OAI21_X1 U5842 ( .B1(n6922), .B2(n5175), .A(n5174), .ZN(U3121) );
  INV_X1 U5843 ( .A(n5182), .ZN(n5176) );
  NAND3_X1 U5844 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5904), .A3(n6967), .ZN(n5747) );
  INV_X1 U5845 ( .A(n5747), .ZN(n5179) );
  OAI21_X1 U5846 ( .B1(n5182), .B2(n7535), .A(n7599), .ZN(n5180) );
  INV_X1 U5847 ( .A(n5180), .ZN(n5177) );
  INV_X1 U5848 ( .A(n5795), .ZN(n5750) );
  NOR2_X1 U5849 ( .A1(n6784), .A2(n5747), .ZN(n6849) );
  AOI21_X1 U5850 ( .B1(n5680), .B2(n5750), .A(n6849), .ZN(n5181) );
  NAND2_X1 U5851 ( .A1(n5177), .A2(n5181), .ZN(n5178) );
  OAI211_X1 U5852 ( .C1(n7599), .C2(n5179), .A(n7602), .B(n5178), .ZN(n6848)
         );
  OAI22_X1 U5853 ( .A1(n5181), .A2(n5180), .B1(n7200), .B2(n5747), .ZN(n6847)
         );
  AOI22_X1 U5854 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6848), .B1(n6805), 
        .B2(n6847), .ZN(n5184) );
  AOI22_X1 U5855 ( .A1(n6895), .A2(n7617), .B1(n6849), .B2(n7616), .ZN(n5183)
         );
  OAI211_X1 U5856 ( .C1(n6852), .C2(n6723), .A(n5184), .B(n5183), .ZN(U3094)
         );
  AOI22_X1 U5857 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6848), .B1(n6820), 
        .B2(n6847), .ZN(n5186) );
  AOI22_X1 U5858 ( .A1(n6895), .A2(n7641), .B1(n6849), .B2(n7640), .ZN(n5185)
         );
  OAI211_X1 U5859 ( .C1(n6852), .C2(n6742), .A(n5186), .B(n5185), .ZN(U3098)
         );
  AOI22_X1 U5860 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6848), .B1(n6798), 
        .B2(n6847), .ZN(n5188) );
  AOI22_X1 U5861 ( .A1(n6895), .A2(n7606), .B1(n7596), .B2(n6849), .ZN(n5187)
         );
  OAI211_X1 U5862 ( .C1(n6714), .C2(n6852), .A(n5188), .B(n5187), .ZN(U3092)
         );
  AOI22_X1 U5863 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6848), .B1(n6816), 
        .B2(n6847), .ZN(n5190) );
  AOI22_X1 U5864 ( .A1(n6895), .A2(n7635), .B1(n6849), .B2(n7634), .ZN(n5189)
         );
  OAI211_X1 U5865 ( .C1(n6852), .C2(n6737), .A(n5190), .B(n5189), .ZN(U3097)
         );
  AOI22_X1 U5866 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6848), .B1(n6809), 
        .B2(n6847), .ZN(n5192) );
  AOI22_X1 U5867 ( .A1(n6895), .A2(n7624), .B1(n6849), .B2(n7622), .ZN(n5191)
         );
  OAI211_X1 U5868 ( .C1(n6852), .C2(n6728), .A(n5192), .B(n5191), .ZN(U3095)
         );
  AOI22_X1 U5869 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6848), .B1(n6825), 
        .B2(n6847), .ZN(n5194) );
  AOI22_X1 U5870 ( .A1(n6895), .A2(n7648), .B1(n6849), .B2(n7647), .ZN(n5193)
         );
  OAI211_X1 U5871 ( .C1(n6852), .C2(n6749), .A(n5194), .B(n5193), .ZN(U3099)
         );
  NAND2_X1 U5872 ( .A1(n5893), .A2(DATAI_8_), .ZN(n5869) );
  INV_X1 U5873 ( .A(n5197), .ZN(n5198) );
  AOI22_X1 U5874 ( .A1(n5894), .A2(EAX_REG_24__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U5875 ( .A1(n5869), .A2(n5200), .ZN(U2932) );
  NAND2_X1 U5876 ( .A1(n5893), .A2(DATAI_7_), .ZN(n5867) );
  AOI22_X1 U5877 ( .A1(n5894), .A2(EAX_REG_23__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5878 ( .A1(n5867), .A2(n5201), .ZN(U2931) );
  NAND2_X1 U5879 ( .A1(n5893), .A2(DATAI_6_), .ZN(n5865) );
  AOI22_X1 U5880 ( .A1(n5894), .A2(EAX_REG_22__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U5881 ( .A1(n5865), .A2(n5202), .ZN(U2930) );
  NAND2_X1 U5882 ( .A1(n5893), .A2(DATAI_9_), .ZN(n5885) );
  AOI22_X1 U5883 ( .A1(n5894), .A2(EAX_REG_25__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U5884 ( .A1(n5885), .A2(n5203), .ZN(U2933) );
  NAND2_X1 U5885 ( .A1(n5893), .A2(DATAI_11_), .ZN(n5863) );
  AOI22_X1 U5886 ( .A1(n5933), .A2(EAX_REG_27__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U5887 ( .A1(n5863), .A2(n5204), .ZN(U2935) );
  NAND2_X1 U5888 ( .A1(n5893), .A2(DATAI_10_), .ZN(n5887) );
  AOI22_X1 U5889 ( .A1(n5933), .A2(EAX_REG_26__SCAN_IN), .B1(n5860), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U5890 ( .A1(n5887), .A2(n5205), .ZN(U2934) );
  NOR2_X1 U5891 ( .A1(n5050), .A2(n4085), .ZN(n7588) );
  NAND2_X1 U5892 ( .A1(n7588), .A2(n5206), .ZN(n5213) );
  OR2_X1 U5893 ( .A1(n5213), .A2(n7535), .ZN(n5207) );
  AND2_X1 U5894 ( .A1(n5207), .A2(n7599), .ZN(n5209) );
  INV_X1 U5895 ( .A(n7589), .ZN(n5246) );
  NAND2_X1 U5896 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6706), .ZN(n7591) );
  OR2_X1 U5897 ( .A1(n7591), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5210)
         );
  NOR2_X1 U5898 ( .A1(n6784), .A2(n5210), .ZN(n6780) );
  AOI21_X1 U5899 ( .B1(n5246), .B2(n5679), .A(n6780), .ZN(n5212) );
  AOI22_X1 U5900 ( .A1(n5209), .A2(n5212), .B1(n7587), .B2(n5210), .ZN(n5208)
         );
  NAND2_X1 U5901 ( .A1(n7602), .A2(n5208), .ZN(n6779) );
  INV_X1 U5902 ( .A(n5209), .ZN(n5211) );
  OAI22_X1 U5903 ( .A1(n5212), .A2(n5211), .B1(n7200), .B2(n5210), .ZN(n6778)
         );
  AOI22_X1 U5904 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6779), .B1(n6825), 
        .B2(n6778), .ZN(n5215) );
  AOI22_X1 U5905 ( .A1(n6827), .A2(n7648), .B1(n7647), .B2(n6780), .ZN(n5214)
         );
  OAI211_X1 U5906 ( .C1(n6749), .C2(n6783), .A(n5215), .B(n5214), .ZN(U3067)
         );
  AOI22_X1 U5907 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6779), .B1(n6809), 
        .B2(n6778), .ZN(n5217) );
  AOI22_X1 U5908 ( .A1(n6827), .A2(n7624), .B1(n7622), .B2(n6780), .ZN(n5216)
         );
  OAI211_X1 U5909 ( .C1(n6728), .C2(n6783), .A(n5217), .B(n5216), .ZN(U3063)
         );
  AOI22_X1 U5910 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6779), .B1(n6816), 
        .B2(n6778), .ZN(n5219) );
  AOI22_X1 U5911 ( .A1(n6827), .A2(n7635), .B1(n7634), .B2(n6780), .ZN(n5218)
         );
  OAI211_X1 U5912 ( .C1(n6737), .C2(n6783), .A(n5219), .B(n5218), .ZN(U3065)
         );
  AOI22_X1 U5913 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6779), .B1(n6805), 
        .B2(n6778), .ZN(n5221) );
  AOI22_X1 U5914 ( .A1(n6827), .A2(n7617), .B1(n7616), .B2(n6780), .ZN(n5220)
         );
  OAI211_X1 U5915 ( .C1(n6723), .C2(n6783), .A(n5221), .B(n5220), .ZN(U3062)
         );
  AOI22_X1 U5916 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6779), .B1(n6798), 
        .B2(n6778), .ZN(n5223) );
  AOI22_X1 U5917 ( .A1(n6827), .A2(n7606), .B1(n7596), .B2(n6780), .ZN(n5222)
         );
  OAI211_X1 U5918 ( .C1(n6714), .C2(n6783), .A(n5223), .B(n5222), .ZN(U3060)
         );
  AOI22_X1 U5919 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6779), .B1(n6820), 
        .B2(n6778), .ZN(n5225) );
  AOI22_X1 U5920 ( .A1(n6827), .A2(n7641), .B1(n7640), .B2(n6780), .ZN(n5224)
         );
  OAI211_X1 U5921 ( .C1(n6742), .C2(n6783), .A(n5225), .B(n5224), .ZN(U3066)
         );
  NOR2_X1 U5922 ( .A1(n4935), .A2(n5226), .ZN(n5227) );
  NAND2_X1 U5923 ( .A1(n7564), .A2(n5230), .ZN(n6356) );
  INV_X1 U5924 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7021) );
  INV_X1 U5925 ( .A(n5230), .ZN(n5231) );
  OAI222_X1 U5926 ( .A1(n6346), .A2(n6356), .B1(n7564), .B2(n7021), .C1(n6354), 
        .C2(n5232), .ZN(U2891) );
  INV_X1 U5927 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7025) );
  INV_X1 U5928 ( .A(n5233), .ZN(n5235) );
  NAND3_X1 U5929 ( .A1(n5235), .A2(n5234), .A3(n4965), .ZN(n5236) );
  NAND2_X1 U5930 ( .A1(n5236), .A2(n5020), .ZN(n7126) );
  OAI222_X1 U5931 ( .A1(n6356), .A2(n5237), .B1(n7564), .B2(n7025), .C1(n6354), 
        .C2(n7126), .ZN(U2889) );
  INV_X1 U5932 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7027) );
  OAI222_X1 U5933 ( .A1(n7566), .A2(n6356), .B1(n7564), .B2(n7027), .C1(n6354), 
        .C2(n5944), .ZN(U2888) );
  INV_X1 U5934 ( .A(DATAI_1_), .ZN(n7559) );
  INV_X1 U5935 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7023) );
  OAI222_X1 U5936 ( .A1(n7559), .A2(n6356), .B1(n7564), .B2(n7023), .C1(n6354), 
        .C2(n5987), .ZN(U2890) );
  OAI222_X1 U5937 ( .A1(n7341), .A2(n6354), .B1(n6356), .B2(n5238), .C1(n7564), 
        .C2(n4299), .ZN(U2886) );
  INV_X1 U5938 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7029) );
  INV_X1 U5939 ( .A(DATAI_4_), .ZN(n6680) );
  INV_X1 U5940 ( .A(n5239), .ZN(n5240) );
  XNOR2_X1 U5941 ( .A(n5022), .B(n5240), .ZN(n7330) );
  INV_X1 U5942 ( .A(n7330), .ZN(n5241) );
  OAI222_X1 U5943 ( .A1(n7564), .A2(n7029), .B1(n6356), .B2(n6680), .C1(n6354), 
        .C2(n5241), .ZN(U2887) );
  INV_X1 U5944 ( .A(n5242), .ZN(n5672) );
  AND2_X1 U5945 ( .A1(n5050), .A2(n5052), .ZN(n5243) );
  INV_X1 U5946 ( .A(n5251), .ZN(n5244) );
  OR2_X1 U5947 ( .A1(n5251), .A2(n7535), .ZN(n5245) );
  AND2_X1 U5948 ( .A1(n5245), .A2(n7599), .ZN(n5248) );
  NAND2_X1 U5949 ( .A1(n6090), .A2(n6665), .ZN(n6712) );
  INV_X1 U5950 ( .A(n6712), .ZN(n5903) );
  NOR2_X1 U5951 ( .A1(n7592), .A2(n5789), .ZN(n6759) );
  AOI21_X1 U5952 ( .B1(n5246), .B2(n5903), .A(n6759), .ZN(n5250) );
  OR2_X1 U5953 ( .A1(n6967), .A2(n5789), .ZN(n6704) );
  AOI22_X1 U5954 ( .A1(n5248), .A2(n5250), .B1(n7587), .B2(n6704), .ZN(n5247)
         );
  NAND2_X1 U5955 ( .A1(n7602), .A2(n5247), .ZN(n6758) );
  INV_X1 U5956 ( .A(n5248), .ZN(n5249) );
  OAI22_X1 U5957 ( .A1(n5250), .A2(n5249), .B1(n7200), .B2(n6704), .ZN(n6757)
         );
  AOI22_X1 U5958 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6758), .B1(n6798), 
        .B2(n6757), .ZN(n5253) );
  AOI22_X1 U5959 ( .A1(n6760), .A2(n7597), .B1(n7596), .B2(n6759), .ZN(n5252)
         );
  OAI211_X1 U5960 ( .C1(n6865), .C2(n6772), .A(n5253), .B(n5252), .ZN(U3044)
         );
  AOI22_X1 U5961 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6758), .B1(n6816), 
        .B2(n6757), .ZN(n5255) );
  AOI22_X1 U5962 ( .A1(n6760), .A2(n7636), .B1(n7634), .B2(n6759), .ZN(n5254)
         );
  OAI211_X1 U5963 ( .C1(n6883), .C2(n6772), .A(n5255), .B(n5254), .ZN(U3049)
         );
  AOI22_X1 U5964 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6758), .B1(n6825), 
        .B2(n6757), .ZN(n5257) );
  AOI22_X1 U5965 ( .A1(n6760), .A2(n7651), .B1(n7647), .B2(n6759), .ZN(n5256)
         );
  OAI211_X1 U5966 ( .C1(n6893), .C2(n6772), .A(n5257), .B(n5256), .ZN(U3051)
         );
  AOI22_X1 U5967 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6758), .B1(n6809), 
        .B2(n6757), .ZN(n5259) );
  AOI22_X1 U5968 ( .A1(n6760), .A2(n7623), .B1(n7622), .B2(n6759), .ZN(n5258)
         );
  OAI211_X1 U5969 ( .C1(n6876), .C2(n6772), .A(n5259), .B(n5258), .ZN(U3047)
         );
  AOI22_X1 U5970 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6758), .B1(n6820), 
        .B2(n6757), .ZN(n5261) );
  AOI22_X1 U5971 ( .A1(n6760), .A2(n7642), .B1(n7640), .B2(n6759), .ZN(n5260)
         );
  OAI211_X1 U5972 ( .C1(n6887), .C2(n6772), .A(n5261), .B(n5260), .ZN(U3050)
         );
  AOI22_X1 U5973 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6758), .B1(n6805), 
        .B2(n6757), .ZN(n5263) );
  AOI22_X1 U5974 ( .A1(n6760), .A2(n7618), .B1(n7616), .B2(n6759), .ZN(n5262)
         );
  OAI211_X1 U5975 ( .C1(n6872), .C2(n6772), .A(n5263), .B(n5262), .ZN(U3046)
         );
  OR2_X1 U5976 ( .A1(n6962), .A2(n3750), .ZN(n5266) );
  NAND2_X1 U5977 ( .A1(n6962), .A2(n5264), .ZN(n5265) );
  INV_X1 U5978 ( .A(n6969), .ZN(n5277) );
  OR2_X1 U5979 ( .A1(n6962), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5276)
         );
  INV_X1 U5980 ( .A(n5267), .ZN(n6664) );
  XNOR2_X1 U5981 ( .A(n5268), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5273)
         );
  XNOR2_X1 U5982 ( .A(n5269), .B(n3744), .ZN(n5270) );
  NAND2_X1 U5983 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  OAI21_X1 U5984 ( .B1(n5273), .B2(n6661), .A(n5272), .ZN(n5274) );
  AOI21_X1 U5985 ( .B1(n6703), .B2(n6664), .A(n5274), .ZN(n7511) );
  NAND2_X1 U5986 ( .A1(n6962), .A2(n7511), .ZN(n5275) );
  NAND3_X1 U5987 ( .A1(n5277), .A2(n6957), .A3(n6667), .ZN(n5281) );
  NOR2_X1 U5988 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6667), .ZN(n5278) );
  NAND2_X1 U5989 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  MUX2_X1 U5990 ( .A(n6962), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5283) );
  INV_X1 U5991 ( .A(n5283), .ZN(n5290) );
  INV_X1 U5992 ( .A(n5284), .ZN(n5285) );
  OR2_X1 U5993 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  XNOR2_X1 U5994 ( .A(n5287), .B(n7520), .ZN(n7514) );
  OR2_X1 U5995 ( .A1(n4904), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5288) );
  NOR2_X1 U5996 ( .A1(n7514), .A2(n5288), .ZN(n5289) );
  AOI21_X1 U5997 ( .B1(n5290), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n5289), 
        .ZN(n6983) );
  OAI21_X1 U5998 ( .B1(n6984), .B2(n5282), .A(n6983), .ZN(n6991) );
  OR2_X1 U5999 ( .A1(n6991), .A2(FLUSH_REG_SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6000 ( .A1(n5291), .A2(n7199), .ZN(n5292) );
  NAND2_X1 U6001 ( .A1(n5292), .A2(n6679), .ZN(n7015) );
  NOR2_X1 U6002 ( .A1(n6082), .A2(n7587), .ZN(n6079) );
  INV_X1 U6003 ( .A(n6079), .ZN(n5821) );
  OAI21_X1 U6004 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6667), .A(n7015), .ZN(
        n6085) );
  INV_X1 U6005 ( .A(n6085), .ZN(n5674) );
  INV_X1 U6006 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7502) );
  OAI21_X1 U6007 ( .B1(n7502), .B2(n7531), .A(n6679), .ZN(n5293) );
  NAND2_X1 U6008 ( .A1(n5293), .A2(n7526), .ZN(n5294) );
  OAI22_X1 U6009 ( .A1(n7015), .A2(n6784), .B1(n6991), .B2(n5294), .ZN(n5295)
         );
  AOI21_X1 U6010 ( .B1(n5674), .B2(n5905), .A(n5295), .ZN(n5296) );
  OAI21_X1 U6011 ( .B1(n5821), .B2(n5057), .A(n5296), .ZN(U3465) );
  INV_X1 U6012 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7013) );
  XNOR2_X1 U6013 ( .A(n7013), .B(keyinput_254), .ZN(n5667) );
  XOR2_X1 U6014 ( .A(DATAI_30_), .B(keyinput_129), .Z(n5299) );
  XOR2_X1 U6015 ( .A(DATAI_31_), .B(keyinput_128), .Z(n5298) );
  XOR2_X1 U6016 ( .A(DATAI_29_), .B(keyinput_130), .Z(n5297) );
  NAND3_X1 U6017 ( .A1(n5299), .A2(n5298), .A3(n5297), .ZN(n5302) );
  XNOR2_X1 U6018 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n5301) );
  XNOR2_X1 U6019 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n5300) );
  NAND3_X1 U6020 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n5305) );
  XNOR2_X1 U6021 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n5304) );
  XNOR2_X1 U6022 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n5303) );
  NAND3_X1 U6023 ( .A1(n5305), .A2(n5304), .A3(n5303), .ZN(n5309) );
  XOR2_X1 U6024 ( .A(DATAI_22_), .B(keyinput_137), .Z(n5308) );
  XOR2_X1 U6025 ( .A(DATAI_24_), .B(keyinput_135), .Z(n5307) );
  XNOR2_X1 U6026 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n5306) );
  NAND4_X1 U6027 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n5312)
         );
  XNOR2_X1 U6028 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n5311) );
  XOR2_X1 U6029 ( .A(DATAI_20_), .B(keyinput_139), .Z(n5310) );
  AOI21_X1 U6030 ( .B1(n5312), .B2(n5311), .A(n5310), .ZN(n5327) );
  XOR2_X1 U6031 ( .A(DATAI_19_), .B(keyinput_140), .Z(n5326) );
  INV_X1 U6032 ( .A(DATAI_13_), .ZN(n6355) );
  INV_X1 U6033 ( .A(DATAI_18_), .ZN(n5313) );
  NAND2_X1 U6034 ( .A1(n5313), .A2(keyinput_141), .ZN(n5318) );
  INV_X1 U6035 ( .A(DATAI_15_), .ZN(n6347) );
  INV_X1 U6036 ( .A(DATAI_17_), .ZN(n5319) );
  OAI22_X1 U6037 ( .A1(n6347), .A2(keyinput_144), .B1(n5319), .B2(keyinput_142), .ZN(n5316) );
  OAI22_X1 U6038 ( .A1(n6355), .A2(keyinput_146), .B1(keyinput_145), .B2(
        DATAI_14_), .ZN(n5315) );
  OAI22_X1 U6039 ( .A1(n5313), .A2(keyinput_141), .B1(keyinput_147), .B2(
        DATAI_12_), .ZN(n5314) );
  NOR3_X1 U6040 ( .A1(n5316), .A2(n5315), .A3(n5314), .ZN(n5317) );
  NAND2_X1 U6041 ( .A1(n5318), .A2(n5317), .ZN(n5323) );
  AOI22_X1 U6042 ( .A1(keyinput_144), .A2(n6347), .B1(n5319), .B2(keyinput_142), .ZN(n5321) );
  AOI22_X1 U6043 ( .A1(DATAI_14_), .A2(keyinput_145), .B1(DATAI_12_), .B2(
        keyinput_147), .ZN(n5320) );
  NAND2_X1 U6044 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  AOI211_X1 U6045 ( .C1(keyinput_146), .C2(n6355), .A(n5323), .B(n5322), .ZN(
        n5325) );
  XNOR2_X1 U6046 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n5324) );
  OAI211_X1 U6047 ( .C1(n5327), .C2(n5326), .A(n5325), .B(n5324), .ZN(n5330)
         );
  XOR2_X1 U6048 ( .A(DATAI_11_), .B(keyinput_148), .Z(n5329) );
  XOR2_X1 U6049 ( .A(DATAI_10_), .B(keyinput_149), .Z(n5328) );
  AOI21_X1 U6050 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(n5333) );
  XOR2_X1 U6051 ( .A(DATAI_8_), .B(keyinput_151), .Z(n5332) );
  XNOR2_X1 U6052 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n5331) );
  NOR3_X1 U6053 ( .A1(n5333), .A2(n5332), .A3(n5331), .ZN(n5337) );
  XNOR2_X1 U6054 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n5336) );
  XNOR2_X1 U6055 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n5335) );
  XNOR2_X1 U6056 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n5334) );
  NOR4_X1 U6057 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n5341)
         );
  XOR2_X1 U6058 ( .A(DATAI_3_), .B(keyinput_156), .Z(n5340) );
  XOR2_X1 U6059 ( .A(DATAI_4_), .B(keyinput_155), .Z(n5339) );
  XNOR2_X1 U6060 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n5338) );
  NOR4_X1 U6061 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n5345)
         );
  XOR2_X1 U6062 ( .A(DATAI_1_), .B(keyinput_158), .Z(n5344) );
  XOR2_X1 U6063 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .Z(n5343) );
  XNOR2_X1 U6064 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n5342) );
  OAI211_X1 U6065 ( .C1(n5345), .C2(n5344), .A(n5343), .B(n5342), .ZN(n5348)
         );
  XOR2_X1 U6066 ( .A(NA_N), .B(keyinput_161), .Z(n5347) );
  INV_X1 U6067 ( .A(BS16_N), .ZN(n6999) );
  XNOR2_X1 U6068 ( .A(n6999), .B(keyinput_162), .ZN(n5346) );
  AOI21_X1 U6069 ( .B1(n5348), .B2(n5347), .A(n5346), .ZN(n5351) );
  XNOR2_X1 U6070 ( .A(READY_N), .B(keyinput_163), .ZN(n5350) );
  XNOR2_X1 U6071 ( .A(HOLD), .B(keyinput_164), .ZN(n5349) );
  NOR3_X1 U6072 ( .A1(n5351), .A2(n5350), .A3(n5349), .ZN(n5354) );
  INV_X1 U6073 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7017) );
  XNOR2_X1 U6074 ( .A(n7017), .B(keyinput_166), .ZN(n5353) );
  XNOR2_X1 U6075 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .ZN(n5352)
         );
  NOR3_X1 U6076 ( .A1(n5354), .A2(n5353), .A3(n5352), .ZN(n5357) );
  XNOR2_X1 U6077 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_168), .ZN(n5356) );
  XNOR2_X1 U6078 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_167), .ZN(n5355) );
  NOR3_X1 U6079 ( .A1(n5357), .A2(n5356), .A3(n5355), .ZN(n5361) );
  XNOR2_X1 U6080 ( .A(n7535), .B(keyinput_171), .ZN(n5360) );
  XOR2_X1 U6081 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .Z(n5359)
         );
  XOR2_X1 U6082 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_169), .Z(n5358) );
  NOR4_X1 U6083 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n5364)
         );
  XOR2_X1 U6084 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .Z(n5363) );
  XNOR2_X1 U6085 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .ZN(n5362) );
  NOR3_X1 U6086 ( .A1(n5364), .A2(n5363), .A3(n5362), .ZN(n5377) );
  XNOR2_X1 U6087 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .ZN(n5376) );
  AOI22_X1 U6088 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_177), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_175), .ZN(n5365) );
  OAI221_X1 U6089 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_177), .C1(
        BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_175), .A(n5365), .ZN(n5368)
         );
  XNOR2_X1 U6090 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n5367) );
  XNOR2_X1 U6091 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .ZN(n5366) );
  NOR3_X1 U6092 ( .A1(n5368), .A2(n5367), .A3(n5366), .ZN(n5375) );
  INV_X1 U6093 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7101) );
  AOI22_X1 U6094 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_176), .B1(
        n7101), .B2(keyinput_178), .ZN(n5369) );
  OAI221_X1 U6095 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_176), .C1(
        n7101), .C2(keyinput_178), .A(n5369), .ZN(n5373) );
  XNOR2_X1 U6096 ( .A(n7094), .B(keyinput_181), .ZN(n5372) );
  XNOR2_X1 U6097 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n5371) );
  XNOR2_X1 U6098 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .ZN(n5370) );
  NOR4_X1 U6099 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n5374)
         );
  OAI211_X1 U6100 ( .C1(n5377), .C2(n5376), .A(n5375), .B(n5374), .ZN(n5380)
         );
  XOR2_X1 U6101 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .Z(n5379) );
  XNOR2_X1 U6102 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .ZN(n5378) );
  AOI21_X1 U6103 ( .B1(n5380), .B2(n5379), .A(n5378), .ZN(n5383) );
  XNOR2_X1 U6104 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n5382) );
  XNOR2_X1 U6105 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .ZN(n5381) );
  OAI21_X1 U6106 ( .B1(n5383), .B2(n5382), .A(n5381), .ZN(n5386) );
  XNOR2_X1 U6107 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n5385) );
  XNOR2_X1 U6108 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .ZN(n5384) );
  AOI21_X1 U6109 ( .B1(n5386), .B2(n5385), .A(n5384), .ZN(n5390) );
  XOR2_X1 U6110 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .Z(n5389) );
  XOR2_X1 U6111 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n5388) );
  XNOR2_X1 U6112 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .ZN(n5387) );
  OAI211_X1 U6113 ( .C1(n5390), .C2(n5389), .A(n5388), .B(n5387), .ZN(n5393)
         );
  XOR2_X1 U6114 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .Z(n5392) );
  XOR2_X1 U6115 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .Z(n5391) );
  AOI21_X1 U6116 ( .B1(n5393), .B2(n5392), .A(n5391), .ZN(n5411) );
  INV_X1 U6117 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7113) );
  XNOR2_X1 U6118 ( .A(n7113), .B(keyinput_196), .ZN(n5397) );
  XNOR2_X1 U6119 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_197), .ZN(n5396) );
  XNOR2_X1 U6120 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_195), .ZN(n5395) );
  XNOR2_X1 U6121 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_198), .ZN(n5394) );
  NAND4_X1 U6122 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n5410)
         );
  INV_X1 U6123 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7081) );
  INV_X1 U6124 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7097) );
  INV_X1 U6125 ( .A(keyinput_199), .ZN(n5403) );
  INV_X1 U6126 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7085) );
  INV_X1 U6127 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7093) );
  AOI22_X1 U6128 ( .A1(n7085), .A2(keyinput_204), .B1(n7093), .B2(keyinput_200), .ZN(n5401) );
  AOI22_X1 U6129 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(keyinput_201), .B1(n7081), 
        .B2(keyinput_206), .ZN(n5400) );
  AOI22_X1 U6130 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_203), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_205), .ZN(n5399) );
  AOI22_X1 U6131 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_202), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(keyinput_199), .ZN(n5398) );
  NAND4_X1 U6132 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n5402)
         );
  AOI21_X1 U6133 ( .B1(n7097), .B2(n5403), .A(n5402), .ZN(n5404) );
  OAI21_X1 U6134 ( .B1(keyinput_206), .B2(n7081), .A(n5404), .ZN(n5408) );
  OAI22_X1 U6135 ( .A1(n7093), .A2(keyinput_200), .B1(ADDRESS_REG_27__SCAN_IN), 
        .B2(keyinput_201), .ZN(n5407) );
  OAI22_X1 U6136 ( .A1(n7085), .A2(keyinput_204), .B1(ADDRESS_REG_26__SCAN_IN), 
        .B2(keyinput_202), .ZN(n5406) );
  OAI22_X1 U6137 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_203), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(keyinput_205), .ZN(n5405) );
  NOR4_X1 U6138 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n5409)
         );
  OAI21_X1 U6139 ( .B1(n5411), .B2(n5410), .A(n5409), .ZN(n5414) );
  XOR2_X1 U6140 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_207), .Z(n5413) );
  XNOR2_X1 U6141 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_208), .ZN(n5412)
         );
  AOI21_X1 U6142 ( .B1(n5414), .B2(n5413), .A(n5412), .ZN(n5420) );
  INV_X1 U6143 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7077) );
  XNOR2_X1 U6144 ( .A(n7077), .B(keyinput_209), .ZN(n5416) );
  INV_X1 U6145 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7076) );
  XNOR2_X1 U6146 ( .A(n7076), .B(keyinput_210), .ZN(n5415) );
  NAND2_X1 U6147 ( .A1(n5416), .A2(n5415), .ZN(n5419) );
  XOR2_X1 U6148 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_211), .Z(n5418) );
  XNOR2_X1 U6149 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_212), .ZN(n5417)
         );
  OAI211_X1 U6150 ( .C1(n5420), .C2(n5419), .A(n5418), .B(n5417), .ZN(n5426)
         );
  XNOR2_X1 U6151 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_213), .ZN(n5425)
         );
  XOR2_X1 U6152 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .Z(n5423) );
  XOR2_X1 U6153 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_214), .Z(n5422) );
  XNOR2_X1 U6154 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_215), .ZN(n5421)
         );
  NAND3_X1 U6155 ( .A1(n5423), .A2(n5422), .A3(n5421), .ZN(n5424) );
  AOI21_X1 U6156 ( .B1(n5426), .B2(n5425), .A(n5424), .ZN(n5434) );
  XNOR2_X1 U6157 ( .A(ADDRESS_REG_7__SCAN_IN), .B(keyinput_221), .ZN(n5433) );
  XNOR2_X1 U6158 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_217), .ZN(n5432)
         );
  XNOR2_X1 U6159 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_218), .ZN(n5430)
         );
  XNOR2_X1 U6160 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n5429) );
  XNOR2_X1 U6161 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_220), .ZN(n5428) );
  XNOR2_X1 U6162 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_222), .ZN(n5427) );
  NAND4_X1 U6163 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n5431)
         );
  NOR4_X1 U6164 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n5443)
         );
  INV_X1 U6165 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7058) );
  XNOR2_X1 U6166 ( .A(n7058), .B(keyinput_223), .ZN(n5442) );
  XOR2_X1 U6167 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_224), .Z(n5440) );
  XOR2_X1 U6168 ( .A(keyinput_227), .B(ADDRESS_REG_1__SCAN_IN), .Z(n5439) );
  XNOR2_X1 U6169 ( .A(keyinput_228), .B(ADDRESS_REG_0__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U6170 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_225), .ZN(n5436) );
  XNOR2_X1 U6171 ( .A(keyinput_226), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n5435) );
  NAND3_X1 U6172 ( .A1(n5437), .A2(n5436), .A3(n5435), .ZN(n5438) );
  NOR3_X1 U6173 ( .A1(n5440), .A2(n5439), .A3(n5438), .ZN(n5441) );
  OAI21_X1 U6174 ( .B1(n5443), .B2(n5442), .A(n5441), .ZN(n5454) );
  XNOR2_X1 U6175 ( .A(n6998), .B(keyinput_229), .ZN(n5453) );
  XNOR2_X1 U6176 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_235), .ZN(n5445)
         );
  XNOR2_X1 U6177 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_234), .ZN(n5444)
         );
  NOR2_X1 U6178 ( .A1(n5445), .A2(n5444), .ZN(n5451) );
  XNOR2_X1 U6179 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .ZN(n5447)
         );
  XNOR2_X1 U6180 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_231), .ZN(n5446) );
  NOR2_X1 U6181 ( .A1(n5447), .A2(n5446), .ZN(n5450) );
  XNOR2_X1 U6182 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_230), .ZN(n5449) );
  XNOR2_X1 U6183 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_232), .ZN(n5448)
         );
  NAND4_X1 U6184 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n5452)
         );
  AOI21_X1 U6185 ( .B1(n5454), .B2(n5453), .A(n5452), .ZN(n5457) );
  INV_X1 U6186 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7002) );
  XNOR2_X1 U6187 ( .A(n7002), .B(keyinput_237), .ZN(n5456) );
  XNOR2_X1 U6188 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_236), .ZN(n5455)
         );
  NOR3_X1 U6189 ( .A1(n5457), .A2(n5456), .A3(n5455), .ZN(n5465) );
  INV_X1 U6190 ( .A(keyinput_240), .ZN(n5458) );
  XNOR2_X1 U6191 ( .A(n5458), .B(DATAWIDTH_REG_8__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U6192 ( .A(DATAWIDTH_REG_6__SCAN_IN), .B(keyinput_238), .ZN(n5461)
         );
  XNOR2_X1 U6193 ( .A(DATAWIDTH_REG_9__SCAN_IN), .B(keyinput_241), .ZN(n5460)
         );
  XNOR2_X1 U6194 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_239), .ZN(n5459)
         );
  NAND4_X1 U6195 ( .A1(n5462), .A2(n5461), .A3(n5460), .A4(n5459), .ZN(n5464)
         );
  XOR2_X1 U6196 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_242), .Z(n5463)
         );
  OAI21_X1 U6197 ( .B1(n5465), .B2(n5464), .A(n5463), .ZN(n5477) );
  INV_X1 U6198 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7008) );
  XNOR2_X1 U6199 ( .A(n7008), .B(keyinput_246), .ZN(n5469) );
  INV_X1 U6200 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7007) );
  XNOR2_X1 U6201 ( .A(n7007), .B(keyinput_245), .ZN(n5468) );
  INV_X1 U6202 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7006) );
  XNOR2_X1 U6203 ( .A(n7006), .B(keyinput_243), .ZN(n5467) );
  XNOR2_X1 U6204 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_244), .ZN(n5466)
         );
  NOR4_X1 U6205 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n5476)
         );
  INV_X1 U6206 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7010) );
  AOI22_X1 U6207 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput_247), .B1(
        n7010), .B2(keyinput_250), .ZN(n5470) );
  OAI221_X1 U6208 ( .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput_247), .C1(
        n7010), .C2(keyinput_250), .A(n5470), .ZN(n5474) );
  INV_X1 U6209 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U6210 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(keyinput_249), .B1(
        n7011), .B2(keyinput_251), .ZN(n5471) );
  OAI221_X1 U6211 ( .B1(DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_249), .C1(
        n7011), .C2(keyinput_251), .A(n5471), .ZN(n5473) );
  XNOR2_X1 U6212 ( .A(DATAWIDTH_REG_16__SCAN_IN), .B(keyinput_248), .ZN(n5472)
         );
  OR3_X1 U6213 ( .A1(n5474), .A2(n5473), .A3(n5472), .ZN(n5475) );
  AOI21_X1 U6214 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5480) );
  XNOR2_X1 U6215 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_252), .ZN(n5479)
         );
  XNOR2_X1 U6216 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_253), .ZN(n5478)
         );
  OAI21_X1 U6217 ( .B1(n5480), .B2(n5479), .A(n5478), .ZN(n5666) );
  XNOR2_X1 U6218 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .ZN(n5665)
         );
  XOR2_X1 U6219 ( .A(DATAI_30_), .B(keyinput_1), .Z(n5483) );
  XOR2_X1 U6220 ( .A(DATAI_31_), .B(keyinput_0), .Z(n5482) );
  XNOR2_X1 U6221 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n5481) );
  NAND3_X1 U6222 ( .A1(n5483), .A2(n5482), .A3(n5481), .ZN(n5486) );
  XOR2_X1 U6223 ( .A(DATAI_27_), .B(keyinput_4), .Z(n5485) );
  XOR2_X1 U6224 ( .A(DATAI_28_), .B(keyinput_3), .Z(n5484) );
  NAND3_X1 U6225 ( .A1(n5486), .A2(n5485), .A3(n5484), .ZN(n5489) );
  XNOR2_X1 U6226 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n5488) );
  XNOR2_X1 U6227 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n5487) );
  NAND3_X1 U6228 ( .A1(n5489), .A2(n5488), .A3(n5487), .ZN(n5493) );
  XOR2_X1 U6229 ( .A(DATAI_24_), .B(keyinput_7), .Z(n5492) );
  XNOR2_X1 U6230 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n5491) );
  XNOR2_X1 U6231 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n5490) );
  NAND4_X1 U6232 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n5496)
         );
  XOR2_X1 U6233 ( .A(DATAI_21_), .B(keyinput_10), .Z(n5495) );
  XOR2_X1 U6234 ( .A(DATAI_20_), .B(keyinput_11), .Z(n5494) );
  AOI21_X1 U6235 ( .B1(n5496), .B2(n5495), .A(n5494), .ZN(n5509) );
  XNOR2_X1 U6236 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n5508) );
  INV_X1 U6237 ( .A(DATAI_16_), .ZN(n5497) );
  INV_X1 U6238 ( .A(DATAI_14_), .ZN(n6350) );
  OAI22_X1 U6239 ( .A1(keyinput_15), .A2(n5497), .B1(n6350), .B2(keyinput_17), 
        .ZN(n5505) );
  OAI22_X1 U6240 ( .A1(DATAI_13_), .A2(keyinput_18), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n5504) );
  INV_X1 U6241 ( .A(DATAI_12_), .ZN(n6327) );
  NOR2_X1 U6242 ( .A1(n6327), .A2(keyinput_19), .ZN(n5503) );
  AOI22_X1 U6243 ( .A1(n5497), .A2(keyinput_15), .B1(n6327), .B2(keyinput_19), 
        .ZN(n5500) );
  AOI22_X1 U6244 ( .A1(DATAI_17_), .A2(keyinput_14), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n5499) );
  AOI22_X1 U6245 ( .A1(DATAI_13_), .A2(keyinput_18), .B1(n6350), .B2(
        keyinput_17), .ZN(n5498) );
  AND3_X1 U6246 ( .A1(n5500), .A2(n5499), .A3(n5498), .ZN(n5501) );
  OAI21_X1 U6247 ( .B1(DATAI_17_), .B2(keyinput_14), .A(n5501), .ZN(n5502) );
  NOR4_X1 U6248 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n5507)
         );
  XNOR2_X1 U6249 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n5506) );
  OAI211_X1 U6250 ( .C1(n5509), .C2(n5508), .A(n5507), .B(n5506), .ZN(n5512)
         );
  XNOR2_X1 U6251 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n5511) );
  XNOR2_X1 U6252 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n5510) );
  AOI21_X1 U6253 ( .B1(n5512), .B2(n5511), .A(n5510), .ZN(n5515) );
  XOR2_X1 U6254 ( .A(DATAI_9_), .B(keyinput_22), .Z(n5514) );
  XNOR2_X1 U6255 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n5513) );
  NOR3_X1 U6256 ( .A1(n5515), .A2(n5514), .A3(n5513), .ZN(n5519) );
  XOR2_X1 U6257 ( .A(DATAI_6_), .B(keyinput_25), .Z(n5518) );
  XOR2_X1 U6258 ( .A(DATAI_5_), .B(keyinput_26), .Z(n5517) );
  XNOR2_X1 U6259 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n5516) );
  NOR4_X1 U6260 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .ZN(n5523)
         );
  XOR2_X1 U6261 ( .A(DATAI_2_), .B(keyinput_29), .Z(n5522) );
  XNOR2_X1 U6262 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n5521) );
  XNOR2_X1 U6263 ( .A(DATAI_3_), .B(keyinput_28), .ZN(n5520) );
  NOR4_X1 U6264 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n5527)
         );
  XOR2_X1 U6265 ( .A(DATAI_1_), .B(keyinput_30), .Z(n5526) );
  XNOR2_X1 U6266 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_32), .ZN(n5525) );
  XNOR2_X1 U6267 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n5524) );
  OAI211_X1 U6268 ( .C1(n5527), .C2(n5526), .A(n5525), .B(n5524), .ZN(n5530)
         );
  XNOR2_X1 U6269 ( .A(NA_N), .B(keyinput_33), .ZN(n5529) );
  XNOR2_X1 U6270 ( .A(BS16_N), .B(keyinput_34), .ZN(n5528) );
  AOI21_X1 U6271 ( .B1(n5530), .B2(n5529), .A(n5528), .ZN(n5533) );
  XNOR2_X1 U6272 ( .A(n7546), .B(keyinput_35), .ZN(n5532) );
  XNOR2_X1 U6273 ( .A(HOLD), .B(keyinput_36), .ZN(n5531) );
  NOR3_X1 U6274 ( .A1(n5533), .A2(n5532), .A3(n5531), .ZN(n5536) );
  XNOR2_X1 U6275 ( .A(n7017), .B(keyinput_38), .ZN(n5535) );
  XOR2_X1 U6276 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_37), .Z(n5534) );
  NOR3_X1 U6277 ( .A1(n5536), .A2(n5535), .A3(n5534), .ZN(n5539) );
  XOR2_X1 U6278 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_39), .Z(n5538) );
  XNOR2_X1 U6279 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_40), .ZN(n5537) );
  NOR3_X1 U6280 ( .A1(n5539), .A2(n5538), .A3(n5537), .ZN(n5543) );
  XNOR2_X1 U6281 ( .A(n7535), .B(keyinput_43), .ZN(n5542) );
  XNOR2_X1 U6282 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_42), .ZN(n5541)
         );
  XNOR2_X1 U6283 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n5540) );
  NOR4_X1 U6284 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n5546)
         );
  XOR2_X1 U6285 ( .A(MORE_REG_SCAN_IN), .B(keyinput_44), .Z(n5545) );
  XNOR2_X1 U6286 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_45), .ZN(n5544) );
  NOR3_X1 U6287 ( .A1(n5546), .A2(n5545), .A3(n5544), .ZN(n5560) );
  INV_X1 U6288 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7193) );
  XNOR2_X1 U6289 ( .A(n7193), .B(keyinput_46), .ZN(n5559) );
  OAI22_X1 U6290 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_54), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_47), .ZN(n5548) );
  AND2_X1 U6291 ( .A1(keyinput_47), .A2(BYTEENABLE_REG_0__SCAN_IN), .ZN(n5547)
         );
  AOI211_X1 U6292 ( .C1(REIP_REG_28__SCAN_IN), .C2(keyinput_54), .A(n5548), 
        .B(n5547), .ZN(n5552) );
  XOR2_X1 U6293 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_50), .Z(n5551) );
  XNOR2_X1 U6294 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .ZN(n5550) );
  XNOR2_X1 U6295 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .ZN(n5549) );
  NAND4_X1 U6296 ( .A1(n5552), .A2(n5551), .A3(n5550), .A4(n5549), .ZN(n5557)
         );
  INV_X1 U6297 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7121) );
  AOI22_X1 U6298 ( .A1(n7121), .A2(keyinput_48), .B1(n7096), .B2(keyinput_52), 
        .ZN(n5553) );
  OAI221_X1 U6299 ( .B1(n7121), .B2(keyinput_48), .C1(n7096), .C2(keyinput_52), 
        .A(n5553), .ZN(n5556) );
  XNOR2_X1 U6300 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n5555) );
  XNOR2_X1 U6301 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_49), .ZN(n5554)
         );
  NOR4_X1 U6302 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n5558)
         );
  OAI21_X1 U6303 ( .B1(n5560), .B2(n5559), .A(n5558), .ZN(n5563) );
  XNOR2_X1 U6304 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n5562) );
  XNOR2_X1 U6305 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .ZN(n5561) );
  AOI21_X1 U6306 ( .B1(n5563), .B2(n5562), .A(n5561), .ZN(n5566) );
  XOR2_X1 U6307 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .Z(n5565) );
  XOR2_X1 U6308 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .Z(n5564) );
  OAI21_X1 U6309 ( .B1(n5566), .B2(n5565), .A(n5564), .ZN(n5569) );
  XNOR2_X1 U6310 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .ZN(n5568) );
  XNOR2_X1 U6311 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n5567) );
  AOI21_X1 U6312 ( .B1(n5569), .B2(n5568), .A(n5567), .ZN(n5573) );
  XOR2_X1 U6313 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .Z(n5572) );
  XOR2_X1 U6314 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .Z(n5571) );
  XNOR2_X1 U6315 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .ZN(n5570) );
  OAI211_X1 U6316 ( .C1(n5573), .C2(n5572), .A(n5571), .B(n5570), .ZN(n5576)
         );
  XOR2_X1 U6317 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_65), .Z(n5575) );
  XNOR2_X1 U6318 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .ZN(n5574) );
  AOI21_X1 U6319 ( .B1(n5576), .B2(n5575), .A(n5574), .ZN(n5594) );
  INV_X1 U6320 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7122) );
  XNOR2_X1 U6321 ( .A(n7122), .B(keyinput_70), .ZN(n5580) );
  INV_X1 U6322 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7100) );
  XNOR2_X1 U6323 ( .A(n7100), .B(keyinput_67), .ZN(n5579) );
  INV_X1 U6324 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7118) );
  XNOR2_X1 U6325 ( .A(n7118), .B(keyinput_69), .ZN(n5578) );
  XNOR2_X1 U6326 ( .A(BE_N_REG_2__SCAN_IN), .B(keyinput_68), .ZN(n5577) );
  NAND4_X1 U6327 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n5593)
         );
  INV_X1 U6328 ( .A(keyinput_76), .ZN(n5586) );
  AOI22_X1 U6329 ( .A1(n7081), .A2(keyinput_78), .B1(keyinput_72), .B2(n7093), 
        .ZN(n5584) );
  INV_X1 U6330 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7084) );
  AOI22_X1 U6331 ( .A1(n7097), .A2(keyinput_71), .B1(keyinput_77), .B2(n7084), 
        .ZN(n5583) );
  AOI22_X1 U6332 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput_76), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput_75), .ZN(n5582) );
  AOI22_X1 U6333 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(keyinput_73), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(keyinput_74), .ZN(n5581) );
  NAND4_X1 U6334 ( .A1(n5584), .A2(n5583), .A3(n5582), .A4(n5581), .ZN(n5585)
         );
  AOI21_X1 U6335 ( .B1(n7085), .B2(n5586), .A(n5585), .ZN(n5587) );
  OAI21_X1 U6336 ( .B1(keyinput_71), .B2(n7097), .A(n5587), .ZN(n5591) );
  OAI22_X1 U6337 ( .A1(keyinput_78), .A2(n7081), .B1(n7084), .B2(keyinput_77), 
        .ZN(n5590) );
  OAI22_X1 U6338 ( .A1(n7093), .A2(keyinput_72), .B1(ADDRESS_REG_26__SCAN_IN), 
        .B2(keyinput_74), .ZN(n5589) );
  OAI22_X1 U6339 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_75), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(keyinput_73), .ZN(n5588) );
  NOR4_X1 U6340 ( .A1(n5591), .A2(n5590), .A3(n5589), .A4(n5588), .ZN(n5592)
         );
  OAI21_X1 U6341 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n5597) );
  XOR2_X1 U6342 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_79), .Z(n5596) );
  XNOR2_X1 U6343 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_80), .ZN(n5595) );
  AOI21_X1 U6344 ( .B1(n5597), .B2(n5596), .A(n5595), .ZN(n5600) );
  XNOR2_X1 U6345 ( .A(n7076), .B(keyinput_82), .ZN(n5599) );
  XNOR2_X1 U6346 ( .A(n7077), .B(keyinput_81), .ZN(n5598) );
  NOR3_X1 U6347 ( .A1(n5600), .A2(n5599), .A3(n5598), .ZN(n5603) );
  XNOR2_X1 U6348 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_83), .ZN(n5602) );
  XNOR2_X1 U6349 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_84), .ZN(n5601) );
  NOR3_X1 U6350 ( .A1(n5603), .A2(n5602), .A3(n5601), .ZN(n5609) );
  INV_X1 U6351 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7072) );
  XNOR2_X1 U6352 ( .A(n7072), .B(keyinput_85), .ZN(n5608) );
  XNOR2_X1 U6353 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_87), .ZN(n5606) );
  XNOR2_X1 U6354 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_88), .ZN(n5605) );
  XNOR2_X1 U6355 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_86), .ZN(n5604) );
  NOR3_X1 U6356 ( .A1(n5606), .A2(n5605), .A3(n5604), .ZN(n5607) );
  OAI21_X1 U6357 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5617) );
  XOR2_X1 U6358 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_89), .Z(n5616) );
  XOR2_X1 U6359 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .Z(n5615) );
  INV_X1 U6360 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7062) );
  XNOR2_X1 U6361 ( .A(n7062), .B(keyinput_92), .ZN(n5613) );
  XNOR2_X1 U6362 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_94), .ZN(n5612) );
  XNOR2_X1 U6363 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_91), .ZN(n5611) );
  XNOR2_X1 U6364 ( .A(ADDRESS_REG_7__SCAN_IN), .B(keyinput_93), .ZN(n5610) );
  NOR4_X1 U6365 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5614)
         );
  NAND4_X1 U6366 ( .A1(n5617), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(n5619)
         );
  XNOR2_X1 U6367 ( .A(n7058), .B(keyinput_95), .ZN(n5618) );
  NAND2_X1 U6368 ( .A1(n5619), .A2(n5618), .ZN(n5625) );
  OAI22_X1 U6369 ( .A1(ADDRESS_REG_0__SCAN_IN), .A2(keyinput_100), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(keyinput_98), .ZN(n5620) );
  AOI221_X1 U6370 ( .B1(ADDRESS_REG_0__SCAN_IN), .B2(keyinput_100), .C1(
        keyinput_98), .C2(ADDRESS_REG_2__SCAN_IN), .A(n5620), .ZN(n5624) );
  XOR2_X1 U6371 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_96), .Z(n5623) );
  INV_X1 U6372 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7053) );
  OAI22_X1 U6373 ( .A1(n7053), .A2(keyinput_99), .B1(ADDRESS_REG_3__SCAN_IN), 
        .B2(keyinput_97), .ZN(n5621) );
  AOI221_X1 U6374 ( .B1(n7053), .B2(keyinput_99), .C1(keyinput_97), .C2(
        ADDRESS_REG_3__SCAN_IN), .A(n5621), .ZN(n5622) );
  NAND4_X1 U6375 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n5635)
         );
  XNOR2_X1 U6376 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .ZN(n5634) );
  XOR2_X1 U6377 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_104), .Z(n5629) );
  XNOR2_X1 U6378 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_107), .ZN(n5628)
         );
  XNOR2_X1 U6379 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .ZN(n5627)
         );
  XNOR2_X1 U6380 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_106), .ZN(n5626)
         );
  NOR4_X1 U6381 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n5632)
         );
  XOR2_X1 U6382 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .Z(n5631) );
  XNOR2_X1 U6383 ( .A(n7547), .B(keyinput_103), .ZN(n5630) );
  NAND3_X1 U6384 ( .A1(n5632), .A2(n5631), .A3(n5630), .ZN(n5633) );
  AOI21_X1 U6385 ( .B1(n5635), .B2(n5634), .A(n5633), .ZN(n5638) );
  INV_X1 U6386 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7001) );
  XNOR2_X1 U6387 ( .A(n7001), .B(keyinput_108), .ZN(n5637) );
  XNOR2_X1 U6388 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_109), .ZN(n5636)
         );
  NOR3_X1 U6389 ( .A1(n5638), .A2(n5637), .A3(n5636), .ZN(n5645) );
  XOR2_X1 U6390 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_112), .Z(n5642) );
  INV_X1 U6391 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7005) );
  XNOR2_X1 U6392 ( .A(n7005), .B(keyinput_113), .ZN(n5641) );
  INV_X1 U6393 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7003) );
  XNOR2_X1 U6394 ( .A(n7003), .B(keyinput_110), .ZN(n5640) );
  INV_X1 U6395 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7004) );
  XNOR2_X1 U6396 ( .A(n7004), .B(keyinput_111), .ZN(n5639) );
  NAND4_X1 U6397 ( .A1(n5642), .A2(n5641), .A3(n5640), .A4(n5639), .ZN(n5644)
         );
  XNOR2_X1 U6398 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_114), .ZN(n5643)
         );
  OAI21_X1 U6399 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5657) );
  XNOR2_X1 U6400 ( .A(n7007), .B(keyinput_117), .ZN(n5649) );
  XNOR2_X1 U6401 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_118), .ZN(n5648)
         );
  XNOR2_X1 U6402 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_115), .ZN(n5647)
         );
  XNOR2_X1 U6403 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_116), .ZN(n5646)
         );
  NOR4_X1 U6404 ( .A1(n5649), .A2(n5648), .A3(n5647), .A4(n5646), .ZN(n5656)
         );
  OAI22_X1 U6405 ( .A1(n7010), .A2(keyinput_122), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_123), .ZN(n5650) );
  AOI221_X1 U6406 ( .B1(n7010), .B2(keyinput_122), .C1(keyinput_123), .C2(
        DATAWIDTH_REG_19__SCAN_IN), .A(n5650), .ZN(n5654) );
  INV_X1 U6407 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7009) );
  OAI22_X1 U6408 ( .A1(n7009), .A2(keyinput_119), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput_120), .ZN(n5651) );
  AOI221_X1 U6409 ( .B1(n7009), .B2(keyinput_119), .C1(keyinput_120), .C2(
        DATAWIDTH_REG_16__SCAN_IN), .A(n5651), .ZN(n5653) );
  XOR2_X1 U6410 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_121), .Z(n5652)
         );
  NAND3_X1 U6411 ( .A1(n5654), .A2(n5653), .A3(n5652), .ZN(n5655) );
  AOI21_X1 U6412 ( .B1(n5657), .B2(n5656), .A(n5655), .ZN(n5660) );
  XNOR2_X1 U6413 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_124), .ZN(n5659)
         );
  XNOR2_X1 U6414 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .ZN(n5658)
         );
  OAI21_X1 U6415 ( .B1(n5660), .B2(n5659), .A(n5658), .ZN(n5663) );
  XNOR2_X1 U6416 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_126), .ZN(n5662)
         );
  XNOR2_X1 U6417 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_127), .ZN(n5661)
         );
  AOI21_X1 U6418 ( .B1(n5663), .B2(n5662), .A(n5661), .ZN(n5664) );
  AOI211_X1 U6419 ( .C1(n5667), .C2(n5666), .A(n5665), .B(n5664), .ZN(n5669)
         );
  INV_X1 U6420 ( .A(n7095), .ZN(n7068) );
  NOR2_X1 U6421 ( .A1(n7553), .A2(STATE_REG_2__SCAN_IN), .ZN(n7069) );
  AOI222_X1 U6422 ( .A1(n7553), .A2(ADDRESS_REG_10__SCAN_IN), .B1(n7068), .B2(
        REIP_REG_11__SCAN_IN), .C1(REIP_REG_12__SCAN_IN), .C2(n7069), .ZN(
        n5668) );
  XNOR2_X1 U6423 ( .A(n5669), .B(n5668), .ZN(U3194) );
  NAND2_X1 U6424 ( .A1(n7588), .A2(n5052), .ZN(n6786) );
  INV_X1 U6425 ( .A(n6786), .ZN(n5671) );
  NOR2_X1 U6426 ( .A1(n5678), .A2(n7535), .ZN(n5681) );
  AOI211_X1 U6427 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5671), .A(n5909), .B(
        n5681), .ZN(n5677) );
  NOR3_X1 U6428 ( .A1(n6082), .A2(n5672), .A3(n6853), .ZN(n5673) );
  AOI21_X1 U6429 ( .B1(n6082), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n5673), 
        .ZN(n5676) );
  NAND2_X1 U6430 ( .A1(n5674), .A2(n6703), .ZN(n5675) );
  OAI211_X1 U6431 ( .C1(n5677), .C2(n5821), .A(n5676), .B(n5675), .ZN(U3462)
         );
  NOR2_X1 U6432 ( .A1(n6784), .A2(n5684), .ZN(n6928) );
  AOI21_X1 U6433 ( .B1(n5680), .B2(n5679), .A(n6928), .ZN(n5686) );
  NOR2_X1 U6434 ( .A1(n5681), .A2(n7587), .ZN(n5683) );
  AOI22_X1 U6435 ( .A1(n5686), .A2(n5683), .B1(n7587), .B2(n5684), .ZN(n5682)
         );
  NAND2_X1 U6436 ( .A1(n7602), .A2(n5682), .ZN(n6927) );
  INV_X1 U6437 ( .A(n5683), .ZN(n5685) );
  OAI22_X1 U6438 ( .A1(n5686), .A2(n5685), .B1(n7200), .B2(n5684), .ZN(n6926)
         );
  AOI22_X1 U6439 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6927), .B1(n6809), 
        .B2(n6926), .ZN(n5688) );
  AOI22_X1 U6440 ( .A1(n6929), .A2(n7623), .B1(n7622), .B2(n6928), .ZN(n5687)
         );
  OAI211_X1 U6441 ( .C1(n6876), .C2(n6932), .A(n5688), .B(n5687), .ZN(U3127)
         );
  AOI22_X1 U6442 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6927), .B1(n6816), 
        .B2(n6926), .ZN(n5690) );
  AOI22_X1 U6443 ( .A1(n6929), .A2(n7636), .B1(n7634), .B2(n6928), .ZN(n5689)
         );
  OAI211_X1 U6444 ( .C1(n6883), .C2(n6932), .A(n5690), .B(n5689), .ZN(U3129)
         );
  AOI22_X1 U6445 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6927), .B1(n6798), 
        .B2(n6926), .ZN(n5692) );
  AOI22_X1 U6446 ( .A1(n6929), .A2(n7597), .B1(n7596), .B2(n6928), .ZN(n5691)
         );
  OAI211_X1 U6447 ( .C1(n6865), .C2(n6932), .A(n5692), .B(n5691), .ZN(U3124)
         );
  AOI22_X1 U6448 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6927), .B1(n6805), 
        .B2(n6926), .ZN(n5694) );
  AOI22_X1 U6449 ( .A1(n6929), .A2(n7618), .B1(n7616), .B2(n6928), .ZN(n5693)
         );
  OAI211_X1 U6450 ( .C1(n6872), .C2(n6932), .A(n5694), .B(n5693), .ZN(U3126)
         );
  AOI22_X1 U6451 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6927), .B1(n6825), 
        .B2(n6926), .ZN(n5696) );
  AOI22_X1 U6452 ( .A1(n6929), .A2(n7651), .B1(n7647), .B2(n6928), .ZN(n5695)
         );
  OAI211_X1 U6453 ( .C1(n6893), .C2(n6932), .A(n5696), .B(n5695), .ZN(U3131)
         );
  AOI22_X1 U6454 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6927), .B1(n6820), 
        .B2(n6926), .ZN(n5698) );
  AOI22_X1 U6455 ( .A1(n6929), .A2(n7642), .B1(n7640), .B2(n6928), .ZN(n5697)
         );
  OAI211_X1 U6456 ( .C1(n6887), .C2(n6932), .A(n5698), .B(n5697), .ZN(U3130)
         );
  OR2_X1 U6457 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  AND2_X1 U6458 ( .A1(n5699), .A2(n5702), .ZN(n7371) );
  INV_X1 U6459 ( .A(n7371), .ZN(n5705) );
  INV_X1 U6460 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5703) );
  OAI21_X1 U6461 ( .B1(n3682), .B2(n3740), .A(n5994), .ZN(n7369) );
  OAI222_X1 U6462 ( .A1(n5705), .A2(n7127), .B1(n5703), .B2(n7143), .C1(n6304), 
        .C2(n7369), .ZN(U2852) );
  OAI222_X1 U6463 ( .A1(n5705), .A2(n6354), .B1(n6356), .B2(n5704), .C1(n7564), 
        .C2(n4314), .ZN(U2884) );
  INV_X1 U6464 ( .A(n6853), .ZN(n5707) );
  NAND2_X1 U6465 ( .A1(n7590), .A2(n7599), .ZN(n6787) );
  AOI211_X1 U6466 ( .C1(n6797), .C2(n6787), .A(n6951), .B(n6939), .ZN(n5706)
         );
  AOI21_X1 U6467 ( .B1(n7590), .B2(n5707), .A(n5706), .ZN(n5711) );
  NOR2_X1 U6468 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5708), .ZN(n6938)
         );
  INV_X1 U6469 ( .A(n6938), .ZN(n5709) );
  AND2_X1 U6470 ( .A1(n6707), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6855)
         );
  NOR2_X1 U6471 ( .A1(n6855), .A2(n5906), .ZN(n6859) );
  AOI211_X1 U6472 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5709), .A(n6859), .B(
        n6789), .ZN(n5710) );
  INV_X1 U6473 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5715) );
  INV_X1 U6474 ( .A(n6855), .ZN(n5712) );
  OAI22_X1 U6475 ( .A1(n6788), .A2(n7590), .B1(n6796), .B2(n5712), .ZN(n6937)
         );
  AOI22_X1 U6476 ( .A1(n7647), .A2(n6938), .B1(n6825), .B2(n6937), .ZN(n5714)
         );
  AOI22_X1 U6477 ( .A1(n7651), .A2(n6939), .B1(n6951), .B2(n7648), .ZN(n5713)
         );
  OAI211_X1 U6478 ( .C1(n6943), .C2(n5715), .A(n5714), .B(n5713), .ZN(U3139)
         );
  INV_X1 U6479 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5718) );
  AOI22_X1 U6480 ( .A1(n7634), .A2(n6938), .B1(n6816), .B2(n6937), .ZN(n5717)
         );
  AOI22_X1 U6481 ( .A1(n7636), .A2(n6939), .B1(n6951), .B2(n7635), .ZN(n5716)
         );
  OAI211_X1 U6482 ( .C1(n6943), .C2(n5718), .A(n5717), .B(n5716), .ZN(U3137)
         );
  INV_X1 U6483 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5721) );
  AOI22_X1 U6484 ( .A1(n7616), .A2(n6938), .B1(n6805), .B2(n6937), .ZN(n5720)
         );
  AOI22_X1 U6485 ( .A1(n7618), .A2(n6939), .B1(n6951), .B2(n7617), .ZN(n5719)
         );
  OAI211_X1 U6486 ( .C1(n6943), .C2(n5721), .A(n5720), .B(n5719), .ZN(U3134)
         );
  INV_X1 U6487 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5724) );
  AOI22_X1 U6488 ( .A1(n7596), .A2(n6938), .B1(n6798), .B2(n6937), .ZN(n5723)
         );
  AOI22_X1 U6489 ( .A1(n7597), .A2(n6939), .B1(n6951), .B2(n7606), .ZN(n5722)
         );
  OAI211_X1 U6490 ( .C1(n6943), .C2(n5724), .A(n5723), .B(n5722), .ZN(U3132)
         );
  INV_X1 U6491 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5727) );
  AOI22_X1 U6492 ( .A1(n7622), .A2(n6938), .B1(n6809), .B2(n6937), .ZN(n5726)
         );
  AOI22_X1 U6493 ( .A1(n7623), .A2(n6939), .B1(n6951), .B2(n7624), .ZN(n5725)
         );
  OAI211_X1 U6494 ( .C1(n6943), .C2(n5727), .A(n5726), .B(n5725), .ZN(U3135)
         );
  INV_X1 U6495 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5730) );
  AOI22_X1 U6496 ( .A1(n7640), .A2(n6938), .B1(n6820), .B2(n6937), .ZN(n5729)
         );
  AOI22_X1 U6497 ( .A1(n7642), .A2(n6939), .B1(n6951), .B2(n7641), .ZN(n5728)
         );
  OAI211_X1 U6498 ( .C1(n6943), .C2(n5730), .A(n5729), .B(n5728), .ZN(U3138)
         );
  NAND2_X1 U6499 ( .A1(n5733), .A2(n3925), .ZN(n5731) );
  NAND2_X1 U6500 ( .A1(n5733), .A2(n5732), .ZN(n7326) );
  INV_X1 U6501 ( .A(n6215), .ZN(n6245) );
  AOI22_X1 U6502 ( .A1(n7490), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6245), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5738) );
  AND2_X1 U6503 ( .A1(n5734), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5735) );
  INV_X1 U6504 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6505 ( .A1(n7483), .A2(n5736), .ZN(n5737) );
  OAI211_X1 U6506 ( .C1(n7326), .C2(n5047), .A(n5738), .B(n5737), .ZN(n5739)
         );
  AOI21_X1 U6507 ( .B1(n7412), .B2(n4974), .A(n5739), .ZN(n5746) );
  INV_X1 U6508 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7114) );
  NAND3_X1 U6509 ( .A1(n3645), .A2(n6260), .A3(n5740), .ZN(n5741) );
  AND2_X1 U6510 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  AOI22_X1 U6511 ( .A1(n7333), .A2(n7114), .B1(n3617), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5745) );
  OAI211_X1 U6512 ( .C1(n7319), .C2(n5987), .A(n5746), .B(n5745), .ZN(U2826)
         );
  NAND2_X1 U6513 ( .A1(n5795), .A2(n7599), .ZN(n5788) );
  AOI211_X1 U6514 ( .C1(n6797), .C2(n5788), .A(n7649), .B(n6841), .ZN(n5752)
         );
  NOR2_X1 U6515 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5747), .ZN(n6837)
         );
  NOR2_X1 U6516 ( .A1(n6837), .A2(n7533), .ZN(n5751) );
  NAND2_X1 U6517 ( .A1(n5748), .A2(n6796), .ZN(n6860) );
  INV_X1 U6518 ( .A(n6860), .ZN(n5749) );
  NOR4_X2 U6519 ( .A1(n5752), .A2(n5751), .A3(n5791), .A4(n3741), .ZN(n6844)
         );
  INV_X1 U6520 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5757) );
  OAI22_X1 U6521 ( .A1(n6788), .A2(n5795), .B1(n6711), .B2(n5753), .ZN(n6836)
         );
  AOI22_X1 U6522 ( .A1(n7616), .A2(n6837), .B1(n6805), .B2(n6836), .ZN(n5754)
         );
  OAI21_X1 U6523 ( .B1(n6723), .B2(n6839), .A(n5754), .ZN(n5755) );
  AOI21_X1 U6524 ( .B1(n6841), .B2(n7617), .A(n5755), .ZN(n5756) );
  OAI21_X1 U6525 ( .B1(n6844), .B2(n5757), .A(n5756), .ZN(U3086) );
  INV_X1 U6526 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5761) );
  AOI22_X1 U6527 ( .A1(n7622), .A2(n6837), .B1(n6809), .B2(n6836), .ZN(n5758)
         );
  OAI21_X1 U6528 ( .B1(n6728), .B2(n6839), .A(n5758), .ZN(n5759) );
  AOI21_X1 U6529 ( .B1(n6841), .B2(n7624), .A(n5759), .ZN(n5760) );
  OAI21_X1 U6530 ( .B1(n6844), .B2(n5761), .A(n5760), .ZN(U3087) );
  INV_X1 U6531 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5765) );
  AOI22_X1 U6532 ( .A1(n7640), .A2(n6837), .B1(n6820), .B2(n6836), .ZN(n5762)
         );
  OAI21_X1 U6533 ( .B1(n6742), .B2(n6839), .A(n5762), .ZN(n5763) );
  AOI21_X1 U6534 ( .B1(n6841), .B2(n7641), .A(n5763), .ZN(n5764) );
  OAI21_X1 U6535 ( .B1(n6844), .B2(n5765), .A(n5764), .ZN(U3090) );
  INV_X1 U6536 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5769) );
  AOI22_X1 U6537 ( .A1(n7647), .A2(n6837), .B1(n6825), .B2(n6836), .ZN(n5766)
         );
  OAI21_X1 U6538 ( .B1(n6749), .B2(n6839), .A(n5766), .ZN(n5767) );
  AOI21_X1 U6539 ( .B1(n6841), .B2(n7648), .A(n5767), .ZN(n5768) );
  OAI21_X1 U6540 ( .B1(n6844), .B2(n5769), .A(n5768), .ZN(U3091) );
  INV_X1 U6541 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5773) );
  AOI22_X1 U6542 ( .A1(n7634), .A2(n6837), .B1(n6816), .B2(n6836), .ZN(n5770)
         );
  OAI21_X1 U6543 ( .B1(n6737), .B2(n6839), .A(n5770), .ZN(n5771) );
  AOI21_X1 U6544 ( .B1(n6841), .B2(n7635), .A(n5771), .ZN(n5772) );
  OAI21_X1 U6545 ( .B1(n6844), .B2(n5773), .A(n5772), .ZN(U3089) );
  INV_X1 U6546 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5777) );
  AOI22_X1 U6547 ( .A1(n7596), .A2(n6837), .B1(n6798), .B2(n6836), .ZN(n5774)
         );
  OAI21_X1 U6548 ( .B1(n6714), .B2(n6839), .A(n5774), .ZN(n5775) );
  AOI21_X1 U6549 ( .B1(n6841), .B2(n7606), .A(n5775), .ZN(n5776) );
  OAI21_X1 U6550 ( .B1(n6844), .B2(n5777), .A(n5776), .ZN(U3084) );
  INV_X1 U6551 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U6552 ( .A1(n7138), .A2(n5779), .ZN(n5781) );
  NAND2_X1 U6553 ( .A1(n5781), .A2(n5780), .ZN(n5783) );
  NAND2_X1 U6554 ( .A1(n5783), .A2(n5782), .ZN(n7359) );
  INV_X1 U6555 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5785) );
  XOR2_X1 U6556 ( .A(n5028), .B(n5784), .Z(n7354) );
  INV_X1 U6557 ( .A(n7354), .ZN(n5786) );
  OAI222_X1 U6558 ( .A1(n7359), .A2(n6304), .B1(n5785), .B2(n7143), .C1(n7127), 
        .C2(n5786), .ZN(U2853) );
  OAI222_X1 U6559 ( .A1(n5787), .A2(n6356), .B1(n7564), .B2(n4308), .C1(n6354), 
        .C2(n5786), .ZN(U2885) );
  AOI211_X1 U6560 ( .C1(n6788), .C2(n5788), .A(n6952), .B(n6686), .ZN(n5793)
         );
  NOR2_X1 U6561 ( .A1(n5824), .A2(n5789), .ZN(n6682) );
  NOR2_X1 U6562 ( .A1(n7533), .A2(n6682), .ZN(n5792) );
  OAI21_X1 U6563 ( .B1(n5830), .B2(n6707), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n5790) );
  INV_X1 U6564 ( .A(n5790), .ZN(n5826) );
  NOR4_X2 U6565 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5826), .ZN(n6689)
         );
  INV_X1 U6566 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5799) );
  INV_X1 U6567 ( .A(n6711), .ZN(n6856) );
  NAND2_X1 U6568 ( .A1(n6856), .A2(n5831), .ZN(n5794) );
  OAI22_X1 U6569 ( .A1(n6797), .A2(n5795), .B1(n5830), .B2(n5794), .ZN(n6681)
         );
  AOI22_X1 U6570 ( .A1(n7616), .A2(n6682), .B1(n6805), .B2(n6681), .ZN(n5796)
         );
  OAI21_X1 U6571 ( .B1(n6684), .B2(n6723), .A(n5796), .ZN(n5797) );
  AOI21_X1 U6572 ( .B1(n7617), .B2(n6686), .A(n5797), .ZN(n5798) );
  OAI21_X1 U6573 ( .B1(n6689), .B2(n5799), .A(n5798), .ZN(U3022) );
  INV_X1 U6574 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5803) );
  AOI22_X1 U6575 ( .A1(n7596), .A2(n6682), .B1(n6798), .B2(n6681), .ZN(n5800)
         );
  OAI21_X1 U6576 ( .B1(n6684), .B2(n6714), .A(n5800), .ZN(n5801) );
  AOI21_X1 U6577 ( .B1(n7606), .B2(n6686), .A(n5801), .ZN(n5802) );
  OAI21_X1 U6578 ( .B1(n6689), .B2(n5803), .A(n5802), .ZN(U3020) );
  INV_X1 U6579 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5807) );
  AOI22_X1 U6580 ( .A1(n7634), .A2(n6682), .B1(n6816), .B2(n6681), .ZN(n5804)
         );
  OAI21_X1 U6581 ( .B1(n6684), .B2(n6737), .A(n5804), .ZN(n5805) );
  AOI21_X1 U6582 ( .B1(n7635), .B2(n6686), .A(n5805), .ZN(n5806) );
  OAI21_X1 U6583 ( .B1(n6689), .B2(n5807), .A(n5806), .ZN(U3025) );
  INV_X1 U6584 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5811) );
  AOI22_X1 U6585 ( .A1(n7640), .A2(n6682), .B1(n6820), .B2(n6681), .ZN(n5808)
         );
  OAI21_X1 U6586 ( .B1(n6684), .B2(n6742), .A(n5808), .ZN(n5809) );
  AOI21_X1 U6587 ( .B1(n7641), .B2(n6686), .A(n5809), .ZN(n5810) );
  OAI21_X1 U6588 ( .B1(n6689), .B2(n5811), .A(n5810), .ZN(U3026) );
  INV_X1 U6589 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5815) );
  AOI22_X1 U6590 ( .A1(n7647), .A2(n6682), .B1(n6825), .B2(n6681), .ZN(n5812)
         );
  OAI21_X1 U6591 ( .B1(n6684), .B2(n6749), .A(n5812), .ZN(n5813) );
  AOI21_X1 U6592 ( .B1(n7648), .B2(n6686), .A(n5813), .ZN(n5814) );
  OAI21_X1 U6593 ( .B1(n6689), .B2(n5815), .A(n5814), .ZN(U3027) );
  INV_X1 U6594 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5819) );
  AOI22_X1 U6595 ( .A1(n7622), .A2(n6682), .B1(n6809), .B2(n6681), .ZN(n5816)
         );
  OAI21_X1 U6596 ( .B1(n6684), .B2(n6728), .A(n5816), .ZN(n5817) );
  AOI21_X1 U6597 ( .B1(n7624), .B2(n6686), .A(n5817), .ZN(n5818) );
  OAI21_X1 U6598 ( .B1(n6689), .B2(n5819), .A(n5818), .ZN(U3023) );
  XNOR2_X1 U6599 ( .A(n5052), .B(STATEBS16_REG_SCAN_IN), .ZN(n5820) );
  OAI222_X1 U6600 ( .A1(n6085), .A2(n5047), .B1(n5821), .B2(n5820), .C1(n6967), 
        .C2(n7015), .ZN(U3464) );
  INV_X1 U6601 ( .A(n6772), .ZN(n5822) );
  AOI211_X1 U6602 ( .C1(n6788), .C2(n5823), .A(n6769), .B(n5822), .ZN(n5828)
         );
  NOR2_X1 U6603 ( .A1(n5824), .A2(n7591), .ZN(n6768) );
  NOR2_X1 U6604 ( .A1(n7533), .A2(n6768), .ZN(n5827) );
  OR2_X1 U6605 ( .A1(n5829), .A2(n6797), .ZN(n5835) );
  INV_X1 U6606 ( .A(n5830), .ZN(n5833) );
  INV_X1 U6607 ( .A(n6796), .ZN(n5832) );
  NAND3_X1 U6608 ( .A1(n5833), .A2(n5832), .A3(n5831), .ZN(n5834) );
  NAND2_X1 U6609 ( .A1(n5835), .A2(n5834), .ZN(n6767) );
  AOI22_X1 U6610 ( .A1(n7596), .A2(n6768), .B1(n6798), .B2(n6767), .ZN(n5837)
         );
  NAND2_X1 U6611 ( .A1(n6769), .A2(n7606), .ZN(n5836) );
  OAI211_X1 U6612 ( .C1(n6772), .C2(n6714), .A(n5837), .B(n5836), .ZN(n5838)
         );
  AOI21_X1 U6613 ( .B1(n6774), .B2(INSTQUEUE_REG_4__0__SCAN_IN), .A(n5838), 
        .ZN(n5839) );
  INV_X1 U6614 ( .A(n5839), .ZN(U3052) );
  AOI22_X1 U6615 ( .A1(n7640), .A2(n6768), .B1(n6820), .B2(n6767), .ZN(n5841)
         );
  NAND2_X1 U6616 ( .A1(n6769), .A2(n7641), .ZN(n5840) );
  OAI211_X1 U6617 ( .C1(n6772), .C2(n6742), .A(n5841), .B(n5840), .ZN(n5842)
         );
  AOI21_X1 U6618 ( .B1(n6774), .B2(INSTQUEUE_REG_4__6__SCAN_IN), .A(n5842), 
        .ZN(n5843) );
  INV_X1 U6619 ( .A(n5843), .ZN(U3058) );
  AOI22_X1 U6620 ( .A1(n7616), .A2(n6768), .B1(n6805), .B2(n6767), .ZN(n5845)
         );
  NAND2_X1 U6621 ( .A1(n6769), .A2(n7617), .ZN(n5844) );
  OAI211_X1 U6622 ( .C1(n6772), .C2(n6723), .A(n5845), .B(n5844), .ZN(n5846)
         );
  AOI21_X1 U6623 ( .B1(n6774), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n5846), 
        .ZN(n5847) );
  INV_X1 U6624 ( .A(n5847), .ZN(U3054) );
  AOI22_X1 U6625 ( .A1(n7622), .A2(n6768), .B1(n6809), .B2(n6767), .ZN(n5849)
         );
  NAND2_X1 U6626 ( .A1(n6769), .A2(n7624), .ZN(n5848) );
  OAI211_X1 U6627 ( .C1(n6772), .C2(n6728), .A(n5849), .B(n5848), .ZN(n5850)
         );
  AOI21_X1 U6628 ( .B1(n6774), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n5850), 
        .ZN(n5851) );
  INV_X1 U6629 ( .A(n5851), .ZN(U3055) );
  AOI22_X1 U6630 ( .A1(n7647), .A2(n6768), .B1(n6825), .B2(n6767), .ZN(n5853)
         );
  NAND2_X1 U6631 ( .A1(n6769), .A2(n7648), .ZN(n5852) );
  OAI211_X1 U6632 ( .C1(n6772), .C2(n6749), .A(n5853), .B(n5852), .ZN(n5854)
         );
  AOI21_X1 U6633 ( .B1(n6774), .B2(INSTQUEUE_REG_4__7__SCAN_IN), .A(n5854), 
        .ZN(n5855) );
  INV_X1 U6634 ( .A(n5855), .ZN(U3059) );
  AOI22_X1 U6635 ( .A1(n7634), .A2(n6768), .B1(n6816), .B2(n6767), .ZN(n5857)
         );
  NAND2_X1 U6636 ( .A1(n6769), .A2(n7635), .ZN(n5856) );
  OAI211_X1 U6637 ( .C1(n6772), .C2(n6737), .A(n5857), .B(n5856), .ZN(n5858)
         );
  AOI21_X1 U6638 ( .B1(n6774), .B2(INSTQUEUE_REG_4__5__SCAN_IN), .A(n5858), 
        .ZN(n5859) );
  INV_X1 U6639 ( .A(n5859), .ZN(U3057) );
  NAND2_X1 U6640 ( .A1(n5893), .A2(DATAI_0_), .ZN(n5871) );
  AOI22_X1 U6641 ( .A1(n5933), .A2(EAX_REG_16__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U6642 ( .A1(n5871), .A2(n5861), .ZN(U2924) );
  AOI22_X1 U6643 ( .A1(n5933), .A2(EAX_REG_11__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6644 ( .A1(n5863), .A2(n5862), .ZN(U2950) );
  AOI22_X1 U6645 ( .A1(n5933), .A2(EAX_REG_6__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U6646 ( .A1(n5865), .A2(n5864), .ZN(U2945) );
  AOI22_X1 U6647 ( .A1(n5933), .A2(EAX_REG_7__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U6648 ( .A1(n5867), .A2(n5866), .ZN(U2946) );
  AOI22_X1 U6649 ( .A1(n5933), .A2(EAX_REG_8__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6650 ( .A1(n5869), .A2(n5868), .ZN(U2947) );
  AOI22_X1 U6651 ( .A1(n5933), .A2(EAX_REG_0__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6652 ( .A1(n5871), .A2(n5870), .ZN(U2939) );
  NAND2_X1 U6653 ( .A1(n5893), .A2(DATAI_1_), .ZN(n5877) );
  AOI22_X1 U6654 ( .A1(n5933), .A2(EAX_REG_1__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U6655 ( .A1(n5877), .A2(n5872), .ZN(U2940) );
  NAND2_X1 U6656 ( .A1(n5893), .A2(DATAI_2_), .ZN(n5879) );
  AOI22_X1 U6657 ( .A1(n5933), .A2(EAX_REG_2__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6658 ( .A1(n5879), .A2(n5873), .ZN(U2941) );
  NAND2_X1 U6659 ( .A1(n5893), .A2(DATAI_13_), .ZN(n5882) );
  AOI22_X1 U6660 ( .A1(n5933), .A2(EAX_REG_13__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U6661 ( .A1(n5882), .A2(n5874), .ZN(U2952) );
  NAND2_X1 U6662 ( .A1(n5893), .A2(DATAI_3_), .ZN(n5889) );
  AOI22_X1 U6663 ( .A1(n5933), .A2(EAX_REG_3__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6664 ( .A1(n5889), .A2(n5875), .ZN(U2942) );
  AOI22_X1 U6665 ( .A1(n5933), .A2(EAX_REG_17__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6666 ( .A1(n5877), .A2(n5876), .ZN(U2925) );
  AOI22_X1 U6667 ( .A1(n5933), .A2(EAX_REG_18__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6668 ( .A1(n5879), .A2(n5878), .ZN(U2926) );
  NAND2_X1 U6669 ( .A1(n5893), .A2(DATAI_12_), .ZN(n5897) );
  AOI22_X1 U6670 ( .A1(n5933), .A2(EAX_REG_28__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U6671 ( .A1(n5897), .A2(n5880), .ZN(U2936) );
  AOI22_X1 U6672 ( .A1(n5933), .A2(EAX_REG_29__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U6673 ( .A1(n5882), .A2(n5881), .ZN(U2937) );
  NAND2_X1 U6674 ( .A1(n5893), .A2(DATAI_14_), .ZN(n5891) );
  AOI22_X1 U6675 ( .A1(n5933), .A2(EAX_REG_30__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U6676 ( .A1(n5891), .A2(n5883), .ZN(U2938) );
  AOI22_X1 U6677 ( .A1(n5933), .A2(EAX_REG_9__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U6678 ( .A1(n5885), .A2(n5884), .ZN(U2948) );
  AOI22_X1 U6679 ( .A1(n5933), .A2(EAX_REG_10__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U6680 ( .A1(n5887), .A2(n5886), .ZN(U2949) );
  AOI22_X1 U6681 ( .A1(n5933), .A2(EAX_REG_19__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6682 ( .A1(n5889), .A2(n5888), .ZN(U2927) );
  AOI22_X1 U6683 ( .A1(n5933), .A2(EAX_REG_14__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U6684 ( .A1(n5891), .A2(n5890), .ZN(U2953) );
  NAND2_X1 U6685 ( .A1(n5893), .A2(DATAI_4_), .ZN(n5899) );
  AOI22_X1 U6686 ( .A1(n5894), .A2(EAX_REG_20__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U6687 ( .A1(n5899), .A2(n5892), .ZN(U2928) );
  NAND2_X1 U6688 ( .A1(n5893), .A2(DATAI_5_), .ZN(n5901) );
  AOI22_X1 U6689 ( .A1(n5894), .A2(EAX_REG_21__SCAN_IN), .B1(n5932), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6690 ( .A1(n5901), .A2(n5895), .ZN(U2929) );
  AOI22_X1 U6691 ( .A1(n5933), .A2(EAX_REG_12__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6692 ( .A1(n5897), .A2(n5896), .ZN(U2951) );
  AOI22_X1 U6693 ( .A1(n5933), .A2(EAX_REG_4__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6694 ( .A1(n5899), .A2(n5898), .ZN(U2943) );
  AOI22_X1 U6695 ( .A1(n5933), .A2(EAX_REG_5__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U6696 ( .A1(n5901), .A2(n5900), .ZN(U2944) );
  INV_X1 U6697 ( .A(n5909), .ZN(n5902) );
  OAI21_X1 U6698 ( .B1(n5052), .B2(n7587), .A(n6853), .ZN(n7585) );
  AOI21_X1 U6699 ( .B1(n5902), .B2(n7599), .A(n7585), .ZN(n5910) );
  AND2_X1 U6700 ( .A1(n5903), .A2(n6703), .ZN(n6858) );
  NAND3_X1 U6701 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5904), .ZN(n6857) );
  NOR2_X1 U6702 ( .A1(n6784), .A2(n6857), .ZN(n6903) );
  AOI21_X1 U6703 ( .B1(n6858), .B2(n5905), .A(n6903), .ZN(n5912) );
  OAI22_X1 U6704 ( .A1(n5910), .A2(n5912), .B1(n6857), .B2(n5906), .ZN(n5907)
         );
  INV_X1 U6705 ( .A(n6805), .ZN(n7621) );
  AND2_X1 U6706 ( .A1(n5052), .A2(n5057), .ZN(n5908) );
  INV_X1 U6707 ( .A(n5910), .ZN(n5911) );
  AOI22_X1 U6708 ( .A1(n5912), .A2(n5911), .B1(n6857), .B2(n7587), .ZN(n5913)
         );
  NAND2_X1 U6709 ( .A1(n7602), .A2(n5913), .ZN(n6902) );
  AOI22_X1 U6710 ( .A1(n7616), .A2(n6903), .B1(INSTQUEUE_REG_11__2__SCAN_IN), 
        .B2(n6902), .ZN(n5914) );
  OAI21_X1 U6711 ( .B1(n6723), .B2(n6905), .A(n5914), .ZN(n5915) );
  AOI21_X1 U6712 ( .B1(n7617), .B2(n6919), .A(n5915), .ZN(n5916) );
  OAI21_X1 U6713 ( .B1(n6909), .B2(n7621), .A(n5916), .ZN(U3110) );
  INV_X1 U6714 ( .A(n6820), .ZN(n7645) );
  AOI22_X1 U6715 ( .A1(n7640), .A2(n6903), .B1(INSTQUEUE_REG_11__6__SCAN_IN), 
        .B2(n6902), .ZN(n5917) );
  OAI21_X1 U6716 ( .B1(n6742), .B2(n6905), .A(n5917), .ZN(n5918) );
  AOI21_X1 U6717 ( .B1(n7641), .B2(n6919), .A(n5918), .ZN(n5919) );
  OAI21_X1 U6718 ( .B1(n6909), .B2(n7645), .A(n5919), .ZN(U3114) );
  INV_X1 U6719 ( .A(n6809), .ZN(n7627) );
  AOI22_X1 U6720 ( .A1(n7622), .A2(n6903), .B1(INSTQUEUE_REG_11__3__SCAN_IN), 
        .B2(n6902), .ZN(n5920) );
  OAI21_X1 U6721 ( .B1(n6728), .B2(n6905), .A(n5920), .ZN(n5921) );
  AOI21_X1 U6722 ( .B1(n7624), .B2(n6919), .A(n5921), .ZN(n5922) );
  OAI21_X1 U6723 ( .B1(n6909), .B2(n7627), .A(n5922), .ZN(U3111) );
  INV_X1 U6724 ( .A(n6798), .ZN(n7609) );
  AOI22_X1 U6725 ( .A1(n7596), .A2(n6903), .B1(INSTQUEUE_REG_11__0__SCAN_IN), 
        .B2(n6902), .ZN(n5923) );
  OAI21_X1 U6726 ( .B1(n6714), .B2(n6905), .A(n5923), .ZN(n5924) );
  AOI21_X1 U6727 ( .B1(n7606), .B2(n6919), .A(n5924), .ZN(n5925) );
  OAI21_X1 U6728 ( .B1(n6909), .B2(n7609), .A(n5925), .ZN(U3108) );
  INV_X1 U6729 ( .A(n6825), .ZN(n7655) );
  AOI22_X1 U6730 ( .A1(n7647), .A2(n6903), .B1(INSTQUEUE_REG_11__7__SCAN_IN), 
        .B2(n6902), .ZN(n5926) );
  OAI21_X1 U6731 ( .B1(n6749), .B2(n6905), .A(n5926), .ZN(n5927) );
  AOI21_X1 U6732 ( .B1(n7648), .B2(n6919), .A(n5927), .ZN(n5928) );
  OAI21_X1 U6733 ( .B1(n6909), .B2(n7655), .A(n5928), .ZN(U3115) );
  INV_X1 U6734 ( .A(n6816), .ZN(n7639) );
  AOI22_X1 U6735 ( .A1(n7634), .A2(n6903), .B1(INSTQUEUE_REG_11__5__SCAN_IN), 
        .B2(n6902), .ZN(n5929) );
  OAI21_X1 U6736 ( .B1(n6737), .B2(n6905), .A(n5929), .ZN(n5930) );
  AOI21_X1 U6737 ( .B1(n7635), .B2(n6919), .A(n5930), .ZN(n5931) );
  OAI21_X1 U6738 ( .B1(n6909), .B2(n7639), .A(n5931), .ZN(U3113) );
  AOI22_X1 U6739 ( .A1(n5933), .A2(EAX_REG_15__SCAN_IN), .B1(n5932), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5934) );
  OAI21_X1 U6740 ( .B1(n5935), .B2(n6347), .A(n5934), .ZN(U2954) );
  NAND3_X1 U6741 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        n6215), .ZN(n5937) );
  OAI21_X1 U6742 ( .B1(n7054), .B2(n5937), .A(n6217), .ZN(n7327) );
  AOI22_X1 U6743 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7490), .B1(
        EBX_REG_3__SCAN_IN), .B2(n3617), .ZN(n5936) );
  OAI221_X1 U6744 ( .B1(n7327), .B2(n7054), .C1(n7327), .C2(n5937), .A(n5936), 
        .ZN(n5938) );
  INV_X1 U6745 ( .A(n5938), .ZN(n5943) );
  INV_X1 U6746 ( .A(n6703), .ZN(n5939) );
  OAI22_X1 U6747 ( .A1(n7326), .A2(n5939), .B1(n7491), .B2(n5964), .ZN(n5940)
         );
  AOI21_X1 U6748 ( .B1(n7412), .B2(n5941), .A(n5940), .ZN(n5942) );
  OAI211_X1 U6749 ( .C1(n7319), .C2(n5944), .A(n5943), .B(n5942), .ZN(U2824)
         );
  INV_X1 U6750 ( .A(n5945), .ZN(n5946) );
  OAI21_X1 U6751 ( .B1(n3662), .B2(n5947), .A(n5946), .ZN(n7391) );
  NOR2_X1 U6752 ( .A1(n5993), .A2(n5948), .ZN(n5949) );
  OR2_X1 U6753 ( .A1(n5979), .A2(n5949), .ZN(n7387) );
  INV_X1 U6754 ( .A(n7387), .ZN(n5950) );
  AOI22_X1 U6755 ( .A1(n7139), .A2(n5950), .B1(EBX_REG_9__SCAN_IN), .B2(n6314), 
        .ZN(n5951) );
  OAI21_X1 U6756 ( .B1(n7391), .B2(n7127), .A(n5951), .ZN(U2850) );
  XNOR2_X1 U6757 ( .A(n5952), .B(n5953), .ZN(n5972) );
  NAND2_X1 U6758 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U6759 ( .A1(n5954), .A2(n7227), .ZN(n7238) );
  NAND3_X1 U6760 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n7238), .ZN(n6502) );
  INV_X1 U6761 ( .A(n7256), .ZN(n7296) );
  NOR2_X1 U6762 ( .A1(n7227), .A2(n5955), .ZN(n7223) );
  NAND3_X1 U6763 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n7223), .ZN(n6498) );
  AOI22_X1 U6764 ( .A1(n7298), .A2(n6502), .B1(n7296), .B2(n6498), .ZN(n5956)
         );
  NAND2_X1 U6765 ( .A1(n7300), .A2(n5956), .ZN(n6626) );
  INV_X1 U6766 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7364) );
  OAI22_X1 U6767 ( .A1(n7301), .A2(n7369), .B1(n7364), .B2(n7248), .ZN(n5957)
         );
  AOI21_X1 U6768 ( .B1(n6626), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5957), 
        .ZN(n5959) );
  NOR2_X1 U6769 ( .A1(n7230), .A2(n6502), .ZN(n6039) );
  NAND2_X1 U6770 ( .A1(n6039), .A2(n5990), .ZN(n5958) );
  OAI211_X1 U6771 ( .C1(n5972), .C2(n7240), .A(n5959), .B(n5958), .ZN(U3011)
         );
  INV_X1 U6772 ( .A(DATAI_8_), .ZN(n6338) );
  INV_X1 U6773 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7035) );
  XOR2_X1 U6774 ( .A(n5699), .B(n5960), .Z(n7383) );
  INV_X1 U6775 ( .A(n7383), .ZN(n5961) );
  OAI222_X1 U6776 ( .A1(n6356), .A2(n6338), .B1(n7564), .B2(n7035), .C1(n6354), 
        .C2(n5961), .ZN(U2883) );
  INV_X1 U6777 ( .A(DATAI_9_), .ZN(n5962) );
  INV_X1 U6778 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7037) );
  OAI222_X1 U6779 ( .A1(n6356), .A2(n5962), .B1(n7564), .B2(n7037), .C1(n6354), 
        .C2(n7391), .ZN(U2882) );
  AOI22_X1 U6780 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n7280), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U6781 ( .B1(n7190), .B2(n5964), .A(n5963), .ZN(n5965) );
  AOI21_X1 U6782 ( .B1(n5966), .B2(n7185), .A(n5965), .ZN(n5967) );
  OAI21_X1 U6783 ( .B1(n5968), .B2(n7501), .A(n5967), .ZN(U2983) );
  AOI22_X1 U6784 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n7280), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n5969) );
  OAI21_X1 U6785 ( .B1(n7190), .B2(n7374), .A(n5969), .ZN(n5970) );
  AOI21_X1 U6786 ( .B1(n7371), .B2(n7185), .A(n5970), .ZN(n5971) );
  OAI21_X1 U6787 ( .B1(n5972), .B2(n7501), .A(n5971), .ZN(U2979) );
  INV_X1 U6788 ( .A(n5973), .ZN(n5974) );
  NOR2_X1 U6789 ( .A1(n5945), .A2(n5975), .ZN(n5976) );
  OR2_X1 U6790 ( .A1(n5974), .A2(n5976), .ZN(n6239) );
  OR2_X1 U6791 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND2_X1 U6792 ( .A1(n5977), .A2(n5980), .ZN(n6248) );
  INV_X1 U6793 ( .A(n6248), .ZN(n7267) );
  AOI22_X1 U6794 ( .A1(n7139), .A2(n7267), .B1(EBX_REG_10__SCAN_IN), .B2(n6314), .ZN(n5981) );
  OAI21_X1 U6795 ( .B1(n6239), .B2(n7127), .A(n5981), .ZN(U2849) );
  NOR2_X1 U6796 ( .A1(n7190), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5982)
         );
  AOI211_X1 U6797 ( .C1(n7183), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5983), 
        .B(n5982), .ZN(n5986) );
  NAND2_X1 U6798 ( .A1(n5984), .A2(n7186), .ZN(n5985) );
  OAI211_X1 U6799 ( .C1(n7174), .C2(n5987), .A(n5986), .B(n5985), .ZN(U2985)
         );
  XNOR2_X1 U6800 ( .A(n3642), .B(n5989), .ZN(n6032) );
  NOR2_X1 U6801 ( .A1(n5991), .A2(n5990), .ZN(n6497) );
  AOI21_X1 U6802 ( .B1(n5991), .B2(n5990), .A(n6497), .ZN(n5992) );
  AOI22_X1 U6803 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n6626), .B1(n6039), 
        .B2(n5992), .ZN(n5998) );
  AOI21_X1 U6804 ( .B1(n5995), .B2(n5994), .A(n5993), .ZN(n7377) );
  INV_X1 U6805 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5996) );
  NOR2_X1 U6806 ( .A1(n7248), .A2(n5996), .ZN(n6028) );
  AOI21_X1 U6807 ( .B1(n7313), .B2(n7377), .A(n6028), .ZN(n5997) );
  OAI211_X1 U6808 ( .C1(n6032), .C2(n7240), .A(n5998), .B(n5997), .ZN(U3010)
         );
  INV_X1 U6809 ( .A(DATAI_10_), .ZN(n6333) );
  INV_X1 U6810 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7039) );
  OAI222_X1 U6811 ( .A1(n6356), .A2(n6333), .B1(n7564), .B2(n7039), .C1(n6354), 
        .C2(n6239), .ZN(U2881) );
  NOR2_X1 U6812 ( .A1(n5974), .A2(n6001), .ZN(n6002) );
  OR2_X1 U6813 ( .A1(n6000), .A2(n6002), .ZN(n7175) );
  NAND2_X1 U6814 ( .A1(n5977), .A2(n6003), .ZN(n6004) );
  NAND2_X1 U6815 ( .A1(n6021), .A2(n6004), .ZN(n6657) );
  INV_X1 U6816 ( .A(n6657), .ZN(n6005) );
  AOI22_X1 U6817 ( .A1(n7139), .A2(n6005), .B1(EBX_REG_11__SCAN_IN), .B2(n6314), .ZN(n6006) );
  OAI21_X1 U6818 ( .B1(n7175), .B2(n7127), .A(n6006), .ZN(U2848) );
  OAI21_X1 U6819 ( .B1(n7473), .B2(n6007), .A(n6215), .ZN(n7403) );
  OAI21_X1 U6820 ( .B1(n7473), .B2(n6018), .A(n7064), .ZN(n6014) );
  INV_X1 U6821 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6012) );
  OAI22_X1 U6822 ( .A1(n6008), .A2(n7476), .B1(n7493), .B2(n6657), .ZN(n6010)
         );
  NAND2_X1 U6823 ( .A1(n6009), .A2(n6215), .ZN(n7423) );
  AOI211_X1 U6824 ( .C1(n7483), .C2(n7172), .A(n6010), .B(n7449), .ZN(n6011)
         );
  OAI21_X1 U6825 ( .B1(n6012), .B2(n7478), .A(n6011), .ZN(n6013) );
  AOI21_X1 U6826 ( .B1(n7403), .B2(n6014), .A(n6013), .ZN(n6015) );
  OAI21_X1 U6827 ( .B1(n7175), .B2(n7467), .A(n6015), .ZN(U2816) );
  OAI21_X1 U6828 ( .B1(n6000), .B2(n6017), .A(n6016), .ZN(n6489) );
  INV_X1 U6829 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U6830 ( .A1(n7410), .A2(n6019), .ZN(n6020) );
  OAI21_X1 U6831 ( .B1(n6491), .B2(n7491), .A(n6020), .ZN(n6025) );
  INV_X1 U6832 ( .A(n6647), .ZN(n6639) );
  AOI21_X1 U6833 ( .B1(n6022), .B2(n6021), .A(n6639), .ZN(n7278) );
  AOI22_X1 U6834 ( .A1(EBX_REG_12__SCAN_IN), .A2(n3617), .B1(n7412), .B2(n7278), .ZN(n6023) );
  OAI211_X1 U6835 ( .C1(n7478), .C2(n4386), .A(n6023), .B(n7423), .ZN(n6024)
         );
  AOI211_X1 U6836 ( .C1(REIP_REG_12__SCAN_IN), .C2(n7403), .A(n6025), .B(n6024), .ZN(n6026) );
  OAI21_X1 U6837 ( .B1(n6489), .B2(n7467), .A(n6026), .ZN(U2815) );
  AOI22_X1 U6838 ( .A1(n7139), .A2(n7278), .B1(EBX_REG_12__SCAN_IN), .B2(n6314), .ZN(n6027) );
  OAI21_X1 U6839 ( .B1(n6489), .B2(n7127), .A(n6027), .ZN(U2847) );
  INV_X1 U6840 ( .A(DATAI_11_), .ZN(n6330) );
  INV_X1 U6841 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7041) );
  OAI222_X1 U6842 ( .A1(n6356), .A2(n6330), .B1(n7564), .B2(n7041), .C1(n6354), 
        .C2(n7175), .ZN(U2880) );
  AOI21_X1 U6843 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6028), 
        .ZN(n6029) );
  OAI21_X1 U6844 ( .B1(n7190), .B2(n7381), .A(n6029), .ZN(n6030) );
  AOI21_X1 U6845 ( .B1(n7383), .B2(n7185), .A(n6030), .ZN(n6031) );
  OAI21_X1 U6846 ( .B1(n6032), .B2(n7501), .A(n6031), .ZN(U2978) );
  INV_X1 U6847 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7043) );
  OAI222_X1 U6848 ( .A1(n6356), .A2(n6327), .B1(n7564), .B2(n7043), .C1(n6354), 
        .C2(n6489), .ZN(U2879) );
  XOR2_X1 U6849 ( .A(n6033), .B(n6034), .Z(n6040) );
  NAND2_X1 U6850 ( .A1(n6040), .A2(n7186), .ZN(n6038) );
  INV_X1 U6851 ( .A(n7190), .ZN(n6466) );
  INV_X1 U6852 ( .A(n7183), .ZN(n6464) );
  INV_X1 U6853 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U6854 ( .A1(n7280), .A2(REIP_REG_9__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U6855 ( .B1(n6464), .B2(n6035), .A(n6042), .ZN(n6036) );
  AOI21_X1 U6856 ( .B1(n6466), .B2(n7392), .A(n6036), .ZN(n6037) );
  OAI211_X1 U6857 ( .C1(n7174), .C2(n7391), .A(n6038), .B(n6037), .ZN(U2977)
         );
  NAND2_X1 U6858 ( .A1(n6497), .A2(n6039), .ZN(n7273) );
  NAND2_X1 U6859 ( .A1(n6040), .A2(n7314), .ZN(n6045) );
  INV_X1 U6860 ( .A(n6626), .ZN(n6041) );
  OAI21_X1 U6861 ( .B1(n6497), .B2(n6628), .A(n6041), .ZN(n7268) );
  OAI21_X1 U6862 ( .B1(n7301), .B2(n7387), .A(n6042), .ZN(n6043) );
  AOI21_X1 U6863 ( .B1(n7268), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6043), 
        .ZN(n6044) );
  OAI211_X1 U6864 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n7273), .A(n6045), 
        .B(n6044), .ZN(U3009) );
  MUX2_X1 U6865 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .B(n6046), .S(n6444), 
        .Z(n6047) );
  XNOR2_X1 U6866 ( .A(n6048), .B(n6047), .ZN(n7269) );
  NAND2_X1 U6867 ( .A1(n7269), .A2(n7186), .ZN(n6052) );
  INV_X1 U6868 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6049) );
  NOR2_X1 U6869 ( .A1(n7248), .A2(n6049), .ZN(n7266) );
  NOR2_X1 U6870 ( .A1(n7190), .A2(n6247), .ZN(n6050) );
  AOI211_X1 U6871 ( .C1(n7183), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7266), 
        .B(n6050), .ZN(n6051) );
  OAI211_X1 U6872 ( .C1(n7174), .C2(n6239), .A(n6052), .B(n6051), .ZN(U2976)
         );
  XNOR2_X2 U6873 ( .A(n6067), .B(n6054), .ZN(n6319) );
  INV_X1 U6874 ( .A(n6319), .ZN(n6126) );
  INV_X1 U6875 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6059) );
  INV_X1 U6876 ( .A(n6055), .ZN(n6056) );
  OAI22_X1 U6877 ( .A1(n6069), .A2(n4789), .B1(n6056), .B2(n6131), .ZN(n6057)
         );
  OAI222_X1 U6878 ( .A1(n7127), .A2(n6126), .B1(n6059), .B2(n7143), .C1(n6527), 
        .C2(n6304), .ZN(U2829) );
  NAND2_X1 U6879 ( .A1(n6062), .A2(n6061), .ZN(n6065) );
  INV_X1 U6880 ( .A(n3908), .ZN(n6063) );
  AOI22_X1 U6881 ( .A1(n7578), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7581), .ZN(n6064) );
  NAND2_X1 U6882 ( .A1(n6065), .A2(n6064), .ZN(U2860) );
  OAI21_X1 U6883 ( .B1(n6066), .B2(n6068), .A(n6067), .ZN(n6322) );
  AOI21_X1 U6884 ( .B1(n6070), .B2(n6131), .A(n6069), .ZN(n6538) );
  AOI22_X1 U6885 ( .A1(n6538), .A2(n7139), .B1(EBX_REG_29__SCAN_IN), .B2(n6314), .ZN(n6071) );
  OAI21_X1 U6886 ( .B1(n6322), .B2(n7127), .A(n6071), .ZN(U2830) );
  NAND3_X1 U6887 ( .A1(n6135), .A2(REIP_REG_28__SCAN_IN), .A3(n7094), .ZN(
        n6076) );
  INV_X1 U6888 ( .A(n6072), .ZN(n6361) );
  OAI22_X1 U6889 ( .A1(n6073), .A2(n7478), .B1(n7491), .B2(n6361), .ZN(n6074)
         );
  AOI21_X1 U6890 ( .B1(n3617), .B2(EBX_REG_29__SCAN_IN), .A(n6074), .ZN(n6075)
         );
  OAI211_X1 U6891 ( .C1(n6137), .C2(n7094), .A(n6076), .B(n6075), .ZN(n6077)
         );
  AOI21_X1 U6892 ( .B1(n6538), .B2(n7412), .A(n6077), .ZN(n6078) );
  OAI21_X1 U6893 ( .B1(n6322), .B2(n7467), .A(n6078), .ZN(U2798) );
  NAND2_X1 U6894 ( .A1(n7015), .A2(n7585), .ZN(n6081) );
  NAND3_X1 U6895 ( .A1(n6079), .A2(STATEBS16_REG_SCAN_IN), .A3(n5052), .ZN(
        n6080) );
  MUX2_X1 U6896 ( .A(n6081), .B(n6080), .S(n5050), .Z(n6084) );
  NAND2_X1 U6897 ( .A1(n6082), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6083) );
  OAI211_X1 U6898 ( .C1(n6090), .C2(n6085), .A(n6084), .B(n6083), .ZN(U3463)
         );
  OR2_X1 U6899 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  AND2_X1 U6900 ( .A1(n6089), .A2(n6088), .ZN(n7247) );
  INV_X1 U6901 ( .A(n7326), .ZN(n6091) );
  AOI22_X1 U6902 ( .A1(n6091), .A2(n4050), .B1(n3617), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n6097) );
  AOI22_X1 U6903 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7490), .B1(n6245), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U6904 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6092) );
  OAI211_X1 U6905 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n7333), .B(n6092), .ZN(n6095) );
  INV_X1 U6906 ( .A(n7155), .ZN(n6093) );
  NAND2_X1 U6907 ( .A1(n7483), .A2(n6093), .ZN(n6094) );
  NAND4_X1 U6908 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n6098)
         );
  AOI21_X1 U6909 ( .B1(n7412), .B2(n7247), .A(n6098), .ZN(n6099) );
  OAI21_X1 U6910 ( .B1(n7319), .B2(n7126), .A(n6099), .ZN(U2825) );
  XNOR2_X1 U6911 ( .A(n6104), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6531)
         );
  INV_X1 U6912 ( .A(n6105), .ZN(n6119) );
  AND2_X1 U6913 ( .A1(n7280), .A2(REIP_REG_30__SCAN_IN), .ZN(n6525) );
  AOI21_X1 U6914 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6525), 
        .ZN(n6106) );
  OAI21_X1 U6915 ( .B1(n7190), .B2(n6119), .A(n6106), .ZN(n6107) );
  OAI21_X1 U6916 ( .B1(n6531), .B2(n7501), .A(n6108), .ZN(U2956) );
  AND2_X1 U6917 ( .A1(n6109), .A2(n4764), .ZN(n6114) );
  NAND2_X1 U6918 ( .A1(n4772), .A2(n6110), .ZN(n6113) );
  NAND2_X1 U6919 ( .A1(n6115), .A2(n6111), .ZN(n6112) );
  OAI211_X1 U6920 ( .C1(n6115), .C2(n6114), .A(n6113), .B(n6112), .ZN(n6976)
         );
  NAND2_X1 U6921 ( .A1(n6116), .A2(n7194), .ZN(n7202) );
  AND2_X1 U6922 ( .A1(n7202), .A2(n7546), .ZN(n6117) );
  OR2_X1 U6923 ( .A1(n6118), .A2(n6117), .ZN(n6979) );
  AND2_X1 U6924 ( .A1(n6979), .A2(n7522), .ZN(n7503) );
  MUX2_X1 U6925 ( .A(MORE_REG_SCAN_IN), .B(n6976), .S(n7503), .Z(U3471) );
  OAI22_X1 U6926 ( .A1(n6120), .A2(n7478), .B1(n7491), .B2(n6119), .ZN(n6121)
         );
  AOI21_X1 U6927 ( .B1(EBX_REG_30__SCAN_IN), .B2(n3617), .A(n6121), .ZN(n6122)
         );
  OAI21_X1 U6928 ( .B1(n6123), .B2(REIP_REG_30__SCAN_IN), .A(n6122), .ZN(n6124) );
  INV_X1 U6929 ( .A(n6127), .ZN(n6142) );
  INV_X1 U6930 ( .A(n6372), .ZN(n6263) );
  NAND2_X1 U6931 ( .A1(n6146), .A2(n6129), .ZN(n6130) );
  NAND2_X1 U6932 ( .A1(n6131), .A2(n6130), .ZN(n6261) );
  INV_X1 U6933 ( .A(n6261), .ZN(n6547) );
  INV_X1 U6934 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7092) );
  INV_X1 U6935 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6262) );
  NOR2_X1 U6936 ( .A1(n7476), .A2(n6262), .ZN(n6134) );
  OAI22_X1 U6937 ( .A1(n6132), .A2(n7478), .B1(n7491), .B2(n6370), .ZN(n6133)
         );
  AOI211_X1 U6938 ( .C1(n6135), .C2(n7092), .A(n6134), .B(n6133), .ZN(n6136)
         );
  OAI21_X1 U6939 ( .B1(n7092), .B2(n6137), .A(n6136), .ZN(n6138) );
  AOI21_X1 U6940 ( .B1(n6547), .B2(n7412), .A(n6138), .ZN(n6139) );
  OAI21_X1 U6941 ( .B1(n6263), .B2(n7467), .A(n6139), .ZN(U2799) );
  OR2_X1 U6943 ( .A1(n6164), .A2(n6144), .ZN(n6145) );
  NAND2_X1 U6944 ( .A1(n6146), .A2(n6145), .ZN(n6550) );
  OAI22_X1 U6945 ( .A1(n6147), .A2(n7478), .B1(n7491), .B2(n6380), .ZN(n6149)
         );
  NOR3_X1 U6946 ( .A1(n6159), .A2(REIP_REG_27__SCAN_IN), .A3(n7088), .ZN(n6148) );
  AOI211_X1 U6947 ( .C1(EBX_REG_27__SCAN_IN), .C2(n3617), .A(n6149), .B(n6148), 
        .ZN(n6151) );
  NAND3_X1 U6948 ( .A1(n6217), .A2(REIP_REG_27__SCAN_IN), .A3(n6160), .ZN(
        n6150) );
  OAI211_X1 U6949 ( .C1(n6550), .C2(n7493), .A(n6151), .B(n6150), .ZN(n6152)
         );
  AOI21_X1 U6950 ( .B1(n6382), .B2(n7496), .A(n6152), .ZN(n6153) );
  INV_X1 U6951 ( .A(n6153), .ZN(U2800) );
  INV_X1 U6952 ( .A(n6141), .ZN(n6155) );
  AOI21_X1 U6953 ( .B1(n6156), .B2(n6154), .A(n6155), .ZN(n6390) );
  INV_X1 U6954 ( .A(n6390), .ZN(n6267) );
  INV_X1 U6955 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6157) );
  OAI22_X1 U6956 ( .A1(n6158), .A2(n7478), .B1(n6157), .B2(n7476), .ZN(n6163)
         );
  NAND2_X1 U6957 ( .A1(n6159), .A2(n7088), .ZN(n6161) );
  AND3_X1 U6958 ( .A1(n6217), .A2(n6161), .A3(n6160), .ZN(n6162) );
  AOI211_X1 U6959 ( .C1(n7483), .C2(n6386), .A(n6163), .B(n6162), .ZN(n6167)
         );
  AOI21_X1 U6960 ( .B1(n6165), .B2(n6170), .A(n6164), .ZN(n6566) );
  NAND2_X1 U6961 ( .A1(n6566), .A2(n7412), .ZN(n6166) );
  OAI211_X1 U6962 ( .C1(n6267), .C2(n7467), .A(n6167), .B(n6166), .ZN(U2801)
         );
  OAI21_X1 U6963 ( .B1(n6168), .B2(n6169), .A(n6154), .ZN(n6394) );
  INV_X1 U6964 ( .A(n6170), .ZN(n6171) );
  AOI21_X1 U6965 ( .B1(n6172), .B2(n6184), .A(n6171), .ZN(n6575) );
  AOI211_X1 U6966 ( .C1(n6174), .C2(n7086), .A(n6173), .B(n7473), .ZN(n6175)
         );
  AOI21_X1 U6967 ( .B1(EBX_REG_25__SCAN_IN), .B2(n3617), .A(n6175), .ZN(n6177)
         );
  AOI22_X1 U6968 ( .A1(n7490), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6245), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n6176) );
  OAI211_X1 U6969 ( .C1(n6396), .C2(n7491), .A(n6177), .B(n6176), .ZN(n6178)
         );
  AOI21_X1 U6970 ( .B1(n6575), .B2(n7412), .A(n6178), .ZN(n6179) );
  OAI21_X1 U6971 ( .B1(n6394), .B2(n7467), .A(n6179), .ZN(U2802) );
  INV_X1 U6972 ( .A(n6180), .ZN(n6183) );
  INV_X1 U6973 ( .A(n6181), .ZN(n6182) );
  AOI21_X1 U6974 ( .B1(n6183), .B2(n6182), .A(n6168), .ZN(n6409) );
  INV_X1 U6975 ( .A(n6409), .ZN(n6271) );
  AOI21_X1 U6976 ( .B1(n6185), .B2(n3650), .A(n3688), .ZN(n6582) );
  INV_X1 U6977 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6270) );
  INV_X1 U6978 ( .A(n6407), .ZN(n6191) );
  INV_X1 U6979 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7083) );
  INV_X1 U6980 ( .A(n6186), .ZN(n6188) );
  OAI21_X1 U6981 ( .B1(n6245), .B2(n6188), .A(n6217), .ZN(n7499) );
  OAI22_X1 U6982 ( .A1(n6187), .A2(n7478), .B1(n7083), .B2(n7499), .ZN(n6190)
         );
  NOR3_X1 U6983 ( .A1(n7473), .A2(REIP_REG_24__SCAN_IN), .A3(n6188), .ZN(n6189) );
  AOI211_X1 U6984 ( .C1(n7483), .C2(n6191), .A(n6190), .B(n6189), .ZN(n6192)
         );
  OAI21_X1 U6985 ( .B1(n7476), .B2(n6270), .A(n6192), .ZN(n6193) );
  AOI21_X1 U6986 ( .B1(n6582), .B2(n7412), .A(n6193), .ZN(n6194) );
  OAI21_X1 U6987 ( .B1(n6271), .B2(n7467), .A(n6194), .ZN(U2803) );
  NOR2_X1 U6988 ( .A1(n6196), .A2(n6197), .ZN(n6198) );
  OR2_X1 U6989 ( .A1(n6195), .A2(n6198), .ZN(n6441) );
  NAND4_X1 U6990 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .A4(n7410), .ZN(n7439) );
  OAI21_X1 U6991 ( .B1(n6199), .B2(n7439), .A(n7078), .ZN(n6208) );
  INV_X1 U6992 ( .A(n7461), .ZN(n6200) );
  NAND2_X1 U6993 ( .A1(n7333), .A2(n6200), .ZN(n6201) );
  AND2_X1 U6994 ( .A1(n6201), .A2(n6215), .ZN(n7464) );
  INV_X1 U6995 ( .A(n7464), .ZN(n7475) );
  NAND2_X1 U6996 ( .A1(n6295), .A2(n6202), .ZN(n6203) );
  AND2_X1 U6997 ( .A1(n6287), .A2(n6203), .ZN(n7212) );
  INV_X1 U6998 ( .A(n7212), .ZN(n6206) );
  INV_X1 U6999 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6290) );
  OAI22_X1 U7000 ( .A1(n6436), .A2(n7478), .B1(n6290), .B2(n7476), .ZN(n6204)
         );
  AOI21_X1 U7001 ( .B1(n7483), .B2(n6438), .A(n6204), .ZN(n6205) );
  OAI21_X1 U7002 ( .B1(n6206), .B2(n7493), .A(n6205), .ZN(n6207) );
  AOI21_X1 U7003 ( .B1(n6208), .B2(n7475), .A(n6207), .ZN(n6209) );
  OAI21_X1 U7004 ( .B1(n6441), .B2(n7467), .A(n6209), .ZN(U2807) );
  OAI21_X1 U7005 ( .B1(n3723), .B2(n3735), .A(n6211), .ZN(n6453) );
  NOR3_X1 U7006 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6212), .A3(n7439), .ZN(n7457) );
  INV_X1 U7007 ( .A(n6217), .ZN(n7348) );
  INV_X1 U7008 ( .A(n6212), .ZN(n6218) );
  INV_X1 U7009 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7010 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  NAND2_X1 U7011 ( .A1(n6217), .A2(n6216), .ZN(n7415) );
  OAI21_X1 U7012 ( .B1(n7348), .B2(n6218), .A(n7415), .ZN(n7456) );
  AOI22_X1 U7013 ( .A1(EBX_REG_18__SCAN_IN), .A2(n3617), .B1(
        REIP_REG_18__SCAN_IN), .B2(n7456), .ZN(n6219) );
  OAI211_X1 U7014 ( .C1(n7478), .C2(n6220), .A(n6219), .B(n7423), .ZN(n6225)
         );
  AOI21_X1 U7015 ( .B1(n6222), .B2(n3648), .A(n6221), .ZN(n7312) );
  INV_X1 U7016 ( .A(n7312), .ZN(n6298) );
  INV_X1 U7017 ( .A(n6450), .ZN(n6223) );
  OAI22_X1 U7018 ( .A1(n6298), .A2(n7493), .B1(n6223), .B2(n7491), .ZN(n6224)
         );
  NOR3_X1 U7019 ( .A1(n7457), .A2(n6225), .A3(n6224), .ZN(n6226) );
  OAI21_X1 U7020 ( .B1(n6453), .B2(n7467), .A(n6226), .ZN(U2809) );
  AOI21_X1 U7021 ( .B1(n6230), .B2(n6228), .A(n6229), .ZN(n6343) );
  INV_X1 U7022 ( .A(n6343), .ZN(n6460) );
  AOI21_X1 U7023 ( .B1(n6231), .B2(n6313), .A(n3664), .ZN(n7287) );
  AOI22_X1 U7024 ( .A1(n6232), .A2(n7483), .B1(EBX_REG_16__SCAN_IN), .B2(n3617), .ZN(n6233) );
  OAI211_X1 U7025 ( .C1(n7478), .C2(n6234), .A(n6233), .B(n7423), .ZN(n6236)
         );
  INV_X1 U7026 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7071) );
  INV_X1 U7027 ( .A(n7439), .ZN(n7446) );
  AND3_X1 U7028 ( .A1(n7071), .A2(REIP_REG_15__SCAN_IN), .A3(n7446), .ZN(n6235) );
  AOI211_X1 U7029 ( .C1(n7287), .C2(n7412), .A(n6236), .B(n6235), .ZN(n6238)
         );
  NOR2_X1 U7030 ( .A1(REIP_REG_15__SCAN_IN), .A2(n7439), .ZN(n7426) );
  INV_X1 U7031 ( .A(n7415), .ZN(n7428) );
  OAI21_X1 U7032 ( .B1(n7426), .B2(n7428), .A(REIP_REG_16__SCAN_IN), .ZN(n6237) );
  OAI211_X1 U7033 ( .C1(n6460), .C2(n7467), .A(n6238), .B(n6237), .ZN(U2811)
         );
  INV_X1 U7034 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7035 ( .A1(n6240), .A2(n7496), .ZN(n6259) );
  INV_X1 U7036 ( .A(n6241), .ZN(n6242) );
  NOR2_X1 U7037 ( .A1(n7473), .A2(n6242), .ZN(n7350) );
  AND2_X1 U7038 ( .A1(n7350), .A2(REIP_REG_5__SCAN_IN), .ZN(n7361) );
  INV_X1 U7039 ( .A(n7361), .ZN(n7375) );
  NOR3_X1 U7040 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6243), .A3(n7375), .ZN(n7389)
         );
  INV_X1 U7041 ( .A(n6243), .ZN(n6246) );
  NOR2_X1 U7042 ( .A1(n6245), .A2(n6244), .ZN(n7349) );
  AOI21_X1 U7043 ( .B1(n6246), .B2(n7349), .A(n7348), .ZN(n7390) );
  OAI21_X1 U7044 ( .B1(n7389), .B2(n7390), .A(REIP_REG_10__SCAN_IN), .ZN(n6258) );
  INV_X1 U7045 ( .A(n6247), .ZN(n6251) );
  OAI22_X1 U7046 ( .A1(n6249), .A2(n7476), .B1(n7493), .B2(n6248), .ZN(n6250)
         );
  AOI21_X1 U7047 ( .B1(n7483), .B2(n6251), .A(n6250), .ZN(n6257) );
  NAND3_X1 U7048 ( .A1(n7333), .A2(n6252), .A3(n6049), .ZN(n6253) );
  OAI211_X1 U7049 ( .C1(n7478), .C2(n6254), .A(n7423), .B(n6253), .ZN(n6255)
         );
  INV_X1 U7050 ( .A(n6255), .ZN(n6256) );
  NAND4_X1 U7051 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(U2817)
         );
  OAI22_X1 U7052 ( .A1(n6496), .A2(n6304), .B1(n7143), .B2(n6260), .ZN(U2828)
         );
  OAI222_X1 U7053 ( .A1(n7127), .A2(n6263), .B1(n6262), .B2(n7143), .C1(n6261), 
        .C2(n6304), .ZN(U2831) );
  INV_X1 U7054 ( .A(n6382), .ZN(n6265) );
  INV_X1 U7055 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6264) );
  OAI222_X1 U7056 ( .A1(n7127), .A2(n6265), .B1(n6264), .B2(n7143), .C1(n6550), 
        .C2(n6304), .ZN(U2832) );
  AOI22_X1 U7057 ( .A1(n6566), .A2(n7139), .B1(EBX_REG_26__SCAN_IN), .B2(n6314), .ZN(n6266) );
  OAI21_X1 U7058 ( .B1(n6267), .B2(n7127), .A(n6266), .ZN(U2833) );
  AOI22_X1 U7059 ( .A1(n6575), .A2(n7139), .B1(EBX_REG_25__SCAN_IN), .B2(n6314), .ZN(n6268) );
  OAI21_X1 U7060 ( .B1(n6394), .B2(n7127), .A(n6268), .ZN(U2834) );
  INV_X1 U7061 ( .A(n6582), .ZN(n6269) );
  OAI222_X1 U7062 ( .A1(n7127), .A2(n6271), .B1(n6270), .B2(n7143), .C1(n6269), 
        .C2(n6304), .ZN(U2835) );
  AND2_X1 U7063 ( .A1(n6272), .A2(n6273), .ZN(n6274) );
  OR2_X1 U7064 ( .A1(n6274), .A2(n6181), .ZN(n6417) );
  INV_X1 U7065 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7066 ( .A1(n6283), .A2(n6275), .ZN(n6276) );
  NAND2_X1 U7067 ( .A1(n3650), .A2(n6276), .ZN(n7494) );
  OAI222_X1 U7068 ( .A1(n7127), .A2(n6417), .B1(n6277), .B2(n7143), .C1(n7494), 
        .C2(n6304), .ZN(U2836) );
  INV_X1 U7069 ( .A(n6272), .ZN(n6279) );
  AOI21_X1 U7070 ( .B1(n6280), .B2(n6278), .A(n6279), .ZN(n7575) );
  INV_X1 U7071 ( .A(n7575), .ZN(n6284) );
  INV_X1 U7072 ( .A(EBX_REG_22__SCAN_IN), .ZN(n7477) );
  NOR2_X1 U7073 ( .A1(n6286), .A2(n6281), .ZN(n6282) );
  OR2_X1 U7074 ( .A1(n6283), .A2(n6282), .ZN(n7487) );
  OAI222_X1 U7075 ( .A1(n7127), .A2(n6284), .B1(n7143), .B2(n7477), .C1(n7487), 
        .C2(n6304), .ZN(U2837) );
  OAI21_X1 U7076 ( .B1(n6195), .B2(n6285), .A(n6278), .ZN(n7571) );
  AOI21_X1 U7077 ( .B1(n6288), .B2(n6287), .A(n6286), .ZN(n7465) );
  AOI22_X1 U7078 ( .A1(n7465), .A2(n7139), .B1(EBX_REG_21__SCAN_IN), .B2(n6314), .ZN(n6289) );
  OAI21_X1 U7079 ( .B1(n7571), .B2(n7127), .A(n6289), .ZN(U2838) );
  NOR2_X1 U7080 ( .A1(n7143), .A2(n6290), .ZN(n6291) );
  AOI21_X1 U7081 ( .B1(n7212), .B2(n7139), .A(n6291), .ZN(n6292) );
  OAI21_X1 U7082 ( .B1(n6441), .B2(n7127), .A(n6292), .ZN(U2839) );
  AND2_X1 U7083 ( .A1(n6211), .A2(n6293), .ZN(n6294) );
  OR2_X1 U7084 ( .A1(n6294), .A2(n6196), .ZN(n7184) );
  INV_X1 U7085 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6297) );
  OAI21_X1 U7086 ( .B1(n6221), .B2(n6296), .A(n6295), .ZN(n7460) );
  OAI222_X1 U7087 ( .A1(n7184), .A2(n7127), .B1(n6297), .B2(n7143), .C1(n6304), 
        .C2(n7460), .ZN(U2840) );
  INV_X1 U7088 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6299) );
  OAI222_X1 U7089 ( .A1(n6453), .A2(n7127), .B1(n6299), .B2(n7143), .C1(n6304), 
        .C2(n6298), .ZN(U2841) );
  OR2_X1 U7090 ( .A1(n6229), .A2(n6300), .ZN(n6301) );
  AND2_X1 U7091 ( .A1(n6210), .A2(n6301), .ZN(n7557) );
  INV_X1 U7092 ( .A(n7557), .ZN(n6306) );
  INV_X1 U7093 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6305) );
  INV_X1 U7094 ( .A(n6302), .ZN(n6303) );
  OAI21_X1 U7095 ( .B1(n3664), .B2(n6303), .A(n3648), .ZN(n7444) );
  OAI222_X1 U7096 ( .A1(n6306), .A2(n7127), .B1(n6305), .B2(n7143), .C1(n6304), 
        .C2(n7444), .ZN(U2842) );
  AOI22_X1 U7097 ( .A1(n7287), .A2(n7139), .B1(EBX_REG_16__SCAN_IN), .B2(n6314), .ZN(n6307) );
  OAI21_X1 U7098 ( .B1(n6460), .B2(n7127), .A(n6307), .ZN(U2843) );
  NAND2_X1 U7099 ( .A1(n6308), .A2(n6309), .ZN(n6310) );
  NAND2_X1 U7100 ( .A1(n6228), .A2(n6310), .ZN(n7430) );
  OR2_X1 U7101 ( .A1(n6640), .A2(n6311), .ZN(n6312) );
  NAND2_X1 U7102 ( .A1(n6313), .A2(n6312), .ZN(n7434) );
  INV_X1 U7103 ( .A(n7434), .ZN(n6315) );
  AOI22_X1 U7104 ( .A1(n6315), .A2(n7139), .B1(EBX_REG_15__SCAN_IN), .B2(n6314), .ZN(n6316) );
  OAI21_X1 U7105 ( .B1(n7430), .B2(n7127), .A(n6316), .ZN(U2844) );
  AND2_X1 U7106 ( .A1(n6317), .A2(n3900), .ZN(n6318) );
  NAND2_X1 U7107 ( .A1(n6319), .A2(n7579), .ZN(n6321) );
  AOI22_X1 U7108 ( .A1(n7578), .A2(DATAI_30_), .B1(n7581), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6320) );
  OAI211_X1 U7109 ( .C1(n7567), .C2(n6350), .A(n6321), .B(n6320), .ZN(U2861)
         );
  INV_X1 U7110 ( .A(n6322), .ZN(n6363) );
  NAND2_X1 U7111 ( .A1(n6363), .A2(n7579), .ZN(n6324) );
  AOI22_X1 U7112 ( .A1(n7578), .A2(DATAI_29_), .B1(n7581), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6323) );
  OAI211_X1 U7113 ( .C1(n7567), .C2(n6355), .A(n6324), .B(n6323), .ZN(U2862)
         );
  NAND2_X1 U7114 ( .A1(n6372), .A2(n7579), .ZN(n6326) );
  AOI22_X1 U7115 ( .A1(n7578), .A2(DATAI_28_), .B1(n7581), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U7116 ( .C1(n7567), .C2(n6327), .A(n6326), .B(n6325), .ZN(U2863)
         );
  NAND2_X1 U7117 ( .A1(n6382), .A2(n7579), .ZN(n6329) );
  AOI22_X1 U7118 ( .A1(n7578), .A2(DATAI_27_), .B1(n7581), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6328) );
  OAI211_X1 U7119 ( .C1(n7567), .C2(n6330), .A(n6329), .B(n6328), .ZN(U2864)
         );
  NAND2_X1 U7120 ( .A1(n6390), .A2(n7579), .ZN(n6332) );
  AOI22_X1 U7121 ( .A1(n7578), .A2(DATAI_26_), .B1(n7581), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6331) );
  OAI211_X1 U7122 ( .C1(n7567), .C2(n6333), .A(n6332), .B(n6331), .ZN(U2865)
         );
  AOI22_X1 U7123 ( .A1(n7578), .A2(DATAI_25_), .B1(n7581), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7124 ( .A1(n7582), .A2(DATAI_9_), .ZN(n6334) );
  OAI211_X1 U7125 ( .C1(n6394), .C2(n6354), .A(n6335), .B(n6334), .ZN(U2866)
         );
  NAND2_X1 U7126 ( .A1(n6409), .A2(n7579), .ZN(n6337) );
  AOI22_X1 U7127 ( .A1(n7578), .A2(DATAI_24_), .B1(n7581), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6336) );
  OAI211_X1 U7128 ( .C1(n7567), .C2(n6338), .A(n6337), .B(n6336), .ZN(U2867)
         );
  AOI22_X1 U7129 ( .A1(n7578), .A2(DATAI_20_), .B1(n7581), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7130 ( .A1(n7582), .A2(DATAI_4_), .ZN(n6339) );
  OAI211_X1 U7131 ( .C1(n6441), .C2(n6354), .A(n6340), .B(n6339), .ZN(U2871)
         );
  AOI22_X1 U7132 ( .A1(n7578), .A2(DATAI_18_), .B1(n7581), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7133 ( .A1(n7582), .A2(DATAI_2_), .ZN(n6341) );
  OAI211_X1 U7134 ( .C1(n6453), .C2(n6354), .A(n6342), .B(n6341), .ZN(U2873)
         );
  NAND2_X1 U7135 ( .A1(n6343), .A2(n7579), .ZN(n6345) );
  AOI22_X1 U7136 ( .A1(n7578), .A2(DATAI_16_), .B1(n7581), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6344) );
  OAI211_X1 U7137 ( .C1(n7567), .C2(n6346), .A(n6345), .B(n6344), .ZN(U2875)
         );
  INV_X1 U7138 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7051) );
  OAI222_X1 U7139 ( .A1(n6347), .A2(n6356), .B1(n7564), .B2(n7051), .C1(n6354), 
        .C2(n7430), .ZN(U2876) );
  INV_X1 U7140 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7047) );
  XOR2_X1 U7141 ( .A(n6348), .B(n3660), .Z(n7419) );
  INV_X1 U7142 ( .A(n7419), .ZN(n6349) );
  OAI222_X1 U7143 ( .A1(n6356), .A2(n6350), .B1(n7564), .B2(n7047), .C1(n6354), 
        .C2(n6349), .ZN(U2877) );
  XOR2_X1 U7144 ( .A(n6352), .B(n6351), .Z(n7402) );
  INV_X1 U7145 ( .A(n7402), .ZN(n6353) );
  OAI222_X1 U7146 ( .A1(n6356), .A2(n6355), .B1(n6354), .B2(n6353), .C1(n7045), 
        .C2(n7564), .ZN(U2878) );
  AOI22_X1 U7147 ( .A1(n6366), .A2(n6357), .B1(n3618), .B2(n6545), .ZN(n6358)
         );
  AND2_X1 U7148 ( .A1(n7280), .A2(REIP_REG_29__SCAN_IN), .ZN(n6537) );
  AOI21_X1 U7149 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6537), 
        .ZN(n6360) );
  OAI21_X1 U7150 ( .B1(n7190), .B2(n6361), .A(n6360), .ZN(n6362) );
  AOI21_X1 U7151 ( .B1(n6363), .B2(n7185), .A(n6362), .ZN(n6364) );
  OAI21_X1 U7152 ( .B1(n7501), .B2(n3653), .A(n6364), .ZN(U2957) );
  NAND2_X1 U7153 ( .A1(n6366), .A2(n6365), .ZN(n6368) );
  XNOR2_X1 U7154 ( .A(n3618), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6367)
         );
  XNOR2_X1 U7155 ( .A(n6368), .B(n6367), .ZN(n6549) );
  AND2_X1 U7156 ( .A1(n7280), .A2(REIP_REG_28__SCAN_IN), .ZN(n6542) );
  AOI21_X1 U7157 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6542), 
        .ZN(n6369) );
  OAI21_X1 U7158 ( .B1(n7190), .B2(n6370), .A(n6369), .ZN(n6371) );
  AOI21_X1 U7159 ( .B1(n6372), .B2(n7185), .A(n6371), .ZN(n6373) );
  OAI21_X1 U7160 ( .B1(n6549), .B2(n7501), .A(n6373), .ZN(U2958) );
  NAND2_X1 U7161 ( .A1(n6374), .A2(n6562), .ZN(n6375) );
  AND2_X1 U7162 ( .A1(n7280), .A2(REIP_REG_27__SCAN_IN), .ZN(n6551) );
  AOI21_X1 U7163 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6551), 
        .ZN(n6379) );
  OAI21_X1 U7164 ( .B1(n7190), .B2(n6380), .A(n6379), .ZN(n6381) );
  AOI21_X1 U7165 ( .B1(n6382), .B2(n7185), .A(n6381), .ZN(n6383) );
  OAI21_X1 U7166 ( .B1(n7501), .B2(n6559), .A(n6383), .ZN(U2959) );
  XNOR2_X1 U7167 ( .A(n3618), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6385)
         );
  XNOR2_X1 U7168 ( .A(n6384), .B(n6385), .ZN(n6569) );
  INV_X1 U7169 ( .A(n6386), .ZN(n6388) );
  AND2_X1 U7170 ( .A1(n7280), .A2(REIP_REG_26__SCAN_IN), .ZN(n6564) );
  AOI21_X1 U7171 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6564), 
        .ZN(n6387) );
  OAI21_X1 U7172 ( .B1(n7190), .B2(n6388), .A(n6387), .ZN(n6389) );
  AOI21_X1 U7173 ( .B1(n6390), .B2(n7185), .A(n6389), .ZN(n6391) );
  OAI21_X1 U7174 ( .B1(n6569), .B2(n7501), .A(n6391), .ZN(U2960) );
  XNOR2_X1 U7175 ( .A(n6392), .B(n6393), .ZN(n6577) );
  INV_X1 U7176 ( .A(n6394), .ZN(n6398) );
  AND2_X1 U7177 ( .A1(n7280), .A2(REIP_REG_25__SCAN_IN), .ZN(n6570) );
  AOI21_X1 U7178 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6570), 
        .ZN(n6395) );
  OAI21_X1 U7179 ( .B1(n7190), .B2(n6396), .A(n6395), .ZN(n6397) );
  AOI21_X1 U7180 ( .B1(n6398), .B2(n7185), .A(n6397), .ZN(n6399) );
  OAI21_X1 U7181 ( .B1(n6577), .B2(n7501), .A(n6399), .ZN(U2961) );
  XNOR2_X1 U7182 ( .A(n6483), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6616)
         );
  NAND2_X2 U7183 ( .A1(n6617), .A2(n6616), .ZN(n6615) );
  NOR2_X1 U7184 ( .A1(n6444), .A2(n6433), .ZN(n6400) );
  OAI22_X2 U7185 ( .A1(n6615), .A2(n6400), .B1(n6443), .B2(n7217), .ZN(n6427)
         );
  XNOR2_X1 U7186 ( .A(n6483), .B(n6609), .ZN(n6426) );
  NAND3_X1 U7187 ( .A1(n6483), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6404) );
  NOR2_X1 U7188 ( .A1(n3618), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6411)
         );
  NAND3_X1 U7189 ( .A1(n6411), .A2(n6412), .A3(n6402), .ZN(n6403) );
  OAI22_X1 U7190 ( .A1(n6422), .A2(n6404), .B1(n6615), .B2(n6403), .ZN(n6405)
         );
  XNOR2_X1 U7191 ( .A(n6405), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6584)
         );
  NAND2_X1 U7192 ( .A1(n7280), .A2(REIP_REG_24__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U7193 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6406)
         );
  OAI211_X1 U7194 ( .C1(n7190), .C2(n6407), .A(n6578), .B(n6406), .ZN(n6408)
         );
  AOI21_X1 U7195 ( .B1(n6409), .B2(n7185), .A(n6408), .ZN(n6410) );
  OAI21_X1 U7196 ( .B1(n6584), .B2(n7501), .A(n6410), .ZN(U2962) );
  INV_X1 U7197 ( .A(n6411), .ZN(n6432) );
  INV_X1 U7198 ( .A(n6412), .ZN(n6600) );
  NOR2_X1 U7199 ( .A1(n6432), .A2(n6600), .ZN(n6415) );
  NOR2_X1 U7200 ( .A1(n6443), .A2(n6413), .ZN(n6414) );
  MUX2_X1 U7201 ( .A(n6415), .B(n6414), .S(n6615), .Z(n6416) );
  XNOR2_X1 U7202 ( .A(n6416), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6592)
         );
  NAND2_X1 U7203 ( .A1(n7280), .A2(REIP_REG_23__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U7204 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6418)
         );
  OAI211_X1 U7205 ( .C1(n7190), .C2(n7492), .A(n6586), .B(n6418), .ZN(n6419)
         );
  AOI21_X1 U7206 ( .B1(n7580), .B2(n7185), .A(n6419), .ZN(n6420) );
  OAI21_X1 U7207 ( .B1(n7501), .B2(n6592), .A(n6420), .ZN(U2963) );
  XNOR2_X1 U7208 ( .A(n3618), .B(n6594), .ZN(n6421) );
  NAND2_X1 U7209 ( .A1(n6466), .A2(n7484), .ZN(n6423) );
  NAND2_X1 U7210 ( .A1(n7280), .A2(REIP_REG_22__SCAN_IN), .ZN(n6595) );
  OAI211_X1 U7211 ( .C1(n6464), .C2(n7479), .A(n6423), .B(n6595), .ZN(n6424)
         );
  AOI21_X1 U7212 ( .B1(n7575), .B2(n7185), .A(n6424), .ZN(n6425) );
  OAI21_X1 U7213 ( .B1(n6596), .B2(n7501), .A(n6425), .ZN(U2964) );
  NAND2_X1 U7214 ( .A1(n6427), .A2(n6426), .ZN(n6602) );
  NAND2_X1 U7215 ( .A1(n7280), .A2(REIP_REG_21__SCAN_IN), .ZN(n6604) );
  INV_X1 U7216 ( .A(n6604), .ZN(n6429) );
  NOR2_X1 U7217 ( .A1(n7190), .A2(n7471), .ZN(n6428) );
  AOI211_X1 U7218 ( .C1(n7183), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n6429), 
        .B(n6428), .ZN(n6430) );
  OAI211_X1 U7219 ( .C1(n7174), .C2(n7571), .A(n6431), .B(n6430), .ZN(U2965)
         );
  OAI21_X1 U7220 ( .B1(n6443), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6615), 
        .ZN(n6435) );
  OAI21_X1 U7221 ( .B1(n6443), .B2(n6433), .A(n6432), .ZN(n6434) );
  XNOR2_X1 U7222 ( .A(n6435), .B(n6434), .ZN(n7213) );
  NAND2_X1 U7223 ( .A1(n7213), .A2(n7186), .ZN(n6440) );
  OAI22_X1 U7224 ( .A1(n6464), .A2(n6436), .B1(n7248), .B2(n7078), .ZN(n6437)
         );
  AOI21_X1 U7225 ( .B1(n6466), .B2(n6438), .A(n6437), .ZN(n6439) );
  OAI211_X1 U7226 ( .C1(n7174), .C2(n6441), .A(n6440), .B(n6439), .ZN(U2966)
         );
  INV_X1 U7227 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U7228 ( .A1(n6443), .A2(n7302), .ZN(n6447) );
  NAND2_X1 U7229 ( .A1(n6444), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6445) );
  OAI22_X1 U7230 ( .A1(n6442), .A2(n6447), .B1(n6446), .B2(n6445), .ZN(n6448)
         );
  XOR2_X1 U7231 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n6448), .Z(n7315) );
  NAND2_X1 U7232 ( .A1(n7315), .A2(n7186), .ZN(n6452) );
  OAI22_X1 U7233 ( .A1(n6464), .A2(n6220), .B1(n7248), .B2(n7074), .ZN(n6449)
         );
  AOI21_X1 U7234 ( .B1(n6466), .B2(n6450), .A(n6449), .ZN(n6451) );
  OAI211_X1 U7235 ( .C1(n7174), .C2(n6453), .A(n6452), .B(n6451), .ZN(U2968)
         );
  XNOR2_X1 U7236 ( .A(n3618), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6455)
         );
  XNOR2_X1 U7237 ( .A(n6454), .B(n6455), .ZN(n7289) );
  NAND2_X1 U7238 ( .A1(n7289), .A2(n7186), .ZN(n6459) );
  AND2_X1 U7239 ( .A1(n7280), .A2(REIP_REG_16__SCAN_IN), .ZN(n7286) );
  NOR2_X1 U7240 ( .A1(n7190), .A2(n6456), .ZN(n6457) );
  AOI211_X1 U7241 ( .C1(n7183), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7286), 
        .B(n6457), .ZN(n6458) );
  OAI211_X1 U7242 ( .C1(n7174), .C2(n6460), .A(n6459), .B(n6458), .ZN(U2970)
         );
  OAI21_X1 U7243 ( .B1(n6463), .B2(n6462), .A(n6461), .ZN(n6625) );
  NAND2_X1 U7244 ( .A1(n6625), .A2(n7186), .ZN(n6468) );
  INV_X1 U7245 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U7246 ( .A1(n7280), .A2(REIP_REG_15__SCAN_IN), .ZN(n6630) );
  OAI21_X1 U7247 ( .B1(n6464), .B2(n7425), .A(n6630), .ZN(n6465) );
  AOI21_X1 U7248 ( .B1(n7432), .B2(n6466), .A(n6465), .ZN(n6467) );
  OAI211_X1 U7249 ( .C1(n7174), .C2(n7430), .A(n6468), .B(n6467), .ZN(U2971)
         );
  OAI21_X1 U7250 ( .B1(n6469), .B2(n6471), .A(n6470), .ZN(n6644) );
  INV_X1 U7251 ( .A(n6644), .ZN(n6475) );
  AOI22_X1 U7252 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n7280), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n6472) );
  OAI21_X1 U7253 ( .B1(n7190), .B2(n7417), .A(n6472), .ZN(n6473) );
  AOI21_X1 U7254 ( .B1(n7419), .B2(n7185), .A(n6473), .ZN(n6474) );
  OAI21_X1 U7255 ( .B1(n6475), .B2(n7501), .A(n6474), .ZN(U2972) );
  XOR2_X1 U7256 ( .A(n6476), .B(n6477), .Z(n6653) );
  INV_X1 U7257 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U7258 ( .A1(n7248), .A2(n6478), .ZN(n6651) );
  AOI21_X1 U7259 ( .B1(n7183), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6651), 
        .ZN(n6479) );
  OAI21_X1 U7260 ( .B1(n7190), .B2(n7400), .A(n6479), .ZN(n6480) );
  AOI21_X1 U7261 ( .B1(n7402), .B2(n7185), .A(n6480), .ZN(n6481) );
  OAI21_X1 U7262 ( .B1(n6653), .B2(n7501), .A(n6481), .ZN(U2973) );
  OAI21_X1 U7263 ( .B1(n6046), .B2(n6483), .A(n6482), .ZN(n6656) );
  XNOR2_X1 U7264 ( .A(n6483), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6655)
         );
  NAND2_X1 U7265 ( .A1(n6656), .A2(n6655), .ZN(n6654) );
  OAI21_X1 U7266 ( .B1(n6484), .B2(n6444), .A(n6654), .ZN(n6488) );
  OAI21_X1 U7267 ( .B1(n6486), .B2(n6483), .A(n6485), .ZN(n6487) );
  XNOR2_X1 U7268 ( .A(n6488), .B(n6487), .ZN(n7279) );
  INV_X1 U7269 ( .A(n7279), .ZN(n6495) );
  INV_X1 U7270 ( .A(n6489), .ZN(n6493) );
  AOI22_X1 U7271 ( .A1(n7183), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n7280), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6490) );
  OAI21_X1 U7272 ( .B1(n7190), .B2(n6491), .A(n6490), .ZN(n6492) );
  AOI21_X1 U7273 ( .B1(n6493), .B2(n7185), .A(n6492), .ZN(n6494) );
  OAI21_X1 U7274 ( .B1(n6495), .B2(n7501), .A(n6494), .ZN(U2974) );
  NOR2_X1 U7275 ( .A1(n6496), .A2(n7301), .ZN(n6520) );
  NAND2_X1 U7276 ( .A1(n6509), .A2(n7252), .ZN(n6511) );
  NAND3_X1 U7277 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6497), .ZN(n6627) );
  NOR2_X1 U7278 ( .A1(n6498), .A2(n6627), .ZN(n6611) );
  NAND3_X1 U7279 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6635) );
  NOR2_X1 U7280 ( .A1(n6499), .A2(n6635), .ZN(n6629) );
  NAND3_X1 U7281 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6629), .ZN(n6501) );
  INV_X1 U7282 ( .A(n6501), .ZN(n7294) );
  NAND2_X1 U7283 ( .A1(n6611), .A2(n7294), .ZN(n7295) );
  NOR2_X1 U7284 ( .A1(n6500), .A2(n7295), .ZN(n6618) );
  AND2_X1 U7285 ( .A1(n6618), .A2(n7217), .ZN(n6505) );
  OAI21_X1 U7286 ( .B1(n7256), .B2(n6505), .A(n7300), .ZN(n6504) );
  INV_X1 U7287 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6614) );
  NOR2_X1 U7288 ( .A1(n7302), .A2(n6501), .ZN(n6613) );
  NOR2_X1 U7289 ( .A1(n6627), .A2(n6502), .ZN(n6612) );
  NAND2_X1 U7290 ( .A1(n6613), .A2(n6612), .ZN(n7297) );
  NOR2_X1 U7291 ( .A1(n6614), .A2(n7297), .ZN(n6620) );
  AND2_X1 U7292 ( .A1(n6620), .A2(n7217), .ZN(n6506) );
  NOR2_X1 U7293 ( .A1(n7252), .A2(n6506), .ZN(n6503) );
  NOR2_X1 U7294 ( .A1(n6504), .A2(n6503), .ZN(n6610) );
  INV_X1 U7295 ( .A(n6505), .ZN(n6508) );
  INV_X1 U7296 ( .A(n6506), .ZN(n6507) );
  OAI22_X1 U7297 ( .A1(n6509), .A2(n6508), .B1(n7252), .B2(n6507), .ZN(n6603)
         );
  INV_X1 U7298 ( .A(n6514), .ZN(n6510) );
  NAND2_X1 U7299 ( .A1(n6603), .A2(n6510), .ZN(n6593) );
  NAND2_X1 U7300 ( .A1(n6610), .A2(n6593), .ZN(n6590) );
  AOI21_X1 U7301 ( .B1(n6515), .B2(n6511), .A(n6590), .ZN(n6580) );
  NOR2_X1 U7302 ( .A1(n6562), .A2(n6573), .ZN(n6561) );
  NAND2_X1 U7303 ( .A1(n6580), .A2(n6561), .ZN(n6540) );
  NAND2_X1 U7304 ( .A1(n6580), .A2(n6628), .ZN(n6541) );
  OAI21_X1 U7305 ( .B1(n6540), .B2(n6523), .A(n6541), .ZN(n6535) );
  INV_X1 U7306 ( .A(n6541), .ZN(n6513) );
  AOI211_X1 U7307 ( .C1(n6535), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6513), .B(n6512), .ZN(n6519) );
  NAND2_X1 U7308 ( .A1(n6571), .A2(n6561), .ZN(n6532) );
  INV_X1 U7309 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6516) );
  NOR4_X1 U7310 ( .A1(n6532), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6516), 
        .A4(n6523), .ZN(n6517) );
  NOR4_X2 U7311 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n6521)
         );
  OAI21_X1 U7312 ( .B1(n6522), .B2(n7240), .A(n6521), .ZN(U2987) );
  INV_X1 U7313 ( .A(n6535), .ZN(n6526) );
  NOR3_X1 U7314 ( .A1(n6532), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6523), 
        .ZN(n6524) );
  AOI211_X1 U7315 ( .C1(n6526), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6525), .B(n6524), .ZN(n6530) );
  INV_X1 U7316 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U7317 ( .A1(n6528), .A2(n7313), .ZN(n6529) );
  OAI211_X1 U7318 ( .C1(n6531), .C2(n7240), .A(n6530), .B(n6529), .ZN(U2988)
         );
  INV_X1 U7319 ( .A(n6532), .ZN(n6552) );
  AOI21_X1 U7320 ( .B1(n6552), .B2(n6533), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n6534) );
  NOR2_X1 U7321 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  AOI211_X1 U7322 ( .C1(n6538), .C2(n7313), .A(n6537), .B(n6536), .ZN(n6539)
         );
  OAI21_X1 U7323 ( .B1(n3653), .B2(n7240), .A(n6539), .ZN(U2989) );
  NAND2_X1 U7324 ( .A1(n6541), .A2(n6540), .ZN(n6555) );
  XNOR2_X1 U7325 ( .A(n6554), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6543)
         );
  AOI21_X1 U7326 ( .B1(n6552), .B2(n6543), .A(n6542), .ZN(n6544) );
  OAI21_X1 U7327 ( .B1(n6555), .B2(n6545), .A(n6544), .ZN(n6546) );
  AOI21_X1 U7328 ( .B1(n6547), .B2(n7313), .A(n6546), .ZN(n6548) );
  OAI21_X1 U7329 ( .B1(n6549), .B2(n7240), .A(n6548), .ZN(U2990) );
  INV_X1 U7330 ( .A(n6550), .ZN(n6557) );
  AOI21_X1 U7331 ( .B1(n6552), .B2(n6554), .A(n6551), .ZN(n6553) );
  OAI21_X1 U7332 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(n6556) );
  AOI21_X1 U7333 ( .B1(n6557), .B2(n7313), .A(n6556), .ZN(n6558) );
  OAI21_X1 U7334 ( .B1(n6559), .B2(n7240), .A(n6558), .ZN(U2991) );
  INV_X1 U7335 ( .A(n6580), .ZN(n6565) );
  INV_X1 U7336 ( .A(n6571), .ZN(n6560) );
  AOI211_X1 U7337 ( .C1(n6573), .C2(n6562), .A(n6561), .B(n6560), .ZN(n6563)
         );
  AOI211_X1 U7338 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n6565), .A(n6564), .B(n6563), .ZN(n6568) );
  NAND2_X1 U7339 ( .A1(n6566), .A2(n7313), .ZN(n6567) );
  OAI211_X1 U7340 ( .C1(n6569), .C2(n7240), .A(n6568), .B(n6567), .ZN(U2992)
         );
  AOI21_X1 U7341 ( .B1(n6571), .B2(n6573), .A(n6570), .ZN(n6572) );
  OAI21_X1 U7342 ( .B1(n6580), .B2(n6573), .A(n6572), .ZN(n6574) );
  AOI21_X1 U7343 ( .B1(n6575), .B2(n7313), .A(n6574), .ZN(n6576) );
  OAI21_X1 U7344 ( .B1(n6577), .B2(n7240), .A(n6576), .ZN(U2993) );
  AOI21_X1 U7345 ( .B1(n6585), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6579) );
  OAI21_X1 U7346 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(n6581) );
  AOI21_X1 U7347 ( .B1(n6582), .B2(n7313), .A(n6581), .ZN(n6583) );
  OAI21_X1 U7348 ( .B1(n6584), .B2(n7240), .A(n6583), .ZN(U2994) );
  INV_X1 U7349 ( .A(n6585), .ZN(n6587) );
  OAI21_X1 U7350 ( .B1(n6587), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6586), 
        .ZN(n6589) );
  NOR2_X1 U7351 ( .A1(n7494), .A2(n7301), .ZN(n6588) );
  AOI211_X1 U7352 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n6590), .A(n6589), .B(n6588), .ZN(n6591) );
  OAI21_X1 U7353 ( .B1(n6592), .B2(n7240), .A(n6591), .ZN(U2995) );
  OAI21_X1 U7354 ( .B1(n6610), .B2(n6594), .A(n6593), .ZN(n6599) );
  OAI21_X1 U7355 ( .B1(n7487), .B2(n7301), .A(n6595), .ZN(n6598) );
  NOR2_X1 U7356 ( .A1(n6596), .A2(n7240), .ZN(n6597) );
  INV_X1 U7357 ( .A(n6601), .ZN(U2996) );
  INV_X1 U7358 ( .A(n6603), .ZN(n6605) );
  OAI21_X1 U7359 ( .B1(n6605), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6604), 
        .ZN(n6606) );
  AOI21_X1 U7360 ( .B1(n7465), .B2(n7313), .A(n6606), .ZN(n6607) );
  OAI211_X1 U7361 ( .C1(n6610), .C2(n6609), .A(n6608), .B(n6607), .ZN(U2997)
         );
  NAND2_X1 U7362 ( .A1(n7260), .A2(n6611), .ZN(n7310) );
  INV_X1 U7363 ( .A(n7307), .ZN(n7277) );
  NAND2_X1 U7364 ( .A1(n6613), .A2(n7277), .ZN(n7318) );
  NOR2_X1 U7365 ( .A1(n6614), .A2(n7318), .ZN(n7210) );
  INV_X1 U7366 ( .A(n7210), .ZN(n6624) );
  OAI21_X1 U7367 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(n7187) );
  NAND2_X1 U7368 ( .A1(n7187), .A2(n7314), .ZN(n6623) );
  OR2_X1 U7369 ( .A1(n7256), .A2(n6618), .ZN(n6619) );
  OAI211_X1 U7370 ( .C1(n6620), .C2(n7252), .A(n7300), .B(n6619), .ZN(n7211)
         );
  INV_X1 U7371 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7445) );
  OAI22_X1 U7372 ( .A1(n7460), .A2(n7301), .B1(n7248), .B2(n7445), .ZN(n6621)
         );
  AOI21_X1 U7373 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n7211), .A(n6621), 
        .ZN(n6622) );
  OAI211_X1 U7374 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6624), .A(n6623), .B(n6622), .ZN(U2999) );
  NAND2_X1 U7375 ( .A1(n6629), .A2(n7277), .ZN(n7293) );
  NAND2_X1 U7376 ( .A1(n6625), .A2(n7314), .ZN(n6633) );
  AOI21_X1 U7377 ( .B1(n6627), .B2(n7226), .A(n6626), .ZN(n6634) );
  OAI21_X1 U7378 ( .B1(n6629), .B2(n6628), .A(n6634), .ZN(n7288) );
  OAI21_X1 U7379 ( .B1(n7301), .B2(n7434), .A(n6630), .ZN(n6631) );
  AOI21_X1 U7380 ( .B1(n7288), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6631), 
        .ZN(n6632) );
  OAI211_X1 U7381 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n7293), .A(n6633), .B(n6632), .ZN(U3003) );
  NOR2_X1 U7382 ( .A1(n7307), .A2(n6635), .ZN(n6637) );
  INV_X1 U7383 ( .A(n6634), .ZN(n7274) );
  AOI21_X1 U7384 ( .B1(n6635), .B2(n7226), .A(n7274), .ZN(n6636) );
  INV_X1 U7385 ( .A(n6636), .ZN(n6648) );
  MUX2_X1 U7386 ( .A(n6637), .B(n6648), .S(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .Z(n6643) );
  AOI21_X1 U7387 ( .B1(n6639), .B2(n6646), .A(n6638), .ZN(n6641) );
  OR2_X1 U7388 ( .A1(n6641), .A2(n6640), .ZN(n7133) );
  INV_X1 U7389 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7414) );
  OAI22_X1 U7390 ( .A1(n7301), .A2(n7133), .B1(n7414), .B2(n7248), .ZN(n6642)
         );
  AOI211_X1 U7391 ( .C1(n6644), .C2(n7314), .A(n6643), .B(n6642), .ZN(n6645)
         );
  INV_X1 U7392 ( .A(n6645), .ZN(U3004) );
  XNOR2_X1 U7393 ( .A(n6647), .B(n6646), .ZN(n7399) );
  NAND2_X1 U7394 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7276) );
  NOR2_X1 U7395 ( .A1(n7307), .A2(n7276), .ZN(n6649) );
  MUX2_X1 U7396 ( .A(n6649), .B(n6648), .S(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .Z(n6650) );
  AOI211_X1 U7397 ( .C1(n7313), .C2(n7399), .A(n6651), .B(n6650), .ZN(n6652)
         );
  OAI21_X1 U7398 ( .B1(n6653), .B2(n7240), .A(n6652), .ZN(U3005) );
  OAI21_X1 U7399 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(n7179) );
  OAI22_X1 U7400 ( .A1(n7301), .A2(n6657), .B1(n7064), .B2(n7248), .ZN(n6658)
         );
  AOI21_X1 U7401 ( .B1(n7274), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6658), 
        .ZN(n6660) );
  OR2_X1 U7402 ( .A1(n7307), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6659)
         );
  OAI211_X1 U7403 ( .C1(n7179), .C2(n7240), .A(n6660), .B(n6659), .ZN(U3007)
         );
  NOR2_X1 U7404 ( .A1(n6661), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6663)
         );
  NOR3_X1 U7405 ( .A1(n4437), .A2(n4939), .A3(n5282), .ZN(n6662) );
  AOI211_X1 U7406 ( .C1(n6665), .C2(n6664), .A(n6663), .B(n6662), .ZN(n6963)
         );
  INV_X1 U7407 ( .A(n7517), .ZN(n7510) );
  INV_X1 U7408 ( .A(n5282), .ZN(n6670) );
  NOR2_X1 U7409 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  AOI22_X1 U7410 ( .A1(n6671), .A2(n6670), .B1(n6669), .B2(n6668), .ZN(n6672)
         );
  OAI21_X1 U7411 ( .B1(n6963), .B2(n7510), .A(n6672), .ZN(n6673) );
  MUX2_X1 U7412 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6673), .S(n7521), 
        .Z(U3460) );
  INV_X1 U7413 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U7414 ( .A1(n7185), .A2(DATAI_25_), .ZN(n6899) );
  NOR2_X2 U7415 ( .A1(n6678), .A2(n3907), .ZN(n7610) );
  NOR2_X2 U7416 ( .A1(n7559), .A2(n6679), .ZN(n6944) );
  AOI22_X1 U7417 ( .A1(n7610), .A2(n6682), .B1(n6944), .B2(n6681), .ZN(n6674)
         );
  OAI21_X1 U7418 ( .B1(n6684), .B2(n6899), .A(n6674), .ZN(n6675) );
  AOI21_X1 U7419 ( .B1(n7611), .B2(n6686), .A(n6675), .ZN(n6676) );
  OAI21_X1 U7420 ( .B1(n6689), .B2(n6677), .A(n6676), .ZN(U3021) );
  INV_X1 U7421 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U7422 ( .A1(n7185), .A2(DATAI_28_), .ZN(n6906) );
  NOR2_X2 U7423 ( .A1(n6678), .A2(n3920), .ZN(n7628) );
  NOR2_X2 U7424 ( .A1(n6680), .A2(n6679), .ZN(n6949) );
  AOI22_X1 U7425 ( .A1(n7628), .A2(n6682), .B1(n6949), .B2(n6681), .ZN(n6683)
         );
  OAI21_X1 U7426 ( .B1(n6684), .B2(n6906), .A(n6683), .ZN(n6685) );
  AOI21_X1 U7427 ( .B1(n7629), .B2(n6686), .A(n6685), .ZN(n6687) );
  OAI21_X1 U7428 ( .B1(n6689), .B2(n6688), .A(n6687), .ZN(U3024) );
  INV_X1 U7429 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6693) );
  AOI22_X1 U7430 ( .A1(n7610), .A2(n6695), .B1(n6944), .B2(n6694), .ZN(n6690)
         );
  OAI21_X1 U7431 ( .B1(n6899), .B2(n6697), .A(n6690), .ZN(n6691) );
  AOI21_X1 U7432 ( .B1(n7611), .B2(n6710), .A(n6691), .ZN(n6692) );
  OAI21_X1 U7433 ( .B1(n6701), .B2(n6693), .A(n6692), .ZN(U3029) );
  INV_X1 U7434 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6700) );
  AOI22_X1 U7435 ( .A1(n7628), .A2(n6695), .B1(n6949), .B2(n6694), .ZN(n6696)
         );
  OAI21_X1 U7436 ( .B1(n6906), .B2(n6697), .A(n6696), .ZN(n6698) );
  AOI21_X1 U7437 ( .B1(n7629), .B2(n6710), .A(n6698), .ZN(n6699) );
  OAI21_X1 U7438 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(U3032) );
  OAI21_X1 U7439 ( .B1(n6760), .B2(n6710), .A(n6853), .ZN(n6702) );
  OAI21_X1 U7440 ( .B1(n6703), .B2(n6712), .A(n6702), .ZN(n6705) );
  NOR2_X1 U7441 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6704), .ZN(n6747)
         );
  AOI21_X1 U7442 ( .B1(n6705), .B2(n7533), .A(n6747), .ZN(n6709) );
  NAND2_X1 U7443 ( .A1(n6707), .A2(n6706), .ZN(n6795) );
  NAND2_X1 U7444 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6795), .ZN(n6792) );
  INV_X1 U7445 ( .A(n6792), .ZN(n6708) );
  NOR3_X2 U7446 ( .A1(n6709), .A2(n6860), .A3(n6708), .ZN(n6754) );
  INV_X1 U7447 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6717) );
  OAI22_X1 U7448 ( .A1(n6797), .A2(n6712), .B1(n6795), .B2(n6711), .ZN(n6746)
         );
  AOI22_X1 U7449 ( .A1(n7596), .A2(n6747), .B1(n6798), .B2(n6746), .ZN(n6713)
         );
  OAI21_X1 U7450 ( .B1(n6750), .B2(n6714), .A(n6713), .ZN(n6715) );
  AOI21_X1 U7451 ( .B1(n7606), .B2(n6760), .A(n6715), .ZN(n6716) );
  OAI21_X1 U7452 ( .B1(n6754), .B2(n6717), .A(n6716), .ZN(U3036) );
  INV_X1 U7453 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7454 ( .A1(n7610), .A2(n6747), .B1(n6944), .B2(n6746), .ZN(n6718)
         );
  OAI21_X1 U7455 ( .B1(n6750), .B2(n6899), .A(n6718), .ZN(n6719) );
  AOI21_X1 U7456 ( .B1(n7611), .B2(n6760), .A(n6719), .ZN(n6720) );
  OAI21_X1 U7457 ( .B1(n6754), .B2(n6721), .A(n6720), .ZN(U3037) );
  INV_X1 U7458 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U7459 ( .A1(n7616), .A2(n6747), .B1(n6805), .B2(n6746), .ZN(n6722)
         );
  OAI21_X1 U7460 ( .B1(n6750), .B2(n6723), .A(n6722), .ZN(n6724) );
  AOI21_X1 U7461 ( .B1(n7617), .B2(n6760), .A(n6724), .ZN(n6725) );
  OAI21_X1 U7462 ( .B1(n6754), .B2(n6726), .A(n6725), .ZN(U3038) );
  INV_X1 U7463 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U7464 ( .A1(n7622), .A2(n6747), .B1(n6809), .B2(n6746), .ZN(n6727)
         );
  OAI21_X1 U7465 ( .B1(n6750), .B2(n6728), .A(n6727), .ZN(n6729) );
  AOI21_X1 U7466 ( .B1(n7624), .B2(n6760), .A(n6729), .ZN(n6730) );
  OAI21_X1 U7467 ( .B1(n6754), .B2(n6731), .A(n6730), .ZN(U3039) );
  INV_X1 U7468 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7469 ( .A1(n7628), .A2(n6747), .B1(n6949), .B2(n6746), .ZN(n6732)
         );
  OAI21_X1 U7470 ( .B1(n6750), .B2(n6906), .A(n6732), .ZN(n6733) );
  AOI21_X1 U7471 ( .B1(n7629), .B2(n6760), .A(n6733), .ZN(n6734) );
  OAI21_X1 U7472 ( .B1(n6754), .B2(n6735), .A(n6734), .ZN(U3040) );
  INV_X1 U7473 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7474 ( .A1(n7634), .A2(n6747), .B1(n6816), .B2(n6746), .ZN(n6736)
         );
  OAI21_X1 U7475 ( .B1(n6750), .B2(n6737), .A(n6736), .ZN(n6738) );
  AOI21_X1 U7476 ( .B1(n7635), .B2(n6760), .A(n6738), .ZN(n6739) );
  OAI21_X1 U7477 ( .B1(n6754), .B2(n6740), .A(n6739), .ZN(U3041) );
  INV_X1 U7478 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7479 ( .A1(n7640), .A2(n6747), .B1(n6820), .B2(n6746), .ZN(n6741)
         );
  OAI21_X1 U7480 ( .B1(n6750), .B2(n6742), .A(n6741), .ZN(n6743) );
  AOI21_X1 U7481 ( .B1(n7641), .B2(n6760), .A(n6743), .ZN(n6744) );
  OAI21_X1 U7482 ( .B1(n6754), .B2(n6745), .A(n6744), .ZN(U3042) );
  INV_X1 U7483 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7484 ( .A1(n7647), .A2(n6747), .B1(n6825), .B2(n6746), .ZN(n6748)
         );
  OAI21_X1 U7485 ( .B1(n6750), .B2(n6749), .A(n6748), .ZN(n6751) );
  AOI21_X1 U7486 ( .B1(n7648), .B2(n6760), .A(n6751), .ZN(n6752) );
  OAI21_X1 U7487 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(U3043) );
  INV_X1 U7488 ( .A(n7611), .ZN(n6925) );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6758), .B1(n6944), 
        .B2(n6757), .ZN(n6756) );
  INV_X1 U7490 ( .A(n6899), .ZN(n7612) );
  AOI22_X1 U7491 ( .A1(n6760), .A2(n7612), .B1(n7610), .B2(n6759), .ZN(n6755)
         );
  OAI211_X1 U7492 ( .C1(n6925), .C2(n6772), .A(n6756), .B(n6755), .ZN(U3045)
         );
  INV_X1 U7493 ( .A(n7629), .ZN(n6933) );
  AOI22_X1 U7494 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6758), .B1(n6949), 
        .B2(n6757), .ZN(n6762) );
  INV_X1 U7495 ( .A(n6906), .ZN(n7630) );
  AOI22_X1 U7496 ( .A1(n6760), .A2(n7630), .B1(n7628), .B2(n6759), .ZN(n6761)
         );
  OAI211_X1 U7497 ( .C1(n6933), .C2(n6772), .A(n6762), .B(n6761), .ZN(U3048)
         );
  AOI22_X1 U7498 ( .A1(n7610), .A2(n6768), .B1(n6944), .B2(n6767), .ZN(n6764)
         );
  NAND2_X1 U7499 ( .A1(n6769), .A2(n7611), .ZN(n6763) );
  OAI211_X1 U7500 ( .C1(n6772), .C2(n6899), .A(n6764), .B(n6763), .ZN(n6765)
         );
  AOI21_X1 U7501 ( .B1(n6774), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n6765), 
        .ZN(n6766) );
  INV_X1 U7502 ( .A(n6766), .ZN(U3053) );
  AOI22_X1 U7503 ( .A1(n7628), .A2(n6768), .B1(n6949), .B2(n6767), .ZN(n6771)
         );
  NAND2_X1 U7504 ( .A1(n6769), .A2(n7629), .ZN(n6770) );
  OAI211_X1 U7505 ( .C1(n6772), .C2(n6906), .A(n6771), .B(n6770), .ZN(n6773)
         );
  AOI21_X1 U7506 ( .B1(n6774), .B2(INSTQUEUE_REG_4__4__SCAN_IN), .A(n6773), 
        .ZN(n6775) );
  INV_X1 U7507 ( .A(n6775), .ZN(U3056) );
  AOI22_X1 U7508 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6779), .B1(n6944), 
        .B2(n6778), .ZN(n6777) );
  AOI22_X1 U7509 ( .A1(n6827), .A2(n7611), .B1(n7610), .B2(n6780), .ZN(n6776)
         );
  OAI211_X1 U7510 ( .C1(n6899), .C2(n6783), .A(n6777), .B(n6776), .ZN(U3061)
         );
  AOI22_X1 U7511 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6779), .B1(n6949), 
        .B2(n6778), .ZN(n6782) );
  AOI22_X1 U7512 ( .A1(n6827), .A2(n7629), .B1(n7628), .B2(n6780), .ZN(n6781)
         );
  OAI211_X1 U7513 ( .C1(n6906), .C2(n6783), .A(n6782), .B(n6781), .ZN(U3064)
         );
  NOR2_X1 U7514 ( .A1(n6967), .A2(n7591), .ZN(n7598) );
  AND2_X1 U7515 ( .A1(n6784), .A2(n7598), .ZN(n6826) );
  NOR2_X2 U7516 ( .A1(n6786), .A2(n6785), .ZN(n7652) );
  OAI21_X1 U7517 ( .B1(n7652), .B2(n6827), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6791) );
  NAND2_X1 U7518 ( .A1(n6788), .A2(n6787), .ZN(n6790) );
  AOI21_X1 U7519 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6793) );
  OAI211_X1 U7520 ( .C1(n6826), .C2(n7533), .A(n6793), .B(n6792), .ZN(n6794)
         );
  INV_X1 U7521 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6801) );
  OAI22_X1 U7522 ( .A1(n6797), .A2(n7590), .B1(n6796), .B2(n6795), .ZN(n6824)
         );
  AOI22_X1 U7523 ( .A1(n7596), .A2(n6826), .B1(n6798), .B2(n6824), .ZN(n6800)
         );
  AOI22_X1 U7524 ( .A1(n7597), .A2(n6827), .B1(n7652), .B2(n7606), .ZN(n6799)
         );
  OAI211_X1 U7525 ( .C1(n6831), .C2(n6801), .A(n6800), .B(n6799), .ZN(U3068)
         );
  INV_X1 U7526 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6804) );
  AOI22_X1 U7527 ( .A1(n7610), .A2(n6826), .B1(n6944), .B2(n6824), .ZN(n6803)
         );
  AOI22_X1 U7528 ( .A1(n7612), .A2(n6827), .B1(n7652), .B2(n7611), .ZN(n6802)
         );
  OAI211_X1 U7529 ( .C1(n6831), .C2(n6804), .A(n6803), .B(n6802), .ZN(U3069)
         );
  INV_X1 U7530 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7531 ( .A1(n7616), .A2(n6826), .B1(n6805), .B2(n6824), .ZN(n6807)
         );
  AOI22_X1 U7532 ( .A1(n7618), .A2(n6827), .B1(n7652), .B2(n7617), .ZN(n6806)
         );
  OAI211_X1 U7533 ( .C1(n6831), .C2(n6808), .A(n6807), .B(n6806), .ZN(U3070)
         );
  INV_X1 U7534 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6812) );
  AOI22_X1 U7535 ( .A1(n7622), .A2(n6826), .B1(n6809), .B2(n6824), .ZN(n6811)
         );
  AOI22_X1 U7536 ( .A1(n7623), .A2(n6827), .B1(n7652), .B2(n7624), .ZN(n6810)
         );
  OAI211_X1 U7537 ( .C1(n6831), .C2(n6812), .A(n6811), .B(n6810), .ZN(U3071)
         );
  INV_X1 U7538 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7539 ( .A1(n7628), .A2(n6826), .B1(n6949), .B2(n6824), .ZN(n6814)
         );
  AOI22_X1 U7540 ( .A1(n7630), .A2(n6827), .B1(n7652), .B2(n7629), .ZN(n6813)
         );
  OAI211_X1 U7541 ( .C1(n6831), .C2(n6815), .A(n6814), .B(n6813), .ZN(U3072)
         );
  INV_X1 U7542 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7543 ( .A1(n7634), .A2(n6826), .B1(n6816), .B2(n6824), .ZN(n6818)
         );
  AOI22_X1 U7544 ( .A1(n7636), .A2(n6827), .B1(n7652), .B2(n7635), .ZN(n6817)
         );
  OAI211_X1 U7545 ( .C1(n6831), .C2(n6819), .A(n6818), .B(n6817), .ZN(U3073)
         );
  INV_X1 U7546 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U7547 ( .A1(n7640), .A2(n6826), .B1(n6820), .B2(n6824), .ZN(n6822)
         );
  AOI22_X1 U7548 ( .A1(n7642), .A2(n6827), .B1(n7652), .B2(n7641), .ZN(n6821)
         );
  OAI211_X1 U7549 ( .C1(n6831), .C2(n6823), .A(n6822), .B(n6821), .ZN(U3074)
         );
  INV_X1 U7550 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6830) );
  AOI22_X1 U7551 ( .A1(n7647), .A2(n6826), .B1(n6825), .B2(n6824), .ZN(n6829)
         );
  AOI22_X1 U7552 ( .A1(n7651), .A2(n6827), .B1(n7652), .B2(n7648), .ZN(n6828)
         );
  OAI211_X1 U7553 ( .C1(n6831), .C2(n6830), .A(n6829), .B(n6828), .ZN(U3075)
         );
  INV_X1 U7554 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7555 ( .A1(n7610), .A2(n6837), .B1(n6944), .B2(n6836), .ZN(n6832)
         );
  OAI21_X1 U7556 ( .B1(n6899), .B2(n6839), .A(n6832), .ZN(n6833) );
  AOI21_X1 U7557 ( .B1(n6841), .B2(n7611), .A(n6833), .ZN(n6834) );
  OAI21_X1 U7558 ( .B1(n6844), .B2(n6835), .A(n6834), .ZN(U3085) );
  INV_X1 U7559 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U7560 ( .A1(n7628), .A2(n6837), .B1(n6949), .B2(n6836), .ZN(n6838)
         );
  OAI21_X1 U7561 ( .B1(n6906), .B2(n6839), .A(n6838), .ZN(n6840) );
  AOI21_X1 U7562 ( .B1(n6841), .B2(n7629), .A(n6840), .ZN(n6842) );
  OAI21_X1 U7563 ( .B1(n6844), .B2(n6843), .A(n6842), .ZN(U3088) );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6848), .B1(n6944), 
        .B2(n6847), .ZN(n6846) );
  AOI22_X1 U7565 ( .A1(n6895), .A2(n7611), .B1(n6849), .B2(n7610), .ZN(n6845)
         );
  OAI211_X1 U7566 ( .C1(n6852), .C2(n6899), .A(n6846), .B(n6845), .ZN(U3093)
         );
  AOI22_X1 U7567 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6848), .B1(n6949), 
        .B2(n6847), .ZN(n6851) );
  AOI22_X1 U7568 ( .A1(n6895), .A2(n7629), .B1(n6849), .B2(n7628), .ZN(n6850)
         );
  OAI211_X1 U7569 ( .C1(n6852), .C2(n6906), .A(n6851), .B(n6850), .ZN(U3096)
         );
  NAND2_X1 U7570 ( .A1(n6905), .A2(n7599), .ZN(n6854) );
  OAI21_X1 U7571 ( .B1(n6895), .B2(n6854), .A(n6853), .ZN(n6862) );
  NOR2_X1 U7572 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6857), .ZN(n6891)
         );
  INV_X1 U7573 ( .A(n6858), .ZN(n6861) );
  AOI211_X1 U7574 ( .C1(n6862), .C2(n6861), .A(n6860), .B(n6859), .ZN(n6863)
         );
  OAI21_X1 U7575 ( .B1(n6891), .B2(n7533), .A(n6863), .ZN(n6890) );
  AOI22_X1 U7576 ( .A1(n7596), .A2(n6891), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n6890), .ZN(n6864) );
  OAI21_X1 U7577 ( .B1(n6865), .B2(n6905), .A(n6864), .ZN(n6866) );
  AOI21_X1 U7578 ( .B1(n7597), .B2(n6895), .A(n6866), .ZN(n6867) );
  OAI21_X1 U7579 ( .B1(n6897), .B2(n7609), .A(n6867), .ZN(U3100) );
  INV_X1 U7580 ( .A(n6944), .ZN(n7615) );
  AOI22_X1 U7581 ( .A1(n7610), .A2(n6891), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n6890), .ZN(n6868) );
  OAI21_X1 U7582 ( .B1(n6925), .B2(n6905), .A(n6868), .ZN(n6869) );
  AOI21_X1 U7583 ( .B1(n6895), .B2(n7612), .A(n6869), .ZN(n6870) );
  OAI21_X1 U7584 ( .B1(n6897), .B2(n7615), .A(n6870), .ZN(U3101) );
  AOI22_X1 U7585 ( .A1(n7616), .A2(n6891), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n6890), .ZN(n6871) );
  OAI21_X1 U7586 ( .B1(n6872), .B2(n6905), .A(n6871), .ZN(n6873) );
  AOI21_X1 U7587 ( .B1(n6895), .B2(n7618), .A(n6873), .ZN(n6874) );
  OAI21_X1 U7588 ( .B1(n6897), .B2(n7621), .A(n6874), .ZN(U3102) );
  AOI22_X1 U7589 ( .A1(n7622), .A2(n6891), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n6890), .ZN(n6875) );
  OAI21_X1 U7590 ( .B1(n6876), .B2(n6905), .A(n6875), .ZN(n6877) );
  AOI21_X1 U7591 ( .B1(n6895), .B2(n7623), .A(n6877), .ZN(n6878) );
  OAI21_X1 U7592 ( .B1(n6897), .B2(n7627), .A(n6878), .ZN(U3103) );
  INV_X1 U7593 ( .A(n6949), .ZN(n7633) );
  AOI22_X1 U7594 ( .A1(n7628), .A2(n6891), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n6890), .ZN(n6879) );
  OAI21_X1 U7595 ( .B1(n6933), .B2(n6905), .A(n6879), .ZN(n6880) );
  AOI21_X1 U7596 ( .B1(n6895), .B2(n7630), .A(n6880), .ZN(n6881) );
  OAI21_X1 U7597 ( .B1(n6897), .B2(n7633), .A(n6881), .ZN(U3104) );
  AOI22_X1 U7598 ( .A1(n7634), .A2(n6891), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n6890), .ZN(n6882) );
  OAI21_X1 U7599 ( .B1(n6883), .B2(n6905), .A(n6882), .ZN(n6884) );
  AOI21_X1 U7600 ( .B1(n6895), .B2(n7636), .A(n6884), .ZN(n6885) );
  OAI21_X1 U7601 ( .B1(n6897), .B2(n7639), .A(n6885), .ZN(U3105) );
  AOI22_X1 U7602 ( .A1(n7640), .A2(n6891), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n6890), .ZN(n6886) );
  OAI21_X1 U7603 ( .B1(n6887), .B2(n6905), .A(n6886), .ZN(n6888) );
  AOI21_X1 U7604 ( .B1(n6895), .B2(n7642), .A(n6888), .ZN(n6889) );
  OAI21_X1 U7605 ( .B1(n6897), .B2(n7645), .A(n6889), .ZN(U3106) );
  AOI22_X1 U7606 ( .A1(n7647), .A2(n6891), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n6890), .ZN(n6892) );
  OAI21_X1 U7607 ( .B1(n6893), .B2(n6905), .A(n6892), .ZN(n6894) );
  AOI21_X1 U7608 ( .B1(n6895), .B2(n7651), .A(n6894), .ZN(n6896) );
  OAI21_X1 U7609 ( .B1(n6897), .B2(n7655), .A(n6896), .ZN(U3107) );
  AOI22_X1 U7610 ( .A1(n7610), .A2(n6903), .B1(INSTQUEUE_REG_11__1__SCAN_IN), 
        .B2(n6902), .ZN(n6898) );
  OAI21_X1 U7611 ( .B1(n6899), .B2(n6905), .A(n6898), .ZN(n6900) );
  AOI21_X1 U7612 ( .B1(n7611), .B2(n6919), .A(n6900), .ZN(n6901) );
  OAI21_X1 U7613 ( .B1(n6909), .B2(n7615), .A(n6901), .ZN(U3109) );
  AOI22_X1 U7614 ( .A1(n7628), .A2(n6903), .B1(INSTQUEUE_REG_11__4__SCAN_IN), 
        .B2(n6902), .ZN(n6904) );
  OAI21_X1 U7615 ( .B1(n6906), .B2(n6905), .A(n6904), .ZN(n6907) );
  AOI21_X1 U7616 ( .B1(n7629), .B2(n6919), .A(n6907), .ZN(n6908) );
  OAI21_X1 U7617 ( .B1(n6909), .B2(n7633), .A(n6908), .ZN(U3112) );
  INV_X1 U7618 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7619 ( .A1(n7610), .A2(n6915), .B1(n6944), .B2(n6914), .ZN(n6910)
         );
  OAI21_X1 U7620 ( .B1(n6917), .B2(n6925), .A(n6910), .ZN(n6911) );
  AOI21_X1 U7621 ( .B1(n7612), .B2(n6919), .A(n6911), .ZN(n6912) );
  OAI21_X1 U7622 ( .B1(n6922), .B2(n6913), .A(n6912), .ZN(U3117) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U7624 ( .A1(n7628), .A2(n6915), .B1(n6949), .B2(n6914), .ZN(n6916)
         );
  OAI21_X1 U7625 ( .B1(n6917), .B2(n6933), .A(n6916), .ZN(n6918) );
  AOI21_X1 U7626 ( .B1(n7630), .B2(n6919), .A(n6918), .ZN(n6920) );
  OAI21_X1 U7627 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(U3120) );
  AOI22_X1 U7628 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6927), .B1(n6944), 
        .B2(n6926), .ZN(n6924) );
  AOI22_X1 U7629 ( .A1(n6929), .A2(n7612), .B1(n7610), .B2(n6928), .ZN(n6923)
         );
  OAI211_X1 U7630 ( .C1(n6925), .C2(n6932), .A(n6924), .B(n6923), .ZN(U3125)
         );
  AOI22_X1 U7631 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6927), .B1(n6949), 
        .B2(n6926), .ZN(n6931) );
  AOI22_X1 U7632 ( .A1(n6929), .A2(n7630), .B1(n7628), .B2(n6928), .ZN(n6930)
         );
  OAI211_X1 U7633 ( .C1(n6933), .C2(n6932), .A(n6931), .B(n6930), .ZN(U3128)
         );
  INV_X1 U7634 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7635 ( .A1(n7610), .A2(n6938), .B1(n6944), .B2(n6937), .ZN(n6935)
         );
  AOI22_X1 U7636 ( .A1(n7612), .A2(n6939), .B1(n6951), .B2(n7611), .ZN(n6934)
         );
  OAI211_X1 U7637 ( .C1(n6943), .C2(n6936), .A(n6935), .B(n6934), .ZN(U3133)
         );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U7639 ( .A1(n7628), .A2(n6938), .B1(n6949), .B2(n6937), .ZN(n6941)
         );
  AOI22_X1 U7640 ( .A1(n7630), .A2(n6939), .B1(n6951), .B2(n7629), .ZN(n6940)
         );
  OAI211_X1 U7641 ( .C1(n6943), .C2(n6942), .A(n6941), .B(n6940), .ZN(U3136)
         );
  INV_X1 U7642 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6947) );
  AOI22_X1 U7643 ( .A1(n7610), .A2(n6950), .B1(n6944), .B2(n6948), .ZN(n6946)
         );
  AOI22_X1 U7644 ( .A1(n7611), .A2(n6952), .B1(n6951), .B2(n7612), .ZN(n6945)
         );
  OAI211_X1 U7645 ( .C1(n6956), .C2(n6947), .A(n6946), .B(n6945), .ZN(U3141)
         );
  INV_X1 U7646 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7647 ( .A1(n7628), .A2(n6950), .B1(n6949), .B2(n6948), .ZN(n6954)
         );
  AOI22_X1 U7648 ( .A1(n7629), .A2(n6952), .B1(n6951), .B2(n7630), .ZN(n6953)
         );
  OAI211_X1 U7649 ( .C1(n6956), .C2(n6955), .A(n6954), .B(n6953), .ZN(U3144)
         );
  INV_X1 U7650 ( .A(n6957), .ZN(n6974) );
  NAND2_X1 U7651 ( .A1(n6958), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U7652 ( .A1(n6959), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6960) );
  NOR2_X1 U7653 ( .A1(n6961), .A2(n6960), .ZN(n6965) );
  INV_X1 U7654 ( .A(n6965), .ZN(n6968) );
  INV_X1 U7655 ( .A(n6962), .ZN(n6964) );
  OAI22_X1 U7656 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6965), .B1(n6964), .B2(n6963), .ZN(n6966) );
  OAI21_X1 U7657 ( .B1(n6968), .B2(n6967), .A(n6966), .ZN(n6970) );
  AOI222_X1 U7658 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6970), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6969), .C1(n6970), .C2(n6969), 
        .ZN(n6971) );
  INV_X1 U7659 ( .A(n6971), .ZN(n6972) );
  AND2_X1 U7660 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6972), .ZN(n6973)
         );
  OAI22_X1 U7661 ( .A1(n6974), .A2(n6973), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6972), .ZN(n6981) );
  NOR2_X1 U7662 ( .A1(MORE_REG_SCAN_IN), .A2(FLUSH_REG_SCAN_IN), .ZN(n6978) );
  NOR2_X1 U7663 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  OAI21_X1 U7664 ( .B1(n6979), .B2(n6978), .A(n6977), .ZN(n6980) );
  AOI21_X1 U7665 ( .B1(n6981), .B2(n7016), .A(n6980), .ZN(n6982) );
  NAND3_X1 U7666 ( .A1(n6984), .A2(n6983), .A3(n6982), .ZN(n6994) );
  OAI22_X1 U7667 ( .A1(n6994), .A2(n6986), .B1(n7546), .B2(n6985), .ZN(n6990)
         );
  OR2_X1 U7668 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  NAND2_X1 U7669 ( .A1(n6990), .A2(n6989), .ZN(n7532) );
  NAND2_X1 U7670 ( .A1(READY_N), .A2(n7200), .ZN(n7196) );
  AOI21_X1 U7671 ( .B1(n7532), .B2(n7196), .A(n4049), .ZN(n7525) );
  INV_X1 U7672 ( .A(n7525), .ZN(n6997) );
  NOR2_X1 U7673 ( .A1(n6991), .A2(n7531), .ZN(n6992) );
  AOI211_X1 U7674 ( .C1(n7522), .C2(n6994), .A(n6993), .B(n6992), .ZN(n6996)
         );
  OAI211_X1 U7675 ( .C1(n7505), .C2(n7203), .A(n7532), .B(n4049), .ZN(n6995)
         );
  NAND3_X1 U7676 ( .A1(n6997), .A2(n6996), .A3(n6995), .ZN(U3148) );
  INV_X1 U7677 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7000) );
  AND2_X1 U7678 ( .A1(n6998), .A2(STATE_REG_1__SCAN_IN), .ZN(n7541) );
  NOR2_X1 U7679 ( .A1(n7547), .A2(n7541), .ZN(n7018) );
  NOR2_X2 U7680 ( .A1(n7556), .A2(n7018), .ZN(n7538) );
  INV_X1 U7681 ( .A(n7538), .ZN(n7014) );
  NAND2_X1 U7682 ( .A1(n6998), .A2(n7547), .ZN(n7192) );
  AOI21_X1 U7683 ( .B1(n6999), .B2(n7192), .A(n7014), .ZN(n7534) );
  AOI21_X1 U7684 ( .B1(n7000), .B2(n7014), .A(n7534), .ZN(U3451) );
  AND2_X1 U7685 ( .A1(n7014), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  AND2_X1 U7686 ( .A1(n7014), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  NOR2_X1 U7687 ( .A1(n7538), .A2(n7001), .ZN(U3178) );
  NOR2_X1 U7688 ( .A1(n7538), .A2(n7002), .ZN(U3177) );
  NOR2_X1 U7689 ( .A1(n7538), .A2(n7003), .ZN(U3176) );
  NOR2_X1 U7690 ( .A1(n7538), .A2(n7004), .ZN(U3175) );
  AND2_X1 U7691 ( .A1(n7014), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  NOR2_X1 U7692 ( .A1(n7538), .A2(n7005), .ZN(U3173) );
  AND2_X1 U7693 ( .A1(n7014), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  NOR2_X1 U7694 ( .A1(n7538), .A2(n7006), .ZN(U3171) );
  AND2_X1 U7695 ( .A1(n7014), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  NOR2_X1 U7696 ( .A1(n7538), .A2(n7007), .ZN(U3169) );
  NOR2_X1 U7697 ( .A1(n7538), .A2(n7008), .ZN(U3168) );
  NOR2_X1 U7698 ( .A1(n7538), .A2(n7009), .ZN(U3167) );
  AND2_X1 U7699 ( .A1(n7014), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7700 ( .A1(n7014), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  NOR2_X1 U7701 ( .A1(n7538), .A2(n7010), .ZN(U3164) );
  NOR2_X1 U7702 ( .A1(n7538), .A2(n7011), .ZN(U3163) );
  AND2_X1 U7703 ( .A1(n7014), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  INV_X1 U7704 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U7705 ( .A1(n7538), .A2(n7012), .ZN(U3161) );
  NOR2_X1 U7706 ( .A1(n7538), .A2(n7013), .ZN(U3160) );
  AND2_X1 U7707 ( .A1(n7014), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7708 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7014), .ZN(U3158) );
  AND2_X1 U7709 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7014), .ZN(U3157) );
  AND2_X1 U7710 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7014), .ZN(U3156) );
  AND2_X1 U7711 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7014), .ZN(U3155) );
  AND2_X1 U7712 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7014), .ZN(U3154) );
  AND2_X1 U7713 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7014), .ZN(U3153) );
  AND2_X1 U7714 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7014), .ZN(U3152) );
  AND2_X1 U7715 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7014), .ZN(U3151) );
  NOR2_X1 U7716 ( .A1(n7016), .A2(n7015), .ZN(U3019) );
  AND2_X1 U7717 ( .A1(n7031), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7718 ( .B1(n7018), .B2(n7017), .A(n7556), .ZN(U2789) );
  AOI22_X1 U7719 ( .A1(n7048), .A2(LWORD_REG_0__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n7020) );
  OAI21_X1 U7720 ( .B1(n7021), .B2(n7050), .A(n7020), .ZN(U2923) );
  AOI22_X1 U7721 ( .A1(n7048), .A2(LWORD_REG_1__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U7722 ( .B1(n7023), .B2(n7050), .A(n7022), .ZN(U2922) );
  AOI22_X1 U7723 ( .A1(n7048), .A2(LWORD_REG_2__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n7024) );
  OAI21_X1 U7724 ( .B1(n7025), .B2(n7050), .A(n7024), .ZN(U2921) );
  AOI22_X1 U7725 ( .A1(n7048), .A2(LWORD_REG_3__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7026) );
  OAI21_X1 U7726 ( .B1(n7027), .B2(n7050), .A(n7026), .ZN(U2920) );
  AOI22_X1 U7727 ( .A1(n7048), .A2(LWORD_REG_4__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7028) );
  OAI21_X1 U7728 ( .B1(n7029), .B2(n7050), .A(n7028), .ZN(U2919) );
  AOI22_X1 U7729 ( .A1(n7048), .A2(LWORD_REG_5__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7030) );
  OAI21_X1 U7730 ( .B1(n4299), .B2(n7050), .A(n7030), .ZN(U2918) );
  AOI22_X1 U7731 ( .A1(n7048), .A2(LWORD_REG_6__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7032) );
  OAI21_X1 U7732 ( .B1(n4308), .B2(n7050), .A(n7032), .ZN(U2917) );
  AOI22_X1 U7733 ( .A1(n7048), .A2(LWORD_REG_7__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7033) );
  OAI21_X1 U7734 ( .B1(n4314), .B2(n7050), .A(n7033), .ZN(U2916) );
  AOI22_X1 U7735 ( .A1(n7048), .A2(LWORD_REG_8__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7034) );
  OAI21_X1 U7736 ( .B1(n7035), .B2(n7050), .A(n7034), .ZN(U2915) );
  AOI22_X1 U7737 ( .A1(n7048), .A2(LWORD_REG_9__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7036) );
  OAI21_X1 U7738 ( .B1(n7037), .B2(n7050), .A(n7036), .ZN(U2914) );
  AOI22_X1 U7739 ( .A1(n7048), .A2(LWORD_REG_10__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7038) );
  OAI21_X1 U7740 ( .B1(n7039), .B2(n7050), .A(n7038), .ZN(U2913) );
  AOI22_X1 U7741 ( .A1(n7048), .A2(LWORD_REG_11__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7040) );
  OAI21_X1 U7742 ( .B1(n7041), .B2(n7050), .A(n7040), .ZN(U2912) );
  AOI22_X1 U7743 ( .A1(n7048), .A2(LWORD_REG_12__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7042) );
  OAI21_X1 U7744 ( .B1(n7043), .B2(n7050), .A(n7042), .ZN(U2911) );
  AOI22_X1 U7745 ( .A1(n7048), .A2(LWORD_REG_13__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U7746 ( .B1(n7045), .B2(n7050), .A(n7044), .ZN(U2910) );
  AOI22_X1 U7747 ( .A1(n7048), .A2(LWORD_REG_14__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7046) );
  OAI21_X1 U7748 ( .B1(n7047), .B2(n7050), .A(n7046), .ZN(U2909) );
  AOI22_X1 U7749 ( .A1(n7048), .A2(LWORD_REG_15__SCAN_IN), .B1(n7031), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7049) );
  OAI21_X1 U7750 ( .B1(n7051), .B2(n7050), .A(n7049), .ZN(U2908) );
  INV_X1 U7751 ( .A(n7069), .ZN(n7099) );
  INV_X1 U7752 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7249) );
  INV_X1 U7753 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7052) );
  OAI222_X1 U7754 ( .A1(n7099), .A2(n7249), .B1(n7052), .B2(n7556), .C1(n7114), 
        .C2(n7095), .ZN(U3184) );
  OAI222_X1 U7755 ( .A1(n7099), .A2(n7054), .B1(n7053), .B2(n7556), .C1(n7249), 
        .C2(n7095), .ZN(U3185) );
  INV_X1 U7756 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7055) );
  OAI222_X1 U7757 ( .A1(n7099), .A2(n7328), .B1(n7055), .B2(n7556), .C1(n7054), 
        .C2(n7095), .ZN(U3186) );
  AOI222_X1 U7758 ( .A1(n7069), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7553), .C1(REIP_REG_4__SCAN_IN), .C2(
        n7068), .ZN(n7056) );
  INV_X1 U7759 ( .A(n7056), .ZN(U3187) );
  AOI222_X1 U7760 ( .A1(n7069), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7553), .C1(REIP_REG_5__SCAN_IN), .C2(
        n7068), .ZN(n7057) );
  INV_X1 U7761 ( .A(n7057), .ZN(U3188) );
  INV_X1 U7762 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7365) );
  OAI222_X1 U7763 ( .A1(n7099), .A2(n7364), .B1(n7058), .B2(n7556), .C1(n7365), 
        .C2(n7095), .ZN(U3189) );
  INV_X1 U7764 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7059) );
  OAI222_X1 U7765 ( .A1(n7099), .A2(n5996), .B1(n7059), .B2(n7556), .C1(n7364), 
        .C2(n7095), .ZN(U3190) );
  INV_X1 U7766 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7060) );
  OAI222_X1 U7767 ( .A1(n7099), .A2(n7061), .B1(n7060), .B2(n7556), .C1(n5996), 
        .C2(n7095), .ZN(U3191) );
  OAI222_X1 U7768 ( .A1(n7099), .A2(n6049), .B1(n7062), .B2(n7556), .C1(n7061), 
        .C2(n7095), .ZN(U3192) );
  INV_X1 U7769 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7063) );
  OAI222_X1 U7770 ( .A1(n7099), .A2(n7064), .B1(n7063), .B2(n7556), .C1(n6049), 
        .C2(n7095), .ZN(U3193) );
  AOI222_X1 U7771 ( .A1(n7068), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7553), .C1(REIP_REG_13__SCAN_IN), .C2(
        n7069), .ZN(n7065) );
  INV_X1 U7772 ( .A(n7065), .ZN(U3195) );
  AOI222_X1 U7773 ( .A1(n7069), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7553), .C1(REIP_REG_13__SCAN_IN), .C2(
        n7068), .ZN(n7066) );
  INV_X1 U7774 ( .A(n7066), .ZN(U3196) );
  AOI222_X1 U7775 ( .A1(n7069), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7553), .C1(REIP_REG_14__SCAN_IN), .C2(
        n7068), .ZN(n7067) );
  INV_X1 U7776 ( .A(n7067), .ZN(U3197) );
  AOI222_X1 U7777 ( .A1(n7069), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7553), .C1(REIP_REG_15__SCAN_IN), .C2(
        n7068), .ZN(n7070) );
  INV_X1 U7778 ( .A(n7070), .ZN(U3198) );
  INV_X1 U7779 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7438) );
  OAI222_X1 U7780 ( .A1(n7099), .A2(n7438), .B1(n7072), .B2(n7556), .C1(n7071), 
        .C2(n7095), .ZN(U3199) );
  INV_X1 U7781 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7073) );
  OAI222_X1 U7782 ( .A1(n7099), .A2(n7074), .B1(n7073), .B2(n7556), .C1(n7438), 
        .C2(n7095), .ZN(U3200) );
  INV_X1 U7783 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7075) );
  OAI222_X1 U7784 ( .A1(n7099), .A2(n7445), .B1(n7075), .B2(n7556), .C1(n7074), 
        .C2(n7095), .ZN(U3201) );
  OAI222_X1 U7785 ( .A1(n7095), .A2(n7445), .B1(n7076), .B2(n7556), .C1(n7078), 
        .C2(n7099), .ZN(U3202) );
  INV_X1 U7786 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7463) );
  OAI222_X1 U7787 ( .A1(n7095), .A2(n7078), .B1(n7077), .B2(n7556), .C1(n7463), 
        .C2(n7099), .ZN(U3203) );
  INV_X1 U7788 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7079) );
  OAI222_X1 U7789 ( .A1(n7095), .A2(n7463), .B1(n7079), .B2(n7556), .C1(n7482), 
        .C2(n7099), .ZN(U3204) );
  INV_X1 U7790 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7080) );
  OAI222_X1 U7791 ( .A1(n7099), .A2(n7082), .B1(n7080), .B2(n7556), .C1(n7482), 
        .C2(n7095), .ZN(U3205) );
  OAI222_X1 U7792 ( .A1(n7095), .A2(n7082), .B1(n7081), .B2(n7556), .C1(n7083), 
        .C2(n7099), .ZN(U3206) );
  OAI222_X1 U7793 ( .A1(n7099), .A2(n7086), .B1(n7084), .B2(n7556), .C1(n7083), 
        .C2(n7095), .ZN(U3207) );
  OAI222_X1 U7794 ( .A1(n7095), .A2(n7086), .B1(n7085), .B2(n7556), .C1(n7088), 
        .C2(n7099), .ZN(U3208) );
  INV_X1 U7795 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7087) );
  OAI222_X1 U7796 ( .A1(n7095), .A2(n7088), .B1(n7087), .B2(n7556), .C1(n7090), 
        .C2(n7099), .ZN(U3209) );
  INV_X1 U7797 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7089) );
  OAI222_X1 U7798 ( .A1(n7095), .A2(n7090), .B1(n7089), .B2(n7556), .C1(n7092), 
        .C2(n7099), .ZN(U3210) );
  INV_X1 U7799 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7091) );
  OAI222_X1 U7800 ( .A1(n7095), .A2(n7092), .B1(n7091), .B2(n7556), .C1(n7094), 
        .C2(n7099), .ZN(U3211) );
  OAI222_X1 U7801 ( .A1(n7095), .A2(n7094), .B1(n7093), .B2(n7556), .C1(n7096), 
        .C2(n7099), .ZN(U3212) );
  INV_X1 U7802 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7098) );
  OAI222_X1 U7803 ( .A1(n7099), .A2(n7098), .B1(n7097), .B2(n7556), .C1(n7096), 
        .C2(n7095), .ZN(U3213) );
  AOI22_X1 U7804 ( .A1(n7556), .A2(n7101), .B1(n7100), .B2(n7553), .ZN(U3445)
         );
  AOI221_X1 U7805 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7112) );
  NOR4_X1 U7806 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7105) );
  NOR4_X1 U7807 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n7104) );
  NOR4_X1 U7808 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n7103) );
  NOR4_X1 U7809 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n7102) );
  NAND4_X1 U7810 ( .A1(n7105), .A2(n7104), .A3(n7103), .A4(n7102), .ZN(n7111)
         );
  NOR4_X1 U7811 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(
        n7109) );
  AOI211_X1 U7812 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n7108) );
  NOR4_X1 U7813 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n7107) );
  NOR4_X1 U7814 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7106) );
  NAND4_X1 U7815 ( .A1(n7109), .A2(n7108), .A3(n7107), .A4(n7106), .ZN(n7110)
         );
  NOR2_X1 U7816 ( .A1(n7111), .A2(n7110), .ZN(n7125) );
  MUX2_X1 U7817 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7112), .S(n7125), .Z(
        U2795) );
  INV_X1 U7818 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7117) );
  AOI22_X1 U7819 ( .A1(n7556), .A2(n7117), .B1(n7113), .B2(n7553), .ZN(U3446)
         );
  AOI21_X1 U7820 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7115) );
  OAI221_X1 U7821 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7115), .C1(n7114), .C2(
        REIP_REG_0__SCAN_IN), .A(n7125), .ZN(n7116) );
  OAI21_X1 U7822 ( .B1(n7125), .B2(n7117), .A(n7116), .ZN(U3468) );
  AOI22_X1 U7823 ( .A1(n7556), .A2(n7121), .B1(n7118), .B2(n7553), .ZN(U3447)
         );
  NOR3_X1 U7824 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7119) );
  OAI21_X1 U7825 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7119), .A(n7125), .ZN(n7120)
         );
  OAI21_X1 U7826 ( .B1(n7125), .B2(n7121), .A(n7120), .ZN(U2794) );
  INV_X1 U7827 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7124) );
  AOI22_X1 U7828 ( .A1(n7556), .A2(n7124), .B1(n7122), .B2(n7553), .ZN(U3448)
         );
  OAI21_X1 U7829 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n7125), .ZN(n7123) );
  OAI21_X1 U7830 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(U3469) );
  INV_X1 U7831 ( .A(n7126), .ZN(n7152) );
  INV_X1 U7832 ( .A(n7127), .ZN(n7140) );
  AOI22_X1 U7833 ( .A1(n7152), .A2(n7140), .B1(n7139), .B2(n7247), .ZN(n7128)
         );
  OAI21_X1 U7834 ( .B1(n7143), .B2(n7129), .A(n7128), .ZN(U2857) );
  INV_X1 U7835 ( .A(EBX_REG_8__SCAN_IN), .ZN(n7131) );
  AOI22_X1 U7836 ( .A1(n7383), .A2(n7140), .B1(n7139), .B2(n7377), .ZN(n7130)
         );
  OAI21_X1 U7837 ( .B1(n7143), .B2(n7131), .A(n7130), .ZN(U2851) );
  AOI22_X1 U7838 ( .A1(n7402), .A2(n7140), .B1(n7139), .B2(n7399), .ZN(n7132)
         );
  OAI21_X1 U7839 ( .B1(n7143), .B2(n7396), .A(n7132), .ZN(U2846) );
  INV_X1 U7840 ( .A(n7133), .ZN(n7411) );
  AOI22_X1 U7841 ( .A1(n7419), .A2(n7140), .B1(n7139), .B2(n7411), .ZN(n7134)
         );
  OAI21_X1 U7842 ( .B1(n7143), .B2(n7413), .A(n7134), .ZN(U2845) );
  INV_X1 U7843 ( .A(EBX_REG_4__SCAN_IN), .ZN(n7142) );
  AND2_X1 U7844 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  NOR2_X1 U7845 ( .A1(n7138), .A2(n7137), .ZN(n7334) );
  AOI22_X1 U7846 ( .A1(n7330), .A2(n7140), .B1(n7139), .B2(n7334), .ZN(n7141)
         );
  OAI21_X1 U7847 ( .B1(n7143), .B2(n7142), .A(n7141), .ZN(U2855) );
  INV_X1 U7848 ( .A(n7144), .ZN(n7145) );
  AOI22_X1 U7849 ( .A1(n7186), .A2(n7145), .B1(n7185), .B2(n7323), .ZN(n7149)
         );
  INV_X1 U7850 ( .A(n7146), .ZN(n7147) );
  OAI21_X1 U7851 ( .B1(n7183), .B2(n7147), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n7148) );
  OAI211_X1 U7852 ( .C1(n5016), .C2(n7248), .A(n7149), .B(n7148), .ZN(U2986)
         );
  AOI22_X1 U7853 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7154) );
  XNOR2_X1 U7854 ( .A(n7150), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7151)
         );
  AOI22_X1 U7855 ( .A1(n7257), .A2(n7186), .B1(n7185), .B2(n7152), .ZN(n7153)
         );
  OAI211_X1 U7856 ( .C1(n7190), .C2(n7155), .A(n7154), .B(n7153), .ZN(U2984)
         );
  AOI22_X1 U7857 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n7161) );
  INV_X1 U7858 ( .A(n7158), .ZN(n7159) );
  AOI21_X1 U7859 ( .B1(n7156), .B2(n7157), .A(n7159), .ZN(n7218) );
  AOI22_X1 U7860 ( .A1(n7218), .A2(n7186), .B1(n7185), .B2(n7330), .ZN(n7160)
         );
  OAI211_X1 U7861 ( .C1(n7190), .C2(n7340), .A(n7161), .B(n7160), .ZN(U2982)
         );
  AOI22_X1 U7862 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n7166) );
  OAI22_X1 U7863 ( .A1(n7241), .A2(n7501), .B1(n7174), .B2(n7341), .ZN(n7164)
         );
  INV_X1 U7864 ( .A(n7164), .ZN(n7165) );
  OAI211_X1 U7865 ( .C1(n7190), .C2(n7353), .A(n7166), .B(n7165), .ZN(U2981)
         );
  AOI22_X1 U7866 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n7171) );
  XNOR2_X1 U7867 ( .A(n7167), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7168)
         );
  XNOR2_X1 U7868 ( .A(n7169), .B(n7168), .ZN(n7232) );
  AOI22_X1 U7869 ( .A1(n7232), .A2(n7186), .B1(n7185), .B2(n7354), .ZN(n7170)
         );
  OAI211_X1 U7870 ( .C1(n7190), .C2(n7363), .A(n7171), .B(n7170), .ZN(U2980)
         );
  AOI22_X1 U7871 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n7178) );
  INV_X1 U7872 ( .A(n7172), .ZN(n7173) );
  OAI22_X1 U7873 ( .A1(n7175), .A2(n7174), .B1(n7190), .B2(n7173), .ZN(n7176)
         );
  INV_X1 U7874 ( .A(n7176), .ZN(n7177) );
  OAI211_X1 U7875 ( .C1(n7501), .C2(n7179), .A(n7178), .B(n7177), .ZN(U2975)
         );
  AOI22_X1 U7876 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n7182) );
  XNOR2_X1 U7877 ( .A(n3618), .B(n7302), .ZN(n7180) );
  XNOR2_X1 U7878 ( .A(n6442), .B(n7180), .ZN(n7304) );
  AOI22_X1 U7879 ( .A1(n7304), .A2(n7186), .B1(n7185), .B2(n7557), .ZN(n7181)
         );
  OAI211_X1 U7880 ( .C1(n7190), .C2(n7435), .A(n7182), .B(n7181), .ZN(U2969)
         );
  AOI22_X1 U7881 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n7183), .B1(n7280), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n7189) );
  AOI22_X1 U7882 ( .A1(n7187), .A2(n7186), .B1(n7185), .B2(n7563), .ZN(n7188)
         );
  OAI211_X1 U7883 ( .C1(n7190), .C2(n7448), .A(n7189), .B(n7188), .ZN(U2967)
         );
  NOR2_X1 U7884 ( .A1(n7556), .A2(D_C_N_REG_SCAN_IN), .ZN(n7191) );
  AOI22_X1 U7885 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7556), .B1(n7192), .B2(
        n7191), .ZN(U2791) );
  AOI22_X1 U7886 ( .A1(n7556), .A2(READREQUEST_REG_SCAN_IN), .B1(n7193), .B2(
        n7553), .ZN(U3470) );
  AND2_X1 U7887 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7540) );
  INV_X1 U7888 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7539) );
  NOR2_X1 U7889 ( .A1(n7547), .A2(n7539), .ZN(n7545) );
  AOI21_X1 U7890 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7545), .ZN(n7195)
         );
  NAND2_X1 U7891 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7551) );
  OAI211_X1 U7892 ( .C1(n7540), .C2(n7195), .A(n7194), .B(n7551), .ZN(U3182)
         );
  OAI221_X1 U7893 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(STATE2_REG_1__SCAN_IN), .A(n7196), 
        .ZN(n7198) );
  OAI21_X1 U7894 ( .B1(n7199), .B2(n7198), .A(n7197), .ZN(U3150) );
  AND2_X1 U7895 ( .A1(n7202), .A2(n7201), .ZN(n7204) );
  OAI21_X1 U7896 ( .B1(n7204), .B2(n4049), .A(n7203), .ZN(n7208) );
  AOI211_X1 U7897 ( .C1(n7048), .C2(n7546), .A(n7206), .B(n7205), .ZN(n7207)
         );
  MUX2_X1 U7898 ( .A(n7208), .B(REQUESTPENDING_REG_SCAN_IN), .S(n7207), .Z(
        U3472) );
  NAND2_X1 U7899 ( .A1(n7210), .A2(n7209), .ZN(n7216) );
  AOI22_X1 U7900 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n7211), .B1(n7280), .B2(REIP_REG_20__SCAN_IN), .ZN(n7215) );
  AOI22_X1 U7901 ( .A1(n7213), .A2(n7314), .B1(n7313), .B2(n7212), .ZN(n7214)
         );
  OAI211_X1 U7902 ( .C1(n7217), .C2(n7216), .A(n7215), .B(n7214), .ZN(U2998)
         );
  AOI22_X1 U7903 ( .A1(n7313), .A2(n7334), .B1(n7280), .B2(REIP_REG_4__SCAN_IN), .ZN(n7222) );
  AOI22_X1 U7904 ( .A1(n7218), .A2(n7314), .B1(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .B2(n7224), .ZN(n7221) );
  OAI211_X1 U7905 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7219), .B(n7227), .ZN(n7220) );
  NAND3_X1 U7906 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(U3014) );
  NAND2_X1 U7907 ( .A1(n7260), .A2(n7223), .ZN(n7236) );
  AOI21_X1 U7908 ( .B1(n7252), .B2(n7236), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n7225) );
  AOI211_X1 U7909 ( .C1(n7227), .C2(n7226), .A(n7225), .B(n7224), .ZN(n7246)
         );
  INV_X1 U7910 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7235) );
  INV_X1 U7911 ( .A(n7359), .ZN(n7228) );
  AOI22_X1 U7912 ( .A1(n7313), .A2(n7228), .B1(n7280), .B2(REIP_REG_6__SCAN_IN), .ZN(n7234) );
  NOR3_X1 U7913 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n7230), .A3(n7229), 
        .ZN(n7231) );
  AOI22_X1 U7914 ( .A1(n7232), .A2(n7314), .B1(n7231), .B2(n7238), .ZN(n7233)
         );
  OAI211_X1 U7915 ( .C1(n7246), .C2(n7235), .A(n7234), .B(n7233), .ZN(U3012)
         );
  INV_X1 U7916 ( .A(n7236), .ZN(n7237) );
  AOI211_X1 U7917 ( .C1(n7298), .C2(n7238), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .B(n7237), .ZN(n7245) );
  OAI22_X1 U7918 ( .A1(n7241), .A2(n7240), .B1(n7239), .B2(n7301), .ZN(n7242)
         );
  INV_X1 U7919 ( .A(n7242), .ZN(n7244) );
  NAND2_X1 U7920 ( .A1(n7280), .A2(REIP_REG_5__SCAN_IN), .ZN(n7243) );
  OAI211_X1 U7921 ( .C1(n7246), .C2(n7245), .A(n7244), .B(n7243), .ZN(U3013)
         );
  INV_X1 U7922 ( .A(n7247), .ZN(n7250) );
  OAI22_X1 U7923 ( .A1(n7301), .A2(n7250), .B1(n7249), .B2(n7248), .ZN(n7254)
         );
  NAND3_X1 U7924 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n7251) );
  NOR2_X1 U7925 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  NOR2_X1 U7926 ( .A1(n7254), .A2(n7253), .ZN(n7264) );
  OAI21_X1 U7927 ( .B1(n7256), .B2(n7255), .A(n7300), .ZN(n7258) );
  AOI22_X1 U7928 ( .A1(n7258), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n7314), 
        .B2(n7257), .ZN(n7263) );
  NAND3_X1 U7929 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7260), .A3(n7259), 
        .ZN(n7261) );
  NAND4_X1 U7930 ( .A1(n7264), .A2(n7263), .A3(n7262), .A4(n7261), .ZN(U3016)
         );
  AOI22_X1 U7931 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n7265), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6046), .ZN(n7272) );
  AOI21_X1 U7932 ( .B1(n7313), .B2(n7267), .A(n7266), .ZN(n7271) );
  AOI22_X1 U7933 ( .A1(n7269), .A2(n7314), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7268), .ZN(n7270) );
  OAI211_X1 U7934 ( .C1(n7273), .C2(n7272), .A(n7271), .B(n7270), .ZN(U3008)
         );
  AOI221_X1 U7935 ( .B1(n7298), .B2(n7276), .C1(n7275), .C2(n7276), .A(n7274), 
        .ZN(n7284) );
  AOI21_X1 U7936 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n7277), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n7283) );
  AOI22_X1 U7937 ( .A1(n7279), .A2(n7314), .B1(n7313), .B2(n7278), .ZN(n7282)
         );
  NAND2_X1 U7938 ( .A1(n7280), .A2(REIP_REG_12__SCAN_IN), .ZN(n7281) );
  OAI211_X1 U7939 ( .C1(n7284), .C2(n7283), .A(n7282), .B(n7281), .ZN(U3006)
         );
  AOI22_X1 U7940 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n7285), .B1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4177), .ZN(n7292) );
  AOI21_X1 U7941 ( .B1(n7287), .B2(n7313), .A(n7286), .ZN(n7291) );
  AOI22_X1 U7942 ( .A1(n7289), .A2(n7314), .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n7288), .ZN(n7290) );
  OAI211_X1 U7943 ( .C1(n7293), .C2(n7292), .A(n7291), .B(n7290), .ZN(U3002)
         );
  NAND2_X1 U7944 ( .A1(n7294), .A2(n7302), .ZN(n7309) );
  AOI22_X1 U7945 ( .A1(n7298), .A2(n7297), .B1(n7296), .B2(n7295), .ZN(n7299)
         );
  AND2_X1 U7946 ( .A1(n7300), .A2(n7299), .ZN(n7308) );
  OAI22_X1 U7947 ( .A1(n7308), .A2(n7302), .B1(n7301), .B2(n7444), .ZN(n7303)
         );
  AOI21_X1 U7948 ( .B1(n7304), .B2(n7314), .A(n7303), .ZN(n7306) );
  NAND2_X1 U7949 ( .A1(n7280), .A2(REIP_REG_17__SCAN_IN), .ZN(n7305) );
  OAI211_X1 U7950 ( .C1(n7307), .C2(n7309), .A(n7306), .B(n7305), .ZN(U3001)
         );
  OAI21_X1 U7951 ( .B1(n7310), .B2(n7309), .A(n7308), .ZN(n7311) );
  AOI22_X1 U7952 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7311), .B1(n7280), .B2(REIP_REG_18__SCAN_IN), .ZN(n7317) );
  AOI22_X1 U7953 ( .A1(n7315), .A2(n7314), .B1(n7313), .B2(n7312), .ZN(n7316)
         );
  OAI211_X1 U7954 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n7318), .A(n7317), .B(n7316), .ZN(U3000) );
  INV_X1 U7955 ( .A(n7319), .ZN(n7346) );
  OAI22_X1 U7956 ( .A1(n7476), .A2(n4779), .B1(n4267), .B2(n7326), .ZN(n7322)
         );
  OAI22_X1 U7957 ( .A1(n7493), .A2(n7320), .B1(n7348), .B2(n5016), .ZN(n7321)
         );
  AOI211_X1 U7958 ( .C1(n7346), .C2(n7323), .A(n7322), .B(n7321), .ZN(n7324)
         );
  OAI221_X1 U7959 ( .B1(n7325), .B2(n7478), .C1(n7325), .C2(n7491), .A(n7324), 
        .ZN(U2827) );
  OAI22_X1 U7960 ( .A1(n7328), .A2(n7327), .B1(n7514), .B2(n7326), .ZN(n7329)
         );
  AOI211_X1 U7961 ( .C1(n7490), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7449), 
        .B(n7329), .ZN(n7339) );
  NAND2_X1 U7962 ( .A1(n7330), .A2(n7346), .ZN(n7337) );
  NOR2_X1 U7963 ( .A1(REIP_REG_4__SCAN_IN), .A2(n7331), .ZN(n7332) );
  AOI22_X1 U7964 ( .A1(n7333), .A2(n7332), .B1(n3617), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n7336) );
  NAND2_X1 U7965 ( .A1(n7412), .A2(n7334), .ZN(n7335) );
  AND3_X1 U7966 ( .A1(n7337), .A2(n7336), .A3(n7335), .ZN(n7338) );
  OAI211_X1 U7967 ( .C1(n7340), .C2(n7491), .A(n7339), .B(n7338), .ZN(U2823)
         );
  INV_X1 U7968 ( .A(n7341), .ZN(n7347) );
  AOI22_X1 U7969 ( .A1(EBX_REG_5__SCAN_IN), .A2(n3617), .B1(n7412), .B2(n7342), 
        .ZN(n7343) );
  OAI211_X1 U7970 ( .C1(n7478), .C2(n7344), .A(n7423), .B(n7343), .ZN(n7345)
         );
  AOI21_X1 U7971 ( .B1(n7347), .B2(n7346), .A(n7345), .ZN(n7352) );
  NOR2_X1 U7972 ( .A1(n7349), .A2(n7348), .ZN(n7367) );
  OAI21_X1 U7973 ( .B1(n7350), .B2(REIP_REG_5__SCAN_IN), .A(n7367), .ZN(n7351)
         );
  OAI211_X1 U7974 ( .C1(n7491), .C2(n7353), .A(n7352), .B(n7351), .ZN(U2822)
         );
  NAND2_X1 U7975 ( .A1(n7354), .A2(n7496), .ZN(n7358) );
  OAI21_X1 U7976 ( .B1(n7478), .B2(n7355), .A(n7423), .ZN(n7356) );
  AOI21_X1 U7977 ( .B1(n3617), .B2(EBX_REG_6__SCAN_IN), .A(n7356), .ZN(n7357)
         );
  OAI211_X1 U7978 ( .C1(n7493), .C2(n7359), .A(n7358), .B(n7357), .ZN(n7360)
         );
  AOI221_X1 U7979 ( .B1(n7367), .B2(REIP_REG_6__SCAN_IN), .C1(n7361), .C2(
        n7365), .A(n7360), .ZN(n7362) );
  OAI21_X1 U7980 ( .B1(n7363), .B2(n7491), .A(n7362), .ZN(U2821) );
  AOI21_X1 U7981 ( .B1(n7365), .B2(n7364), .A(n7375), .ZN(n7366) );
  NAND2_X1 U7982 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n7376) );
  AOI22_X1 U7983 ( .A1(REIP_REG_7__SCAN_IN), .A2(n7367), .B1(n7366), .B2(n7376), .ZN(n7373) );
  AOI22_X1 U7984 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7490), .B1(
        EBX_REG_7__SCAN_IN), .B2(n3617), .ZN(n7368) );
  OAI211_X1 U7985 ( .C1(n7493), .C2(n7369), .A(n7423), .B(n7368), .ZN(n7370)
         );
  AOI21_X1 U7986 ( .B1(n7371), .B2(n7496), .A(n7370), .ZN(n7372) );
  OAI211_X1 U7987 ( .C1(n7374), .C2(n7491), .A(n7373), .B(n7372), .ZN(U2820)
         );
  NOR3_X1 U7988 ( .A1(REIP_REG_8__SCAN_IN), .A2(n7376), .A3(n7375), .ZN(n7380)
         );
  AOI22_X1 U7989 ( .A1(EBX_REG_8__SCAN_IN), .A2(n3617), .B1(n7412), .B2(n7377), 
        .ZN(n7378) );
  OAI211_X1 U7990 ( .C1(n7478), .C2(n4329), .A(n7378), .B(n7423), .ZN(n7379)
         );
  AOI211_X1 U7991 ( .C1(n7390), .C2(REIP_REG_8__SCAN_IN), .A(n7380), .B(n7379), 
        .ZN(n7385) );
  INV_X1 U7992 ( .A(n7381), .ZN(n7382) );
  AOI22_X1 U7993 ( .A1(n7383), .A2(n7496), .B1(n7382), .B2(n7483), .ZN(n7384)
         );
  NAND2_X1 U7994 ( .A1(n7385), .A2(n7384), .ZN(U2819) );
  AOI22_X1 U7995 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n7490), .B1(
        EBX_REG_9__SCAN_IN), .B2(n3617), .ZN(n7386) );
  OAI211_X1 U7996 ( .C1(n7493), .C2(n7387), .A(n7386), .B(n7423), .ZN(n7388)
         );
  AOI211_X1 U7997 ( .C1(REIP_REG_9__SCAN_IN), .C2(n7390), .A(n7389), .B(n7388), 
        .ZN(n7395) );
  INV_X1 U7998 ( .A(n7391), .ZN(n7393) );
  AOI22_X1 U7999 ( .A1(n7393), .A2(n7496), .B1(n7483), .B2(n7392), .ZN(n7394)
         );
  NAND2_X1 U8000 ( .A1(n7395), .A2(n7394), .ZN(U2818) );
  OAI22_X1 U8001 ( .A1(n7397), .A2(n7478), .B1(n7396), .B2(n7476), .ZN(n7398)
         );
  AOI211_X1 U8002 ( .C1(n7399), .C2(n7412), .A(n7449), .B(n7398), .ZN(n7407)
         );
  INV_X1 U8003 ( .A(n7400), .ZN(n7401) );
  AOI22_X1 U8004 ( .A1(n7402), .A2(n7496), .B1(n7401), .B2(n7483), .ZN(n7406)
         );
  NAND2_X1 U8005 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7403), .ZN(n7405) );
  NAND2_X1 U8006 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n7408) );
  OAI211_X1 U8007 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n7410), .B(n7408), .ZN(n7404) );
  NAND4_X1 U8008 ( .A1(n7407), .A2(n7406), .A3(n7405), .A4(n7404), .ZN(U2814)
         );
  NOR2_X1 U8009 ( .A1(REIP_REG_14__SCAN_IN), .A2(n7408), .ZN(n7409) );
  AOI22_X1 U8010 ( .A1(n7412), .A2(n7411), .B1(n7410), .B2(n7409), .ZN(n7422)
         );
  OAI22_X1 U8011 ( .A1(n7415), .A2(n7414), .B1(n7413), .B2(n7476), .ZN(n7416)
         );
  AOI211_X1 U8012 ( .C1(n7490), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7449), 
        .B(n7416), .ZN(n7421) );
  INV_X1 U8013 ( .A(n7417), .ZN(n7418) );
  AOI22_X1 U8014 ( .A1(n7419), .A2(n7496), .B1(n7418), .B2(n7483), .ZN(n7420)
         );
  NAND3_X1 U8015 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(U2813) );
  NAND2_X1 U8016 ( .A1(n3617), .A2(EBX_REG_15__SCAN_IN), .ZN(n7424) );
  OAI211_X1 U8017 ( .C1(n7478), .C2(n7425), .A(n7424), .B(n7423), .ZN(n7427)
         );
  AOI211_X1 U8018 ( .C1(n7428), .C2(REIP_REG_15__SCAN_IN), .A(n7427), .B(n7426), .ZN(n7429) );
  OAI21_X1 U8019 ( .B1(n7430), .B2(n7467), .A(n7429), .ZN(n7431) );
  AOI21_X1 U8020 ( .B1(n7432), .B2(n7483), .A(n7431), .ZN(n7433) );
  OAI21_X1 U8021 ( .B1(n7493), .B2(n7434), .A(n7433), .ZN(U2812) );
  INV_X1 U8022 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7436) );
  OAI22_X1 U8023 ( .A1(n7436), .A2(n7478), .B1(n7435), .B2(n7491), .ZN(n7437)
         );
  AOI211_X1 U8024 ( .C1(n3617), .C2(EBX_REG_17__SCAN_IN), .A(n7449), .B(n7437), 
        .ZN(n7443) );
  NAND2_X1 U8025 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n7440) );
  OAI21_X1 U8026 ( .B1(n7440), .B2(n7439), .A(n7438), .ZN(n7441) );
  AOI22_X1 U8027 ( .A1(n7557), .A2(n7496), .B1(n7441), .B2(n7456), .ZN(n7442)
         );
  OAI211_X1 U8028 ( .C1(n7493), .C2(n7444), .A(n7443), .B(n7442), .ZN(U2810)
         );
  AND3_X1 U8029 ( .A1(n7447), .A2(n7446), .A3(n7445), .ZN(n7455) );
  INV_X1 U8030 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U8031 ( .A1(n3617), .A2(EBX_REG_19__SCAN_IN), .ZN(n7452) );
  INV_X1 U8032 ( .A(n7448), .ZN(n7450) );
  AOI21_X1 U8033 ( .B1(n7483), .B2(n7450), .A(n7449), .ZN(n7451) );
  OAI211_X1 U8034 ( .C1(n7453), .C2(n7478), .A(n7452), .B(n7451), .ZN(n7454)
         );
  AOI211_X1 U8035 ( .C1(n7563), .C2(n7496), .A(n7455), .B(n7454), .ZN(n7459)
         );
  OAI21_X1 U8036 ( .B1(n7457), .B2(n7456), .A(REIP_REG_19__SCAN_IN), .ZN(n7458) );
  OAI211_X1 U8037 ( .C1(n7460), .C2(n7493), .A(n7459), .B(n7458), .ZN(U2808)
         );
  NOR2_X1 U8038 ( .A1(n7473), .A2(REIP_REG_21__SCAN_IN), .ZN(n7474) );
  AOI22_X1 U8039 ( .A1(EBX_REG_21__SCAN_IN), .A2(n3617), .B1(n7461), .B2(n7474), .ZN(n7462) );
  OAI21_X1 U8040 ( .B1(n7464), .B2(n7463), .A(n7462), .ZN(n7469) );
  INV_X1 U8041 ( .A(n7465), .ZN(n7466) );
  OAI22_X1 U8042 ( .A1(n7571), .A2(n7467), .B1(n7493), .B2(n7466), .ZN(n7468)
         );
  AOI211_X1 U8043 ( .C1(PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n7490), .A(n7469), 
        .B(n7468), .ZN(n7470) );
  OAI21_X1 U8044 ( .B1(n7471), .B2(n7491), .A(n7470), .ZN(U2806) );
  NOR2_X1 U8045 ( .A1(n7473), .A2(n7472), .ZN(n7488) );
  OR2_X1 U8046 ( .A1(n7475), .A2(n7474), .ZN(n7481) );
  OAI22_X1 U8047 ( .A1(n7479), .A2(n7478), .B1(n7477), .B2(n7476), .ZN(n7480)
         );
  AOI221_X1 U8048 ( .B1(n7488), .B2(n7482), .C1(n7481), .C2(
        REIP_REG_22__SCAN_IN), .A(n7480), .ZN(n7486) );
  AOI22_X1 U8049 ( .A1(n7575), .A2(n7496), .B1(n7484), .B2(n7483), .ZN(n7485)
         );
  OAI211_X1 U8050 ( .C1(n7487), .C2(n7493), .A(n7486), .B(n7485), .ZN(U2805)
         );
  AOI21_X1 U8051 ( .B1(REIP_REG_22__SCAN_IN), .B2(n7488), .A(
        REIP_REG_23__SCAN_IN), .ZN(n7500) );
  AOI22_X1 U8052 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n7490), .B1(
        EBX_REG_23__SCAN_IN), .B2(n3617), .ZN(n7498) );
  OAI22_X1 U8053 ( .A1(n7494), .A2(n7493), .B1(n7492), .B2(n7491), .ZN(n7495)
         );
  AOI21_X1 U8054 ( .B1(n7580), .B2(n7496), .A(n7495), .ZN(n7497) );
  OAI211_X1 U8055 ( .C1(n7500), .C2(n7499), .A(n7498), .B(n7497), .ZN(U2804)
         );
  OAI21_X1 U8056 ( .B1(n7503), .B2(n7502), .A(n7501), .ZN(U2793) );
  INV_X1 U8057 ( .A(n7504), .ZN(n7508) );
  INV_X1 U8058 ( .A(n7505), .ZN(n7506) );
  OAI211_X1 U8059 ( .C1(n7508), .C2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n7507), .B(n7506), .ZN(n7509) );
  OAI21_X1 U8060 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7513) );
  MUX2_X1 U8061 ( .A(n7513), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n7512), 
        .Z(U3456) );
  INV_X1 U8062 ( .A(n4904), .ZN(n7516) );
  INV_X1 U8063 ( .A(n7514), .ZN(n7515) );
  NAND4_X1 U8064 ( .A1(n7518), .A2(n7517), .A3(n7516), .A4(n7515), .ZN(n7519)
         );
  OAI21_X1 U8065 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(U3455) );
  INV_X1 U8066 ( .A(n7532), .ZN(n7530) );
  AOI21_X1 U8067 ( .B1(n7523), .B2(n7546), .A(n7522), .ZN(n7529) );
  AOI21_X1 U8068 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7525), .A(n7524), .ZN(
        n7528) );
  NAND2_X1 U8069 ( .A1(n7530), .A2(n7526), .ZN(n7527) );
  OAI211_X1 U8070 ( .C1(n7530), .C2(n7529), .A(n7528), .B(n7527), .ZN(U3149)
         );
  OAI221_X1 U8071 ( .B1(n7533), .B2(STATE2_REG_0__SCAN_IN), .C1(n7533), .C2(
        n7532), .A(n7531), .ZN(U3453) );
  INV_X1 U8072 ( .A(n7534), .ZN(n7536) );
  OAI21_X1 U8073 ( .B1(n7538), .B2(n7535), .A(n7536), .ZN(U2792) );
  INV_X1 U8074 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7537) );
  OAI21_X1 U8075 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(U3452) );
  AOI211_X1 U8076 ( .C1(STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n7540), .B(n7539), 
        .ZN(n7543) );
  INV_X1 U8077 ( .A(NA_N), .ZN(n7544) );
  AOI221_X1 U8078 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7544), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7549) );
  AOI21_X1 U8079 ( .B1(n7541), .B2(READY_N), .A(n7549), .ZN(n7542) );
  OAI21_X1 U8080 ( .B1(n7556), .B2(n7543), .A(n7542), .ZN(U3181) );
  AOI21_X1 U8081 ( .B1(n7545), .B2(n7544), .A(STATE_REG_2__SCAN_IN), .ZN(n7552) );
  AOI221_X1 U8082 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7546), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7548) );
  AOI221_X1 U8083 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7548), .C2(HOLD), .A(n7547), .ZN(n7550) );
  OAI22_X1 U8084 ( .A1(n7552), .A2(n7551), .B1(n7550), .B2(n7549), .ZN(U3183)
         );
  INV_X1 U8085 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7554) );
  AOI22_X1 U8086 ( .A1(n7556), .A2(n7555), .B1(n7554), .B2(n7553), .ZN(U3473)
         );
  AOI22_X1 U8087 ( .A1(n7557), .A2(n7579), .B1(n7578), .B2(DATAI_17_), .ZN(
        n7562) );
  OAI22_X1 U8088 ( .A1(n7567), .A2(n7559), .B1(n7558), .B2(n7564), .ZN(n7560)
         );
  INV_X1 U8089 ( .A(n7560), .ZN(n7561) );
  NAND2_X1 U8090 ( .A1(n7562), .A2(n7561), .ZN(U2874) );
  AOI22_X1 U8091 ( .A1(n7563), .A2(n7579), .B1(n7578), .B2(DATAI_19_), .ZN(
        n7570) );
  OAI22_X1 U8092 ( .A1(n7567), .A2(n7566), .B1(n7565), .B2(n7564), .ZN(n7568)
         );
  INV_X1 U8093 ( .A(n7568), .ZN(n7569) );
  NAND2_X1 U8094 ( .A1(n7570), .A2(n7569), .ZN(U2872) );
  INV_X1 U8095 ( .A(n7571), .ZN(n7572) );
  AOI22_X1 U8096 ( .A1(n7572), .A2(n7579), .B1(n7578), .B2(DATAI_21_), .ZN(
        n7574) );
  AOI22_X1 U8097 ( .A1(n7582), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7581), .ZN(n7573) );
  NAND2_X1 U8098 ( .A1(n7574), .A2(n7573), .ZN(U2870) );
  AOI22_X1 U8099 ( .A1(n7575), .A2(n7579), .B1(n7578), .B2(DATAI_22_), .ZN(
        n7577) );
  AOI22_X1 U8100 ( .A1(n7582), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7581), .ZN(n7576) );
  NAND2_X1 U8101 ( .A1(n7577), .A2(n7576), .ZN(U2869) );
  AOI22_X1 U8102 ( .A1(n7580), .A2(n7579), .B1(n7578), .B2(DATAI_23_), .ZN(
        n7584) );
  AOI22_X1 U8103 ( .A1(n7582), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n7581), .ZN(n7583) );
  NAND2_X1 U8104 ( .A1(n7584), .A2(n7583), .ZN(U2868) );
  INV_X1 U8105 ( .A(n7585), .ZN(n7586) );
  OAI21_X1 U8106 ( .B1(n7588), .B2(n7587), .A(n7586), .ZN(n7601) );
  OR2_X1 U8107 ( .A1(n7590), .A2(n7589), .ZN(n7594) );
  NOR2_X1 U8108 ( .A1(n7592), .A2(n7591), .ZN(n7646) );
  INV_X1 U8109 ( .A(n7646), .ZN(n7593) );
  INV_X1 U8110 ( .A(n7600), .ZN(n7595) );
  AOI22_X1 U8111 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7598), .B1(n7601), .B2(
        n7595), .ZN(n7656) );
  AOI22_X1 U8112 ( .A1(n7652), .A2(n7597), .B1(n7596), .B2(n7646), .ZN(n7608)
         );
  OR2_X1 U8113 ( .A1(n7599), .A2(n7598), .ZN(n7605) );
  NAND2_X1 U8114 ( .A1(n7601), .A2(n7600), .ZN(n7603) );
  AND2_X1 U8115 ( .A1(n7603), .A2(n7602), .ZN(n7604) );
  NAND2_X1 U8116 ( .A1(n7605), .A2(n7604), .ZN(n7650) );
  AOI22_X1 U8117 ( .A1(n7649), .A2(n7606), .B1(INSTQUEUE_REG_7__0__SCAN_IN), 
        .B2(n7650), .ZN(n7607) );
  OAI211_X1 U8118 ( .C1(n7656), .C2(n7609), .A(n7608), .B(n7607), .ZN(U3076)
         );
  AOI22_X1 U8119 ( .A1(n7649), .A2(n7611), .B1(n7610), .B2(n7646), .ZN(n7614)
         );
  AOI22_X1 U8120 ( .A1(n7652), .A2(n7612), .B1(INSTQUEUE_REG_7__1__SCAN_IN), 
        .B2(n7650), .ZN(n7613) );
  OAI211_X1 U8121 ( .C1(n7656), .C2(n7615), .A(n7614), .B(n7613), .ZN(U3077)
         );
  AOI22_X1 U8122 ( .A1(n7649), .A2(n7617), .B1(n7616), .B2(n7646), .ZN(n7620)
         );
  AOI22_X1 U8123 ( .A1(n7652), .A2(n7618), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n7650), .ZN(n7619) );
  OAI211_X1 U8124 ( .C1(n7656), .C2(n7621), .A(n7620), .B(n7619), .ZN(U3078)
         );
  AOI22_X1 U8125 ( .A1(n7652), .A2(n7623), .B1(n7622), .B2(n7646), .ZN(n7626)
         );
  AOI22_X1 U8126 ( .A1(n7649), .A2(n7624), .B1(INSTQUEUE_REG_7__3__SCAN_IN), 
        .B2(n7650), .ZN(n7625) );
  OAI211_X1 U8127 ( .C1(n7656), .C2(n7627), .A(n7626), .B(n7625), .ZN(U3079)
         );
  AOI22_X1 U8128 ( .A1(n7649), .A2(n7629), .B1(n7628), .B2(n7646), .ZN(n7632)
         );
  AOI22_X1 U8129 ( .A1(n7652), .A2(n7630), .B1(INSTQUEUE_REG_7__4__SCAN_IN), 
        .B2(n7650), .ZN(n7631) );
  OAI211_X1 U8130 ( .C1(n7656), .C2(n7633), .A(n7632), .B(n7631), .ZN(U3080)
         );
  AOI22_X1 U8131 ( .A1(n7649), .A2(n7635), .B1(n7634), .B2(n7646), .ZN(n7638)
         );
  AOI22_X1 U8132 ( .A1(n7652), .A2(n7636), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n7650), .ZN(n7637) );
  OAI211_X1 U8133 ( .C1(n7656), .C2(n7639), .A(n7638), .B(n7637), .ZN(U3081)
         );
  AOI22_X1 U8134 ( .A1(n7649), .A2(n7641), .B1(n7640), .B2(n7646), .ZN(n7644)
         );
  AOI22_X1 U8135 ( .A1(n7652), .A2(n7642), .B1(INSTQUEUE_REG_7__6__SCAN_IN), 
        .B2(n7650), .ZN(n7643) );
  OAI211_X1 U8136 ( .C1(n7656), .C2(n7645), .A(n7644), .B(n7643), .ZN(U3082)
         );
  AOI22_X1 U8137 ( .A1(n7649), .A2(n7648), .B1(n7647), .B2(n7646), .ZN(n7654)
         );
  AOI22_X1 U8138 ( .A1(n7652), .A2(n7651), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n7650), .ZN(n7653) );
  OAI211_X1 U8139 ( .C1(n7656), .C2(n7655), .A(n7654), .B(n7653), .ZN(U3083)
         );
  AND2_X2 U4330 ( .A1(n3751), .A2(n4939), .ZN(n4420) );
  INV_X1 U4460 ( .A(n3926), .ZN(n5069) );
  CLKBUF_X2 U3653 ( .A(n4420), .Z(n4701) );
  CLKBUF_X1 U3669 ( .A(n6140), .Z(n6141) );
  CLKBUF_X1 U6942 ( .A(n5860), .Z(n5932) );
endmodule

