

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2956, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621;

  OR2_X1 U3404 ( .A1(n4273), .A2(n3010), .ZN(n4211) );
  AND2_X1 U3405 ( .A1(n5159), .A2(n3650), .ZN(n4228) );
  NAND2_X1 U3406 ( .A1(n3605), .A2(n3604), .ZN(n4681) );
  NAND2_X4 U3408 ( .A1(n3433), .A2(n3432), .ZN(n3439) );
  INV_X1 U3409 ( .A(n4167), .ZN(n4156) );
  BUF_X1 U3410 ( .A(n3577), .Z(n2964) );
  NAND2_X1 U3411 ( .A1(n3346), .A2(n3345), .ZN(n3347) );
  CLKBUF_X2 U3412 ( .A(n3571), .Z(n2962) );
  XNOR2_X1 U3413 ( .A(n3242), .B(n3297), .ZN(n3702) );
  CLKBUF_X2 U3414 ( .A(n3207), .Z(n4036) );
  NAND2_X1 U3415 ( .A1(n3536), .A2(n4491), .ZN(n5664) );
  CLKBUF_X2 U3416 ( .A(n3131), .Z(n4098) );
  NOR2_X1 U3417 ( .A1(n3226), .A2(n3227), .ZN(n3536) );
  BUF_X2 U3418 ( .A(n3331), .Z(n4097) );
  CLKBUF_X2 U3419 ( .A(n3132), .Z(n4105) );
  CLKBUF_X2 U3420 ( .A(n3123), .Z(n3276) );
  CLKBUF_X2 U3421 ( .A(n3121), .Z(n4094) );
  CLKBUF_X2 U3422 ( .A(n3171), .Z(n4103) );
  BUF_X2 U3423 ( .A(n3324), .Z(n4018) );
  BUF_X2 U3424 ( .A(n3172), .Z(n4095) );
  CLKBUF_X2 U3425 ( .A(n3124), .Z(n4106) );
  CLKBUF_X2 U3426 ( .A(n3129), .Z(n4104) );
  BUF_X2 U3427 ( .A(n3326), .Z(n3282) );
  INV_X1 U3428 ( .A(n3148), .ZN(n4500) );
  AND4_X1 U3429 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3116)
         );
  AND4_X1 U3430 ( .A1(n3031), .A2(n3030), .A3(n3029), .A4(n3028), .ZN(n3032)
         );
  AND2_X2 U3431 ( .A1(n5089), .A2(n4394), .ZN(n3324) );
  AND2_X2 U3432 ( .A1(n3027), .A2(n4389), .ZN(n3122) );
  AND2_X2 U3433 ( .A1(n5089), .A2(n4390), .ZN(n3207) );
  AND2_X2 U3434 ( .A1(n5087), .A2(n4391), .ZN(n3326) );
  AND2_X2 U3435 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4391) );
  CLKBUF_X1 U3436 ( .A(n5799), .Z(n2956) );
  NOR2_X1 U3437 ( .A1(n4267), .A2(n4178), .ZN(n5799) );
  INV_X1 U3439 ( .A(n6621), .ZN(n2958) );
  AOI22_X1 U3440 ( .A1(n6536), .A2(keyinput16), .B1(keyinput3), .B2(n6535), 
        .ZN(n6534) );
  OAI221_X1 U3441 ( .B1(n6536), .B2(keyinput16), .C1(n6535), .C2(keyinput3), 
        .A(n6534), .ZN(n6537) );
  XNOR2_X1 U3442 ( .A(n3347), .B(n6102), .ZN(n6016) );
  AND4_X1 U3443 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3115)
         );
  NAND2_X1 U3444 ( .A1(n3148), .A2(n3117), .ZN(n3571) );
  INV_X1 U34450 ( .A(n2963), .ZN(n3580) );
  INV_X1 U34460 ( .A(n3155), .ZN(n4296) );
  CLKBUF_X3 U34470 ( .A(n3439), .Z(n2965) );
  INV_X1 U34480 ( .A(n4530), .ZN(n3605) );
  CLKBUF_X2 U3449 ( .A(n3122), .Z(n4396) );
  INV_X1 U3450 ( .A(n5804), .ZN(n5790) );
  INV_X1 U34510 ( .A(n4314), .ZN(n6030) );
  INV_X1 U34520 ( .A(n5770), .ZN(n5780) );
  OR2_X1 U34530 ( .A1(n5861), .A2(n4466), .ZN(n5858) );
  XNOR2_X1 U3454 ( .A(n5122), .B(n5121), .ZN(n5341) );
  AND2_X2 U34550 ( .A1(n3027), .A2(n4389), .ZN(n2959) );
  NOR2_X2 U3457 ( .A1(n3141), .A2(n3532), .ZN(n3225) );
  NAND2_X2 U3458 ( .A1(n3467), .A2(n3466), .ZN(n4222) );
  NAND2_X2 U34590 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  NAND2_X2 U34600 ( .A1(n3460), .A2(n3459), .ZN(n5311) );
  NAND2_X2 U34610 ( .A1(n2972), .A2(n2968), .ZN(n3653) );
  AND4_X2 U34620 ( .A1(n3049), .A2(n3048), .A3(n3047), .A4(n3046), .ZN(n3055)
         );
  AND4_X2 U34630 ( .A1(n3053), .A2(n3052), .A3(n3051), .A4(n3050), .ZN(n3054)
         );
  NOR2_X2 U34640 ( .A1(n3158), .A2(n4510), .ZN(n3526) );
  NAND2_X2 U3466 ( .A1(n3306), .A2(n3305), .ZN(n3349) );
  NOR2_X2 U3467 ( .A1(n4208), .A2(n5379), .ZN(n5290) );
  NAND2_X1 U34680 ( .A1(n3169), .A2(n3168), .ZN(n3238) );
  AND2_X1 U34690 ( .A1(n3152), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3267) );
  OR2_X1 U34700 ( .A1(n2969), .A2(n4491), .ZN(n3163) );
  NAND2_X1 U34710 ( .A1(n3710), .A2(n3056), .ZN(n3147) );
  CLKBUF_X2 U34730 ( .A(n3146), .Z(n4505) );
  INV_X1 U34740 ( .A(n3710), .ZN(n2960) );
  NAND4_X1 U3475 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3117)
         );
  INV_X2 U3476 ( .A(n4946), .ZN(n2961) );
  AOI22_X1 U3477 ( .A1(n3324), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3050) );
  CLKBUF_X2 U3478 ( .A(n3130), .Z(n4096) );
  AND2_X1 U3479 ( .A1(n4218), .A2(n4217), .ZN(n2998) );
  AND2_X1 U3480 ( .A1(n5290), .A2(n2970), .ZN(n4273) );
  OR2_X1 U3481 ( .A1(n4215), .A2(n4314), .ZN(n4216) );
  AND2_X1 U3482 ( .A1(n5312), .A2(n3463), .ZN(n5417) );
  AND2_X1 U3483 ( .A1(n5217), .A2(n5216), .ZN(n5594) );
  CLKBUF_X1 U3484 ( .A(n5281), .Z(n5392) );
  NAND2_X1 U3485 ( .A1(n3458), .A2(n4219), .ZN(n3459) );
  NAND2_X1 U3486 ( .A1(n3005), .A2(n3004), .ZN(n5320) );
  NAND2_X1 U3487 ( .A1(n3691), .A2(n3690), .ZN(n4529) );
  XNOR2_X1 U3488 ( .A(n3433), .B(n3423), .ZN(n3684) );
  AND2_X1 U3489 ( .A1(n3315), .A2(n3314), .ZN(n6017) );
  NAND2_X1 U3490 ( .A1(n3339), .A2(n3338), .ZN(n4449) );
  NAND2_X1 U3491 ( .A1(n4381), .A2(n6530), .ZN(n3339) );
  NAND2_X1 U3492 ( .A1(n3206), .A2(n3205), .ZN(n3294) );
  CLKBUF_X1 U3493 ( .A(n4381), .Z(n5812) );
  NAND2_X1 U3494 ( .A1(n3250), .A2(n3197), .ZN(n3254) );
  XNOR2_X1 U3495 ( .A(n3316), .B(n6167), .ZN(n4381) );
  NAND2_X1 U3496 ( .A1(n3204), .A2(n3251), .ZN(n3206) );
  NAND2_X1 U3497 ( .A1(n3266), .A2(n3265), .ZN(n3275) );
  CLKBUF_X1 U3498 ( .A(n3711), .Z(n3712) );
  NAND2_X1 U3499 ( .A1(n3322), .A2(n3321), .ZN(n6167) );
  INV_X1 U3500 ( .A(n3238), .ZN(n3264) );
  NAND2_X1 U3501 ( .A1(n3273), .A2(n3272), .ZN(n3274) );
  OR2_X1 U3502 ( .A1(n3317), .A2(n4415), .ZN(n3322) );
  OR2_X1 U3503 ( .A1(n3317), .A2(n5106), .ZN(n3273) );
  NAND2_X1 U3504 ( .A1(n3154), .A2(n3153), .ZN(n3169) );
  CLKBUF_X1 U3505 ( .A(n3536), .Z(n4286) );
  NAND2_X1 U3506 ( .A1(n3203), .A2(n3202), .ZN(n3251) );
  NOR2_X1 U3507 ( .A1(n3198), .A2(n6530), .ZN(n3431) );
  AND2_X1 U3508 ( .A1(n3147), .A2(n4505), .ZN(n3118) );
  OR2_X1 U3509 ( .A1(n3194), .A2(n3193), .ZN(n3255) );
  OR2_X1 U3510 ( .A1(n3182), .A2(n3181), .ZN(n3436) );
  INV_X1 U3511 ( .A(n3653), .ZN(n4495) );
  INV_X2 U3512 ( .A(n3117), .ZN(n4491) );
  AND2_X2 U3513 ( .A1(n3033), .A2(n3032), .ZN(n3532) );
  CLKBUF_X2 U3514 ( .A(n3120), .Z(n3200) );
  AND4_X1 U3515 ( .A1(n3026), .A2(n3025), .A3(n3024), .A4(n3023), .ZN(n3033)
         );
  NAND3_X1 U3516 ( .A1(n3066), .A2(n3061), .A3(n3065), .ZN(n3120) );
  AND4_X1 U3517 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3104)
         );
  AND4_X1 U3518 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3042)
         );
  AND4_X1 U3519 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3083)
         );
  AND4_X1 U3520 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3084)
         );
  AND4_X1 U3521 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3105)
         );
  AND4_X1 U3522 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3085)
         );
  AND2_X1 U3523 ( .A1(n3045), .A2(n3044), .ZN(n3049) );
  AND2_X1 U3524 ( .A1(n3020), .A2(n3019), .ZN(n3026) );
  AND4_X1 U3525 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3043)
         );
  AND3_X1 U3526 ( .A1(n3064), .A2(n3063), .A3(n3062), .ZN(n3065) );
  AND4_X1 U3527 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .ZN(n3086)
         );
  AND4_X1 U3528 ( .A1(n3060), .A2(n3059), .A3(n3058), .A4(n3057), .ZN(n3066)
         );
  AND4_X1 U3529 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3103)
         );
  OR2_X2 U3530 ( .A1(n6355), .A2(n6238), .ZN(n4314) );
  NAND2_X1 U3531 ( .A1(n3532), .A2(n3685), .ZN(n3710) );
  AND2_X4 U3532 ( .A1(n3021), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3027)
         );
  OAI22_X2 U3533 ( .A1(n5116), .A2(n3580), .B1(n5208), .B2(n5220), .ZN(n5213)
         );
  OR2_X2 U3534 ( .A1(n5220), .A2(n5209), .ZN(n5116) );
  NAND2_X2 U3535 ( .A1(n3254), .A2(n3253), .ZN(n3709) );
  AOI21_X2 U3536 ( .B1(n4446), .B2(n3533), .A(n3310), .ZN(n6027) );
  BUF_X4 U3537 ( .A(n3571), .Z(n2963) );
  NAND2_X2 U3538 ( .A1(n5175), .A2(n5176), .ZN(n5256) );
  NOR2_X4 U3539 ( .A1(n5075), .A2(n5179), .ZN(n5175) );
  NOR2_X2 U3540 ( .A1(n4681), .A2(n4682), .ZN(n4896) );
  AND2_X2 U3541 ( .A1(n4871), .A2(n2992), .ZN(n4958) );
  NOR2_X4 U3542 ( .A1(n4608), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U3543 ( .A1(n4500), .A2(n4946), .ZN(n3577) );
  AND2_X2 U3544 ( .A1(n5251), .A2(n2991), .ZN(n4190) );
  NOR2_X4 U3545 ( .A1(n5256), .A2(n5255), .ZN(n5251) );
  XNOR2_X2 U3546 ( .A(n4262), .B(n4261), .ZN(n4215) );
  NAND2_X1 U3547 ( .A1(n2984), .A2(n2983), .ZN(n4608) );
  NOR2_X1 U3548 ( .A1(n4370), .A2(n2974), .ZN(n2983) );
  INV_X1 U3549 ( .A(n4610), .ZN(n2986) );
  NAND2_X1 U3550 ( .A1(n5520), .A2(n3004), .ZN(n3003) );
  INV_X1 U3551 ( .A(n3156), .ZN(n2996) );
  INV_X1 U3552 ( .A(n2978), .ZN(n3457) );
  AND2_X1 U3553 ( .A1(n5522), .A2(n5323), .ZN(n3004) );
  NAND2_X1 U3554 ( .A1(n3396), .A2(n3395), .ZN(n3418) );
  AND2_X1 U3555 ( .A1(n4946), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3490) );
  INV_X1 U3556 ( .A(n3504), .ZN(n3513) );
  AOI22_X1 U3557 ( .A1(n3207), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3030) );
  AOI22_X1 U3558 ( .A1(n3172), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3129), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3029) );
  AOI22_X1 U3559 ( .A1(n3121), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3025) );
  OR2_X1 U3560 ( .A1(n4123), .A2(n3323), .ZN(n3503) );
  NAND2_X1 U3561 ( .A1(n5108), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4124) );
  INV_X1 U3562 ( .A(n3510), .ZN(n3533) );
  NAND2_X1 U3563 ( .A1(n4131), .A2(n3560), .ZN(n3510) );
  NAND2_X1 U3564 ( .A1(n3490), .A2(n3200), .ZN(n3504) );
  AND2_X1 U3565 ( .A1(n4430), .A2(n4429), .ZN(n6324) );
  INV_X1 U3566 ( .A(n3225), .ZN(n4130) );
  INV_X1 U3567 ( .A(n3838), .ZN(n4263) );
  INV_X1 U3568 ( .A(n4124), .ZN(n4264) );
  INV_X1 U3569 ( .A(n4369), .ZN(n2985) );
  AND2_X1 U3570 ( .A1(n4438), .A2(n6329), .ZN(n4305) );
  AND2_X1 U3571 ( .A1(n2965), .A2(n5465), .ZN(n3456) );
  AOI22_X1 U3572 ( .A1(n3184), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3059) );
  OR2_X1 U3573 ( .A1(n3217), .A2(n3216), .ZN(n3244) );
  INV_X1 U3574 ( .A(n3200), .ZN(n2997) );
  NAND2_X1 U3575 ( .A1(n3184), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3044)
         );
  NAND2_X1 U3576 ( .A1(n3132), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3045) );
  OR2_X1 U3577 ( .A1(n3504), .A2(n3545), .ZN(n3485) );
  OAI22_X1 U3578 ( .A1(n3515), .A2(n3514), .B1(n3513), .B2(n3540), .ZN(n3516)
         );
  AND2_X1 U3579 ( .A1(n4432), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3482)
         );
  AOI21_X1 U3580 ( .B1(n3509), .B2(n3507), .A(n3478), .ZN(n3483) );
  NOR2_X1 U3581 ( .A1(n3551), .A2(n2961), .ZN(n4139) );
  AOI22_X1 U3582 ( .A1(n3184), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3035) );
  OR2_X1 U3583 ( .A1(n4120), .A2(n5532), .ZN(n4137) );
  OR2_X1 U3584 ( .A1(n3288), .A2(n3287), .ZN(n3340) );
  NOR2_X1 U3585 ( .A1(n3439), .A2(n2979), .ZN(n3006) );
  AOI21_X1 U3586 ( .B1(n3457), .B2(n3004), .A(n2980), .ZN(n3002) );
  NAND2_X1 U3587 ( .A1(n3274), .A2(n6530), .ZN(n3009) );
  INV_X1 U3588 ( .A(n4650), .ZN(n4729) );
  INV_X1 U3589 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6309) );
  AOI22_X1 U3590 ( .A1(n3331), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3023) );
  OAI21_X1 U3591 ( .B1(n6453), .B2(n4439), .A(n6338), .ZN(n4478) );
  AND2_X1 U3592 ( .A1(n4406), .A2(n3657), .ZN(n4388) );
  NOR2_X2 U3593 ( .A1(n5790), .A2(n6326), .ZN(n5123) );
  INV_X1 U3594 ( .A(n4532), .ZN(n3598) );
  INV_X1 U3595 ( .A(n4531), .ZN(n3599) );
  AND2_X1 U3596 ( .A1(n3603), .A2(n3602), .ZN(n4471) );
  NAND2_X1 U3597 ( .A1(n3224), .A2(n3223), .ZN(n4382) );
  INV_X1 U3598 ( .A(n4255), .ZN(n4093) );
  NAND2_X1 U3599 ( .A1(n4053), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4120)
         );
  AND2_X1 U3600 ( .A1(n5153), .A2(n5252), .ZN(n2991) );
  NAND2_X1 U3601 ( .A1(n3787), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3811)
         );
  CLKBUF_X1 U3602 ( .A(n4608), .Z(n4609) );
  AOI21_X1 U3603 ( .B1(n4264), .B2(EAX_REG_7__SCAN_IN), .A(n3689), .ZN(n3690)
         );
  AOI211_X1 U3604 ( .C1(n3743), .C2(n3852), .A(n3742), .B(n3741), .ZN(n4370)
         );
  NAND2_X1 U3605 ( .A1(n3698), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3697)
         );
  XNOR2_X1 U3606 ( .A(n3439), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5391)
         );
  NAND2_X1 U3607 ( .A1(n3462), .A2(n3461), .ZN(n5312) );
  INV_X1 U3608 ( .A(n5314), .ZN(n3461) );
  NAND2_X1 U3609 ( .A1(n5640), .A2(n5641), .ZN(n3454) );
  NOR2_X1 U3610 ( .A1(n5059), .A2(n3666), .ZN(n6068) );
  INV_X1 U3611 ( .A(n5056), .ZN(n3666) );
  AND2_X1 U3612 ( .A1(n3556), .A2(n3555), .ZN(n3665) );
  CLKBUF_X1 U3613 ( .A(n4454), .Z(n4455) );
  INV_X1 U3614 ( .A(n6347), .ZN(n6329) );
  OAI21_X1 U3615 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n4193), .A(n4729), 
        .ZN(n6237) );
  NAND2_X1 U3616 ( .A1(n6530), .A2(n4478), .ZN(n4650) );
  AND3_X1 U3617 ( .A1(n6325), .A2(n6324), .A3(n6323), .ZN(n6330) );
  NAND2_X1 U3618 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  OAI21_X1 U3619 ( .B1(n3521), .B2(n3544), .A(n3520), .ZN(n3525) );
  INV_X1 U3620 ( .A(n3544), .ZN(n3522) );
  INV_X2 U3621 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6326) );
  OR2_X1 U3622 ( .A1(n5861), .A2(n4130), .ZN(n5857) );
  CLKBUF_X1 U3623 ( .A(n4132), .Z(n5867) );
  INV_X1 U3624 ( .A(n5857), .ZN(n5864) );
  INV_X1 U3625 ( .A(n5892), .ZN(n6450) );
  NAND2_X1 U3626 ( .A1(n4305), .A2(n4128), .ZN(n5945) );
  NOR2_X1 U3627 ( .A1(n4408), .A2(READY_N), .ZN(n4128) );
  AND2_X1 U3628 ( .A1(n4305), .A2(n6316), .ZN(n6029) );
  INV_X2 U3629 ( .A(n5315), .ZN(n6025) );
  XNOR2_X1 U3630 ( .A(n3470), .B(n4206), .ZN(n4189) );
  AND2_X1 U3631 ( .A1(n5441), .A2(n3678), .ZN(n5414) );
  INV_X1 U3632 ( .A(n6120), .ZN(n6106) );
  INV_X1 U3633 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6490) );
  AND2_X1 U3634 ( .A1(n4943), .A2(n3488), .ZN(n3511) );
  OR2_X1 U3635 ( .A1(n3406), .A2(n3405), .ZN(n3424) );
  OR2_X1 U3636 ( .A1(n3361), .A2(n3360), .ZN(n3386) );
  AND2_X1 U3637 ( .A1(n3535), .A2(n3534), .ZN(n3661) );
  NAND2_X1 U3638 ( .A1(n3118), .A2(n2999), .ZN(n3535) );
  INV_X1 U3639 ( .A(n2996), .ZN(n2999) );
  OR2_X1 U3640 ( .A1(n3337), .A2(n3336), .ZN(n3364) );
  NAND2_X1 U3641 ( .A1(n2990), .A2(n5224), .ZN(n2989) );
  INV_X1 U3642 ( .A(n5229), .ZN(n2990) );
  NOR2_X1 U3643 ( .A1(n3983), .A2(n5569), .ZN(n4000) );
  NAND2_X1 U3644 ( .A1(n4190), .A2(n4192), .ZN(n4191) );
  NAND2_X1 U3645 ( .A1(n2988), .A2(n2976), .ZN(n5075) );
  INV_X1 U3646 ( .A(n5039), .ZN(n2988) );
  INV_X1 U3647 ( .A(n5077), .ZN(n2987) );
  AND2_X1 U3648 ( .A1(n4167), .A2(n2962), .ZN(n3646) );
  NAND2_X1 U3649 ( .A1(n3420), .A2(n3419), .ZN(n3433) );
  INV_X1 U3650 ( .A(n3646), .ZN(n4153) );
  NAND2_X1 U3651 ( .A1(n3152), .A2(n2977), .ZN(n3154) );
  OAI211_X1 U3652 ( .C1(n3504), .C2(n3220), .A(n3219), .B(n3218), .ZN(n3298)
         );
  AND2_X1 U3653 ( .A1(n3222), .A2(n3148), .ZN(n2994) );
  INV_X1 U3654 ( .A(n3267), .ZN(n3317) );
  AND2_X1 U3655 ( .A1(n3485), .A2(n3484), .ZN(n3517) );
  AOI21_X1 U3656 ( .B1(n3521), .B2(n3533), .A(n3545), .ZN(n3518) );
  NAND2_X1 U3657 ( .A1(n3481), .A2(n3480), .ZN(n3544) );
  INV_X1 U3658 ( .A(n3482), .ZN(n3480) );
  NOR2_X1 U3659 ( .A1(n3504), .A2(n3510), .ZN(n3523) );
  AND2_X1 U3660 ( .A1(n4286), .A2(n4141), .ZN(n4282) );
  CLKBUF_X1 U3661 ( .A(n4139), .Z(n4140) );
  INV_X1 U3662 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5712) );
  INV_X1 U3663 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5728) );
  AND2_X1 U3664 ( .A1(n3645), .A2(n3644), .ZN(n5157) );
  NOR2_X2 U3665 ( .A1(n5247), .A2(n5157), .ZN(n5159) );
  CLKBUF_X1 U3666 ( .A(n3243), .Z(n4131) );
  NAND2_X1 U3667 ( .A1(n3708), .A2(n3707), .ZN(n4319) );
  NAND2_X1 U3668 ( .A1(n4319), .A2(n4318), .ZN(n4321) );
  NAND2_X1 U3669 ( .A1(n4140), .A2(n4305), .ZN(n4293) );
  XNOR2_X1 U3670 ( .A(n4138), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4267)
         );
  OR2_X1 U3671 ( .A1(n5540), .A2(n4092), .ZN(n4072) );
  NOR2_X1 U3672 ( .A1(n4016), .A2(n5140), .ZN(n4017) );
  NAND2_X1 U3673 ( .A1(n4017), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4052)
         );
  NOR2_X2 U3674 ( .A1(n4191), .A2(n4243), .ZN(n5136) );
  INV_X1 U3675 ( .A(n5146), .ZN(n4245) );
  NOR2_X1 U3676 ( .A1(n3940), .A2(n5308), .ZN(n3941) );
  AND2_X1 U3677 ( .A1(n3939), .A2(n3938), .ZN(n5252) );
  NOR2_X1 U3678 ( .A1(n3910), .A2(n5171), .ZN(n3911) );
  NAND2_X1 U3679 ( .A1(n3884), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3910)
         );
  NAND2_X1 U3680 ( .A1(n3869), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3883)
         );
  CLKBUF_X1 U3681 ( .A(n5075), .Z(n5076) );
  NAND2_X1 U3682 ( .A1(n3842), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3843)
         );
  NOR2_X1 U3683 ( .A1(n6536), .A2(n3843), .ZN(n3869) );
  CLKBUF_X1 U3684 ( .A(n5039), .Z(n5040) );
  NOR2_X1 U3685 ( .A1(n3839), .A2(n5712), .ZN(n3842) );
  NAND2_X1 U3686 ( .A1(n3814), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3839)
         );
  CLKBUF_X1 U3687 ( .A(n4985), .Z(n4986) );
  NOR2_X1 U3688 ( .A1(n4959), .A2(n2993), .ZN(n2992) );
  INV_X1 U3689 ( .A(n4875), .ZN(n2993) );
  NOR2_X1 U3690 ( .A1(n3811), .A2(n5728), .ZN(n3814) );
  INV_X1 U3691 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U3692 ( .A1(n3759), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3784)
         );
  INV_X1 U3693 ( .A(n3758), .ZN(n3759) );
  NOR2_X1 U3694 ( .A1(n3739), .A2(n3686), .ZN(n3687) );
  INV_X1 U3695 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3686) );
  NAND2_X1 U3696 ( .A1(n3687), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3758)
         );
  NAND2_X1 U3697 ( .A1(n3733), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3739)
         );
  INV_X1 U3698 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5791) );
  NOR2_X1 U3699 ( .A1(n3697), .A2(n5791), .ZN(n3733) );
  AOI21_X1 U3700 ( .B1(n4448), .B2(n3852), .A(n3701), .ZN(n4474) );
  NAND2_X1 U3701 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U3702 ( .A1(n5227), .A2(n5218), .ZN(n5220) );
  AND2_X1 U3703 ( .A1(n5234), .A2(n5225), .ZN(n5227) );
  NOR2_X2 U3704 ( .A1(n5232), .A2(n5231), .ZN(n5234) );
  NAND2_X1 U3705 ( .A1(n4228), .A2(n4227), .ZN(n5131) );
  AND2_X1 U3706 ( .A1(n4237), .A2(n4236), .ZN(n5383) );
  NAND2_X1 U3707 ( .A1(n3003), .A2(n3002), .ZN(n3458) );
  CLKBUF_X1 U3708 ( .A(n5320), .Z(n5321) );
  XNOR2_X1 U3709 ( .A(n2965), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5641)
         );
  CLKBUF_X1 U3710 ( .A(n5962), .Z(n5963) );
  INV_X1 U3711 ( .A(n4374), .ZN(n3590) );
  INV_X1 U3712 ( .A(n5808), .ZN(n3591) );
  OR2_X1 U3713 ( .A1(n3665), .A2(n4414), .ZN(n4888) );
  NAND2_X1 U3714 ( .A1(n4949), .A2(n4167), .ZN(n4328) );
  NAND2_X1 U3715 ( .A1(n2964), .A2(n2962), .ZN(n5120) );
  OAI211_X1 U3716 ( .C1(n3275), .C2(n3009), .A(n3007), .B(n3289), .ZN(n3293)
         );
  INV_X1 U3717 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6296) );
  INV_X1 U3718 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3018) );
  CLKBUF_X1 U3719 ( .A(n3526), .Z(n3527) );
  CLKBUF_X1 U3720 ( .A(n4389), .Z(n5096) );
  INV_X1 U3721 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4415) );
  NAND3_X1 U3722 ( .A1(n3225), .A2(n2961), .A3(n4500), .ZN(n3227) );
  AND2_X1 U3723 ( .A1(n4905), .A2(n4612), .ZN(n4615) );
  AND2_X1 U3724 ( .A1(n5481), .A2(n4901), .ZN(n6134) );
  AND2_X1 U3725 ( .A1(n4479), .A2(n4455), .ZN(n6169) );
  AND2_X1 U3726 ( .A1(n4446), .A2(n4450), .ZN(n4999) );
  NOR2_X1 U3727 ( .A1(n6235), .A2(n4447), .ZN(n4541) );
  AND2_X1 U3728 ( .A1(n6131), .A2(n4448), .ZN(n4781) );
  NOR2_X1 U3729 ( .A1(n4416), .A2(n4455), .ZN(n4763) );
  BUF_X1 U3730 ( .A(n3532), .Z(n4515) );
  NOR2_X1 U3731 ( .A1(n4481), .A2(n4447), .ZN(n4685) );
  INV_X1 U3732 ( .A(n3709), .ZN(n4906) );
  NOR2_X1 U3733 ( .A1(n4481), .A2(n4903), .ZN(n4487) );
  INV_X1 U3734 ( .A(n6238), .ZN(n6233) );
  INV_X1 U3735 ( .A(n6237), .ZN(n6175) );
  NAND2_X1 U3736 ( .A1(n4293), .A2(n5527), .ZN(n6448) );
  INV_X1 U3737 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5190) );
  NOR2_X1 U3738 ( .A1(n5693), .A2(n5198), .ZN(n5189) );
  INV_X1 U3739 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6536) );
  AND2_X1 U3740 ( .A1(n4267), .A2(n4177), .ZN(n5770) );
  INV_X1 U3741 ( .A(n5820), .ZN(n5834) );
  NAND2_X2 U3742 ( .A1(n4169), .A2(n4168), .ZN(n5817) );
  AND2_X1 U3743 ( .A1(n4184), .A2(n5123), .ZN(n5821) );
  INV_X1 U3744 ( .A(n5799), .ZN(n5835) );
  NAND2_X1 U3745 ( .A1(n4167), .A2(n4166), .ZN(n5824) );
  INV_X1 U3746 ( .A(n5824), .ZN(n5831) );
  AND2_X1 U3747 ( .A1(n5852), .A2(n5108), .ZN(n5849) );
  OR2_X1 U3748 ( .A1(n4327), .A2(n4326), .ZN(n5852) );
  INV_X1 U3749 ( .A(n3685), .ZN(n5108) );
  INV_X1 U3750 ( .A(n5858), .ZN(n5865) );
  INV_X1 U3751 ( .A(n5861), .ZN(n5109) );
  INV_X2 U3752 ( .A(n5888), .ZN(n5895) );
  INV_X1 U3753 ( .A(n5890), .ZN(n5897) );
  NAND2_X1 U3754 ( .A1(n4305), .A2(n4292), .ZN(n5951) );
  INV_X1 U3755 ( .A(n6334), .ZN(n4292) );
  INV_X1 U3756 ( .A(n5945), .ZN(n5949) );
  OR2_X1 U3757 ( .A1(n6029), .A2(n4195), .ZN(n5315) );
  NOR2_X1 U3758 ( .A1(n4370), .A2(n4469), .ZN(n2982) );
  AND2_X1 U3759 ( .A1(n5315), .A2(n4310), .ZN(n6012) );
  INV_X1 U3760 ( .A(n6029), .ZN(n5675) );
  XNOR2_X1 U3761 ( .A(n3000), .B(n5088), .ZN(n5331) );
  NAND2_X1 U3762 ( .A1(n3001), .A2(n2971), .ZN(n3000) );
  NAND2_X1 U3763 ( .A1(n5290), .A2(n2981), .ZN(n3001) );
  AOI21_X1 U3764 ( .B1(n4252), .B2(n5279), .A(n2973), .ZN(n4253) );
  AND2_X1 U3765 ( .A1(n5414), .A2(n4232), .ZN(n5332) );
  AND2_X1 U3767 ( .A1(n3672), .A2(n3671), .ZN(n5412) );
  CLKBUF_X1 U3768 ( .A(n5449), .Z(n5450) );
  CLKBUF_X1 U3769 ( .A(n5520), .Z(n5521) );
  CLKBUF_X1 U3770 ( .A(n5048), .Z(n5049) );
  CLKBUF_X1 U3771 ( .A(n4963), .Z(n4964) );
  OR2_X1 U3772 ( .A1(n5429), .A2(n4972), .ZN(n6037) );
  CLKBUF_X1 U3773 ( .A(n4880), .Z(n4881) );
  OR2_X1 U3774 ( .A1(n4194), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6071) );
  CLKBUF_X1 U3775 ( .A(n5988), .Z(n5989) );
  CLKBUF_X1 U3776 ( .A(n6007), .Z(n6008) );
  INV_X1 U3777 ( .A(n6070), .ZN(n6122) );
  OR2_X1 U3778 ( .A1(n3665), .A2(n3568), .ZN(n6120) );
  NOR2_X1 U3779 ( .A1(n3665), .A2(n5092), .ZN(n5059) );
  INV_X1 U3780 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4997) );
  NOR2_X1 U3781 ( .A1(n4903), .A2(n4534), .ZN(n6232) );
  INV_X1 U3782 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U3783 ( .B1(n4440), .B2(n6428), .A(n4650), .ZN(n6130) );
  INV_X1 U3784 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6513) );
  INV_X1 U3785 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3017) );
  NOR2_X1 U3786 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5665) );
  NAND2_X1 U3787 ( .A1(n4615), .A2(n3709), .ZN(n4757) );
  INV_X1 U3788 ( .A(n6164), .ZN(n6152) );
  OAI21_X1 U3789 ( .B1(n6139), .B2(n6136), .A(n6135), .ZN(n6161) );
  OR2_X1 U3790 ( .A1(n5484), .A2(n3709), .ZN(n6164) );
  INV_X1 U3791 ( .A(n5485), .ZN(n5514) );
  AND2_X1 U3792 ( .A1(n4999), .A2(n4998), .ZN(n6204) );
  INV_X1 U3793 ( .A(n4811), .ZN(n4565) );
  NAND2_X1 U3794 ( .A1(n4541), .A2(n4906), .ZN(n4811) );
  NAND2_X1 U3795 ( .A1(n4781), .A2(n4998), .ZN(n6294) );
  INV_X1 U3796 ( .A(n6278), .ZN(n6286) );
  INV_X1 U3797 ( .A(n6244), .ZN(n6181) );
  INV_X1 U3798 ( .A(n6250), .ZN(n6185) );
  INV_X1 U3799 ( .A(n6262), .ZN(n6193) );
  INV_X1 U3800 ( .A(n6268), .ZN(n6196) );
  INV_X1 U3801 ( .A(n6275), .ZN(n6199) );
  INV_X1 U3802 ( .A(n6282), .ZN(n6203) );
  NOR2_X1 U3803 ( .A1(n5923), .A2(n4650), .ZN(n6250) );
  NOR2_X1 U3804 ( .A1(n5925), .A2(n4650), .ZN(n6256) );
  NOR2_X1 U3805 ( .A1(n4477), .A2(n4650), .ZN(n6262) );
  NOR2_X1 U3806 ( .A1(n4298), .A2(n4650), .ZN(n6275) );
  NOR2_X1 U3807 ( .A1(n5931), .A2(n4650), .ZN(n6282) );
  NAND2_X1 U3808 ( .A1(n4487), .A2(n3709), .ZN(n4715) );
  NAND2_X1 U3809 ( .A1(n4487), .A2(n4906), .ZN(n4756) );
  AND2_X1 U3810 ( .A1(n6336), .A2(n6335), .ZN(n6345) );
  CLKBUF_X1 U3811 ( .A(n6447), .Z(n6418) );
  INV_X1 U3812 ( .A(n6416), .ZN(n6419) );
  NOR2_X1 U3813 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6363), .ZN(n6458) );
  AND2_X1 U3814 ( .A1(n4134), .A2(n4133), .ZN(n4135) );
  OAI21_X1 U3815 ( .B1(n5276), .B2(n4314), .A(n4248), .ZN(n4249) );
  INV_X1 U3816 ( .A(n4202), .ZN(n4203) );
  OAI21_X1 U3817 ( .B1(n5578), .B2(n4314), .A(n4201), .ZN(n4202) );
  AND2_X1 U3818 ( .A1(n3680), .A2(n3679), .ZN(n3681) );
  NAND2_X1 U3819 ( .A1(n4189), .A2(n6126), .ZN(n3682) );
  OR2_X1 U3820 ( .A1(n5135), .A2(n2989), .ZN(n2967) );
  OAI22_X1 U3821 ( .A1(n5311), .A2(n3006), .B1(n4205), .B2(n4219), .ZN(n5281)
         );
  AND4_X1 U3822 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n2968)
         );
  AND4_X1 U3823 ( .A1(n2995), .A2(n3149), .A3(n3147), .A4(n3148), .ZN(n2969)
         );
  INV_X1 U3824 ( .A(n4446), .ZN(n6131) );
  NAND2_X1 U3825 ( .A1(n4871), .A2(n4875), .ZN(n4874) );
  AND2_X1 U3826 ( .A1(n5363), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n2970)
         );
  NAND2_X1 U3827 ( .A1(n5281), .A2(n5391), .ZN(n4271) );
  INV_X1 U3828 ( .A(n3120), .ZN(n3146) );
  AND2_X1 U3829 ( .A1(n3005), .A2(n5522), .ZN(n5322) );
  NOR2_X1 U3830 ( .A1(n5039), .A2(n5072), .ZN(n5071) );
  OR3_X1 U3831 ( .A1(n4271), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4272), 
        .ZN(n2971) );
  AND4_X1 U3832 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n2972)
         );
  NOR2_X1 U3833 ( .A1(n5135), .A2(n5229), .ZN(n5223) );
  AND2_X1 U3834 ( .A1(n5290), .A2(n5363), .ZN(n2973) );
  AND2_X1 U3835 ( .A1(n5251), .A2(n5252), .ZN(n5152) );
  NAND2_X1 U3836 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  NOR2_X1 U3838 ( .A1(n4985), .A2(n5036), .ZN(n5035) );
  NOR2_X1 U3839 ( .A1(n4369), .A2(n4370), .ZN(n4528) );
  OR2_X1 U3840 ( .A1(n4469), .A2(n2986), .ZN(n2974) );
  AND2_X1 U3841 ( .A1(n2984), .A2(n2982), .ZN(n2975) );
  NOR2_X1 U3842 ( .A1(n5072), .A2(n2987), .ZN(n2976) );
  AND2_X1 U3843 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2977) );
  OAI21_X1 U3844 ( .B1(n3275), .B2(n3274), .A(n3316), .ZN(n4416) );
  INV_X1 U3845 ( .A(n6083), .ZN(n6126) );
  NAND2_X1 U3846 ( .A1(n4528), .A2(n4529), .ZN(n4468) );
  NAND2_X1 U3847 ( .A1(n3730), .A2(n3729), .ZN(n4355) );
  OR2_X1 U3848 ( .A1(n3439), .A2(n5656), .ZN(n2978) );
  NAND2_X1 U3849 ( .A1(n3599), .A2(n3598), .ZN(n4530) );
  NAND2_X1 U3850 ( .A1(n2961), .A2(n4491), .ZN(n4943) );
  INV_X1 U3851 ( .A(n4943), .ZN(n3224) );
  AND4_X1 U3852 ( .A1(n5421), .A2(n5400), .A3(n4225), .A4(n4206), .ZN(n2979)
         );
  NAND2_X1 U3853 ( .A1(n5433), .A2(n5438), .ZN(n2980) );
  AND2_X1 U3854 ( .A1(n2970), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n2981)
         );
  INV_X1 U3855 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5354) );
  AND2_X2 U3856 ( .A1(n4529), .A2(n2985), .ZN(n2984) );
  NOR3_X2 U3857 ( .A1(n5135), .A2(n5215), .A3(n2989), .ZN(n4254) );
  AND2_X2 U3858 ( .A1(n4254), .A2(n4093), .ZN(n4262) );
  NAND2_X1 U3859 ( .A1(n4958), .A2(n4987), .ZN(n4985) );
  NAND4_X1 U3860 ( .A1(n2995), .A2(n3149), .A3(n3147), .A4(n2994), .ZN(n3551)
         );
  NAND2_X2 U3861 ( .A1(n2996), .A2(n2997), .ZN(n2995) );
  NAND2_X1 U3862 ( .A1(n2995), .A2(n3147), .ZN(n3528) );
  NAND2_X1 U3863 ( .A1(n4216), .A2(n2998), .ZN(U2956) );
  XNOR2_X2 U3864 ( .A(n3349), .B(n4449), .ZN(n4448) );
  OR2_X2 U3865 ( .A1(n5520), .A2(n3457), .ZN(n3005) );
  NAND2_X1 U3866 ( .A1(n3275), .A2(n3274), .ZN(n3316) );
  INV_X1 U3867 ( .A(n3274), .ZN(n3008) );
  NAND3_X1 U3868 ( .A1(n3275), .A2(n3008), .A3(n6530), .ZN(n3007) );
  OAI21_X2 U3869 ( .B1(n4963), .B2(n4967), .A(n4965), .ZN(n5640) );
  OAI21_X2 U3870 ( .B1(n5953), .B2(n3451), .A(n3450), .ZN(n4963) );
  XNOR2_X1 U3871 ( .A(n3418), .B(n3419), .ZN(n3743) );
  NAND2_X1 U3872 ( .A1(n4463), .A2(n4464), .ZN(n4369) );
  AOI21_X1 U3873 ( .B1(n4255), .B2(n5217), .A(n4262), .ZN(n5207) );
  AOI22_X1 U3874 ( .A1(n3123), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3875 ( .A1(n3684), .A2(n3852), .ZN(n3691) );
  NAND2_X1 U3876 ( .A1(n3249), .A2(n3251), .ZN(n3250) );
  CLKBUF_X1 U3877 ( .A(n4191), .Z(n4244) );
  NAND2_X1 U3878 ( .A1(n5342), .A2(n6029), .ZN(n4218) );
  CLKBUF_X1 U3879 ( .A(n6016), .Z(n6019) );
  OAI21_X2 U3880 ( .B1(n5048), .B2(n3456), .A(n3455), .ZN(n5520) );
  AND2_X1 U3881 ( .A1(n5279), .A2(n4209), .ZN(n3010) );
  AND2_X1 U3882 ( .A1(n4188), .A2(n4187), .ZN(n3011) );
  AND2_X2 U3883 ( .A1(n4129), .A2(n5945), .ZN(n5861) );
  NOR2_X1 U3884 ( .A1(n6229), .A2(n6490), .ZN(n3012) );
  INV_X1 U3885 ( .A(n5900), .ZN(n6614) );
  AND2_X1 U3886 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3013) );
  NAND2_X1 U3887 ( .A1(n6326), .A2(n4193), .ZN(n6238) );
  NOR2_X1 U3888 ( .A1(n6229), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3014)
         );
  OR2_X1 U3889 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4092) );
  INV_X1 U3890 ( .A(n4092), .ZN(n4121) );
  INV_X1 U3891 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4432) );
  OR2_X1 U3892 ( .A1(n4894), .A2(n4876), .ZN(n3015) );
  BUF_X1 U3893 ( .A(n4208), .Z(n5279) );
  NAND2_X1 U3894 ( .A1(n5988), .A2(n5991), .ZN(n5990) );
  INV_X2 U3895 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6530) );
  INV_X1 U3896 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3471) );
  INV_X1 U3897 ( .A(n3551), .ZN(n3552) );
  INV_X1 U3898 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4193) );
  OR2_X1 U3899 ( .A1(n3234), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3016)
         );
  AND2_X1 U3900 ( .A1(n5852), .A2(n3685), .ZN(n5850) );
  OR2_X1 U3901 ( .A1(n3487), .A2(n3486), .ZN(n3474) );
  AND2_X1 U3902 ( .A1(n4495), .A2(n4491), .ZN(n3137) );
  INV_X1 U3903 ( .A(n3234), .ZN(n3235) );
  NAND2_X1 U3904 ( .A1(n6309), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3476) );
  AND2_X1 U3905 ( .A1(n3476), .A2(n3475), .ZN(n3502) );
  INV_X1 U3906 ( .A(n3431), .ZN(n3205) );
  NAND2_X1 U3907 ( .A1(n3477), .A2(n3476), .ZN(n3509) );
  OR2_X1 U3908 ( .A1(n3383), .A2(n3382), .ZN(n3409) );
  NOR2_X1 U3909 ( .A1(n4946), .A2(n6530), .ZN(n3323) );
  AOI22_X1 U3910 ( .A1(n3326), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3911 ( .A1(n3324), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3038) );
  INV_X1 U3912 ( .A(n4323), .ZN(n3223) );
  INV_X1 U3913 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U3914 ( .A1(n5999), .A2(n5998), .ZN(n5997) );
  AOI22_X1 U3915 ( .A1(n3324), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U3916 ( .A1(n3326), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3047) );
  NOR2_X1 U3917 ( .A1(n3200), .A2(n6530), .ZN(n4123) );
  NOR2_X1 U3918 ( .A1(n4052), .A2(n5288), .ZN(n4053) );
  INV_X1 U3919 ( .A(n3688), .ZN(n3689) );
  NAND2_X1 U3920 ( .A1(n3439), .A2(n4220), .ZN(n4221) );
  NAND2_X1 U3921 ( .A1(n4880), .A2(n4879), .ZN(n5953) );
  NAND2_X1 U3922 ( .A1(n3702), .A2(n3533), .ZN(n3248) );
  INV_X1 U3923 ( .A(n3503), .ZN(n3521) );
  AND4_X1 U3924 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3106)
         );
  OR2_X1 U3925 ( .A1(n4137), .A2(n4136), .ZN(n4138) );
  OR2_X1 U3926 ( .A1(n3995), .A2(n3994), .ZN(n4011) );
  NAND2_X1 U3927 ( .A1(n4946), .A2(n4491), .ZN(n3155) );
  AND2_X1 U3928 ( .A1(n3527), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4086) );
  NAND2_X1 U3929 ( .A1(n3726), .A2(n4321), .ZN(n4357) );
  INV_X1 U3930 ( .A(n4471), .ZN(n3604) );
  NAND2_X1 U3931 ( .A1(n5806), .A2(n5805), .ZN(n5808) );
  NOR2_X1 U3932 ( .A1(n3558), .A2(n4943), .ZN(n4411) );
  INV_X1 U3933 ( .A(n4936), .ZN(n4907) );
  OAI21_X1 U3934 ( .B1(n5517), .B2(n4193), .A(n5491), .ZN(n5513) );
  NOR2_X1 U3935 ( .A1(n4570), .A2(n4447), .ZN(n4580) );
  INV_X1 U3936 ( .A(n4781), .ZN(n6235) );
  INV_X1 U3937 ( .A(n4768), .ZN(n4833) );
  NAND2_X1 U3938 ( .A1(n6513), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U3939 ( .A1(n3941), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3983)
         );
  OR2_X1 U3940 ( .A1(n4175), .A2(n5817), .ZN(n5693) );
  AND2_X1 U3941 ( .A1(n5804), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4177) );
  INV_X1 U3942 ( .A(n4177), .ZN(n4178) );
  OR2_X1 U3943 ( .A1(n4125), .A2(n4124), .ZN(n4324) );
  NAND2_X1 U3944 ( .A1(n4000), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4016)
         );
  INV_X1 U3945 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5171) );
  NOR2_X1 U3946 ( .A1(n3784), .A2(n3783), .ZN(n3787) );
  NOR2_X2 U3947 ( .A1(n3683), .A2(n6326), .ZN(n3852) );
  NOR2_X1 U3948 ( .A1(n3558), .A2(n3557), .ZN(n6316) );
  INV_X1 U3949 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4210) );
  OR2_X1 U3950 ( .A1(n5398), .A2(n5361), .ZN(n5371) );
  NOR2_X1 U3951 ( .A1(n2965), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5297)
         );
  NAND2_X1 U3952 ( .A1(n3591), .A2(n3590), .ZN(n4460) );
  OR2_X1 U3953 ( .A1(n6068), .A2(n6121), .ZN(n6112) );
  OR2_X1 U3954 ( .A1(n3665), .A2(n3663), .ZN(n5056) );
  INV_X1 U3955 ( .A(n4447), .ZN(n4903) );
  NAND2_X1 U3956 ( .A1(n3525), .A2(n3524), .ZN(n4438) );
  AND2_X1 U3957 ( .A1(n3230), .A2(n3269), .ZN(n4724) );
  NAND2_X1 U3958 ( .A1(n4580), .A2(n4906), .ZN(n5030) );
  NAND2_X1 U3959 ( .A1(n4685), .A2(n4906), .ZN(n4835) );
  NAND2_X1 U3960 ( .A1(n5086), .A2(n4478), .ZN(n4520) );
  OR2_X1 U3961 ( .A1(n6328), .A2(n6530), .ZN(n6347) );
  INV_X1 U3962 ( .A(n6339), .ZN(n6453) );
  NOR2_X1 U3963 ( .A1(n6404), .A2(n5592), .ZN(n5160) );
  NOR2_X1 U3964 ( .A1(n6399), .A2(n5181), .ZN(n5174) );
  AND3_X1 U3965 ( .A1(n4181), .A2(EBX_REG_31__SCAN_IN), .A3(n5123), .ZN(n4166)
         );
  OR2_X1 U3966 ( .A1(n6448), .A2(n4145), .ZN(n5804) );
  OR2_X2 U3967 ( .A1(n5131), .A2(n5132), .ZN(n5232) );
  NOR2_X2 U3968 ( .A1(n5065), .A2(n3623), .ZN(n5081) );
  INV_X1 U3969 ( .A(n5852), .ZN(n5261) );
  AOI211_X1 U3970 ( .C1(n4245), .C2(n4121), .A(n3999), .B(n3998), .ZN(n4243)
         );
  AND2_X1 U3971 ( .A1(n5109), .A2(n4466), .ZN(n5042) );
  NOR2_X1 U3972 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6352), .ZN(n5883) );
  AND2_X1 U3973 ( .A1(n4307), .A2(n4407), .ZN(n5890) );
  INV_X1 U3974 ( .A(n5951), .ZN(n6613) );
  NAND2_X1 U3975 ( .A1(n3911), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3940)
         );
  NOR2_X1 U3976 ( .A1(n3883), .A2(n5190), .ZN(n3884) );
  INV_X1 U3977 ( .A(n3721), .ZN(n3698) );
  INV_X1 U3978 ( .A(n4222), .ZN(n5304) );
  INV_X1 U3979 ( .A(n4888), .ZN(n6107) );
  NAND2_X1 U3980 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4438), .ZN(n6338) );
  OAI21_X1 U3981 ( .B1(n4733), .B2(n4732), .A(n4731), .ZN(n4755) );
  OAI221_X1 U3982 ( .B1(n4938), .B2(n4193), .C1(n4938), .C2(n4911), .A(n4910), 
        .ZN(n4935) );
  INV_X1 U3983 ( .A(n6155), .ZN(n6159) );
  INV_X1 U3984 ( .A(n6227), .ZN(n6207) );
  AND2_X1 U3985 ( .A1(n6166), .A2(n6233), .ZN(n6174) );
  NAND2_X1 U3986 ( .A1(n4854), .A2(n4853), .ZN(n6224) );
  AND2_X1 U3987 ( .A1(n4541), .A2(n3709), .ZN(n6222) );
  OAI211_X1 U3988 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6326), .A(n4910), .B(n4788), .ZN(n4810) );
  AND2_X1 U3989 ( .A1(n4447), .A2(n4906), .ZN(n4850) );
  AND2_X1 U3990 ( .A1(n4447), .A2(n3709), .ZN(n4998) );
  OR2_X1 U3991 ( .A1(n4653), .A2(n4652), .ZN(n4675) );
  OAI211_X1 U3992 ( .C1(n4692), .C2(n4691), .A(n5005), .B(n4690), .ZN(n4714)
         );
  NOR2_X1 U3993 ( .A1(n5921), .A2(n4650), .ZN(n6244) );
  NOR2_X1 U3994 ( .A1(n5928), .A2(n4650), .ZN(n6268) );
  NOR2_X1 U3995 ( .A1(n5933), .A2(n4650), .ZN(n6290) );
  NOR2_X1 U3996 ( .A1(n6513), .A2(n6326), .ZN(n4439) );
  INV_X1 U3997 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6514) );
  INV_X1 U3998 ( .A(n6458), .ZN(n6447) );
  INV_X1 U3999 ( .A(n5782), .ZN(n5793) );
  INV_X1 U4000 ( .A(n5821), .ZN(n5836) );
  OR2_X1 U4001 ( .A1(n5213), .A2(n5212), .ZN(n5529) );
  INV_X1 U4002 ( .A(n5849), .ZN(n5267) );
  INV_X1 U4003 ( .A(n5042), .ZN(n4841) );
  OR2_X1 U4004 ( .A1(n5890), .A2(n6450), .ZN(n5888) );
  INV_X1 U4005 ( .A(n5883), .ZN(n5892) );
  INV_X1 U4006 ( .A(n4297), .ZN(n5900) );
  INV_X1 U4007 ( .A(n4270), .ZN(n4275) );
  INV_X1 U4008 ( .A(n4249), .ZN(n4250) );
  INV_X1 U4009 ( .A(n6012), .ZN(n6035) );
  AND2_X1 U4010 ( .A1(n4239), .A2(n4238), .ZN(n4240) );
  INV_X1 U4011 ( .A(n6037), .ZN(n5663) );
  OR2_X1 U4012 ( .A1(n4891), .A2(n6093), .ZN(n6064) );
  OR2_X1 U4013 ( .A1(n3665), .A2(n3564), .ZN(n6083) );
  INV_X1 U4014 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6303) );
  INV_X1 U4015 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5106) );
  OR2_X1 U4016 ( .A1(n5484), .A2(n4906), .ZN(n6155) );
  AOI22_X1 U4017 ( .A1(n4576), .A2(n4578), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4575), .ZN(n4607) );
  NAND2_X1 U4018 ( .A1(n4999), .A2(n4850), .ZN(n6227) );
  INV_X1 U4019 ( .A(n6178), .ZN(n6247) );
  NAND2_X1 U4020 ( .A1(n4781), .A2(n4850), .ZN(n6278) );
  INV_X1 U4021 ( .A(n4767), .ZN(n4839) );
  INV_X1 U4022 ( .A(n6256), .ZN(n6189) );
  INV_X1 U4023 ( .A(n6290), .ZN(n6211) );
  INV_X1 U4024 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6363) );
  OR2_X1 U4025 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6418), .ZN(n6416) );
  NOR2_X4 U4026 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4390) );
  AND2_X4 U4027 ( .A1(n3017), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5087)
         );
  AND2_X4 U4028 ( .A1(n4390), .A2(n5087), .ZN(n3132) );
  NAND2_X1 U4029 ( .A1(n3132), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3020) );
  AND2_X4 U4030 ( .A1(n5089), .A2(n4391), .ZN(n3184) );
  NAND2_X1 U4031 ( .A1(n3184), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3019)
         );
  INV_X1 U4032 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3021) );
  AND2_X4 U4033 ( .A1(n5087), .A2(n3027), .ZN(n3121) );
  INV_X1 U4034 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3022) );
  AND2_X4 U4035 ( .A1(n3022), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4394)
         );
  NOR2_X4 U4036 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4431) );
  AND2_X4 U4037 ( .A1(n4394), .A2(n4431), .ZN(n3171) );
  AND2_X4 U4038 ( .A1(n4431), .A2(n4391), .ZN(n4075) );
  AND2_X4 U4039 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4389) );
  AND2_X4 U4040 ( .A1(n4391), .A2(n4389), .ZN(n3131) );
  AOI22_X1 U4041 ( .A1(n4075), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3024) );
  AND2_X4 U4043 ( .A1(n4390), .A2(n4389), .ZN(n3130) );
  AND2_X4 U4044 ( .A1(n4431), .A2(n3027), .ZN(n3123) );
  AOI22_X1 U4045 ( .A1(n3324), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3031) );
  AND2_X2 U4046 ( .A1(n5089), .A2(n3027), .ZN(n3172) );
  AND2_X4 U4047 ( .A1(n4394), .A2(n4389), .ZN(n3129) );
  AND2_X2 U4048 ( .A1(n4431), .A2(n4390), .ZN(n3124) );
  AOI22_X1 U4049 ( .A1(n3326), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        INSTQUEUE_REG_0__6__SCAN_IN), .B2(n3124), .ZN(n3028) );
  AOI22_X1 U4050 ( .A1(n3326), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        INSTQUEUE_REG_0__7__SCAN_IN), .B2(n3124), .ZN(n3037) );
  AOI22_X1 U4051 ( .A1(n3172), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3036) );
  AOI22_X1 U4052 ( .A1(n3129), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3123), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3034) );
  AOI22_X1 U4053 ( .A1(n3171), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3041) );
  AOI22_X1 U4054 ( .A1(n3207), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3040) );
  AOI22_X1 U4055 ( .A1(n3331), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3039) );
  NAND2_X2 U4056 ( .A1(n3043), .A2(n3042), .ZN(n3685) );
  AOI22_X1 U4057 ( .A1(n3331), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3124), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3048) );
  AOI22_X1 U4058 ( .A1(n3207), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3046) );
  AOI22_X1 U4059 ( .A1(n3122), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U4060 ( .A1(n3172), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3129), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3052) );
  NAND2_X2 U4061 ( .A1(n3055), .A2(n3054), .ZN(n3243) );
  NAND2_X1 U4062 ( .A1(n3243), .A2(n3685), .ZN(n3056) );
  AOI22_X1 U4063 ( .A1(n3331), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3124), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3060) );
  AOI22_X1 U4064 ( .A1(n3207), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U4065 ( .A1(n3324), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3061) );
  AOI22_X1 U4066 ( .A1(n3172), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3129), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U4067 ( .A1(n2959), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U4068 ( .A1(n3123), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U4069 ( .A1(n3121), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U4070 ( .A1(n3207), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U4071 ( .A1(n2959), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U4072 ( .A1(n4075), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3067)
         );
  NAND2_X1 U4073 ( .A1(n3184), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3074)
         );
  NAND2_X1 U4074 ( .A1(n3172), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U4075 ( .A1(n3326), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3072)
         );
  NAND2_X1 U4076 ( .A1(n3130), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U4077 ( .A1(n3171), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3078) );
  NAND2_X1 U4078 ( .A1(n3324), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3077)
         );
  NAND2_X1 U4079 ( .A1(n3129), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3076)
         );
  NAND2_X1 U4080 ( .A1(n3123), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U4081 ( .A1(n3132), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U4082 ( .A1(n3331), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U4083 ( .A1(n3124), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U4084 ( .A1(n3131), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3079)
         );
  NAND4_X4 U4085 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n4946)
         );
  NAND2_X1 U4086 ( .A1(n3324), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U4087 ( .A1(n3121), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U4088 ( .A1(n3123), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U4089 ( .A1(n3171), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U4090 ( .A1(n3129), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3094)
         );
  NAND2_X1 U4091 ( .A1(n3172), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U4092 ( .A1(n3122), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U4093 ( .A1(n4075), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U4094 ( .A1(n3207), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U4095 ( .A1(n3132), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U4096 ( .A1(n3184), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3096)
         );
  NAND2_X1 U4097 ( .A1(n3131), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3095)
         );
  NAND2_X1 U4098 ( .A1(n3331), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4099 ( .A1(n3326), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3101)
         );
  NAND2_X1 U4100 ( .A1(n3124), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U4101 ( .A1(n3130), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3099) );
  NAND2_X1 U4102 ( .A1(n3146), .A2(n3243), .ZN(n3138) );
  AOI22_X1 U4103 ( .A1(n3184), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4104 ( .A1(n3172), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3132), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4105 ( .A1(n3331), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3326), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4106 ( .A1(n3121), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3129), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U4107 ( .A1(n3123), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4108 ( .A1(n3207), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4109 ( .A1(n3124), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3112) );
  NAND2_X2 U4110 ( .A1(n3116), .A2(n3115), .ZN(n3148) );
  OAI22_X1 U4111 ( .A1(n3118), .A2(n3155), .B1(n3557), .B2(n3571), .ZN(n3119)
         );
  INV_X1 U4112 ( .A(n3119), .ZN(n3161) );
  NAND2_X1 U4113 ( .A1(n2960), .A2(n3200), .ZN(n3158) );
  INV_X1 U4114 ( .A(n3243), .ZN(n4510) );
  AOI22_X1 U4115 ( .A1(n3121), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4116 ( .A1(n3184), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4117 ( .A1(n3123), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3122), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4118 ( .A1(n3326), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3124), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4119 ( .A1(n3324), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3129), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4120 ( .A1(n3172), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4121 ( .A1(n3331), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4122 ( .A1(n3132), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U4123 ( .A1(n3526), .A2(n3137), .ZN(n3145) );
  INV_X1 U4124 ( .A(n3138), .ZN(n3139) );
  NAND2_X1 U4125 ( .A1(n3139), .A2(n3653), .ZN(n3226) );
  NOR2_X2 U4126 ( .A1(n3653), .A2(n3243), .ZN(n3222) );
  INV_X1 U4127 ( .A(n3222), .ZN(n3140) );
  NAND2_X1 U4128 ( .A1(n3226), .A2(n3140), .ZN(n3143) );
  INV_X1 U4129 ( .A(n3685), .ZN(n3141) );
  AND2_X1 U4130 ( .A1(n3225), .A2(n4500), .ZN(n3142) );
  AOI21_X1 U4131 ( .B1(n3143), .B2(n3142), .A(n4946), .ZN(n3144) );
  NAND2_X1 U4132 ( .A1(n3145), .A2(n3144), .ZN(n3164) );
  NAND2_X2 U4133 ( .A1(n3532), .A2(n3243), .ZN(n3156) );
  NAND2_X1 U4134 ( .A1(n3156), .A2(n3200), .ZN(n3149) );
  INV_X1 U4135 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U4136 ( .A1(n6577), .A2(n6363), .ZN(n6365) );
  INV_X1 U4137 ( .A(n6365), .ZN(n3150) );
  OAI21_X1 U4138 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n3150), .ZN(n3538) );
  NAND2_X1 U4139 ( .A1(n4491), .A2(n3538), .ZN(n3221) );
  AOI21_X1 U4140 ( .B1(n3221), .B2(n4510), .A(n3653), .ZN(n3151) );
  NAND4_X1 U4141 ( .A1(n3161), .A2(n3164), .A3(n2969), .A4(n3151), .ZN(n3152)
         );
  INV_X1 U4142 ( .A(n6328), .ZN(n3319) );
  NAND2_X1 U4143 ( .A1(n5665), .A2(n6530), .ZN(n4194) );
  MUX2_X1 U4144 ( .A(n3319), .B(n4194), .S(n4997), .Z(n3153) );
  INV_X2 U4145 ( .A(n4491), .ZN(n3560) );
  NAND2_X1 U4146 ( .A1(n3156), .A2(n3148), .ZN(n3157) );
  NAND2_X1 U4147 ( .A1(n5665), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6346) );
  AOI21_X1 U4148 ( .B1(n4296), .B2(n3157), .A(n6346), .ZN(n3162) );
  INV_X1 U4149 ( .A(n3158), .ZN(n3160) );
  NAND2_X1 U4150 ( .A1(n4500), .A2(n4495), .ZN(n3658) );
  NOR2_X1 U4151 ( .A1(n3658), .A2(n4946), .ZN(n3159) );
  NAND2_X1 U4152 ( .A1(n3160), .A2(n3159), .ZN(n4417) );
  NAND4_X1 U4153 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n4417), .ZN(n3166)
         );
  NAND2_X1 U4154 ( .A1(n3653), .A2(n4946), .ZN(n3165) );
  NAND2_X1 U4155 ( .A1(n3164), .A2(n3165), .ZN(n3660) );
  NOR2_X1 U4156 ( .A1(n3166), .A2(n3660), .ZN(n3167) );
  INV_X1 U4157 ( .A(n3167), .ZN(n3168) );
  OAI21_X1 U4158 ( .B1(n3169), .B2(n3168), .A(n3238), .ZN(n3711) );
  INV_X1 U4159 ( .A(n3711), .ZN(n3170) );
  NAND2_X1 U4160 ( .A1(n3170), .A2(n6530), .ZN(n3249) );
  AOI22_X1 U4161 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4018), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4162 ( .A1(n3276), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4163 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n4095), .B1(n4104), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3174) );
  CLKBUF_X2 U4164 ( .A(n4075), .Z(n3351) );
  AOI22_X1 U4165 ( .A1(n3122), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3173) );
  NAND4_X1 U4166 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3182)
         );
  AOI22_X1 U4168 ( .A1(n3325), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3180) );
  INV_X1 U4169 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6581) );
  AOI22_X1 U4170 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n4097), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4171 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n3282), .B1(n3130), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4172 ( .A1(n3207), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3131), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3177) );
  NAND4_X1 U4173 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3181)
         );
  INV_X1 U4174 ( .A(n3436), .ZN(n3183) );
  NAND2_X1 U4175 ( .A1(n4123), .A2(n3183), .ZN(n3218) );
  INV_X1 U4176 ( .A(n3218), .ZN(n3196) );
  NAND2_X1 U4177 ( .A1(n4505), .A2(n3436), .ZN(n3198) );
  AOI22_X1 U4178 ( .A1(n4094), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3188) );
  BUF_X1 U4179 ( .A(n3184), .Z(n3281) );
  AOI22_X1 U4180 ( .A1(n3281), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4181 ( .A1(n4097), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4182 ( .A1(n4095), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3185) );
  NAND4_X1 U4183 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3194)
         );
  AOI22_X1 U4184 ( .A1(n4018), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4185 ( .A1(n4104), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4186 ( .A1(n3207), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4187 ( .A1(n4105), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3189) );
  NAND4_X1 U4188 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3193)
         );
  INV_X1 U4189 ( .A(n3255), .ZN(n3195) );
  MUX2_X1 U4190 ( .A(n3196), .B(n3431), .S(n3195), .Z(n3252) );
  INV_X1 U4191 ( .A(n3252), .ZN(n3197) );
  NAND2_X1 U4192 ( .A1(n3249), .A2(n3197), .ZN(n3204) );
  AOI21_X1 U4193 ( .B1(n2961), .B2(n3255), .A(n6530), .ZN(n3199) );
  AND2_X1 U4194 ( .A1(n3199), .A2(n3198), .ZN(n3203) );
  INV_X1 U4195 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3201) );
  OR2_X1 U4196 ( .A1(n3504), .A2(n3201), .ZN(n3202) );
  INV_X1 U4197 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4198 ( .A1(n4018), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4199 ( .A1(n4095), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4200 ( .A1(n4036), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4201 ( .A1(n3281), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3208) );
  NAND4_X1 U4202 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3217)
         );
  AOI22_X1 U4203 ( .A1(n4104), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4204 ( .A1(n4105), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3214) );
  AOI22_X1 U4205 ( .A1(n4097), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4206 ( .A1(n2959), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3212) );
  NAND4_X1 U4207 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3216)
         );
  NAND2_X1 U4208 ( .A1(n3323), .A2(n3244), .ZN(n3219) );
  NAND2_X1 U4210 ( .A1(n4139), .A2(n3221), .ZN(n3228) );
  NAND2_X1 U4211 ( .A1(n3222), .A2(n4500), .ZN(n4323) );
  OR2_X2 U4212 ( .A1(n4382), .A2(n4130), .ZN(n3565) );
  NAND3_X1 U4213 ( .A1(n3228), .A2(n3565), .A3(n5664), .ZN(n3229) );
  NAND2_X1 U4214 ( .A1(n3229), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3237) );
  INV_X1 U4215 ( .A(n3237), .ZN(n3233) );
  INV_X1 U4216 ( .A(n4194), .ZN(n3271) );
  NAND2_X1 U4217 ( .A1(n6303), .A2(n4997), .ZN(n3230) );
  NAND2_X1 U4218 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4219 ( .A1(n3271), .A2(n4724), .ZN(n3232) );
  NAND2_X1 U4220 ( .A1(n6328), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4221 ( .A1(n3232), .A2(n3231), .ZN(n3234) );
  NAND2_X1 U4222 ( .A1(n3233), .A2(n3016), .ZN(n3265) );
  NAND2_X1 U4223 ( .A1(n3267), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3236) );
  NAND3_X1 U4224 ( .A1(n3237), .A2(n3236), .A3(n3235), .ZN(n3263) );
  NAND2_X1 U4225 ( .A1(n3265), .A2(n3263), .ZN(n3239) );
  XNOR2_X1 U4226 ( .A(n3239), .B(n3264), .ZN(n4454) );
  NAND2_X1 U4227 ( .A1(n4454), .A2(n6530), .ZN(n3241) );
  NAND2_X1 U4228 ( .A1(n4123), .A2(n3244), .ZN(n3240) );
  NAND2_X2 U4229 ( .A1(n3241), .A2(n3240), .ZN(n3297) );
  NAND2_X1 U4230 ( .A1(n3244), .A2(n3255), .ZN(n3342) );
  OAI21_X1 U4231 ( .B1(n3255), .B2(n3244), .A(n3342), .ZN(n3245) );
  INV_X1 U4232 ( .A(n4296), .ZN(n6452) );
  OAI211_X1 U4233 ( .C1(n3245), .C2(n6452), .A(n4131), .B(n3148), .ZN(n3246)
         );
  INV_X1 U4234 ( .A(n3246), .ZN(n3247) );
  NAND2_X1 U4235 ( .A1(n3248), .A2(n3247), .ZN(n4363) );
  NAND2_X1 U4236 ( .A1(n3252), .A2(n3251), .ZN(n3253) );
  NAND2_X1 U4237 ( .A1(n2961), .A2(n3148), .ZN(n3308) );
  OAI21_X1 U4238 ( .B1(n6452), .B2(n3255), .A(n3308), .ZN(n3256) );
  INV_X1 U4239 ( .A(n3256), .ZN(n3257) );
  OAI21_X2 U4240 ( .B1(n3709), .B2(n3510), .A(n3257), .ZN(n4309) );
  NAND2_X1 U4241 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3258)
         );
  INV_X1 U4242 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U4243 ( .A1(n3258), .A2(n6507), .ZN(n3260) );
  AND2_X1 U4244 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4245 ( .A1(n4309), .A2(n3259), .ZN(n3261) );
  AND2_X1 U4246 ( .A1(n3260), .A2(n3261), .ZN(n4364) );
  NAND2_X1 U4247 ( .A1(n4363), .A2(n4364), .ZN(n3262) );
  NAND2_X1 U4248 ( .A1(n3262), .A2(n3261), .ZN(n6026) );
  NAND2_X1 U4249 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4250 ( .A1(n3264), .A2(n3263), .ZN(n3266) );
  INV_X1 U4251 ( .A(n3269), .ZN(n3268) );
  NAND2_X1 U4252 ( .A1(n3268), .A2(n6309), .ZN(n6229) );
  NAND2_X1 U4253 ( .A1(n3269), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4254 ( .A1(n6229), .A2(n3270), .ZN(n4649) );
  AOI22_X1 U4255 ( .A1(n3271), .A2(n4649), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6328), .ZN(n3272) );
  AOI22_X1 U4256 ( .A1(n4018), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4257 ( .A1(n3276), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3279) );
  INV_X1 U4258 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6565) );
  AOI22_X1 U4259 ( .A1(n4095), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4260 ( .A1(n3122), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4261 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3288)
         );
  AOI22_X1 U4262 ( .A1(n3281), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4263 ( .A1(n4097), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4264 ( .A1(n3282), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4265 ( .A1(n4036), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4266 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3287)
         );
  NAND2_X1 U4267 ( .A1(n4123), .A2(n3340), .ZN(n3289) );
  INV_X1 U4268 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4269 ( .A1(n3323), .A2(n3340), .ZN(n3290) );
  OAI21_X1 U4270 ( .B1(n3504), .B2(n3291), .A(n3290), .ZN(n3292) );
  XNOR2_X1 U4271 ( .A(n3293), .B(n3292), .ZN(n3304) );
  NAND2_X1 U4272 ( .A1(n3297), .A2(n3298), .ZN(n3296) );
  INV_X1 U4273 ( .A(n3294), .ZN(n3295) );
  NAND2_X1 U4274 ( .A1(n3296), .A2(n3295), .ZN(n3302) );
  INV_X1 U4275 ( .A(n3297), .ZN(n3300) );
  INV_X1 U4276 ( .A(n3298), .ZN(n3299) );
  NAND2_X1 U4277 ( .A1(n3300), .A2(n3299), .ZN(n3301) );
  NAND2_X1 U4278 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  NAND2_X1 U4279 ( .A1(n3304), .A2(n3303), .ZN(n3307) );
  INV_X1 U4280 ( .A(n3303), .ZN(n3306) );
  INV_X1 U4281 ( .A(n3304), .ZN(n3305) );
  AND2_X2 U4282 ( .A1(n3307), .A2(n3349), .ZN(n4446) );
  XNOR2_X1 U4283 ( .A(n3342), .B(n3340), .ZN(n3309) );
  OAI21_X1 U4284 ( .B1(n3309), .B2(n6452), .A(n3308), .ZN(n3310) );
  NAND2_X1 U4285 ( .A1(n3311), .A2(n6027), .ZN(n3315) );
  INV_X1 U4286 ( .A(n6026), .ZN(n3313) );
  INV_X1 U4287 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4288 ( .A1(n3313), .A2(n3312), .ZN(n3314) );
  NOR3_X1 U4289 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6309), .A3(n6303), 
        .ZN(n6177) );
  NAND2_X1 U4290 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6177), .ZN(n6171) );
  NAND2_X1 U4291 ( .A1(n6490), .A2(n6171), .ZN(n3318) );
  NAND3_X1 U4292 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4688) );
  INV_X1 U4293 ( .A(n4688), .ZN(n4485) );
  NAND2_X1 U4294 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4485), .ZN(n4527) );
  NAND2_X1 U4295 ( .A1(n3318), .A2(n4527), .ZN(n4723) );
  OAI22_X1 U4296 ( .A1(n4194), .A2(n4723), .B1(n3319), .B2(n6490), .ZN(n3320)
         );
  INV_X1 U4297 ( .A(n3320), .ZN(n3321) );
  AOI22_X1 U4298 ( .A1(n4018), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4299 ( .A1(n4104), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4300 ( .A1(n3281), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4301 ( .A1(n4036), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4302 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3337)
         );
  AOI22_X1 U4303 ( .A1(n4094), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4304 ( .A1(n4095), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4305 ( .A1(n4097), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4306 ( .A1(n4105), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3332) );
  NAND4_X1 U4307 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3336)
         );
  AOI22_X1 U4308 ( .A1(n3503), .A2(n3364), .B1(n3513), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4309 ( .A1(n4448), .A2(n3533), .ZN(n3346) );
  INV_X1 U4310 ( .A(n3340), .ZN(n3341) );
  NAND2_X1 U4311 ( .A1(n3342), .A2(n3341), .ZN(n3365) );
  INV_X1 U4312 ( .A(n3364), .ZN(n3343) );
  XNOR2_X1 U4313 ( .A(n3365), .B(n3343), .ZN(n3344) );
  NAND2_X1 U4314 ( .A1(n3344), .A2(n4296), .ZN(n3345) );
  INV_X1 U4315 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U4316 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  NAND2_X1 U4317 ( .A1(n3347), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3348)
         );
  NAND2_X1 U4318 ( .A1(n6018), .A2(n3348), .ZN(n6006) );
  INV_X1 U4319 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4320 ( .A1(n3350), .A2(n4449), .ZN(n3371) );
  AOI22_X1 U4321 ( .A1(n4018), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4322 ( .A1(n3276), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4323 ( .A1(n4095), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4324 ( .A1(n3122), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4325 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3361)
         );
  AOI22_X1 U4326 ( .A1(n3281), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4327 ( .A1(n4097), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4328 ( .A1(n3282), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4329 ( .A1(n4036), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3356) );
  NAND4_X1 U4330 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  NAND2_X1 U4331 ( .A1(n3503), .A2(n3386), .ZN(n3363) );
  INV_X1 U4332 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6596) );
  OR2_X1 U4333 ( .A1(n3504), .A2(n6596), .ZN(n3362) );
  NAND2_X1 U4334 ( .A1(n3363), .A2(n3362), .ZN(n3372) );
  XNOR2_X1 U4335 ( .A(n3371), .B(n3372), .ZN(n3696) );
  NAND2_X1 U4336 ( .A1(n3696), .A2(n3533), .ZN(n3368) );
  NAND2_X1 U4337 ( .A1(n3365), .A2(n3364), .ZN(n3388) );
  XNOR2_X1 U4338 ( .A(n3388), .B(n3386), .ZN(n3366) );
  NAND2_X1 U4339 ( .A1(n3366), .A2(n4296), .ZN(n3367) );
  INV_X1 U4340 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6522) );
  XNOR2_X1 U4341 ( .A(n3369), .B(n6522), .ZN(n6009) );
  NAND2_X1 U4342 ( .A1(n6006), .A2(n6009), .ZN(n6007) );
  NAND2_X1 U4343 ( .A1(n3369), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3370)
         );
  NAND2_X1 U4344 ( .A1(n6007), .A2(n3370), .ZN(n5999) );
  INV_X1 U4345 ( .A(n3371), .ZN(n3373) );
  NAND2_X1 U4346 ( .A1(n3373), .A2(n3372), .ZN(n3394) );
  AOI22_X1 U4347 ( .A1(n4018), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4348 ( .A1(n4104), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4349 ( .A1(n4097), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4350 ( .A1(n4036), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3374) );
  NAND4_X1 U4351 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3383)
         );
  AOI22_X1 U4352 ( .A1(n4095), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4353 ( .A1(n3281), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4354 ( .A1(n4396), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4355 ( .A1(n4105), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3378) );
  NAND4_X1 U4356 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3382)
         );
  NAND2_X1 U4357 ( .A1(n3503), .A2(n3409), .ZN(n3385) );
  NAND2_X1 U4358 ( .A1(n3513), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4359 ( .A1(n3385), .A2(n3384), .ZN(n3395) );
  XNOR2_X1 U4360 ( .A(n3394), .B(n3395), .ZN(n3732) );
  NAND2_X1 U4361 ( .A1(n3732), .A2(n3533), .ZN(n3391) );
  INV_X1 U4362 ( .A(n3386), .ZN(n3387) );
  OR2_X1 U4363 ( .A1(n3388), .A2(n3387), .ZN(n3410) );
  XNOR2_X1 U4364 ( .A(n3410), .B(n3409), .ZN(n3389) );
  NAND2_X1 U4365 ( .A1(n3389), .A2(n4296), .ZN(n3390) );
  NAND2_X1 U4366 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  INV_X1 U4367 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6082) );
  XNOR2_X1 U4368 ( .A(n3392), .B(n6082), .ZN(n5998) );
  NAND2_X1 U4369 ( .A1(n3392), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3393)
         );
  NAND2_X1 U4370 ( .A1(n5997), .A2(n3393), .ZN(n5988) );
  INV_X1 U4371 ( .A(n3394), .ZN(n3396) );
  AOI22_X1 U4372 ( .A1(n4018), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4373 ( .A1(n3276), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4374 ( .A1(n4095), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4375 ( .A1(n4396), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4376 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3406)
         );
  AOI22_X1 U4377 ( .A1(n3281), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4378 ( .A1(n4097), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3403) );
  INV_X1 U4379 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U4380 ( .A1(n3282), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4381 ( .A1(n4036), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4382 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3405)
         );
  NAND2_X1 U4383 ( .A1(n3503), .A2(n3424), .ZN(n3408) );
  NAND2_X1 U4384 ( .A1(n3513), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3407) );
  NAND2_X1 U4385 ( .A1(n3408), .A2(n3407), .ZN(n3419) );
  NAND2_X1 U4386 ( .A1(n3743), .A2(n3533), .ZN(n3415) );
  INV_X1 U4387 ( .A(n3409), .ZN(n3411) );
  NOR2_X1 U4388 ( .A1(n3411), .A2(n3410), .ZN(n3425) );
  INV_X1 U4389 ( .A(n3425), .ZN(n3412) );
  XNOR2_X1 U4390 ( .A(n3424), .B(n3412), .ZN(n3413) );
  NAND2_X1 U4391 ( .A1(n4296), .A2(n3413), .ZN(n3414) );
  NAND2_X1 U4392 ( .A1(n3415), .A2(n3414), .ZN(n3416) );
  INV_X1 U4393 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6076) );
  XNOR2_X1 U4394 ( .A(n3416), .B(n6076), .ZN(n5991) );
  NAND2_X1 U4395 ( .A1(n3416), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3417)
         );
  NAND2_X1 U4396 ( .A1(n5990), .A2(n3417), .ZN(n5981) );
  INV_X1 U4397 ( .A(n3418), .ZN(n3420) );
  INV_X1 U4398 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4399 ( .A1(n3503), .A2(n3436), .ZN(n3421) );
  OAI21_X1 U4400 ( .B1(n3504), .B2(n3422), .A(n3421), .ZN(n3423) );
  NAND2_X1 U4401 ( .A1(n3684), .A2(n3533), .ZN(n3428) );
  NAND2_X1 U4402 ( .A1(n3425), .A2(n3424), .ZN(n3434) );
  XNOR2_X1 U4403 ( .A(n3436), .B(n3434), .ZN(n3426) );
  NAND2_X1 U4404 ( .A1(n4296), .A2(n3426), .ZN(n3427) );
  NAND2_X1 U4405 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  INV_X1 U4406 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6050) );
  XNOR2_X1 U4407 ( .A(n3429), .B(n6050), .ZN(n5980) );
  NAND2_X1 U4408 ( .A1(n5981), .A2(n5980), .ZN(n5983) );
  NAND2_X1 U4409 ( .A1(n3429), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3430)
         );
  NAND2_X1 U4410 ( .A1(n5983), .A2(n3430), .ZN(n5962) );
  NOR2_X1 U4411 ( .A1(n3205), .A2(n3510), .ZN(n3432) );
  INV_X1 U4412 ( .A(n3434), .ZN(n3435) );
  NAND2_X1 U4413 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  OR2_X1 U4414 ( .A1(n6452), .A2(n3437), .ZN(n3438) );
  NAND2_X1 U4415 ( .A1(n3439), .A2(n3438), .ZN(n3442) );
  INV_X1 U4416 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6057) );
  XNOR2_X1 U4417 ( .A(n3442), .B(n6057), .ZN(n5972) );
  INV_X1 U4418 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U4419 ( .A1(n2965), .A2(n5965), .ZN(n3441) );
  AND2_X1 U4420 ( .A1(n5972), .A2(n3441), .ZN(n3440) );
  NAND2_X1 U4421 ( .A1(n5962), .A2(n3440), .ZN(n3447) );
  INV_X1 U4422 ( .A(n3441), .ZN(n3445) );
  NAND2_X1 U4423 ( .A1(n3442), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5964)
         );
  NAND2_X1 U4424 ( .A1(n4219), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3443)
         );
  AND2_X1 U4425 ( .A1(n5964), .A2(n3443), .ZN(n3444) );
  OR2_X1 U4426 ( .A1(n3445), .A2(n3444), .ZN(n3446) );
  NAND2_X1 U4427 ( .A1(n3447), .A2(n3446), .ZN(n4880) );
  INV_X1 U4428 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4429 ( .A1(n3439), .A2(n3448), .ZN(n4879) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5955) );
  AND2_X1 U4431 ( .A1(n3439), .A2(n5955), .ZN(n3451) );
  NAND2_X1 U4432 ( .A1(n4219), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U4433 ( .A1(n4219), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3449) );
  AND2_X1 U4434 ( .A1(n5954), .A2(n3449), .ZN(n3450) );
  INV_X1 U4435 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4975) );
  NOR2_X1 U4436 ( .A1(n2965), .A2(n4975), .ZN(n4967) );
  NAND2_X1 U4437 ( .A1(n3439), .A2(n4975), .ZN(n4965) );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4439 ( .A1(n3439), .A2(n3452), .ZN(n3453) );
  NAND2_X1 U4440 ( .A1(n3454), .A2(n3453), .ZN(n5048) );
  NAND2_X1 U4441 ( .A1(n4219), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3455) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U4443 ( .A1(n2965), .A2(n5656), .ZN(n5522) );
  NAND2_X1 U4444 ( .A1(n3439), .A2(n5467), .ZN(n5323) );
  INV_X1 U4445 ( .A(n5320), .ZN(n5449) );
  NAND2_X1 U4446 ( .A1(n5449), .A2(n3013), .ZN(n3460) );
  NOR2_X1 U4447 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5433) );
  INV_X1 U4448 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5438) );
  INV_X1 U4449 ( .A(n5311), .ZN(n3462) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3631) );
  XNOR2_X1 U4451 ( .A(n2965), .B(n3631), .ZN(n5314) );
  NAND2_X1 U4452 ( .A1(n2965), .A2(n3631), .ZN(n3463) );
  INV_X1 U4453 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U4454 ( .A1(n2965), .A2(n5418), .ZN(n3464) );
  NAND2_X1 U4455 ( .A1(n5417), .A2(n3464), .ZN(n3469) );
  AND2_X1 U4456 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U4457 ( .A1(n3439), .A2(n5399), .ZN(n3468) );
  NAND2_X1 U4458 ( .A1(n4219), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3465) );
  NAND2_X1 U4459 ( .A1(n3469), .A2(n3465), .ZN(n5305) );
  INV_X1 U4460 ( .A(n5305), .ZN(n3467) );
  XNOR2_X1 U4461 ( .A(n3439), .B(n4220), .ZN(n5306) );
  INV_X1 U4462 ( .A(n5306), .ZN(n3466) );
  NAND2_X1 U4463 ( .A1(n5304), .A2(n5297), .ZN(n4224) );
  OAI21_X1 U4464 ( .B1(n3469), .B2(n3468), .A(n4224), .ZN(n3470) );
  INV_X1 U4465 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U4466 ( .A1(n6303), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4467 ( .A1(n3471), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U4468 ( .A1(n3473), .A2(n3472), .ZN(n3487) );
  NAND2_X1 U4469 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n4997), .ZN(n3486) );
  NAND2_X1 U4470 ( .A1(n3474), .A2(n3473), .ZN(n3501) );
  NAND2_X1 U4471 ( .A1(n5106), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U4472 ( .A1(n3501), .A2(n3502), .ZN(n3477) );
  XNOR2_X1 U4473 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3507) );
  NOR2_X1 U4474 ( .A1(n4415), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3478)
         );
  NAND2_X1 U4475 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6314), .ZN(n3479) );
  NAND2_X1 U4476 ( .A1(n3483), .A2(n3479), .ZN(n3481) );
  NAND2_X1 U4477 ( .A1(n3483), .A2(n3482), .ZN(n3545) );
  NAND2_X1 U4478 ( .A1(n6530), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3484) );
  AOI21_X1 U4479 ( .B1(n3503), .B2(n3560), .A(n4510), .ZN(n3500) );
  INV_X1 U4480 ( .A(n3486), .ZN(n3489) );
  XNOR2_X1 U4481 ( .A(n3487), .B(n3489), .ZN(n3542) );
  NAND2_X1 U4482 ( .A1(n3542), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U4483 ( .A1(n4491), .A2(n4131), .ZN(n3488) );
  AOI21_X1 U4484 ( .B1(n6296), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n3489), 
        .ZN(n3495) );
  NAND2_X1 U4485 ( .A1(n3557), .A2(n3495), .ZN(n3491) );
  NAND2_X1 U4486 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  AND2_X1 U4487 ( .A1(n3511), .A2(n3492), .ZN(n3493) );
  AOI21_X1 U4488 ( .B1(n3500), .B2(n3499), .A(n3493), .ZN(n3496) );
  INV_X1 U4489 ( .A(n3542), .ZN(n3494) );
  OAI21_X1 U4490 ( .B1(n3496), .B2(n3494), .A(n3523), .ZN(n3498) );
  NAND3_X1 U4491 ( .A1(n3496), .A2(n3495), .A3(n3503), .ZN(n3497) );
  OAI211_X1 U4492 ( .C1(n3500), .C2(n3499), .A(n3498), .B(n3497), .ZN(n3506)
         );
  XOR2_X1 U4493 ( .A(n3502), .B(n3501), .Z(n3541) );
  NAND2_X1 U4494 ( .A1(n3503), .A2(n3541), .ZN(n3512) );
  OAI211_X1 U4495 ( .C1(n3541), .C2(n3504), .A(n3512), .B(n3511), .ZN(n3505)
         );
  AND2_X1 U4496 ( .A1(n3506), .A2(n3505), .ZN(n3515) );
  INV_X1 U4497 ( .A(n3507), .ZN(n3508) );
  XNOR2_X1 U4498 ( .A(n3509), .B(n3508), .ZN(n3540) );
  OAI22_X1 U4499 ( .A1(n3512), .A2(n3511), .B1(n3540), .B2(n3510), .ZN(n3514)
         );
  AOI222_X1 U4500 ( .A1(n3518), .A2(n3517), .B1(n3518), .B2(n3516), .C1(n3517), 
        .C2(n3516), .ZN(n3519) );
  INV_X1 U4501 ( .A(n3519), .ZN(n3520) );
  NAND2_X1 U4502 ( .A1(n3527), .A2(n3560), .ZN(n3549) );
  OR2_X1 U4503 ( .A1(n3527), .A2(n4946), .ZN(n3531) );
  NAND2_X1 U4504 ( .A1(n4495), .A2(n3148), .ZN(n3529) );
  NOR2_X1 U4505 ( .A1(n3528), .A2(n3529), .ZN(n3530) );
  NAND2_X1 U4506 ( .A1(n3531), .A2(n3530), .ZN(n3558) );
  NAND2_X1 U4507 ( .A1(n3533), .A2(n4515), .ZN(n3656) );
  AND2_X1 U4508 ( .A1(n3656), .A2(n4946), .ZN(n3534) );
  INV_X1 U4509 ( .A(n4286), .ZN(n3537) );
  OAI21_X1 U4510 ( .B1(n3558), .B2(n3661), .A(n3537), .ZN(n3655) );
  INV_X1 U4511 ( .A(n3538), .ZN(n3539) );
  NAND2_X1 U4512 ( .A1(n3539), .A2(n6514), .ZN(n6362) );
  NAND2_X1 U4513 ( .A1(n3560), .A2(n6362), .ZN(n3547) );
  NAND3_X1 U4514 ( .A1(n3542), .A2(n3541), .A3(n3540), .ZN(n3543) );
  NAND2_X1 U4515 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  AND2_X1 U4516 ( .A1(n3546), .A2(n3545), .ZN(n4285) );
  NOR2_X1 U4517 ( .A1(READY_N), .A2(n4285), .ZN(n4403) );
  NAND3_X1 U4518 ( .A1(n3547), .A2(n4403), .A3(n3653), .ZN(n3548) );
  OAI211_X1 U4519 ( .C1(n4438), .C2(n3549), .A(n3655), .B(n3548), .ZN(n3550)
         );
  NAND2_X1 U4520 ( .A1(n3550), .A2(n6329), .ZN(n3556) );
  NAND2_X1 U4521 ( .A1(n4491), .A2(n6362), .ZN(n4169) );
  NAND3_X1 U4522 ( .A1(n3552), .A2(n4295), .A3(n4169), .ZN(n3553) );
  NAND3_X1 U4523 ( .A1(n3553), .A2(n4946), .A3(n4130), .ZN(n3554) );
  NAND3_X1 U4524 ( .A1(n4305), .A2(n4495), .A3(n3554), .ZN(n3555) );
  INV_X1 U4525 ( .A(n4411), .ZN(n3563) );
  INV_X1 U4526 ( .A(n6316), .ZN(n3562) );
  OAI21_X1 U4527 ( .B1(n3565), .B2(n4505), .A(n5664), .ZN(n3559) );
  INV_X1 U4528 ( .A(n3559), .ZN(n3561) );
  NAND2_X1 U4529 ( .A1(n4946), .A2(n3560), .ZN(n3584) );
  INV_X2 U4530 ( .A(n3584), .ZN(n4167) );
  NAND2_X1 U4531 ( .A1(n3552), .A2(n4167), .ZN(n4408) );
  AND4_X1 U4532 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n4408), .ZN(n3564)
         );
  NAND2_X1 U4533 ( .A1(n3552), .A2(n4296), .ZN(n6334) );
  INV_X1 U4534 ( .A(n3565), .ZN(n3566) );
  NAND2_X1 U4535 ( .A1(n3566), .A2(n4505), .ZN(n3567) );
  AND2_X1 U4536 ( .A1(n6334), .A2(n3567), .ZN(n3568) );
  NAND2_X1 U4537 ( .A1(n3577), .A2(EBX_REG_0__SCAN_IN), .ZN(n3570) );
  INV_X1 U4538 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U4539 ( .A1(n2962), .A2(n5837), .ZN(n3569) );
  NAND2_X1 U4540 ( .A1(n3570), .A2(n3569), .ZN(n4332) );
  MUX2_X1 U4541 ( .A(n2963), .B(n3577), .S(EBX_REG_1__SCAN_IN), .Z(n3573) );
  NAND2_X1 U4542 ( .A1(n3584), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3572)
         );
  XNOR2_X1 U4543 ( .A(n4332), .B(n3574), .ZN(n4949) );
  INV_X1 U4544 ( .A(n3574), .ZN(n3575) );
  NAND2_X1 U4545 ( .A1(n3575), .A2(n4332), .ZN(n3576) );
  NAND2_X1 U4546 ( .A1(n4328), .A2(n3576), .ZN(n4360) );
  NAND2_X1 U4547 ( .A1(n2964), .A2(n3312), .ZN(n3579) );
  INV_X1 U4548 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3581) );
  NAND2_X1 U4549 ( .A1(n4167), .A2(n3581), .ZN(n3578) );
  NAND3_X1 U4550 ( .A1(n3579), .A2(n2963), .A3(n3578), .ZN(n3583) );
  NAND2_X1 U4551 ( .A1(n3580), .A2(n3581), .ZN(n3582) );
  AND2_X1 U4552 ( .A1(n3583), .A2(n3582), .ZN(n4359) );
  NOR2_X2 U4553 ( .A1(n4360), .A2(n4359), .ZN(n5806) );
  INV_X1 U4554 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U4555 ( .A1(n3646), .A2(n6482), .ZN(n3587) );
  NAND2_X1 U4556 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3585)
         );
  OAI211_X1 U4557 ( .C1(n4156), .C2(EBX_REG_3__SCAN_IN), .A(n2964), .B(n3585), 
        .ZN(n3586) );
  AND2_X1 U4558 ( .A1(n3587), .A2(n3586), .ZN(n5805) );
  MUX2_X1 U4559 ( .A(n2963), .B(n2964), .S(EBX_REG_4__SCAN_IN), .Z(n3589) );
  NAND2_X1 U4560 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3588)
         );
  AND2_X1 U4561 ( .A1(n3589), .A2(n3588), .ZN(n4374) );
  MUX2_X1 U4562 ( .A(n4153), .B(n2963), .S(EBX_REG_5__SCAN_IN), .Z(n3592) );
  OAI21_X1 U4563 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5120), .A(n3592), 
        .ZN(n4459) );
  NOR2_X2 U4564 ( .A1(n4460), .A2(n4459), .ZN(n4462) );
  NAND2_X1 U4565 ( .A1(n2964), .A2(n6076), .ZN(n3594) );
  INV_X1 U4566 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U4567 ( .A1(n4167), .A2(n5773), .ZN(n3593) );
  NAND3_X1 U4568 ( .A1(n3594), .A2(n2963), .A3(n3593), .ZN(n3596) );
  NAND2_X1 U4569 ( .A1(n3580), .A2(n5773), .ZN(n3595) );
  NAND2_X1 U4570 ( .A1(n3596), .A2(n3595), .ZN(n4371) );
  NAND2_X1 U4571 ( .A1(n4462), .A2(n4371), .ZN(n4531) );
  MUX2_X1 U4572 ( .A(n4153), .B(n2963), .S(EBX_REG_7__SCAN_IN), .Z(n3597) );
  OAI21_X1 U4573 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5120), .A(n3597), 
        .ZN(n4532) );
  NAND2_X1 U4574 ( .A1(n2964), .A2(n6057), .ZN(n3601) );
  INV_X1 U4575 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U4576 ( .A1(n4167), .A2(n5756), .ZN(n3600) );
  NAND3_X1 U4577 ( .A1(n3601), .A2(n2963), .A3(n3600), .ZN(n3603) );
  NAND2_X1 U4578 ( .A1(n3580), .A2(n5756), .ZN(n3602) );
  MUX2_X1 U4579 ( .A(n4153), .B(n2963), .S(EBX_REG_9__SCAN_IN), .Z(n3606) );
  OAI21_X1 U4580 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5120), .A(n3606), 
        .ZN(n4682) );
  MUX2_X1 U4581 ( .A(n2962), .B(n2964), .S(EBX_REG_10__SCAN_IN), .Z(n3608) );
  NAND2_X1 U4582 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4583 ( .A1(n3608), .A2(n3607), .ZN(n4895) );
  NAND2_X1 U4584 ( .A1(n4896), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U4585 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3609) );
  OAI211_X1 U4586 ( .C1(n4156), .C2(EBX_REG_11__SCAN_IN), .A(n2964), .B(n3609), 
        .ZN(n3610) );
  OAI21_X1 U4587 ( .B1(n4153), .B2(EBX_REG_11__SCAN_IN), .A(n3610), .ZN(n4876)
         );
  INV_X1 U4588 ( .A(EBX_REG_13__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4589 ( .A1(n3646), .A2(n3611), .ZN(n3614) );
  NAND2_X1 U4590 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3612) );
  OAI211_X1 U4591 ( .C1(n4156), .C2(EBX_REG_13__SCAN_IN), .A(n2964), .B(n3612), 
        .ZN(n3613) );
  AND2_X1 U4592 ( .A1(n3614), .A2(n3613), .ZN(n4988) );
  MUX2_X1 U4593 ( .A(n2962), .B(n2964), .S(EBX_REG_12__SCAN_IN), .Z(n3616) );
  NAND2_X1 U4594 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4595 ( .A1(n3616), .A2(n3615), .ZN(n4989) );
  NAND2_X1 U4596 ( .A1(n4988), .A2(n4989), .ZN(n3617) );
  OR2_X2 U4597 ( .A1(n3015), .A2(n3617), .ZN(n5065) );
  INV_X1 U4598 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U4599 ( .A1(n3646), .A2(n6547), .ZN(n3620) );
  NAND2_X1 U4600 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3618) );
  OAI211_X1 U4601 ( .C1(n4156), .C2(EBX_REG_15__SCAN_IN), .A(n2964), .B(n3618), 
        .ZN(n3619) );
  AND2_X1 U4602 ( .A1(n3620), .A2(n3619), .ZN(n5044) );
  MUX2_X1 U4603 ( .A(n2963), .B(n2964), .S(EBX_REG_14__SCAN_IN), .Z(n3622) );
  NAND2_X1 U4604 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U4605 ( .A1(n3622), .A2(n3621), .ZN(n5064) );
  NAND2_X1 U4606 ( .A1(n5044), .A2(n5064), .ZN(n3623) );
  MUX2_X1 U4607 ( .A(n2963), .B(n2964), .S(EBX_REG_16__SCAN_IN), .Z(n3625) );
  NAND2_X1 U4608 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3624) );
  NAND2_X1 U4609 ( .A1(n3625), .A2(n3624), .ZN(n5080) );
  INV_X1 U4610 ( .A(EBX_REG_17__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4611 ( .A1(n3646), .A2(n3626), .ZN(n3629) );
  NAND2_X1 U4612 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3627) );
  OAI211_X1 U4613 ( .C1(n4156), .C2(EBX_REG_17__SCAN_IN), .A(n2964), .B(n3627), 
        .ZN(n3628) );
  AND2_X1 U4614 ( .A1(n3629), .A2(n3628), .ZN(n5079) );
  AND2_X1 U4615 ( .A1(n5080), .A2(n5079), .ZN(n3630) );
  AND2_X2 U4616 ( .A1(n5081), .A2(n3630), .ZN(n5078) );
  NAND2_X1 U4617 ( .A1(n2964), .A2(n3631), .ZN(n3633) );
  INV_X1 U4618 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4619 ( .A1(n4167), .A2(n3634), .ZN(n3632) );
  NAND3_X1 U4620 ( .A1(n3633), .A2(n2963), .A3(n3632), .ZN(n3636) );
  NAND2_X1 U4621 ( .A1(n3580), .A2(n3634), .ZN(n3635) );
  NAND2_X1 U4622 ( .A1(n3636), .A2(n3635), .ZN(n5167) );
  AND2_X2 U4623 ( .A1(n5078), .A2(n5167), .ZN(n5257) );
  AND2_X1 U4624 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3637)
         );
  AOI21_X1 U4625 ( .B1(n5120), .B2(EBX_REG_18__SCAN_IN), .A(n3637), .ZN(n5258)
         );
  INV_X1 U4626 ( .A(n5258), .ZN(n3638) );
  AND2_X1 U4627 ( .A1(n3638), .A2(n2962), .ZN(n5165) );
  AND2_X1 U4628 ( .A1(n5258), .A2(n3580), .ZN(n5166) );
  OR2_X1 U4629 ( .A1(n5120), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3641)
         );
  INV_X1 U4630 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4631 ( .A1(n4167), .A2(n3639), .ZN(n3640) );
  NAND2_X1 U4632 ( .A1(n3641), .A2(n3640), .ZN(n5259) );
  MUX2_X1 U4633 ( .A(n5165), .B(n5166), .S(n5259), .Z(n3642) );
  NAND2_X1 U4634 ( .A1(n5257), .A2(n3642), .ZN(n5250) );
  MUX2_X1 U4635 ( .A(n4153), .B(n2963), .S(EBX_REG_21__SCAN_IN), .Z(n3643) );
  OAI21_X1 U4636 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5120), .A(n3643), 
        .ZN(n5249) );
  OR2_X2 U4637 ( .A1(n5250), .A2(n5249), .ZN(n5247) );
  MUX2_X1 U4638 ( .A(n2962), .B(n2964), .S(EBX_REG_22__SCAN_IN), .Z(n3645) );
  NAND2_X1 U4639 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3644) );
  INV_X1 U4640 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U4641 ( .A1(n3646), .A2(n6485), .ZN(n3649) );
  NAND2_X1 U4642 ( .A1(n2963), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3647) );
  OAI211_X1 U4643 ( .C1(n4156), .C2(EBX_REG_23__SCAN_IN), .A(n2964), .B(n3647), 
        .ZN(n3648) );
  AND2_X1 U4644 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  NOR2_X1 U4645 ( .A1(n5159), .A2(n3650), .ZN(n3651) );
  OR2_X1 U4646 ( .A1(n4228), .A2(n3651), .ZN(n5241) );
  INV_X1 U4647 ( .A(n5241), .ZN(n5573) );
  INV_X1 U4648 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3652) );
  NOR2_X1 U4649 ( .A1(n6071), .A2(n3652), .ZN(n4200) );
  NAND2_X1 U4650 ( .A1(n2961), .A2(n3560), .ZN(n4278) );
  OR2_X1 U4651 ( .A1(n4278), .A2(n3653), .ZN(n3654) );
  AND2_X1 U4652 ( .A1(n3655), .A2(n3654), .ZN(n4406) );
  INV_X1 U4653 ( .A(n3656), .ZN(n3657) );
  INV_X1 U4654 ( .A(n4388), .ZN(n4414) );
  AOI21_X1 U4655 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6109) );
  NAND2_X1 U4656 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6094) );
  NOR2_X1 U4657 ( .A1(n6109), .A2(n6094), .ZN(n6078) );
  NAND3_X1 U4658 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6078), .ZN(n4891) );
  NAND2_X1 U4659 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U4660 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4889) );
  NOR2_X1 U4661 ( .A1(n4890), .A2(n4889), .ZN(n3668) );
  INV_X1 U4662 ( .A(n3668), .ZN(n4974) );
  NOR2_X1 U4663 ( .A1(n4891), .A2(n4974), .ZN(n4971) );
  INV_X1 U4664 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5451) );
  INV_X1 U4665 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5465) );
  NAND3_X1 U4666 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5466) );
  NOR2_X1 U4667 ( .A1(n5465), .A2(n5466), .ZN(n5463) );
  NAND3_X1 U4668 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5463), .ZN(n5426) );
  NOR2_X1 U4669 ( .A1(n5451), .A2(n5426), .ZN(n5420) );
  NAND2_X1 U4670 ( .A1(n4971), .A2(n5420), .ZN(n3676) );
  OAI21_X1 U4671 ( .B1(n3658), .B2(n4491), .A(n2964), .ZN(n3659) );
  OR2_X1 U4672 ( .A1(n3660), .A2(n3659), .ZN(n4386) );
  INV_X1 U4673 ( .A(n3661), .ZN(n4384) );
  NAND2_X1 U4674 ( .A1(n3528), .A2(n3580), .ZN(n4383) );
  NAND3_X1 U4675 ( .A1(n4384), .A2(n4417), .A3(n4383), .ZN(n3662) );
  NOR2_X1 U4676 ( .A1(n4386), .A2(n3662), .ZN(n3663) );
  NAND2_X1 U4677 ( .A1(n3665), .A2(n6071), .ZN(n6129) );
  OAI21_X1 U4678 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5056), .A(n6129), 
        .ZN(n6066) );
  AOI21_X1 U4679 ( .B1(n6107), .B2(n3676), .A(n6066), .ZN(n5427) );
  AND2_X1 U4680 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5422) );
  AND2_X1 U4681 ( .A1(n5422), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3678)
         );
  INV_X1 U4682 ( .A(n3678), .ZN(n3669) );
  NAND2_X1 U4683 ( .A1(n6107), .A2(n3669), .ZN(n3664) );
  AND2_X1 U4684 ( .A1(n5427), .A2(n3664), .ZN(n3672) );
  NAND2_X1 U4685 ( .A1(n4286), .A2(n3560), .ZN(n5092) );
  NAND2_X1 U4686 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4687 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6080) );
  NOR3_X1 U4688 ( .A1(n6094), .A2(n3667), .A3(n6080), .ZN(n4893) );
  NAND2_X1 U4689 ( .A1(n3668), .A2(n4893), .ZN(n4970) );
  NOR2_X1 U4690 ( .A1(n5426), .A2(n4970), .ZN(n5428) );
  NAND2_X1 U4691 ( .A1(n5428), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3677) );
  NOR2_X1 U4692 ( .A1(n3677), .A2(n3669), .ZN(n3670) );
  OR2_X1 U4693 ( .A1(n6068), .A2(n3670), .ZN(n3671) );
  NAND2_X1 U4694 ( .A1(n6068), .A2(n4888), .ZN(n6070) );
  INV_X1 U4695 ( .A(n5399), .ZN(n3673) );
  NAND2_X1 U4696 ( .A1(n6070), .A2(n3673), .ZN(n3674) );
  AND2_X1 U4697 ( .A1(n5412), .A2(n3674), .ZN(n4237) );
  NOR2_X1 U4698 ( .A1(n4237), .A2(n4206), .ZN(n3675) );
  AOI211_X1 U4699 ( .C1(n6106), .C2(n5573), .A(n4200), .B(n3675), .ZN(n3680)
         );
  NOR2_X1 U4700 ( .A1(n5059), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6121)
         );
  OAI22_X1 U4701 ( .A1(n6112), .A2(n3677), .B1(n3676), .B2(n4888), .ZN(n5441)
         );
  NAND3_X1 U4702 ( .A1(n5414), .A2(n5399), .A3(n4206), .ZN(n3679) );
  NAND2_X1 U4703 ( .A1(n3682), .A2(n3681), .ZN(U2995) );
  INV_X1 U4704 ( .A(n4515), .ZN(n3683) );
  NAND2_X1 U4705 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6326), .ZN(n3838) );
  OAI21_X1 U4706 ( .B1(n3687), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3758), 
        .ZN(n5987) );
  AOI22_X1 U4707 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4263), .B1(n4121), 
        .B2(n5987), .ZN(n3688) );
  AOI21_X1 U4708 ( .B1(n3697), .B2(n5791), .A(n3733), .ZN(n6011) );
  NOR2_X1 U4709 ( .A1(n6011), .A2(n4092), .ZN(n3695) );
  AOI22_X1 U4710 ( .A1(n4264), .A2(EAX_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6326), .ZN(n3693) );
  NAND2_X1 U4711 ( .A1(n3225), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3725) );
  INV_X1 U4712 ( .A(n3725), .ZN(n3716) );
  NAND2_X1 U4713 ( .A1(n3716), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3692) );
  AOI21_X1 U4714 ( .B1(n3693), .B2(n3692), .A(n4121), .ZN(n3694) );
  AOI211_X1 U4715 ( .C1(n3696), .C2(n3852), .A(n3695), .B(n3694), .ZN(n4378)
         );
  OAI21_X1 U4716 ( .B1(n3698), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3697), 
        .ZN(n6024) );
  AOI22_X1 U4717 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4263), .B1(n4121), 
        .B2(n6024), .ZN(n3700) );
  INV_X1 U4718 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4476) );
  OR2_X1 U4719 ( .A1(n4124), .A2(n4476), .ZN(n3699) );
  OAI211_X1 U4720 ( .C1(n3725), .C2(n4415), .A(n3700), .B(n3699), .ZN(n3701)
         );
  NOR2_X1 U4721 ( .A1(n4378), .A2(n4474), .ZN(n3731) );
  AOI21_X1 U4722 ( .B1(n4446), .B2(n3852), .A(n4263), .ZN(n3726) );
  NAND2_X1 U4723 ( .A1(n4447), .A2(n3852), .ZN(n3708) );
  NAND2_X1 U4724 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6326), .ZN(n3705)
         );
  INV_X1 U4725 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3703) );
  OR2_X1 U4726 ( .A1(n4124), .A2(n3703), .ZN(n3704) );
  OAI211_X1 U4727 ( .C1(n3725), .C2(n3471), .A(n3705), .B(n3704), .ZN(n3706)
         );
  INV_X1 U4728 ( .A(n3706), .ZN(n3707) );
  AOI21_X1 U4729 ( .B1(n3709), .B2(n2960), .A(n6326), .ZN(n4313) );
  INV_X1 U4730 ( .A(n3852), .ZN(n3713) );
  OR2_X1 U4731 ( .A1(n3712), .A2(n3713), .ZN(n3718) );
  INV_X1 U4732 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3714) );
  INV_X1 U4733 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5833) );
  OAI22_X1 U4734 ( .A1(n4124), .A2(n3714), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5833), .ZN(n3715) );
  AOI21_X1 U4735 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3716), .A(n3715), 
        .ZN(n3717) );
  NAND2_X1 U4736 ( .A1(n3718), .A2(n3717), .ZN(n4312) );
  NAND2_X1 U4737 ( .A1(n4313), .A2(n4312), .ZN(n4311) );
  INV_X1 U4738 ( .A(n4312), .ZN(n3719) );
  NAND2_X1 U4739 ( .A1(n3719), .A2(n4121), .ZN(n3720) );
  NAND2_X1 U4740 ( .A1(n4311), .A2(n3720), .ZN(n4318) );
  OAI21_X1 U4741 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3721), .ZN(n6034) );
  AOI22_X1 U4742 ( .A1(n6034), .A2(n4121), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n4263), .ZN(n3724) );
  INV_X1 U4743 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3722) );
  OR2_X1 U4744 ( .A1(n4124), .A2(n3722), .ZN(n3723) );
  OAI211_X1 U4745 ( .C1(n3725), .C2(n5106), .A(n3724), .B(n3723), .ZN(n4356)
         );
  NAND2_X1 U4746 ( .A1(n4357), .A2(n4356), .ZN(n3730) );
  INV_X1 U4747 ( .A(n3726), .ZN(n3728) );
  INV_X1 U4748 ( .A(n4321), .ZN(n3727) );
  NAND2_X1 U4749 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  AND2_X2 U4750 ( .A1(n3731), .A2(n4355), .ZN(n4463) );
  NAND2_X1 U4751 ( .A1(n3732), .A2(n3852), .ZN(n3738) );
  INV_X1 U4752 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3735) );
  OAI21_X1 U4753 ( .B1(n3733), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3739), 
        .ZN(n6005) );
  AOI22_X1 U4754 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4263), .B1(n4121), 
        .B2(n6005), .ZN(n3734) );
  OAI21_X1 U4755 ( .B1(n4124), .B2(n3735), .A(n3734), .ZN(n3736) );
  INV_X1 U4756 ( .A(n3736), .ZN(n3737) );
  NAND2_X1 U4757 ( .A1(n3738), .A2(n3737), .ZN(n4464) );
  XNOR2_X1 U4758 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3739), .ZN(n5993) );
  NOR2_X1 U4759 ( .A1(n5993), .A2(n4092), .ZN(n3742) );
  AOI22_X1 U4760 ( .A1(n4264), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6326), .ZN(n3740) );
  NOR2_X1 U4761 ( .A1(n3740), .A2(n4121), .ZN(n3741) );
  INV_X1 U4762 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4763 ( .A1(n3281), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4764 ( .A1(n4104), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4765 ( .A1(n4396), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4766 ( .A1(n4105), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3744) );
  NAND4_X1 U4767 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3753)
         );
  AOI22_X1 U4768 ( .A1(n4018), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4769 ( .A1(n4095), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4770 ( .A1(n3282), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4771 ( .A1(n4036), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4772 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OAI21_X1 U4773 ( .B1(n3753), .B2(n3752), .A(n3852), .ZN(n3754) );
  OAI21_X1 U4774 ( .B1(n3838), .B2(n3755), .A(n3754), .ZN(n3757) );
  XNOR2_X1 U4775 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3758), .ZN(n5975) );
  NOR2_X1 U4776 ( .A1(n5975), .A2(n4092), .ZN(n3756) );
  AOI211_X1 U4777 ( .C1(n4264), .C2(EAX_REG_8__SCAN_IN), .A(n3757), .B(n3756), 
        .ZN(n4469) );
  XNOR2_X1 U4778 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3784), .ZN(n5968) );
  AOI22_X1 U4779 ( .A1(n4264), .A2(EAX_REG_9__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n4263), .ZN(n3771) );
  AOI22_X1 U4780 ( .A1(n4018), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4781 ( .A1(n3281), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4036), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4782 ( .A1(n4104), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4783 ( .A1(n3282), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4784 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4785 ( .A1(n4095), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4786 ( .A1(n4396), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4787 ( .A1(n4097), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4788 ( .A1(n4105), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4789 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  OAI21_X1 U4790 ( .B1(n3769), .B2(n3768), .A(n3852), .ZN(n3770) );
  OAI211_X1 U4791 ( .C1(n5968), .C2(n4092), .A(n3771), .B(n3770), .ZN(n4610)
         );
  INV_X1 U4792 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4884) );
  AOI22_X1 U4793 ( .A1(n4094), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4794 ( .A1(n3276), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4795 ( .A1(n3281), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4796 ( .A1(n4097), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4797 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3781)
         );
  AOI22_X1 U4798 ( .A1(n4018), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4799 ( .A1(n4036), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4800 ( .A1(n3282), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4801 ( .A1(n4095), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4802 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  OAI21_X1 U4803 ( .B1(n3781), .B2(n3780), .A(n3852), .ZN(n3782) );
  OAI21_X1 U4804 ( .B1(n3838), .B2(n4884), .A(n3782), .ZN(n3786) );
  XOR2_X1 U4805 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3787), .Z(n5740) );
  NOR2_X1 U4806 ( .A1(n5740), .A2(n4092), .ZN(n3785) );
  AOI211_X1 U4807 ( .C1(n4264), .C2(EAX_REG_10__SCAN_IN), .A(n3786), .B(n3785), 
        .ZN(n4872) );
  XNOR2_X1 U4808 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3811), .ZN(n5958)
         );
  AOI22_X1 U4809 ( .A1(n4264), .A2(EAX_REG_11__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n4263), .ZN(n3799) );
  AOI22_X1 U4810 ( .A1(n4018), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4811 ( .A1(n4104), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4812 ( .A1(n3282), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4813 ( .A1(n3281), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4814 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4815 ( .A1(n3276), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4816 ( .A1(n4095), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4817 ( .A1(n4097), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4818 ( .A1(n4036), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4819 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  OAI21_X1 U4820 ( .B1(n3797), .B2(n3796), .A(n3852), .ZN(n3798) );
  OAI211_X1 U4821 ( .C1(n5958), .C2(n4092), .A(n3799), .B(n3798), .ZN(n4875)
         );
  INV_X1 U4822 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U4823 ( .A1(n4018), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4824 ( .A1(n4396), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4825 ( .A1(n4097), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4826 ( .A1(n3282), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4827 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3809)
         );
  AOI22_X1 U4828 ( .A1(n4104), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4829 ( .A1(n3281), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4830 ( .A1(n4095), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4831 ( .A1(n4036), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4832 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  OAI21_X1 U4833 ( .B1(n3809), .B2(n3808), .A(n3852), .ZN(n3810) );
  OAI21_X1 U4834 ( .B1(n3838), .B2(n4980), .A(n3810), .ZN(n3813) );
  XOR2_X1 U4835 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3814), .Z(n5724) );
  NOR2_X1 U4836 ( .A1(n5724), .A2(n4092), .ZN(n3812) );
  AOI211_X1 U4837 ( .C1(n4264), .C2(EAX_REG_12__SCAN_IN), .A(n3813), .B(n3812), 
        .ZN(n4959) );
  XNOR2_X1 U4838 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3839), .ZN(n5715)
         );
  AOI22_X1 U4839 ( .A1(n4264), .A2(EAX_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4263), .ZN(n3826) );
  AOI22_X1 U4840 ( .A1(n3276), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4841 ( .A1(n3281), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4842 ( .A1(n4104), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4843 ( .A1(n4097), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4844 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3824)
         );
  AOI22_X1 U4845 ( .A1(n4018), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4846 ( .A1(n4095), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4847 ( .A1(n3282), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4848 ( .A1(n4036), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4849 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3823)
         );
  OAI21_X1 U4850 ( .B1(n3824), .B2(n3823), .A(n3852), .ZN(n3825) );
  OAI211_X1 U4851 ( .C1(n5715), .C2(n4092), .A(n3826), .B(n3825), .ZN(n4987)
         );
  INV_X1 U4852 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5052) );
  AOI22_X1 U4853 ( .A1(n4094), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4854 ( .A1(n4095), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4855 ( .A1(n4105), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4856 ( .A1(n4036), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3827) );
  NAND4_X1 U4857 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3827), .ZN(n3836)
         );
  AOI22_X1 U4858 ( .A1(n4018), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4859 ( .A1(n4104), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4860 ( .A1(n3281), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4861 ( .A1(n4097), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4862 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3835)
         );
  OAI21_X1 U4863 ( .B1(n3836), .B2(n3835), .A(n3852), .ZN(n3837) );
  OAI21_X1 U4864 ( .B1(n3838), .B2(n5052), .A(n3837), .ZN(n3841) );
  XOR2_X1 U4865 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3842), .Z(n5704) );
  NOR2_X1 U4866 ( .A1(n5704), .A2(n4092), .ZN(n3840) );
  AOI211_X1 U4867 ( .C1(n4264), .C2(EAX_REG_14__SCAN_IN), .A(n3841), .B(n3840), 
        .ZN(n5036) );
  AOI21_X1 U4868 ( .B1(n6536), .B2(n3843), .A(n3869), .ZN(n5697) );
  AOI22_X1 U4869 ( .A1(n4264), .A2(EAX_REG_15__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n4263), .ZN(n3856) );
  AOI22_X1 U4870 ( .A1(n4018), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4871 ( .A1(n3325), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4872 ( .A1(n4396), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4873 ( .A1(n4105), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3844) );
  NAND4_X1 U4874 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3854)
         );
  AOI22_X1 U4875 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n4094), .B1(n3276), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4876 ( .A1(n4095), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4877 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n4097), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4878 ( .A1(n4036), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4879 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3853)
         );
  OAI21_X1 U4880 ( .B1(n3854), .B2(n3853), .A(n3852), .ZN(n3855) );
  OAI211_X1 U4881 ( .C1(n5697), .C2(n4092), .A(n3856), .B(n3855), .ZN(n5041)
         );
  NAND2_X1 U4882 ( .A1(n5035), .A2(n5041), .ZN(n5039) );
  AOI22_X1 U4883 ( .A1(n4018), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4884 ( .A1(n4095), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4885 ( .A1(n3351), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4886 ( .A1(n4106), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4887 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3868)
         );
  AOI22_X1 U4888 ( .A1(n3276), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4889 ( .A1(n4036), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4890 ( .A1(n3325), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4891 ( .A1(n4097), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4892 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3867)
         );
  XOR2_X1 U4893 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3869), .Z(n5326) );
  AOI22_X1 U4894 ( .A1(n4264), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n4263), .ZN(n3865) );
  OAI21_X1 U4895 ( .B1(n5326), .B2(n4092), .A(n3865), .ZN(n3866) );
  AOI221_X1 U4896 ( .B1(n3868), .B2(n4086), .C1(n3867), .C2(n4086), .A(n3866), 
        .ZN(n5072) );
  XNOR2_X1 U4897 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n3883), .ZN(n5636)
         );
  AOI22_X1 U4898 ( .A1(n4018), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4899 ( .A1(n3276), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4900 ( .A1(n4095), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4901 ( .A1(n4396), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4902 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4903 ( .A1(n3281), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4904 ( .A1(n4097), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4905 ( .A1(n3282), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4906 ( .A1(n4036), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4907 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  OR2_X1 U4908 ( .A1(n3879), .A2(n3878), .ZN(n3880) );
  AOI22_X1 U4909 ( .A1(n4086), .A2(n3880), .B1(n4264), .B2(EAX_REG_17__SCAN_IN), .ZN(n3882) );
  OAI21_X1 U4910 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4534), .A(n6326), 
        .ZN(n3881) );
  AOI22_X1 U4911 ( .A1(n4121), .A2(n5636), .B1(n3882), .B2(n3881), .ZN(n5077)
         );
  OAI21_X1 U4912 ( .B1(n3884), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n3910), 
        .ZN(n5635) );
  INV_X1 U4913 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6488) );
  AOI22_X1 U4914 ( .A1(n4094), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4915 ( .A1(n3282), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4916 ( .A1(n4105), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4917 ( .A1(n4036), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4918 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3894)
         );
  AOI22_X1 U4919 ( .A1(n4018), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4920 ( .A1(n3281), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4921 ( .A1(n4095), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4922 ( .A1(n4396), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4923 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  OAI21_X1 U4924 ( .B1(n3894), .B2(n3893), .A(n4086), .ZN(n3896) );
  OAI21_X1 U4925 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4534), .A(n6326), 
        .ZN(n3895) );
  OAI211_X1 U4926 ( .C1(n6488), .C2(n4124), .A(n3896), .B(n3895), .ZN(n3897)
         );
  OAI21_X1 U4927 ( .B1(n5635), .B2(n4092), .A(n3897), .ZN(n5179) );
  XNOR2_X1 U4928 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3910), .ZN(n5317)
         );
  AOI22_X1 U4929 ( .A1(n4264), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6326), .ZN(n3909) );
  AOI22_X1 U4930 ( .A1(n4104), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4931 ( .A1(n3325), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4932 ( .A1(n3282), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4933 ( .A1(n4396), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4934 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3907)
         );
  AOI22_X1 U4935 ( .A1(n4018), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4936 ( .A1(n4095), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4937 ( .A1(n4036), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4938 ( .A1(n4097), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4939 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  AOI221_X1 U4940 ( .B1(n3907), .B2(n4086), .C1(n3906), .C2(n4086), .A(n4121), 
        .ZN(n3908) );
  AOI22_X1 U4941 ( .A1(n4121), .A2(n5317), .B1(n3909), .B2(n3908), .ZN(n5176)
         );
  OAI21_X1 U4942 ( .B1(n3911), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3940), 
        .ZN(n5631) );
  AOI22_X1 U4943 ( .A1(n4264), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6326), .ZN(n3923) );
  AOI22_X1 U4944 ( .A1(n4018), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4945 ( .A1(n3325), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4946 ( .A1(n3276), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4947 ( .A1(n4036), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4948 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3921)
         );
  AOI22_X1 U4949 ( .A1(n4104), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4950 ( .A1(n4095), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4951 ( .A1(n3282), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4952 ( .A1(n4105), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4953 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  OAI21_X1 U4954 ( .B1(n3921), .B2(n3920), .A(n4086), .ZN(n3922) );
  NAND3_X1 U4955 ( .A1(n4092), .A2(n3923), .A3(n3922), .ZN(n3924) );
  OAI21_X1 U4956 ( .B1(n4092), .B2(n5631), .A(n3924), .ZN(n5255) );
  INV_X1 U4957 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U4958 ( .A1(n4018), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4959 ( .A1(n3276), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4095), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4960 ( .A1(n4098), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4036), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4961 ( .A1(n4097), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4962 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3934)
         );
  AOI22_X1 U4963 ( .A1(n4104), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4964 ( .A1(n4396), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4965 ( .A1(n3325), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4966 ( .A1(n4106), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4967 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3933)
         );
  AOI221_X1 U4968 ( .B1(n3934), .B2(n4086), .C1(n3933), .C2(n4086), .A(n4121), 
        .ZN(n3935) );
  INV_X1 U4969 ( .A(n3935), .ZN(n3936) );
  AOI21_X1 U4970 ( .B1(n6326), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3936), 
        .ZN(n3937) );
  OAI21_X1 U4971 ( .B1(n4124), .B2(n4299), .A(n3937), .ZN(n3939) );
  XNOR2_X1 U4972 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3940), .ZN(n5580)
         );
  NAND2_X1 U4973 ( .A1(n4121), .A2(n5580), .ZN(n3938) );
  INV_X1 U4974 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5308) );
  OR2_X1 U4975 ( .A1(n3941), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3942)
         );
  NAND2_X1 U4976 ( .A1(n3983), .A2(n3942), .ZN(n5301) );
  INV_X1 U4977 ( .A(n5301), .ZN(n3957) );
  INV_X1 U4978 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4979 ( .A1(n4018), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4980 ( .A1(n4095), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4981 ( .A1(n4396), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4982 ( .A1(n4106), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4983 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3952)
         );
  AOI22_X1 U4984 ( .A1(n4104), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4985 ( .A1(n3351), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4036), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4986 ( .A1(n4105), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4987 ( .A1(n3325), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4988 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  OAI21_X1 U4989 ( .B1(n3952), .B2(n3951), .A(n4086), .ZN(n3953) );
  OAI211_X1 U4990 ( .C1(n3954), .C2(STATE2_REG_2__SCAN_IN), .A(n3953), .B(
        n4092), .ZN(n3955) );
  AOI21_X1 U4991 ( .B1(n4264), .B2(EAX_REG_22__SCAN_IN), .A(n3955), .ZN(n3956)
         );
  AOI21_X1 U4992 ( .B1(n3957), .B2(n4121), .A(n3956), .ZN(n5153) );
  XNOR2_X1 U4993 ( .A(n3983), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5571)
         );
  AOI22_X1 U4994 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4018), .B1(n3276), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4995 ( .A1(n3325), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4996 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4036), .B1(n4396), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4997 ( .A1(n4104), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4998 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3967)
         );
  AOI22_X1 U4999 ( .A1(n4094), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U5000 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3282), .B1(n4106), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U5001 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n4105), .B1(n4096), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U5002 ( .A1(n4095), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U5003 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3966)
         );
  NOR2_X1 U5004 ( .A1(n3967), .A2(n3966), .ZN(n3984) );
  AOI22_X1 U5005 ( .A1(n4018), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U5006 ( .A1(n4104), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U5007 ( .A1(n4105), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U5008 ( .A1(n4097), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3968) );
  NAND4_X1 U5009 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3977)
         );
  AOI22_X1 U5010 ( .A1(n4095), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5011 ( .A1(n4036), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5012 ( .A1(n3282), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5013 ( .A1(n3281), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U5014 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  NOR2_X1 U5015 ( .A1(n3977), .A2(n3976), .ZN(n3985) );
  XOR2_X1 U5016 ( .A(n3984), .B(n3985), .Z(n3981) );
  INV_X1 U5017 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3979) );
  AOI21_X1 U5018 ( .B1(n6326), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4121), 
        .ZN(n3978) );
  OAI21_X1 U5019 ( .B1(n4124), .B2(n3979), .A(n3978), .ZN(n3980) );
  AOI21_X1 U5020 ( .B1(n4086), .B2(n3981), .A(n3980), .ZN(n3982) );
  AOI21_X1 U5021 ( .B1(n5571), .B2(n4121), .A(n3982), .ZN(n4192) );
  INV_X1 U5022 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5569) );
  XOR2_X1 U5023 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .B(n4000), .Z(n5146) );
  NOR2_X1 U5024 ( .A1(n3985), .A2(n3984), .ZN(n4012) );
  AOI22_X1 U5025 ( .A1(n4018), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U5026 ( .A1(n3276), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U5027 ( .A1(n4095), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U5028 ( .A1(n4396), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U5029 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3995)
         );
  AOI22_X1 U5030 ( .A1(n3281), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5031 ( .A1(n4097), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U5032 ( .A1(n3282), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5033 ( .A1(n4036), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U5034 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  OAI21_X1 U5035 ( .B1(n4012), .B2(n4011), .A(n4086), .ZN(n3996) );
  AOI21_X1 U5036 ( .B1(n4012), .B2(n4011), .A(n3996), .ZN(n3999) );
  AOI22_X1 U5037 ( .A1(n4264), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4263), .ZN(n3997) );
  INV_X1 U5038 ( .A(n3997), .ZN(n3998) );
  XNOR2_X1 U5039 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4016), .ZN(n5622)
         );
  AOI22_X1 U5040 ( .A1(n4264), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6326), .ZN(n4015) );
  AOI22_X1 U5041 ( .A1(n4018), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5042 ( .A1(n3276), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5043 ( .A1(n4095), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5044 ( .A1(n4396), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U5045 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U5046 ( .A1(n3325), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5047 ( .A1(n4097), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5048 ( .A1(n3282), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U5049 ( .A1(n4036), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U5050 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  NOR2_X1 U5051 ( .A1(n4010), .A2(n4009), .ZN(n4030) );
  NAND2_X1 U5052 ( .A1(n4012), .A2(n4011), .ZN(n4029) );
  XOR2_X1 U5053 ( .A(n4030), .B(n4029), .Z(n4013) );
  AOI21_X1 U5054 ( .B1(n4013), .B2(n4086), .A(n4121), .ZN(n4014) );
  AOI22_X1 U5055 ( .A1(n4121), .A2(n5622), .B1(n4015), .B2(n4014), .ZN(n5137)
         );
  NAND2_X1 U5056 ( .A1(n5136), .A2(n5137), .ZN(n5135) );
  INV_X1 U5057 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5140) );
  OAI21_X1 U5058 ( .B1(n4017), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n4052), 
        .ZN(n5621) );
  AOI22_X1 U5059 ( .A1(n4018), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5060 ( .A1(n3276), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5061 ( .A1(n4095), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5062 ( .A1(n4396), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U5063 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4028)
         );
  AOI22_X1 U5064 ( .A1(n3325), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5065 ( .A1(n4036), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5066 ( .A1(n4097), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5067 ( .A1(n3282), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U5068 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  OR2_X1 U5069 ( .A1(n4028), .A2(n4027), .ZN(n4034) );
  NOR2_X1 U5070 ( .A1(n4030), .A2(n4029), .ZN(n4035) );
  XNOR2_X1 U5071 ( .A(n4034), .B(n4035), .ZN(n4032) );
  INV_X1 U5072 ( .A(n4086), .ZN(n4118) );
  AOI22_X1 U5073 ( .A1(n4264), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6326), .ZN(n4031) );
  OAI21_X1 U5074 ( .B1(n4032), .B2(n4118), .A(n4031), .ZN(n4033) );
  AOI22_X1 U5075 ( .A1(n4121), .A2(n5621), .B1(n4033), .B2(n4092), .ZN(n5229)
         );
  XNOR2_X1 U5076 ( .A(n4052), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5552)
         );
  NAND2_X1 U5077 ( .A1(n4035), .A2(n4034), .ZN(n4065) );
  AOI22_X1 U5078 ( .A1(n4018), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5079 ( .A1(n3282), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5080 ( .A1(n4095), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4075), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5081 ( .A1(n4036), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U5082 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4046)
         );
  AOI22_X1 U5083 ( .A1(n3276), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5084 ( .A1(n4104), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5085 ( .A1(n3281), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5086 ( .A1(n4097), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5087 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4045)
         );
  NOR2_X1 U5088 ( .A1(n4046), .A2(n4045), .ZN(n4066) );
  XOR2_X1 U5089 ( .A(n4065), .B(n4066), .Z(n4050) );
  INV_X1 U5090 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4048) );
  AOI21_X1 U5091 ( .B1(n6326), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4121), 
        .ZN(n4047) );
  OAI21_X1 U5092 ( .B1(n4124), .B2(n4048), .A(n4047), .ZN(n4049) );
  AOI21_X1 U5093 ( .B1(n4050), .B2(n4086), .A(n4049), .ZN(n4051) );
  AOI21_X1 U5094 ( .B1(n5552), .B2(n4121), .A(n4051), .ZN(n5224) );
  INV_X1 U5095 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5288) );
  OR2_X1 U5096 ( .A1(n4053), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4054)
         );
  NAND2_X1 U5097 ( .A1(n4120), .A2(n4054), .ZN(n5540) );
  AOI22_X1 U5098 ( .A1(n4018), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5099 ( .A1(n3276), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5100 ( .A1(n4095), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5101 ( .A1(n4396), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5102 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U5103 ( .A1(n3281), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5104 ( .A1(n4036), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5105 ( .A1(n4097), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5106 ( .A1(n3282), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5107 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  OR2_X1 U5108 ( .A1(n4064), .A2(n4063), .ZN(n4073) );
  NOR2_X1 U5109 ( .A1(n4066), .A2(n4065), .ZN(n4074) );
  XNOR2_X1 U5110 ( .A(n4073), .B(n4074), .ZN(n4070) );
  INV_X1 U5111 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4067) );
  OAI21_X1 U5112 ( .B1(n4067), .B2(STATE2_REG_2__SCAN_IN), .A(n4092), .ZN(
        n4068) );
  AOI21_X1 U5113 ( .B1(n4264), .B2(EAX_REG_28__SCAN_IN), .A(n4068), .ZN(n4069)
         );
  OAI21_X1 U5114 ( .B1(n4070), .B2(n4118), .A(n4069), .ZN(n4071) );
  NAND2_X1 U5115 ( .A1(n4072), .A2(n4071), .ZN(n5215) );
  XNOR2_X1 U5116 ( .A(n4120), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5530)
         );
  INV_X1 U5117 ( .A(n5530), .ZN(n4257) );
  INV_X1 U5118 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4090) );
  NAND2_X1 U5119 ( .A1(n4074), .A2(n4073), .ZN(n4113) );
  AOI22_X1 U5120 ( .A1(n4094), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5121 ( .A1(n4095), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5122 ( .A1(n3325), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5123 ( .A1(n4075), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4076) );
  NAND4_X1 U5124 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4085)
         );
  AOI22_X1 U5125 ( .A1(n4018), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4104), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5126 ( .A1(n4036), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5127 ( .A1(n4097), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5128 ( .A1(n3282), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U5129 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4084)
         );
  NOR2_X1 U5130 ( .A1(n4085), .A2(n4084), .ZN(n4114) );
  XOR2_X1 U5131 ( .A(n4113), .B(n4114), .Z(n4087) );
  NAND2_X1 U5132 ( .A1(n4087), .A2(n4086), .ZN(n4089) );
  AOI21_X1 U5133 ( .B1(n6326), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4121), 
        .ZN(n4088) );
  OAI211_X1 U5134 ( .C1(n4124), .C2(n4090), .A(n4089), .B(n4088), .ZN(n4091)
         );
  OAI21_X1 U5135 ( .B1(n4257), .B2(n4092), .A(n4091), .ZN(n4255) );
  AOI22_X1 U5136 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4018), .B1(n4094), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5137 ( .A1(n4095), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3351), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5138 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4097), .B1(n4096), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5139 ( .A1(n3281), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4098), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5140 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4112)
         );
  AOI22_X1 U5141 ( .A1(n3276), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4103), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5142 ( .A1(n4104), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4396), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5143 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n4036), .B1(n4105), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5144 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n3282), .B1(n4106), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5145 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4111)
         );
  NOR2_X1 U5146 ( .A1(n4112), .A2(n4111), .ZN(n4116) );
  NOR2_X1 U5147 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  XOR2_X1 U5148 ( .A(n4116), .B(n4115), .Z(n4119) );
  AOI22_X1 U5149 ( .A1(n4264), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6326), .ZN(n4117) );
  OAI21_X1 U5150 ( .B1(n4119), .B2(n4118), .A(n4117), .ZN(n4122) );
  INV_X1 U5151 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5532) );
  XOR2_X1 U5152 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4137), .Z(n4213) );
  MUX2_X1 U5153 ( .A(n4122), .B(n4213), .S(n4121), .Z(n4261) );
  NAND2_X1 U5154 ( .A1(n6329), .A2(n4403), .ZN(n4126) );
  NAND3_X1 U5155 ( .A1(n4123), .A2(n3683), .A3(n6513), .ZN(n4125) );
  OAI22_X1 U5156 ( .A1(n5664), .A2(n4126), .B1(n4382), .B2(n4324), .ZN(n4127)
         );
  AOI21_X1 U5157 ( .B1(n4305), .B2(n4411), .A(n4127), .ZN(n4129) );
  AND2_X1 U5158 ( .A1(n3685), .A2(n3156), .ZN(n4466) );
  NAND2_X1 U5159 ( .A1(n5864), .A2(DATAI_30_), .ZN(n4134) );
  NOR3_X1 U5160 ( .A1(n5861), .A2(n5108), .A3(n4131), .ZN(n4132) );
  AOI22_X1 U5161 ( .A1(n5867), .A2(DATAI_14_), .B1(n5861), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4133) );
  OAI21_X1 U5162 ( .B1(n4215), .B2(n5858), .A(n4135), .ZN(U2861) );
  INV_X1 U5163 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4136) );
  INV_X1 U5164 ( .A(n4285), .ZN(n4141) );
  NAND2_X1 U5165 ( .A1(n4282), .A2(n6329), .ZN(n5527) );
  NAND2_X1 U5166 ( .A1(n6513), .A2(n6326), .ZN(n6339) );
  NOR3_X1 U5167 ( .A1(n6530), .A2(n4193), .A3(n6339), .ZN(n6343) );
  NOR2_X1 U5168 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), .ZN(
        n6344) );
  INV_X1 U5169 ( .A(n6344), .ZN(n4142) );
  NOR3_X1 U5170 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4142), .A3(n6513), .ZN(
        n6349) );
  INV_X1 U5171 ( .A(n6349), .ZN(n4143) );
  NAND2_X1 U5172 ( .A1(n6071), .A2(n4143), .ZN(n4144) );
  OR2_X1 U5173 ( .A1(n6343), .A2(n4144), .ZN(n4145) );
  MUX2_X1 U5174 ( .A(n2962), .B(n2964), .S(EBX_REG_24__SCAN_IN), .Z(n4147) );
  NAND2_X1 U5175 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U5176 ( .A1(n4147), .A2(n4146), .ZN(n4227) );
  MUX2_X1 U5177 ( .A(n4153), .B(n2962), .S(EBX_REG_25__SCAN_IN), .Z(n4148) );
  OAI21_X1 U5178 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5120), .A(n4148), 
        .ZN(n5132) );
  INV_X1 U5179 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5180 ( .A1(n2964), .A2(n5385), .ZN(n4150) );
  INV_X1 U5181 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U5182 ( .A1(n4167), .A2(n5237), .ZN(n4149) );
  NAND3_X1 U5183 ( .A1(n4150), .A2(n2963), .A3(n4149), .ZN(n4152) );
  NAND2_X1 U5184 ( .A1(n3580), .A2(n5237), .ZN(n4151) );
  AND2_X1 U5185 ( .A1(n4152), .A2(n4151), .ZN(n5231) );
  MUX2_X1 U5186 ( .A(n4153), .B(n2962), .S(EBX_REG_27__SCAN_IN), .Z(n4155) );
  OR2_X1 U5187 ( .A1(n5120), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4154)
         );
  AND2_X1 U5188 ( .A1(n4155), .A2(n4154), .ZN(n5225) );
  MUX2_X1 U5189 ( .A(n2963), .B(n2964), .S(EBX_REG_28__SCAN_IN), .Z(n4158) );
  NAND2_X1 U5190 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U5191 ( .A1(n4158), .A2(n4157), .ZN(n5218) );
  OR2_X1 U5192 ( .A1(n5120), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4160)
         );
  INV_X1 U5193 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U5194 ( .A1(n4167), .A2(n5214), .ZN(n4159) );
  NAND2_X1 U5195 ( .A1(n4160), .A2(n4159), .ZN(n5209) );
  INV_X1 U5196 ( .A(n5220), .ZN(n4162) );
  AND2_X1 U5197 ( .A1(n4156), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4161)
         );
  AOI21_X1 U5198 ( .B1(n5120), .B2(EBX_REG_30__SCAN_IN), .A(n4161), .ZN(n5117)
         );
  AOI21_X1 U5199 ( .B1(n5116), .B2(n4162), .A(n5117), .ZN(n4165) );
  NAND2_X1 U5200 ( .A1(n5116), .A2(n2962), .ZN(n5118) );
  INV_X1 U5201 ( .A(n5117), .ZN(n4163) );
  AOI21_X1 U5202 ( .B1(n5220), .B2(n3580), .A(n4163), .ZN(n4164) );
  AOI22_X1 U5203 ( .A1(n4165), .A2(n5118), .B1(n4164), .B2(n5116), .ZN(n5349)
         );
  NOR2_X1 U5204 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4179) );
  INV_X1 U5205 ( .A(n4179), .ZN(n4181) );
  NAND2_X1 U5206 ( .A1(n5349), .A2(n5831), .ZN(n4188) );
  INV_X1 U5207 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6571) );
  INV_X1 U5208 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5545) );
  INV_X1 U5209 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6413) );
  NOR2_X1 U5210 ( .A1(n5545), .A2(n6413), .ZN(n4174) );
  AND3_X1 U5211 ( .A1(n4946), .A2(n5123), .A3(n4179), .ZN(n4168) );
  NAND3_X1 U5212 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4176) );
  NAND2_X1 U5213 ( .A1(n5804), .A2(n5817), .ZN(n5832) );
  INV_X1 U5214 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6598) );
  INV_X1 U5215 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5155) );
  NOR3_X1 U5216 ( .A1(n3652), .A2(n6598), .A3(n5155), .ZN(n4173) );
  AND3_X1 U5217 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4171) );
  INV_X1 U5218 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6392) );
  INV_X1 U5219 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6388) );
  INV_X1 U5220 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6385) );
  INV_X1 U5221 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6379) );
  INV_X1 U5222 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6377) );
  NAND3_X1 U5223 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5794) );
  OR2_X1 U5224 ( .A1(n6377), .A2(n5794), .ZN(n5758) );
  NOR2_X1 U5225 ( .A1(n6379), .A2(n5758), .ZN(n5763) );
  NAND4_X1 U5226 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5763), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U5227 ( .A1(n6385), .A2(n5742), .ZN(n5743) );
  NAND2_X1 U5228 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5743), .ZN(n5731) );
  NOR2_X1 U5229 ( .A1(n6388), .A2(n5731), .ZN(n5716) );
  NAND2_X1 U5230 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5716), .ZN(n5709) );
  NOR2_X1 U5231 ( .A1(n6392), .A2(n5709), .ZN(n5703) );
  NAND2_X1 U5232 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5703), .ZN(n4175) );
  NOR2_X1 U5233 ( .A1(n5790), .A2(n4175), .ZN(n5199) );
  NAND4_X1 U5234 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5199), .ZN(n5168) );
  INV_X1 U5235 ( .A(n5168), .ZN(n4170) );
  NAND2_X1 U5236 ( .A1(n4171), .A2(n4170), .ZN(n4172) );
  NAND2_X1 U5237 ( .A1(n5832), .A2(n4172), .ZN(n5593) );
  OAI21_X1 U5238 ( .B1(n4173), .B2(n5817), .A(n5593), .ZN(n5574) );
  AOI21_X1 U5239 ( .B1(n4176), .B2(n5832), .A(n5574), .ZN(n5563) );
  OAI21_X1 U5240 ( .B1(n4174), .B2(n5817), .A(n5563), .ZN(n5541) );
  NOR2_X1 U5241 ( .A1(n6571), .A2(n5541), .ZN(n5533) );
  INV_X1 U5242 ( .A(n5832), .ZN(n5200) );
  AOI21_X1 U5243 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5533), .A(n5200), .ZN(n5114) );
  INV_X1 U5244 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6404) );
  INV_X1 U5245 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U5246 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5198) );
  NAND2_X1 U5247 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5189), .ZN(n5181) );
  NAND2_X1 U5248 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5174), .ZN(n5592) );
  NAND4_X1 U5249 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5160), .ZN(n5143) );
  NOR2_X1 U5250 ( .A1(n5143), .A2(n4176), .ZN(n5555) );
  NAND3_X1 U5251 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5555), .ZN(n5534) );
  NOR2_X1 U5252 ( .A1(n6571), .A2(n5534), .ZN(n5112) );
  INV_X1 U5253 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6422) );
  INV_X1 U5254 ( .A(n6362), .ZN(n4407) );
  NAND2_X1 U5255 ( .A1(n4407), .A2(n4179), .ZN(n6333) );
  INV_X1 U5256 ( .A(n6333), .ZN(n4180) );
  OR2_X1 U5257 ( .A1(n6452), .A2(n4180), .ZN(n5124) );
  INV_X1 U5258 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4182) );
  NAND3_X1 U5259 ( .A1(n4946), .A2(n4182), .A3(n4181), .ZN(n4183) );
  NAND2_X1 U5260 ( .A1(n5124), .A2(n4183), .ZN(n4184) );
  NOR2_X2 U5261 ( .A1(n5790), .A2(n4193), .ZN(n5820) );
  AOI22_X1 U5262 ( .A1(EBX_REG_30__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5820), .ZN(n4185) );
  OAI21_X1 U5263 ( .B1(n4213), .B2(n5835), .A(n4185), .ZN(n4186) );
  AOI221_X1 U5264 ( .B1(n5114), .B2(REIP_REG_30__SCAN_IN), .C1(n5112), .C2(
        n6422), .A(n4186), .ZN(n4187) );
  OAI21_X1 U5265 ( .B1(n4215), .B2(n5780), .A(n3011), .ZN(U2797) );
  NAND2_X1 U5266 ( .A1(n4189), .A2(n6029), .ZN(n4204) );
  OAI21_X1 U5267 ( .B1(n4190), .B2(n4192), .A(n4244), .ZN(n5578) );
  NAND3_X1 U5268 ( .A1(n6530), .A2(STATE2_REG_1__SCAN_IN), .A3(
        STATEBS16_REG_SCAN_IN), .ZN(n6355) );
  NAND2_X1 U5269 ( .A1(n4194), .A2(n6238), .ZN(n6449) );
  AND2_X1 U5270 ( .A1(n6449), .A2(n6530), .ZN(n4195) );
  NAND2_X1 U5271 ( .A1(n6530), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4197) );
  INV_X1 U5272 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n4534) );
  NAND2_X1 U5273 ( .A1(n4534), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4196) );
  NAND2_X1 U5274 ( .A1(n4197), .A2(n4196), .ZN(n4310) );
  INV_X1 U5275 ( .A(n5571), .ZN(n4198) );
  NOR2_X1 U5276 ( .A1(n6035), .A2(n4198), .ZN(n4199) );
  AOI211_X1 U5277 ( .C1(PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n6025), .A(n4200), 
        .B(n4199), .ZN(n4201) );
  NAND2_X1 U5278 ( .A1(n4204), .A2(n4203), .ZN(U2963) );
  AND2_X1 U5279 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4233) );
  AND3_X1 U5280 ( .A1(n5399), .A2(n5422), .A3(n4233), .ZN(n4205) );
  NOR2_X1 U5281 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5421) );
  NOR2_X1 U5282 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5400) );
  INV_X1 U5283 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4225) );
  INV_X1 U5284 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U5285 ( .A1(n3439), .A2(n5386), .ZN(n4207) );
  NAND2_X1 U5286 ( .A1(n4271), .A2(n4207), .ZN(n4208) );
  NAND2_X1 U5287 ( .A1(n2965), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5379) );
  AND2_X1 U5288 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5363) );
  NOR2_X1 U5289 ( .A1(n2965), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5381)
         );
  NOR2_X1 U5290 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5364) );
  AND2_X1 U5291 ( .A1(n5381), .A2(n5364), .ZN(n4252) );
  NAND2_X1 U5292 ( .A1(n4252), .A2(n5354), .ZN(n4272) );
  INV_X1 U5293 ( .A(n4272), .ZN(n4209) );
  XNOR2_X2 U5294 ( .A(n4211), .B(n4210), .ZN(n5342) );
  INV_X2 U5295 ( .A(n6071), .ZN(n6104) );
  NAND2_X1 U5296 ( .A1(n6104), .A2(REIP_REG_30__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U5297 ( .A1(n6025), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4212)
         );
  OAI211_X1 U5298 ( .C1(n4213), .C2(n6035), .A(n5345), .B(n4212), .ZN(n4214)
         );
  INV_X1 U5299 ( .A(n4214), .ZN(n4217) );
  NAND2_X1 U5300 ( .A1(n4222), .A2(n4221), .ZN(n5296) );
  NAND3_X1 U5301 ( .A1(n2965), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4223) );
  OAI22_X2 U5302 ( .A1(n4224), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5296), .B2(n4223), .ZN(n4226) );
  XNOR2_X1 U5303 ( .A(n4226), .B(n4225), .ZN(n4242) );
  NAND2_X1 U5304 ( .A1(n4242), .A2(n6126), .ZN(n4241) );
  OR2_X1 U5305 ( .A1(n4228), .A2(n4227), .ZN(n4229) );
  NAND2_X1 U5306 ( .A1(n5131), .A2(n4229), .ZN(n5240) );
  INV_X1 U5307 ( .A(n5240), .ZN(n4231) );
  INV_X1 U5308 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4230) );
  NOR2_X1 U5309 ( .A1(n6071), .A2(n4230), .ZN(n4247) );
  AOI21_X1 U5310 ( .B1(n4231), .B2(n6106), .A(n4247), .ZN(n4239) );
  AND2_X1 U5311 ( .A1(n5399), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4232)
         );
  NAND2_X1 U5312 ( .A1(n6112), .A2(n4888), .ZN(n4235) );
  INV_X1 U5313 ( .A(n4233), .ZN(n4234) );
  NAND2_X1 U5314 ( .A1(n4235), .A2(n4234), .ZN(n4236) );
  INV_X1 U5315 ( .A(n5383), .ZN(n5395) );
  OAI21_X1 U5316 ( .B1(n5332), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5395), 
        .ZN(n4238) );
  NAND2_X1 U5317 ( .A1(n4241), .A2(n4240), .ZN(U2994) );
  NAND2_X1 U5318 ( .A1(n4242), .A2(n6029), .ZN(n4251) );
  XNOR2_X1 U5319 ( .A(n4244), .B(n4243), .ZN(n5276) );
  NOR2_X1 U5320 ( .A1(n6035), .A2(n4245), .ZN(n4246) );
  AOI211_X1 U5321 ( .C1(n6025), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4247), 
        .B(n4246), .ZN(n4248) );
  NAND2_X1 U5322 ( .A1(n4251), .A2(n4250), .ZN(U2962) );
  XNOR2_X1 U5323 ( .A(n4253), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5359)
         );
  NAND2_X1 U5324 ( .A1(n5359), .A2(n6029), .ZN(n4260) );
  INV_X1 U5325 ( .A(n4254), .ZN(n5217) );
  NOR2_X1 U5326 ( .A1(n6071), .A2(n6571), .ZN(n5352) );
  AOI21_X1 U5327 ( .B1(n6025), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5352), 
        .ZN(n4256) );
  OAI21_X1 U5328 ( .B1(n4257), .B2(n6035), .A(n4256), .ZN(n4258) );
  AOI21_X1 U5329 ( .B1(n5207), .B2(n6030), .A(n4258), .ZN(n4259) );
  NAND2_X1 U5330 ( .A1(n4260), .A2(n4259), .ZN(U2957) );
  NAND2_X1 U5331 ( .A1(n4262), .A2(n4261), .ZN(n4266) );
  AOI22_X1 U5332 ( .A1(n4264), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4263), .ZN(n4265) );
  XNOR2_X2 U5333 ( .A(n4266), .B(n4265), .ZN(n5130) );
  INV_X1 U5334 ( .A(n4267), .ZN(n4269) );
  NAND2_X1 U5335 ( .A1(n6104), .A2(REIP_REG_31__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U5336 ( .A1(n6025), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4268)
         );
  OAI211_X1 U5337 ( .C1(n4269), .C2(n6035), .A(n5337), .B(n4268), .ZN(n4270)
         );
  NAND2_X1 U5338 ( .A1(n5331), .A2(n6029), .ZN(n4274) );
  OAI211_X1 U5339 ( .C1(n5130), .C2(n4314), .A(n4275), .B(n4274), .ZN(U2955)
         );
  NOR2_X1 U5340 ( .A1(n6238), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5169) );
  INV_X1 U5341 ( .A(n5169), .ZN(n4276) );
  NAND2_X1 U5342 ( .A1(n4293), .A2(n4276), .ZN(n5526) );
  INV_X1 U5343 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n4277) );
  NAND2_X1 U5344 ( .A1(n5527), .A2(n4277), .ZN(n4280) );
  NAND2_X1 U5345 ( .A1(n6452), .A2(n4278), .ZN(n4283) );
  NAND2_X1 U5346 ( .A1(n6448), .A2(n4283), .ZN(n4279) );
  OAI21_X1 U5347 ( .B1(n5526), .B2(n4280), .A(n4279), .ZN(n4281) );
  INV_X1 U5348 ( .A(n4281), .ZN(U3474) );
  OAI22_X1 U5349 ( .A1(n4438), .A2(n3224), .B1(n4140), .B2(n4282), .ZN(n5670)
         );
  AOI21_X1 U5350 ( .B1(n4283), .B2(n6362), .A(READY_N), .ZN(n6451) );
  OR2_X1 U5351 ( .A1(n5670), .A2(n6451), .ZN(n6320) );
  AND2_X1 U5352 ( .A1(n6320), .A2(n6329), .ZN(n5677) );
  INV_X1 U5353 ( .A(MORE_REG_SCAN_IN), .ZN(n4291) );
  OR2_X1 U5354 ( .A1(n4411), .A2(n6316), .ZN(n4284) );
  NOR2_X1 U5355 ( .A1(n4284), .A2(n4140), .ZN(n4289) );
  NAND2_X1 U5356 ( .A1(n4286), .A2(n4285), .ZN(n4288) );
  NAND2_X1 U5357 ( .A1(n4438), .A2(n4388), .ZN(n4287) );
  OAI211_X1 U5358 ( .C1(n4438), .C2(n4289), .A(n4288), .B(n4287), .ZN(n6317)
         );
  NAND2_X1 U5359 ( .A1(n5677), .A2(n6317), .ZN(n4290) );
  OAI21_X1 U5360 ( .B1(n5677), .B2(n4291), .A(n4290), .ZN(U3471) );
  INV_X1 U5361 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6546) );
  INV_X1 U5362 ( .A(READY_N), .ZN(n4295) );
  INV_X1 U5363 ( .A(n4293), .ZN(n4294) );
  OAI21_X1 U5364 ( .B1(n4296), .B2(n4295), .A(n4294), .ZN(n4297) );
  INV_X1 U5365 ( .A(DATAI_5_), .ZN(n4298) );
  OAI222_X1 U5366 ( .A1(n5951), .A2(n4299), .B1(n6546), .B2(n5900), .C1(n5945), 
        .C2(n4298), .ZN(U2929) );
  INV_X1 U5367 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6501) );
  INV_X1 U5368 ( .A(DATAI_12_), .ZN(n4300) );
  NOR2_X1 U5369 ( .A1(n5945), .A2(n4300), .ZN(n5941) );
  AOI21_X1 U5370 ( .B1(n6613), .B2(EAX_REG_28__SCAN_IN), .A(n5941), .ZN(n4301)
         );
  OAI21_X1 U5371 ( .B1(n6501), .B2(n5900), .A(n4301), .ZN(U2936) );
  INV_X1 U5372 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6506) );
  INV_X1 U5373 ( .A(DATAI_11_), .ZN(n4302) );
  NOR2_X1 U5374 ( .A1(n5945), .A2(n4302), .ZN(n5914) );
  AOI21_X1 U5375 ( .B1(n6613), .B2(EAX_REG_11__SCAN_IN), .A(n5914), .ZN(n4303)
         );
  OAI21_X1 U5376 ( .B1(n5900), .B2(n6506), .A(n4303), .ZN(U2950) );
  INV_X1 U5377 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6553) );
  AOI22_X1 U5378 ( .A1(n5949), .A2(DATAI_0_), .B1(n6613), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4304) );
  OAI21_X1 U5379 ( .B1(n5900), .B2(n6553), .A(n4304), .ZN(U2924) );
  INV_X1 U5380 ( .A(n5092), .ZN(n6299) );
  NAND2_X1 U5381 ( .A1(n4305), .A2(n6299), .ZN(n4306) );
  NAND2_X1 U5382 ( .A1(n5951), .A2(n4306), .ZN(n4307) );
  INV_X1 U5383 ( .A(n4439), .ZN(n6352) );
  INV_X1 U5384 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U5385 ( .A1(n5890), .A2(n4946), .ZN(n5870) );
  INV_X1 U5386 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4308) );
  OAI222_X1 U5387 ( .A1(n5888), .A2(n6549), .B1(n5870), .B2(n4308), .C1(n6501), 
        .C2(n5892), .ZN(U2895) );
  INV_X1 U5388 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6550) );
  OAI222_X1 U5389 ( .A1(n5888), .A2(n6550), .B1(n5870), .B2(n4299), .C1(n6546), 
        .C2(n5892), .ZN(U2902) );
  XNOR2_X1 U5390 ( .A(n4309), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4341)
         );
  OAI21_X1 U5391 ( .B1(n6025), .B2(n4310), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4317) );
  OAI21_X1 U5392 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(n5843) );
  INV_X1 U5393 ( .A(n5843), .ZN(n4315) );
  INV_X1 U5394 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6444) );
  NOR2_X1 U5395 ( .A1(n6071), .A2(n6444), .ZN(n4337) );
  AOI21_X1 U5396 ( .B1(n4315), .B2(n6030), .A(n4337), .ZN(n4316) );
  OAI211_X1 U5397 ( .C1(n4341), .C2(n5675), .A(n4317), .B(n4316), .ZN(U2986)
         );
  OR2_X1 U5398 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  NAND2_X1 U5399 ( .A1(n4321), .A2(n4320), .ZN(n4957) );
  NAND2_X1 U5400 ( .A1(n4388), .A2(n6329), .ZN(n4322) );
  NOR2_X1 U5401 ( .A1(n4438), .A2(n4322), .ZN(n4327) );
  OR2_X1 U5402 ( .A1(n4323), .A2(n4156), .ZN(n4325) );
  NOR2_X1 U5403 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  INV_X2 U5404 ( .A(n5850), .ZN(n5264) );
  INV_X1 U5405 ( .A(n4949), .ZN(n4330) );
  INV_X1 U5406 ( .A(n4328), .ZN(n4329) );
  AOI21_X1 U5407 ( .B1(n4330), .B2(n4156), .A(n4329), .ZN(n6119) );
  INV_X1 U5408 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4331) );
  OAI222_X1 U5409 ( .A1(n4957), .A2(n5264), .B1(n5267), .B2(n6119), .C1(n5852), 
        .C2(n4331), .ZN(U2858) );
  INV_X1 U5410 ( .A(n5120), .ZN(n4335) );
  INV_X1 U5411 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4334) );
  INV_X1 U5412 ( .A(n4332), .ZN(n4333) );
  AOI21_X1 U5413 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n5830) );
  NAND2_X1 U5414 ( .A1(n5056), .A2(n4888), .ZN(n5058) );
  NAND2_X1 U5415 ( .A1(n5058), .A2(n4334), .ZN(n6128) );
  INV_X1 U5416 ( .A(n6128), .ZN(n4336) );
  AOI211_X1 U5417 ( .C1(n6106), .C2(n5830), .A(n4337), .B(n4336), .ZN(n4340)
         );
  INV_X1 U5418 ( .A(n6129), .ZN(n4338) );
  OAI21_X1 U5419 ( .B1(n5059), .B2(n4338), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4339) );
  OAI211_X1 U5420 ( .C1(n4341), .C2(n6083), .A(n4340), .B(n4339), .ZN(U3018)
         );
  INV_X1 U5421 ( .A(n5830), .ZN(n4342) );
  OAI222_X1 U5422 ( .A1(n5843), .A2(n5264), .B1(n5852), .B2(n5837), .C1(n4342), 
        .C2(n5267), .ZN(U2859) );
  INV_X1 U5423 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5919) );
  AOI22_X1 U5424 ( .A1(n6450), .A2(UWORD_REG_14__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4343) );
  OAI21_X1 U5425 ( .B1(n5919), .B2(n5870), .A(n4343), .ZN(U2893) );
  AOI22_X1 U5426 ( .A1(n6450), .A2(UWORD_REG_11__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4344) );
  OAI21_X1 U5427 ( .B1(n4048), .B2(n5870), .A(n4344), .ZN(U2896) );
  AOI22_X1 U5428 ( .A1(n6450), .A2(UWORD_REG_13__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4345) );
  OAI21_X1 U5429 ( .B1(n4090), .B2(n5870), .A(n4345), .ZN(U2894) );
  INV_X1 U5430 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5899) );
  AOI22_X1 U5431 ( .A1(n5883), .A2(UWORD_REG_1__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4346) );
  OAI21_X1 U5432 ( .B1(n5899), .B2(n5870), .A(n4346), .ZN(U2906) );
  INV_X1 U5433 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5906) );
  AOI22_X1 U5434 ( .A1(n5883), .A2(UWORD_REG_6__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4347) );
  OAI21_X1 U5435 ( .B1(n5906), .B2(n5870), .A(n4347), .ZN(U2901) );
  AOI22_X1 U5436 ( .A1(n5883), .A2(UWORD_REG_2__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5437 ( .B1(n6488), .B2(n5870), .A(n4348), .ZN(U2905) );
  INV_X1 U5438 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U5439 ( .A1(n5883), .A2(UWORD_REG_9__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5440 ( .B1(n4350), .B2(n5870), .A(n4349), .ZN(U2898) );
  INV_X1 U5441 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5913) );
  AOI22_X1 U5442 ( .A1(n5883), .A2(UWORD_REG_10__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4351) );
  OAI21_X1 U5443 ( .B1(n5913), .B2(n5870), .A(n4351), .ZN(U2897) );
  INV_X1 U5444 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6503) );
  AOI22_X1 U5445 ( .A1(n5883), .A2(UWORD_REG_3__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4352) );
  OAI21_X1 U5446 ( .B1(n6503), .B2(n5870), .A(n4352), .ZN(U2904) );
  INV_X1 U5447 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5904) );
  AOI22_X1 U5448 ( .A1(n5883), .A2(UWORD_REG_4__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5449 ( .B1(n5904), .B2(n5870), .A(n4353), .ZN(U2903) );
  INV_X1 U5450 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5910) );
  AOI22_X1 U5451 ( .A1(n5883), .A2(UWORD_REG_8__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4354) );
  OAI21_X1 U5452 ( .B1(n5910), .B2(n5870), .A(n4354), .ZN(U2899) );
  NOR2_X1 U5453 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  NOR2_X1 U5454 ( .A1(n4355), .A2(n4358), .ZN(n6031) );
  INV_X1 U5455 ( .A(n6031), .ZN(n4840) );
  AND2_X1 U5456 ( .A1(n4360), .A2(n4359), .ZN(n4361) );
  OR2_X1 U5457 ( .A1(n4361), .A2(n5806), .ZN(n5825) );
  INV_X1 U5458 ( .A(n5825), .ZN(n6105) );
  AOI22_X1 U5459 ( .A1(n5849), .A2(n6105), .B1(n5261), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4362) );
  OAI21_X1 U5460 ( .B1(n4840), .B2(n5264), .A(n4362), .ZN(U2857) );
  XOR2_X1 U5461 ( .A(n4363), .B(n4364), .Z(n6125) );
  INV_X1 U5462 ( .A(n6125), .ZN(n4368) );
  NAND2_X1 U5463 ( .A1(n6104), .A2(REIP_REG_1__SCAN_IN), .ZN(n6118) );
  INV_X1 U5464 ( .A(n6118), .ZN(n4366) );
  OAI22_X1 U5465 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6035), .B1(n4314), 
        .B2(n4957), .ZN(n4365) );
  AOI211_X1 U5466 ( .C1(n6025), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4366), 
        .B(n4365), .ZN(n4367) );
  OAI21_X1 U5467 ( .B1(n4368), .B2(n5675), .A(n4367), .ZN(U2985) );
  XNOR2_X1 U5468 ( .A(n4370), .B(n4369), .ZN(n5996) );
  OAI21_X1 U5469 ( .B1(n4462), .B2(n4371), .A(n4531), .ZN(n6072) );
  INV_X1 U5470 ( .A(n6072), .ZN(n4372) );
  AOI22_X1 U5471 ( .A1(n5849), .A2(n4372), .B1(n5261), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4373) );
  OAI21_X1 U5472 ( .B1(n5996), .B2(n5264), .A(n4373), .ZN(U2853) );
  NAND2_X1 U5473 ( .A1(n5808), .A2(n4374), .ZN(n4375) );
  AND2_X1 U5474 ( .A1(n4460), .A2(n4375), .ZN(n6092) );
  INV_X1 U5475 ( .A(n6092), .ZN(n5795) );
  INV_X1 U5476 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4380) );
  INV_X1 U5477 ( .A(n4355), .ZN(n4376) );
  OR2_X1 U5478 ( .A1(n4376), .A2(n4474), .ZN(n4377) );
  AOI21_X1 U5479 ( .B1(n4378), .B2(n4377), .A(n4463), .ZN(n4379) );
  INV_X1 U5480 ( .A(n4379), .ZN(n6015) );
  OAI222_X1 U5481 ( .A1(n5795), .A2(n5267), .B1(n5852), .B2(n4380), .C1(n5264), 
        .C2(n6015), .ZN(U2855) );
  AND2_X1 U5482 ( .A1(n4383), .A2(n4382), .ZN(n4385) );
  NAND4_X1 U5483 ( .A1(n3551), .A2(n4385), .A3(n5664), .A4(n4384), .ZN(n4387)
         );
  NOR2_X1 U5484 ( .A1(n4387), .A2(n4386), .ZN(n4423) );
  INV_X1 U5485 ( .A(n4423), .ZN(n6297) );
  NAND2_X1 U5486 ( .A1(n5812), .A2(n6297), .ZN(n4402) );
  OR2_X1 U5487 ( .A1(n4388), .A2(n4411), .ZN(n4421) );
  MUX2_X1 U5488 ( .A(n4390), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5096), 
        .Z(n4392) );
  NOR2_X1 U5489 ( .A1(n4392), .A2(n4391), .ZN(n4400) );
  NAND2_X1 U5490 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4393) );
  XNOR2_X1 U5491 ( .A(n4415), .B(n4393), .ZN(n4398) );
  INV_X1 U5492 ( .A(n4394), .ZN(n4395) );
  OAI21_X1 U5493 ( .B1(n5096), .B2(n4415), .A(n4395), .ZN(n4397) );
  NOR2_X1 U5494 ( .A1(n4397), .A2(n4396), .ZN(n5476) );
  OAI22_X1 U5495 ( .A1(n5092), .A2(n4398), .B1(n5476), .B2(n4417), .ZN(n4399)
         );
  AOI21_X1 U5496 ( .B1(n4421), .B2(n4400), .A(n4399), .ZN(n4401) );
  AND2_X1 U5497 ( .A1(n4402), .A2(n4401), .ZN(n5477) );
  INV_X1 U5498 ( .A(n4403), .ZN(n4404) );
  OR2_X1 U5499 ( .A1(n5664), .A2(n4404), .ZN(n4405) );
  AND2_X1 U5500 ( .A1(n4406), .A2(n4405), .ZN(n4413) );
  OAI21_X1 U5501 ( .B1(n3552), .B2(n6299), .A(n4407), .ZN(n4409) );
  AOI21_X1 U5502 ( .B1(n4409), .B2(n4408), .A(READY_N), .ZN(n4410) );
  OAI21_X1 U5503 ( .B1(n4411), .B2(n4410), .A(n4438), .ZN(n4412) );
  OAI211_X1 U5504 ( .C1(n4438), .C2(n4414), .A(n4413), .B(n4412), .ZN(n6300)
         );
  MUX2_X1 U5505 ( .A(n4415), .B(n5477), .S(n6300), .Z(n6312) );
  INV_X1 U5506 ( .A(n6312), .ZN(n4428) );
  OR2_X1 U5507 ( .A1(n6300), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4426)
         );
  XNOR2_X1 U5508 ( .A(n5096), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4420)
         );
  XNOR2_X1 U5509 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4418) );
  OAI22_X1 U5510 ( .A1(n5092), .A2(n4418), .B1(n4417), .B2(n4420), .ZN(n4419)
         );
  AOI21_X1 U5511 ( .B1(n4421), .B2(n4420), .A(n4419), .ZN(n4422) );
  OAI21_X1 U5512 ( .B1(n4416), .B2(n4423), .A(n4422), .ZN(n5103) );
  INV_X1 U5513 ( .A(n5103), .ZN(n4424) );
  NAND2_X1 U5514 ( .A1(n6300), .A2(n4424), .ZN(n4425) );
  NAND2_X1 U5515 ( .A1(n4426), .A2(n4425), .ZN(n6307) );
  INV_X1 U5516 ( .A(n6307), .ZN(n4427) );
  NAND3_X1 U5517 ( .A1(n4428), .A2(n4427), .A3(n6513), .ZN(n4430) );
  INV_X1 U5518 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5676) );
  AND2_X1 U5519 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5676), .ZN(n4435) );
  NAND2_X1 U5520 ( .A1(n4391), .A2(n4435), .ZN(n4429) );
  NOR2_X1 U5521 ( .A1(n6324), .A2(n4431), .ZN(n4442) );
  INV_X1 U5522 ( .A(n6167), .ZN(n4572) );
  OR2_X1 U5523 ( .A1(n3316), .A2(n4572), .ZN(n4433) );
  XNOR2_X1 U5524 ( .A(n4433), .B(n4432), .ZN(n5796) );
  OAI22_X1 U5525 ( .A1(n6300), .A2(n4432), .B1(n5664), .B2(n5796), .ZN(n4434)
         );
  NAND2_X1 U5526 ( .A1(n4434), .A2(n6513), .ZN(n4437) );
  NAND2_X1 U5527 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4435), .ZN(n4436) );
  NAND2_X1 U5528 ( .A1(n4437), .A2(n4436), .ZN(n6322) );
  NOR3_X1 U5529 ( .A1(n4442), .A2(n6322), .A3(FLUSH_REG_SCAN_IN), .ZN(n4440)
         );
  NAND2_X1 U5530 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4439), .ZN(n6428) );
  OR2_X1 U5531 ( .A1(n6322), .A2(n6352), .ZN(n4441) );
  OR2_X1 U5532 ( .A1(n4442), .A2(n4441), .ZN(n6327) );
  INV_X1 U5533 ( .A(n6327), .ZN(n4444) );
  AND2_X1 U5534 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4193), .ZN(n5473) );
  OAI22_X1 U5535 ( .A1(n3709), .A2(n6238), .B1(n3712), .B2(n5473), .ZN(n4443)
         );
  OAI21_X1 U5536 ( .B1(n4444), .B2(n4443), .A(n6130), .ZN(n4445) );
  OAI21_X1 U5537 ( .B1(n6130), .B2(n4997), .A(n4445), .ZN(U3465) );
  NAND2_X1 U5538 ( .A1(n4446), .A2(n4449), .ZN(n4481) );
  NAND2_X1 U5539 ( .A1(n4685), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4769) );
  AND2_X1 U5540 ( .A1(n4769), .A2(n6235), .ZN(n6132) );
  INV_X1 U5541 ( .A(n4449), .ZN(n4450) );
  NAND2_X1 U5542 ( .A1(n4999), .A2(n6232), .ZN(n6166) );
  AOI21_X1 U5543 ( .B1(n6132), .B2(n6166), .A(n6238), .ZN(n4452) );
  INV_X1 U5544 ( .A(n4448), .ZN(n4905) );
  OR2_X1 U5545 ( .A1(n6238), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5001) );
  INV_X1 U5546 ( .A(n5812), .ZN(n5481) );
  OAI22_X1 U5547 ( .A1(n4905), .A2(n5001), .B1(n5481), .B2(n5473), .ZN(n4451)
         );
  OAI21_X1 U5548 ( .B1(n4452), .B2(n4451), .A(n6130), .ZN(n4453) );
  OAI21_X1 U5549 ( .B1(n6130), .B2(n6490), .A(n4453), .ZN(U3462) );
  AOI211_X1 U5550 ( .C1(n4903), .C2(n4534), .A(n6238), .B(n6232), .ZN(n4457)
         );
  INV_X1 U5551 ( .A(n4455), .ZN(n4952) );
  NOR2_X1 U5552 ( .A1(n4952), .A2(n5473), .ZN(n4456) );
  OAI21_X1 U5553 ( .B1(n4457), .B2(n4456), .A(n6130), .ZN(n4458) );
  OAI21_X1 U5554 ( .B1(n6130), .B2(n6303), .A(n4458), .ZN(U3464) );
  AND2_X1 U5555 ( .A1(n4460), .A2(n4459), .ZN(n4461) );
  OR2_X1 U5556 ( .A1(n4462), .A2(n4461), .ZN(n5781) );
  XOR2_X1 U5557 ( .A(n4464), .B(n4463), .Z(n6002) );
  INV_X1 U5558 ( .A(n6002), .ZN(n4467) );
  INV_X1 U5559 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4465) );
  OAI222_X1 U5560 ( .A1(n5781), .A2(n5267), .B1(n5264), .B2(n4467), .C1(n5852), 
        .C2(n4465), .ZN(U2854) );
  OAI222_X1 U5561 ( .A1(n5858), .A2(n4467), .B1(n4841), .B2(n4298), .C1(n5109), 
        .C2(n3735), .ZN(U2886) );
  INV_X1 U5562 ( .A(DATAI_1_), .ZN(n5923) );
  OAI222_X1 U5563 ( .A1(n4957), .A2(n5858), .B1(n4841), .B2(n5923), .C1(n5109), 
        .C2(n3703), .ZN(U2890) );
  INV_X1 U5564 ( .A(DATAI_0_), .ZN(n5921) );
  OAI222_X1 U5565 ( .A1(n5843), .A2(n5858), .B1(n4841), .B2(n5921), .C1(n5109), 
        .C2(n3714), .ZN(U2891) );
  INV_X1 U5566 ( .A(DATAI_4_), .ZN(n5928) );
  INV_X1 U5567 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6555) );
  OAI222_X1 U5568 ( .A1(n6015), .A2(n5858), .B1(n4841), .B2(n5928), .C1(n5109), 
        .C2(n6555), .ZN(U2887) );
  XNOR2_X1 U5569 ( .A(n4468), .B(n4469), .ZN(n5979) );
  AOI22_X1 U5570 ( .A1(n5042), .A2(DATAI_8_), .B1(n5861), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5571 ( .B1(n5979), .B2(n5858), .A(n4470), .ZN(U2883) );
  NAND2_X1 U5572 ( .A1(n4530), .A2(n4471), .ZN(n4472) );
  AND2_X1 U5573 ( .A1(n4681), .A2(n4472), .ZN(n5755) );
  AOI22_X1 U5574 ( .A1(n5849), .A2(n5755), .B1(n5261), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4473) );
  OAI21_X1 U5575 ( .B1(n5979), .B2(n5264), .A(n4473), .ZN(U2851) );
  INV_X1 U5576 ( .A(DATAI_3_), .ZN(n4477) );
  XNOR2_X1 U5577 ( .A(n4355), .B(n4474), .ZN(n6021) );
  INV_X1 U5578 ( .A(n6021), .ZN(n4475) );
  OAI222_X1 U5579 ( .A1(n4477), .A2(n4841), .B1(n4476), .B2(n5109), .C1(n4475), 
        .C2(n5858), .ZN(U2888) );
  NOR2_X1 U5580 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4193), .ZN(n5086) );
  INV_X1 U5582 ( .A(n3712), .ZN(n6298) );
  AND2_X1 U5583 ( .A1(n5812), .A2(n6298), .ZN(n4764) );
  INV_X1 U5584 ( .A(n4416), .ZN(n4479) );
  INV_X1 U5585 ( .A(n4527), .ZN(n4480) );
  AOI21_X1 U5586 ( .B1(n4764), .B2(n6169), .A(n4480), .ZN(n4482) );
  OAI22_X1 U5587 ( .A1(n4482), .A2(n6238), .B1(n4688), .B2(n6326), .ZN(n4521)
         );
  NAND2_X1 U5588 ( .A1(n6244), .A2(n4521), .ZN(n4490) );
  OAI21_X1 U5589 ( .B1(n4487), .B2(n4314), .A(n5001), .ZN(n4483) );
  NAND2_X1 U5590 ( .A1(n4483), .A2(n4482), .ZN(n4484) );
  OAI211_X1 U5591 ( .C1(n6233), .C2(n4485), .A(n4484), .B(n6175), .ZN(n4524)
         );
  INV_X1 U5592 ( .A(DATAI_24_), .ZN(n4486) );
  NOR2_X1 U5593 ( .A1(n4314), .A2(n4486), .ZN(n6178) );
  NAND2_X1 U5594 ( .A1(n6030), .A2(DATAI_16_), .ZN(n4918) );
  OAI22_X1 U5595 ( .A1(n6247), .A2(n4715), .B1(n4756), .B2(n4918), .ZN(n4488)
         );
  AOI21_X1 U5596 ( .B1(n4524), .B2(INSTQUEUE_REG_15__0__SCAN_IN), .A(n4488), 
        .ZN(n4489) );
  OAI211_X1 U5597 ( .C1(n6621), .C2(n4527), .A(n4490), .B(n4489), .ZN(U3140)
         );
  NOR2_X2 U5598 ( .A1(n4520), .A2(n4491), .ZN(n6249) );
  INV_X1 U5599 ( .A(n6249), .ZN(n4569) );
  NAND2_X1 U5600 ( .A1(n6250), .A2(n4521), .ZN(n4494) );
  INV_X1 U5601 ( .A(DATAI_25_), .ZN(n5601) );
  NOR2_X1 U5602 ( .A1(n4314), .A2(n5601), .ZN(n6248) );
  INV_X1 U5603 ( .A(n6248), .ZN(n6144) );
  NAND2_X1 U5604 ( .A1(n6030), .A2(DATAI_17_), .ZN(n6253) );
  OAI22_X1 U5605 ( .A1(n6144), .A2(n4715), .B1(n4756), .B2(n6253), .ZN(n4492)
         );
  AOI21_X1 U5606 ( .B1(n4524), .B2(INSTQUEUE_REG_15__1__SCAN_IN), .A(n4492), 
        .ZN(n4493) );
  OAI211_X1 U5607 ( .C1(n4569), .C2(n4527), .A(n4494), .B(n4493), .ZN(U3141)
         );
  NOR2_X2 U5608 ( .A1(n4520), .A2(n4495), .ZN(n6255) );
  INV_X1 U5609 ( .A(n6255), .ZN(n4559) );
  INV_X1 U5610 ( .A(DATAI_2_), .ZN(n5925) );
  NAND2_X1 U5611 ( .A1(n6256), .A2(n4521), .ZN(n4499) );
  NAND2_X1 U5612 ( .A1(n6030), .A2(DATAI_26_), .ZN(n6259) );
  INV_X1 U5613 ( .A(DATAI_18_), .ZN(n4496) );
  NOR2_X1 U5614 ( .A1(n4314), .A2(n4496), .ZN(n6254) );
  INV_X1 U5615 ( .A(n6254), .ZN(n4925) );
  OAI22_X1 U5616 ( .A1(n6259), .A2(n4715), .B1(n4756), .B2(n4925), .ZN(n4497)
         );
  AOI21_X1 U5617 ( .B1(n4524), .B2(INSTQUEUE_REG_15__2__SCAN_IN), .A(n4497), 
        .ZN(n4498) );
  OAI211_X1 U5618 ( .C1(n4559), .C2(n4527), .A(n4499), .B(n4498), .ZN(U3142)
         );
  NOR2_X2 U5619 ( .A1(n4520), .A2(n4500), .ZN(n6261) );
  INV_X1 U5620 ( .A(n6261), .ZN(n4547) );
  NAND2_X1 U5621 ( .A1(n6262), .A2(n4521), .ZN(n4504) );
  INV_X1 U5622 ( .A(DATAI_27_), .ZN(n4501) );
  NOR2_X1 U5623 ( .A1(n4314), .A2(n4501), .ZN(n6190) );
  INV_X1 U5624 ( .A(n6190), .ZN(n6265) );
  NAND2_X1 U5625 ( .A1(n6030), .A2(DATAI_19_), .ZN(n6149) );
  OAI22_X1 U5626 ( .A1(n6265), .A2(n4715), .B1(n4756), .B2(n6149), .ZN(n4502)
         );
  AOI21_X1 U5627 ( .B1(n4524), .B2(INSTQUEUE_REG_15__3__SCAN_IN), .A(n4502), 
        .ZN(n4503) );
  OAI211_X1 U5628 ( .C1(n4547), .C2(n4527), .A(n4504), .B(n4503), .ZN(U3143)
         );
  NOR2_X2 U5629 ( .A1(n4520), .A2(n4505), .ZN(n6267) );
  INV_X1 U5630 ( .A(n6267), .ZN(n4562) );
  NAND2_X1 U5631 ( .A1(n6268), .A2(n4521), .ZN(n4509) );
  INV_X1 U5632 ( .A(DATAI_28_), .ZN(n4506) );
  NOR2_X1 U5633 ( .A1(n4314), .A2(n4506), .ZN(n6266) );
  INV_X1 U5634 ( .A(n6266), .ZN(n6219) );
  NAND2_X1 U5635 ( .A1(n6030), .A2(DATAI_20_), .ZN(n6271) );
  OAI22_X1 U5636 ( .A1(n6219), .A2(n4715), .B1(n4756), .B2(n6271), .ZN(n4507)
         );
  AOI21_X1 U5637 ( .B1(n4524), .B2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n4507), 
        .ZN(n4508) );
  OAI211_X1 U5638 ( .C1(n4562), .C2(n4527), .A(n4509), .B(n4508), .ZN(U3144)
         );
  NOR2_X2 U5639 ( .A1(n4520), .A2(n4510), .ZN(n6274) );
  INV_X1 U5640 ( .A(n6274), .ZN(n4544) );
  NAND2_X1 U5641 ( .A1(n6275), .A2(n4521), .ZN(n4514) );
  NAND2_X1 U5642 ( .A1(n6030), .A2(DATAI_29_), .ZN(n6228) );
  INV_X1 U5643 ( .A(DATAI_21_), .ZN(n4511) );
  NOR2_X1 U5644 ( .A1(n4314), .A2(n4511), .ZN(n6223) );
  INV_X1 U5645 ( .A(n6223), .ZN(n6279) );
  OAI22_X1 U5646 ( .A1(n6228), .A2(n4715), .B1(n4756), .B2(n6279), .ZN(n4512)
         );
  AOI21_X1 U5647 ( .B1(n4524), .B2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4512), 
        .ZN(n4513) );
  OAI211_X1 U5648 ( .C1(n4544), .C2(n4527), .A(n4514), .B(n4513), .ZN(U3145)
         );
  NOR2_X2 U5649 ( .A1(n4520), .A2(n4515), .ZN(n6281) );
  INV_X1 U5650 ( .A(n6281), .ZN(n4553) );
  INV_X1 U5651 ( .A(DATAI_6_), .ZN(n5931) );
  NAND2_X1 U5652 ( .A1(n6282), .A2(n4521), .ZN(n4519) );
  NAND2_X1 U5653 ( .A1(n6030), .A2(DATAI_30_), .ZN(n6285) );
  INV_X1 U5654 ( .A(DATAI_22_), .ZN(n4516) );
  NOR2_X1 U5655 ( .A1(n4314), .A2(n4516), .ZN(n6280) );
  INV_X1 U5656 ( .A(n6280), .ZN(n6158) );
  OAI22_X1 U5657 ( .A1(n6285), .A2(n4715), .B1(n4756), .B2(n6158), .ZN(n4517)
         );
  AOI21_X1 U5658 ( .B1(n4524), .B2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4517), 
        .ZN(n4518) );
  OAI211_X1 U5659 ( .C1(n4553), .C2(n4527), .A(n4519), .B(n4518), .ZN(U3146)
         );
  NOR2_X2 U5660 ( .A1(n4520), .A2(n5108), .ZN(n6288) );
  INV_X1 U5661 ( .A(n6288), .ZN(n4550) );
  INV_X1 U5662 ( .A(DATAI_7_), .ZN(n5933) );
  NAND2_X1 U5663 ( .A1(n6290), .A2(n4521), .ZN(n4526) );
  NAND2_X1 U5664 ( .A1(n6030), .A2(DATAI_31_), .ZN(n6295) );
  INV_X1 U5665 ( .A(DATAI_23_), .ZN(n4522) );
  NOR2_X1 U5666 ( .A1(n4314), .A2(n4522), .ZN(n6287) );
  INV_X1 U5667 ( .A(n6287), .ZN(n6165) );
  OAI22_X1 U5668 ( .A1(n6295), .A2(n4715), .B1(n4756), .B2(n6165), .ZN(n4523)
         );
  AOI21_X1 U5669 ( .B1(n4524), .B2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4523), 
        .ZN(n4525) );
  OAI211_X1 U5670 ( .C1(n4550), .C2(n4527), .A(n4526), .B(n4525), .ZN(U3147)
         );
  XOR2_X1 U5671 ( .A(n4529), .B(n4528), .Z(n5984) );
  INV_X1 U5672 ( .A(n5984), .ZN(n4722) );
  AOI21_X1 U5673 ( .B1(n4532), .B2(n4531), .A(n3605), .ZN(n6059) );
  AOI22_X1 U5674 ( .A1(n5849), .A2(n6059), .B1(n5261), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4533) );
  OAI21_X1 U5675 ( .B1(n4722), .B2(n5264), .A(n4533), .ZN(U2852) );
  NAND3_X1 U5676 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6309), .A3(n6303), .ZN(n4846) );
  NOR2_X1 U5677 ( .A1(n4997), .A2(n4846), .ZN(n4536) );
  INV_X1 U5678 ( .A(n4536), .ZN(n4568) );
  NOR2_X1 U5679 ( .A1(n4447), .A2(n4534), .ZN(n4535) );
  AOI21_X1 U5680 ( .B1(n4781), .B2(n4535), .A(n6238), .ZN(n4538) );
  NAND2_X1 U5681 ( .A1(n4952), .A2(n4416), .ZN(n4852) );
  INV_X1 U5682 ( .A(n4852), .ZN(n4842) );
  AOI21_X1 U5683 ( .B1(n4764), .B2(n4842), .A(n4536), .ZN(n4540) );
  AOI22_X1 U5684 ( .A1(n4538), .A2(n4540), .B1(n6238), .B2(n4846), .ZN(n4537)
         );
  NAND2_X1 U5685 ( .A1(n6175), .A2(n4537), .ZN(n4564) );
  INV_X1 U5686 ( .A(n4538), .ZN(n4539) );
  OAI22_X1 U5687 ( .A1(n4540), .A2(n4539), .B1(n6326), .B2(n4846), .ZN(n4563)
         );
  AOI22_X1 U5688 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4564), .B1(n6275), 
        .B2(n4563), .ZN(n4543) );
  INV_X1 U5689 ( .A(n6228), .ZN(n6272) );
  AOI22_X1 U5690 ( .A1(n4565), .A2(n6223), .B1(n6222), .B2(n6272), .ZN(n4542)
         );
  OAI211_X1 U5691 ( .C1(n4544), .C2(n4568), .A(n4543), .B(n4542), .ZN(U3097)
         );
  AOI22_X1 U5692 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4564), .B1(n6262), 
        .B2(n4563), .ZN(n4546) );
  INV_X1 U5693 ( .A(n6149), .ZN(n6260) );
  AOI22_X1 U5694 ( .A1(n4565), .A2(n6260), .B1(n6222), .B2(n6190), .ZN(n4545)
         );
  OAI211_X1 U5695 ( .C1(n4547), .C2(n4568), .A(n4546), .B(n4545), .ZN(U3095)
         );
  AOI22_X1 U5696 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4564), .B1(n6290), 
        .B2(n4563), .ZN(n4549) );
  INV_X1 U5697 ( .A(n6295), .ZN(n6205) );
  AOI22_X1 U5698 ( .A1(n4565), .A2(n6287), .B1(n6222), .B2(n6205), .ZN(n4548)
         );
  OAI211_X1 U5699 ( .C1(n4550), .C2(n4568), .A(n4549), .B(n4548), .ZN(U3099)
         );
  AOI22_X1 U5700 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4564), .B1(n6282), 
        .B2(n4563), .ZN(n4552) );
  INV_X1 U5701 ( .A(n6285), .ZN(n6200) );
  AOI22_X1 U5702 ( .A1(n4565), .A2(n6280), .B1(n6222), .B2(n6200), .ZN(n4551)
         );
  OAI211_X1 U5703 ( .C1(n4553), .C2(n4568), .A(n4552), .B(n4551), .ZN(U3098)
         );
  AOI22_X1 U5704 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4564), .B1(n6244), 
        .B2(n4563), .ZN(n4555) );
  INV_X1 U5705 ( .A(n4918), .ZN(n6230) );
  AOI22_X1 U5706 ( .A1(n4565), .A2(n6230), .B1(n6222), .B2(n6178), .ZN(n4554)
         );
  OAI211_X1 U5707 ( .C1(n6621), .C2(n4568), .A(n4555), .B(n4554), .ZN(U3092)
         );
  AOI22_X1 U5708 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4564), .B1(n6256), 
        .B2(n4563), .ZN(n4558) );
  INV_X1 U5709 ( .A(n6259), .ZN(n6186) );
  AOI22_X1 U5710 ( .A1(n4565), .A2(n6254), .B1(n6222), .B2(n6186), .ZN(n4557)
         );
  OAI211_X1 U5711 ( .C1(n4559), .C2(n4568), .A(n4558), .B(n4557), .ZN(U3094)
         );
  AOI22_X1 U5712 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4564), .B1(n6268), 
        .B2(n4563), .ZN(n4561) );
  INV_X1 U5713 ( .A(n6271), .ZN(n6216) );
  AOI22_X1 U5714 ( .A1(n4565), .A2(n6216), .B1(n6222), .B2(n6266), .ZN(n4560)
         );
  OAI211_X1 U5715 ( .C1(n4562), .C2(n4568), .A(n4561), .B(n4560), .ZN(U3096)
         );
  AOI22_X1 U5716 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4564), .B1(n6250), 
        .B2(n4563), .ZN(n4567) );
  INV_X1 U5717 ( .A(n6253), .ZN(n6182) );
  AOI22_X1 U5718 ( .A1(n4565), .A2(n6182), .B1(n6222), .B2(n6248), .ZN(n4566)
         );
  OAI211_X1 U5719 ( .C1(n4569), .C2(n4568), .A(n4567), .B(n4566), .ZN(U3093)
         );
  INV_X1 U5720 ( .A(n4999), .ZN(n4570) );
  INV_X1 U5721 ( .A(n4580), .ZN(n4571) );
  OAI21_X1 U5722 ( .B1(n4571), .B2(n4534), .A(n6233), .ZN(n4579) );
  INV_X1 U5723 ( .A(n4579), .ZN(n4576) );
  NAND2_X1 U5724 ( .A1(n4763), .A2(n4572), .ZN(n5487) );
  OR2_X1 U5725 ( .A1(n5487), .A2(n3712), .ZN(n4574) );
  NAND2_X1 U5726 ( .A1(n6303), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4765) );
  OR2_X1 U5727 ( .A1(n4765), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5483)
         );
  NOR2_X1 U5728 ( .A1(n4997), .A2(n5483), .ZN(n4604) );
  INV_X1 U5729 ( .A(n4604), .ZN(n4573) );
  NAND2_X1 U5730 ( .A1(n4574), .A2(n4573), .ZN(n4578) );
  INV_X1 U5731 ( .A(n5483), .ZN(n4575) );
  AOI21_X1 U5732 ( .B1(n6238), .B2(n5483), .A(n6237), .ZN(n4577) );
  OAI21_X1 U5733 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n4603) );
  NAND2_X1 U5734 ( .A1(n4580), .A2(n3709), .ZN(n5485) );
  OAI22_X1 U5735 ( .A1(n6285), .A2(n5485), .B1(n5030), .B2(n6158), .ZN(n4581)
         );
  AOI21_X1 U5736 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(n4603), .A(n4581), 
        .ZN(n4583) );
  NAND2_X1 U5737 ( .A1(n6281), .A2(n4604), .ZN(n4582) );
  OAI211_X1 U5738 ( .C1(n6203), .C2(n4607), .A(n4583), .B(n4582), .ZN(U3066)
         );
  OAI22_X1 U5739 ( .A1(n6265), .A2(n5485), .B1(n5030), .B2(n6149), .ZN(n4584)
         );
  AOI21_X1 U5740 ( .B1(INSTQUEUE_REG_5__3__SCAN_IN), .B2(n4603), .A(n4584), 
        .ZN(n4586) );
  NAND2_X1 U5741 ( .A1(n6261), .A2(n4604), .ZN(n4585) );
  OAI211_X1 U5742 ( .C1(n6193), .C2(n4607), .A(n4586), .B(n4585), .ZN(U3063)
         );
  OAI22_X1 U5743 ( .A1(n6219), .A2(n5485), .B1(n5030), .B2(n6271), .ZN(n4587)
         );
  AOI21_X1 U5744 ( .B1(INSTQUEUE_REG_5__4__SCAN_IN), .B2(n4603), .A(n4587), 
        .ZN(n4589) );
  NAND2_X1 U5745 ( .A1(n6267), .A2(n4604), .ZN(n4588) );
  OAI211_X1 U5746 ( .C1(n6196), .C2(n4607), .A(n4589), .B(n4588), .ZN(U3064)
         );
  OAI22_X1 U5747 ( .A1(n6247), .A2(n5485), .B1(n5030), .B2(n4918), .ZN(n4590)
         );
  AOI21_X1 U5748 ( .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(n4603), .A(n4590), 
        .ZN(n4592) );
  NAND2_X1 U5749 ( .A1(n2958), .A2(n4604), .ZN(n4591) );
  OAI211_X1 U5750 ( .C1(n6181), .C2(n4607), .A(n4592), .B(n4591), .ZN(U3060)
         );
  OAI22_X1 U5751 ( .A1(n6259), .A2(n5485), .B1(n5030), .B2(n4925), .ZN(n4593)
         );
  AOI21_X1 U5752 ( .B1(INSTQUEUE_REG_5__2__SCAN_IN), .B2(n4603), .A(n4593), 
        .ZN(n4595) );
  NAND2_X1 U5753 ( .A1(n6255), .A2(n4604), .ZN(n4594) );
  OAI211_X1 U5754 ( .C1(n6189), .C2(n4607), .A(n4595), .B(n4594), .ZN(U3062)
         );
  OAI22_X1 U5755 ( .A1(n6295), .A2(n5485), .B1(n5030), .B2(n6165), .ZN(n4596)
         );
  AOI21_X1 U5756 ( .B1(INSTQUEUE_REG_5__7__SCAN_IN), .B2(n4603), .A(n4596), 
        .ZN(n4598) );
  NAND2_X1 U5757 ( .A1(n6288), .A2(n4604), .ZN(n4597) );
  OAI211_X1 U5758 ( .C1(n6211), .C2(n4607), .A(n4598), .B(n4597), .ZN(U3067)
         );
  OAI22_X1 U5759 ( .A1(n6228), .A2(n5485), .B1(n5030), .B2(n6279), .ZN(n4599)
         );
  AOI21_X1 U5760 ( .B1(INSTQUEUE_REG_5__5__SCAN_IN), .B2(n4603), .A(n4599), 
        .ZN(n4601) );
  NAND2_X1 U5761 ( .A1(n6274), .A2(n4604), .ZN(n4600) );
  OAI211_X1 U5762 ( .C1(n6199), .C2(n4607), .A(n4601), .B(n4600), .ZN(U3065)
         );
  OAI22_X1 U5763 ( .A1(n6144), .A2(n5485), .B1(n5030), .B2(n6253), .ZN(n4602)
         );
  AOI21_X1 U5764 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(n4603), .A(n4602), 
        .ZN(n4606) );
  NAND2_X1 U5765 ( .A1(n6249), .A2(n4604), .ZN(n4605) );
  OAI211_X1 U5766 ( .C1(n6185), .C2(n4607), .A(n4606), .B(n4605), .ZN(U3061)
         );
  OAI21_X1 U5767 ( .B1(n2975), .B2(n4610), .A(n4609), .ZN(n5971) );
  AOI22_X1 U5768 ( .A1(n5042), .A2(DATAI_9_), .B1(n5861), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4611) );
  OAI21_X1 U5769 ( .B1(n5971), .B2(n5858), .A(n4611), .ZN(U2882) );
  NOR2_X1 U5770 ( .A1(n4446), .A2(n4447), .ZN(n4612) );
  OAI21_X1 U5771 ( .B1(n4615), .B2(n6238), .A(n5001), .ZN(n4617) );
  OR2_X1 U5772 ( .A1(n4852), .A2(n5812), .ZN(n4727) );
  NAND3_X1 U5773 ( .A1(n6490), .A2(n6309), .A3(n6303), .ZN(n4728) );
  NOR2_X1 U5774 ( .A1(n4997), .A2(n4728), .ZN(n4644) );
  INV_X1 U5775 ( .A(n4644), .ZN(n4613) );
  OAI21_X1 U5776 ( .B1(n4727), .B2(n3712), .A(n4613), .ZN(n4616) );
  INV_X1 U5777 ( .A(n4728), .ZN(n4614) );
  AOI22_X1 U5778 ( .A1(n4617), .A2(n4616), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4614), .ZN(n4646) );
  NAND2_X1 U5779 ( .A1(n4615), .A2(n4906), .ZN(n4936) );
  INV_X1 U5780 ( .A(n4616), .ZN(n4618) );
  AOI22_X1 U5781 ( .A1(n4618), .A2(n4617), .B1(n4728), .B2(n6238), .ZN(n4619)
         );
  NAND2_X1 U5782 ( .A1(n6175), .A2(n4619), .ZN(n4641) );
  AOI22_X1 U5783 ( .A1(n4907), .A2(n6230), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n4641), .ZN(n4620) );
  OAI21_X1 U5784 ( .B1(n6247), .B2(n4757), .A(n4620), .ZN(n4621) );
  AOI21_X1 U5785 ( .B1(n2958), .B2(n4644), .A(n4621), .ZN(n4622) );
  OAI21_X1 U5786 ( .B1(n6181), .B2(n4646), .A(n4622), .ZN(U3028) );
  AOI22_X1 U5787 ( .A1(n4907), .A2(n6287), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n4641), .ZN(n4623) );
  OAI21_X1 U5788 ( .B1(n6295), .B2(n4757), .A(n4623), .ZN(n4624) );
  AOI21_X1 U5789 ( .B1(n6288), .B2(n4644), .A(n4624), .ZN(n4625) );
  OAI21_X1 U5790 ( .B1(n6211), .B2(n4646), .A(n4625), .ZN(U3035) );
  AOI22_X1 U5791 ( .A1(n4907), .A2(n6254), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n4641), .ZN(n4626) );
  OAI21_X1 U5792 ( .B1(n6259), .B2(n4757), .A(n4626), .ZN(n4627) );
  AOI21_X1 U5793 ( .B1(n6255), .B2(n4644), .A(n4627), .ZN(n4628) );
  OAI21_X1 U5794 ( .B1(n6189), .B2(n4646), .A(n4628), .ZN(U3030) );
  AOI22_X1 U5795 ( .A1(n4907), .A2(n6280), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n4641), .ZN(n4629) );
  OAI21_X1 U5796 ( .B1(n6285), .B2(n4757), .A(n4629), .ZN(n4630) );
  AOI21_X1 U5797 ( .B1(n6281), .B2(n4644), .A(n4630), .ZN(n4631) );
  OAI21_X1 U5798 ( .B1(n6203), .B2(n4646), .A(n4631), .ZN(U3034) );
  AOI22_X1 U5799 ( .A1(n4907), .A2(n6216), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n4641), .ZN(n4632) );
  OAI21_X1 U5800 ( .B1(n6219), .B2(n4757), .A(n4632), .ZN(n4633) );
  AOI21_X1 U5801 ( .B1(n6267), .B2(n4644), .A(n4633), .ZN(n4634) );
  OAI21_X1 U5802 ( .B1(n6196), .B2(n4646), .A(n4634), .ZN(U3032) );
  AOI22_X1 U5803 ( .A1(n4907), .A2(n6223), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n4641), .ZN(n4635) );
  OAI21_X1 U5804 ( .B1(n6228), .B2(n4757), .A(n4635), .ZN(n4636) );
  AOI21_X1 U5805 ( .B1(n6274), .B2(n4644), .A(n4636), .ZN(n4637) );
  OAI21_X1 U5806 ( .B1(n6199), .B2(n4646), .A(n4637), .ZN(U3033) );
  AOI22_X1 U5807 ( .A1(n4907), .A2(n6182), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n4641), .ZN(n4638) );
  OAI21_X1 U5808 ( .B1(n6144), .B2(n4757), .A(n4638), .ZN(n4639) );
  AOI21_X1 U5809 ( .B1(n6249), .B2(n4644), .A(n4639), .ZN(n4640) );
  OAI21_X1 U5810 ( .B1(n6185), .B2(n4646), .A(n4640), .ZN(U3029) );
  AOI22_X1 U5811 ( .A1(n4907), .A2(n6260), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n4641), .ZN(n4642) );
  OAI21_X1 U5812 ( .B1(n6265), .B2(n4757), .A(n4642), .ZN(n4643) );
  AOI21_X1 U5813 ( .B1(n6261), .B2(n4644), .A(n4643), .ZN(n4645) );
  OAI21_X1 U5814 ( .B1(n6193), .B2(n4646), .A(n4645), .ZN(U3031) );
  INV_X1 U5815 ( .A(n4763), .ZN(n4647) );
  NOR2_X1 U5816 ( .A1(n4647), .A2(n6238), .ZN(n5482) );
  OR2_X1 U5817 ( .A1(n4724), .A2(n4723), .ZN(n4651) );
  INV_X1 U5818 ( .A(n4651), .ZN(n4843) );
  AND2_X1 U5819 ( .A1(n4649), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5479) );
  AOI22_X1 U5820 ( .A1(n5482), .A2(n5812), .B1(n4843), .B2(n5479), .ZN(n4680)
         );
  NAND2_X1 U5821 ( .A1(n4685), .A2(n3709), .ZN(n4768) );
  AOI21_X1 U5822 ( .B1(n4768), .B2(n6278), .A(n4534), .ZN(n4648) );
  AOI211_X1 U5823 ( .C1(n4763), .C2(n6167), .A(n6238), .B(n4648), .ZN(n4653)
         );
  NOR2_X1 U5824 ( .A1(n6490), .A2(n4765), .ZN(n4771) );
  AND2_X1 U5825 ( .A1(n4997), .A2(n4771), .ZN(n4677) );
  OR2_X1 U5826 ( .A1(n4649), .A2(n6326), .ZN(n4687) );
  AOI21_X1 U5827 ( .B1(n4651), .B2(STATE2_REG_2__SCAN_IN), .A(n4650), .ZN(
        n4847) );
  OAI211_X1 U5828 ( .C1(n4193), .C2(n4677), .A(n4687), .B(n4847), .ZN(n4652)
         );
  NAND2_X1 U5829 ( .A1(n4675), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4656)
         );
  OAI22_X1 U5830 ( .A1(n4768), .A2(n4925), .B1(n6278), .B2(n6259), .ZN(n4654)
         );
  AOI21_X1 U5831 ( .B1(n6255), .B2(n4677), .A(n4654), .ZN(n4655) );
  OAI211_X1 U5832 ( .C1(n4680), .C2(n6189), .A(n4656), .B(n4655), .ZN(U3118)
         );
  NAND2_X1 U5833 ( .A1(n4675), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4659)
         );
  OAI22_X1 U5834 ( .A1(n4768), .A2(n6271), .B1(n6278), .B2(n6219), .ZN(n4657)
         );
  AOI21_X1 U5835 ( .B1(n6267), .B2(n4677), .A(n4657), .ZN(n4658) );
  OAI211_X1 U5836 ( .C1(n4680), .C2(n6196), .A(n4659), .B(n4658), .ZN(U3120)
         );
  NAND2_X1 U5837 ( .A1(n4675), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4662)
         );
  OAI22_X1 U5838 ( .A1(n4768), .A2(n6149), .B1(n6278), .B2(n6265), .ZN(n4660)
         );
  AOI21_X1 U5839 ( .B1(n6261), .B2(n4677), .A(n4660), .ZN(n4661) );
  OAI211_X1 U5840 ( .C1(n4680), .C2(n6193), .A(n4662), .B(n4661), .ZN(U3119)
         );
  NAND2_X1 U5841 ( .A1(n4675), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4665)
         );
  OAI22_X1 U5842 ( .A1(n4768), .A2(n4918), .B1(n6278), .B2(n6247), .ZN(n4663)
         );
  AOI21_X1 U5843 ( .B1(n2958), .B2(n4677), .A(n4663), .ZN(n4664) );
  OAI211_X1 U5844 ( .C1(n4680), .C2(n6181), .A(n4665), .B(n4664), .ZN(U3116)
         );
  NAND2_X1 U5845 ( .A1(n4675), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4668)
         );
  OAI22_X1 U5846 ( .A1(n4768), .A2(n6253), .B1(n6278), .B2(n6144), .ZN(n4666)
         );
  AOI21_X1 U5847 ( .B1(n6249), .B2(n4677), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5848 ( .C1(n4680), .C2(n6185), .A(n4668), .B(n4667), .ZN(U3117)
         );
  NAND2_X1 U5849 ( .A1(n4675), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4671)
         );
  OAI22_X1 U5850 ( .A1(n4768), .A2(n6158), .B1(n6278), .B2(n6285), .ZN(n4669)
         );
  AOI21_X1 U5851 ( .B1(n6281), .B2(n4677), .A(n4669), .ZN(n4670) );
  OAI211_X1 U5852 ( .C1(n4680), .C2(n6203), .A(n4671), .B(n4670), .ZN(U3122)
         );
  NAND2_X1 U5853 ( .A1(n4675), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4674)
         );
  OAI22_X1 U5854 ( .A1(n4768), .A2(n6165), .B1(n6278), .B2(n6295), .ZN(n4672)
         );
  AOI21_X1 U5855 ( .B1(n6288), .B2(n4677), .A(n4672), .ZN(n4673) );
  OAI211_X1 U5856 ( .C1(n4680), .C2(n6211), .A(n4674), .B(n4673), .ZN(U3123)
         );
  NAND2_X1 U5857 ( .A1(n4675), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4679)
         );
  OAI22_X1 U5858 ( .A1(n4768), .A2(n6279), .B1(n6278), .B2(n6228), .ZN(n4676)
         );
  AOI21_X1 U5859 ( .B1(n6274), .B2(n4677), .A(n4676), .ZN(n4678) );
  OAI211_X1 U5860 ( .C1(n4680), .C2(n6199), .A(n4679), .B(n4678), .ZN(U3121)
         );
  AOI21_X1 U5861 ( .B1(n4682), .B2(n4681), .A(n4896), .ZN(n6043) );
  INV_X1 U5862 ( .A(n6043), .ZN(n4683) );
  INV_X1 U5863 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5754) );
  OAI222_X1 U5864 ( .A1(n4683), .A2(n5267), .B1(n5852), .B2(n5754), .C1(n5264), 
        .C2(n5971), .ZN(U2850) );
  NAND2_X1 U5865 ( .A1(n6169), .A2(n5812), .ZN(n4686) );
  INV_X1 U5866 ( .A(n4686), .ZN(n4684) );
  INV_X1 U5867 ( .A(n4724), .ZN(n4902) );
  NOR2_X1 U5868 ( .A1(n4902), .A2(n6490), .ZN(n4783) );
  AOI22_X1 U5869 ( .A1(n4684), .A2(n6233), .B1(n4783), .B2(n5479), .ZN(n4720)
         );
  AOI21_X1 U5870 ( .B1(n4835), .B2(n4715), .A(n4534), .ZN(n4692) );
  NAND2_X1 U5871 ( .A1(n4686), .A2(n6233), .ZN(n4691) );
  INV_X1 U5872 ( .A(n4687), .ZN(n5490) );
  OAI21_X1 U5873 ( .B1(n4724), .B2(n6326), .A(n4729), .ZN(n4784) );
  NOR2_X1 U5874 ( .A1(n5490), .A2(n4784), .ZN(n5005) );
  NOR2_X1 U5875 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4688), .ZN(n4717)
         );
  INV_X1 U5876 ( .A(n4717), .ZN(n4689) );
  AOI21_X1 U5877 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4689), .A(n6490), .ZN(
        n4690) );
  NAND2_X1 U5878 ( .A1(n4714), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4695)
         );
  OAI22_X1 U5879 ( .A1(n6219), .A2(n4835), .B1(n4715), .B2(n6271), .ZN(n4693)
         );
  AOI21_X1 U5880 ( .B1(n6267), .B2(n4717), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5881 ( .C1(n4720), .C2(n6196), .A(n4695), .B(n4694), .ZN(U3136)
         );
  NAND2_X1 U5882 ( .A1(n4714), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4698)
         );
  OAI22_X1 U5883 ( .A1(n6247), .A2(n4835), .B1(n4715), .B2(n4918), .ZN(n4696)
         );
  AOI21_X1 U5884 ( .B1(n2958), .B2(n4717), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5885 ( .C1(n4720), .C2(n6181), .A(n4698), .B(n4697), .ZN(U3132)
         );
  NAND2_X1 U5886 ( .A1(n4714), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4701)
         );
  OAI22_X1 U5887 ( .A1(n6285), .A2(n4835), .B1(n4715), .B2(n6158), .ZN(n4699)
         );
  AOI21_X1 U5888 ( .B1(n6281), .B2(n4717), .A(n4699), .ZN(n4700) );
  OAI211_X1 U5889 ( .C1(n4720), .C2(n6203), .A(n4701), .B(n4700), .ZN(U3138)
         );
  NAND2_X1 U5890 ( .A1(n4714), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4704)
         );
  OAI22_X1 U5891 ( .A1(n6295), .A2(n4835), .B1(n4715), .B2(n6165), .ZN(n4702)
         );
  AOI21_X1 U5892 ( .B1(n6288), .B2(n4717), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5893 ( .C1(n4720), .C2(n6211), .A(n4704), .B(n4703), .ZN(U3139)
         );
  NAND2_X1 U5894 ( .A1(n4714), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4707)
         );
  OAI22_X1 U5895 ( .A1(n6259), .A2(n4835), .B1(n4715), .B2(n4925), .ZN(n4705)
         );
  AOI21_X1 U5896 ( .B1(n6255), .B2(n4717), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5897 ( .C1(n4720), .C2(n6189), .A(n4707), .B(n4706), .ZN(U3134)
         );
  NAND2_X1 U5898 ( .A1(n4714), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4710)
         );
  OAI22_X1 U5899 ( .A1(n6144), .A2(n4835), .B1(n4715), .B2(n6253), .ZN(n4708)
         );
  AOI21_X1 U5900 ( .B1(n6249), .B2(n4717), .A(n4708), .ZN(n4709) );
  OAI211_X1 U5901 ( .C1(n4720), .C2(n6185), .A(n4710), .B(n4709), .ZN(U3133)
         );
  NAND2_X1 U5902 ( .A1(n4714), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4713)
         );
  OAI22_X1 U5903 ( .A1(n6228), .A2(n4835), .B1(n4715), .B2(n6279), .ZN(n4711)
         );
  AOI21_X1 U5904 ( .B1(n6274), .B2(n4717), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5905 ( .C1(n4720), .C2(n6199), .A(n4713), .B(n4712), .ZN(U3137)
         );
  NAND2_X1 U5906 ( .A1(n4714), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4719)
         );
  OAI22_X1 U5907 ( .A1(n6265), .A2(n4835), .B1(n4715), .B2(n6149), .ZN(n4716)
         );
  AOI21_X1 U5908 ( .B1(n6261), .B2(n4717), .A(n4716), .ZN(n4718) );
  OAI211_X1 U5909 ( .C1(n4720), .C2(n6193), .A(n4719), .B(n4718), .ZN(U3135)
         );
  AOI22_X1 U5910 ( .A1(n5042), .A2(DATAI_7_), .B1(n5861), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4721) );
  OAI21_X1 U5911 ( .B1(n4722), .B2(n5858), .A(n4721), .ZN(U2884) );
  INV_X1 U5912 ( .A(n4727), .ZN(n4726) );
  INV_X1 U5913 ( .A(n4723), .ZN(n4725) );
  NOR2_X1 U5914 ( .A1(n4725), .A2(n4724), .ZN(n5480) );
  AOI22_X1 U5915 ( .A1(n4726), .A2(n6233), .B1(n5490), .B2(n5480), .ZN(n4762)
         );
  AOI21_X1 U5916 ( .B1(n4757), .B2(n4756), .A(n4534), .ZN(n4733) );
  NAND2_X1 U5917 ( .A1(n4727), .A2(n6233), .ZN(n4732) );
  NOR2_X1 U5918 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4728), .ZN(n4759)
         );
  INV_X1 U5919 ( .A(n4759), .ZN(n4730) );
  OAI21_X1 U5920 ( .B1(n5480), .B2(n6326), .A(n4729), .ZN(n5488) );
  AOI211_X1 U5921 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4730), .A(n5479), .B(
        n5488), .ZN(n4731) );
  NAND2_X1 U5922 ( .A1(n4755), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4736) );
  OAI22_X1 U5923 ( .A1(n4757), .A2(n4918), .B1(n4756), .B2(n6247), .ZN(n4734)
         );
  AOI21_X1 U5924 ( .B1(n2958), .B2(n4759), .A(n4734), .ZN(n4735) );
  OAI211_X1 U5925 ( .C1(n4762), .C2(n6181), .A(n4736), .B(n4735), .ZN(U3020)
         );
  NAND2_X1 U5926 ( .A1(n4755), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4739) );
  OAI22_X1 U5927 ( .A1(n4757), .A2(n6279), .B1(n4756), .B2(n6228), .ZN(n4737)
         );
  AOI21_X1 U5928 ( .B1(n6274), .B2(n4759), .A(n4737), .ZN(n4738) );
  OAI211_X1 U5929 ( .C1(n4762), .C2(n6199), .A(n4739), .B(n4738), .ZN(U3025)
         );
  NAND2_X1 U5930 ( .A1(n4755), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4742) );
  OAI22_X1 U5931 ( .A1(n4757), .A2(n6158), .B1(n4756), .B2(n6285), .ZN(n4740)
         );
  AOI21_X1 U5932 ( .B1(n6281), .B2(n4759), .A(n4740), .ZN(n4741) );
  OAI211_X1 U5933 ( .C1(n4762), .C2(n6203), .A(n4742), .B(n4741), .ZN(U3026)
         );
  NAND2_X1 U5934 ( .A1(n4755), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4745) );
  OAI22_X1 U5935 ( .A1(n4757), .A2(n6253), .B1(n4756), .B2(n6144), .ZN(n4743)
         );
  AOI21_X1 U5936 ( .B1(n6249), .B2(n4759), .A(n4743), .ZN(n4744) );
  OAI211_X1 U5937 ( .C1(n4762), .C2(n6185), .A(n4745), .B(n4744), .ZN(U3021)
         );
  NAND2_X1 U5938 ( .A1(n4755), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4748) );
  OAI22_X1 U5939 ( .A1(n4757), .A2(n4925), .B1(n4756), .B2(n6259), .ZN(n4746)
         );
  AOI21_X1 U5940 ( .B1(n6255), .B2(n4759), .A(n4746), .ZN(n4747) );
  OAI211_X1 U5941 ( .C1(n4762), .C2(n6189), .A(n4748), .B(n4747), .ZN(U3022)
         );
  NAND2_X1 U5942 ( .A1(n4755), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4751) );
  OAI22_X1 U5943 ( .A1(n4757), .A2(n6271), .B1(n4756), .B2(n6219), .ZN(n4749)
         );
  AOI21_X1 U5944 ( .B1(n6267), .B2(n4759), .A(n4749), .ZN(n4750) );
  OAI211_X1 U5945 ( .C1(n4762), .C2(n6196), .A(n4751), .B(n4750), .ZN(U3024)
         );
  NAND2_X1 U5946 ( .A1(n4755), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4754) );
  OAI22_X1 U5947 ( .A1(n4757), .A2(n6149), .B1(n4756), .B2(n6265), .ZN(n4752)
         );
  AOI21_X1 U5948 ( .B1(n6261), .B2(n4759), .A(n4752), .ZN(n4753) );
  OAI211_X1 U5949 ( .C1(n4762), .C2(n6193), .A(n4754), .B(n4753), .ZN(U3023)
         );
  NAND2_X1 U5950 ( .A1(n4755), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4761) );
  OAI22_X1 U5951 ( .A1(n4757), .A2(n6165), .B1(n4756), .B2(n6295), .ZN(n4758)
         );
  AOI21_X1 U5952 ( .B1(n6288), .B2(n4759), .A(n4758), .ZN(n4760) );
  OAI211_X1 U5953 ( .C1(n4762), .C2(n6211), .A(n4761), .B(n4760), .ZN(U3027)
         );
  AND2_X1 U5954 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4771), .ZN(n4837)
         );
  AOI21_X1 U5955 ( .B1(n4764), .B2(n4763), .A(n4837), .ZN(n4770) );
  NAND2_X1 U5956 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4766) );
  OAI22_X1 U5957 ( .A1(n4770), .A2(n6238), .B1(n4766), .B2(n4765), .ZN(n4767)
         );
  NAND2_X1 U5958 ( .A1(n4770), .A2(n4769), .ZN(n4774) );
  INV_X1 U5959 ( .A(n4771), .ZN(n4772) );
  NAND2_X1 U5960 ( .A1(n6238), .A2(n4772), .ZN(n4773) );
  OAI211_X1 U5961 ( .C1(n6238), .C2(n4774), .A(n6175), .B(n4773), .ZN(n4832)
         );
  AOI22_X1 U5962 ( .A1(n4833), .A2(n6190), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4832), .ZN(n4775) );
  OAI21_X1 U5963 ( .B1(n6149), .B2(n4835), .A(n4775), .ZN(n4776) );
  AOI21_X1 U5964 ( .B1(n6261), .B2(n4837), .A(n4776), .ZN(n4777) );
  OAI21_X1 U5965 ( .B1(n6193), .B2(n4839), .A(n4777), .ZN(U3127) );
  AOI22_X1 U5966 ( .A1(n4833), .A2(n6248), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4832), .ZN(n4778) );
  OAI21_X1 U5967 ( .B1(n6253), .B2(n4835), .A(n4778), .ZN(n4779) );
  AOI21_X1 U5968 ( .B1(n6249), .B2(n4837), .A(n4779), .ZN(n4780) );
  OAI21_X1 U5969 ( .B1(n6185), .B2(n4839), .A(n4780), .ZN(U3125) );
  AOI21_X1 U5970 ( .B1(n4811), .B2(n6294), .A(n4534), .ZN(n4782) );
  NOR2_X1 U5971 ( .A1(n4782), .A2(n6238), .ZN(n4787) );
  AND2_X1 U5972 ( .A1(n4416), .A2(n4455), .ZN(n4901) );
  AND2_X1 U5973 ( .A1(n4901), .A2(n5812), .ZN(n6236) );
  AOI22_X1 U5974 ( .A1(n4787), .A2(n6236), .B1(n5490), .B2(n4783), .ZN(n4816)
         );
  NOR2_X1 U5975 ( .A1(n5479), .A2(n4784), .ZN(n4910) );
  INV_X1 U5976 ( .A(n6236), .ZN(n4786) );
  NAND3_X1 U5977 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6309), .ZN(n6241) );
  NOR2_X1 U5978 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6241), .ZN(n4813)
         );
  INV_X1 U5979 ( .A(n4813), .ZN(n4785) );
  AOI22_X1 U5980 ( .A1(n4787), .A2(n4786), .B1(n4785), .B2(
        STATE2_REG_3__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U5981 ( .A1(n4810), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4791)
         );
  OAI22_X1 U5982 ( .A1(n4811), .A2(n6144), .B1(n6294), .B2(n6253), .ZN(n4789)
         );
  AOI21_X1 U5983 ( .B1(n4813), .B2(n6249), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5984 ( .C1(n4816), .C2(n6185), .A(n4791), .B(n4790), .ZN(U3101)
         );
  NAND2_X1 U5985 ( .A1(n4810), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4794)
         );
  OAI22_X1 U5986 ( .A1(n4811), .A2(n6247), .B1(n6294), .B2(n4918), .ZN(n4792)
         );
  AOI21_X1 U5987 ( .B1(n2958), .B2(n4813), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5988 ( .C1(n4816), .C2(n6181), .A(n4794), .B(n4793), .ZN(U3100)
         );
  NAND2_X1 U5989 ( .A1(n4810), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4797)
         );
  OAI22_X1 U5990 ( .A1(n4811), .A2(n6295), .B1(n6294), .B2(n6165), .ZN(n4795)
         );
  AOI21_X1 U5991 ( .B1(n4813), .B2(n6288), .A(n4795), .ZN(n4796) );
  OAI211_X1 U5992 ( .C1(n4816), .C2(n6211), .A(n4797), .B(n4796), .ZN(U3107)
         );
  NAND2_X1 U5993 ( .A1(n4810), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4800)
         );
  OAI22_X1 U5994 ( .A1(n4811), .A2(n6219), .B1(n6294), .B2(n6271), .ZN(n4798)
         );
  AOI21_X1 U5995 ( .B1(n4813), .B2(n6267), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5996 ( .C1(n4816), .C2(n6196), .A(n4800), .B(n4799), .ZN(U3104)
         );
  NAND2_X1 U5997 ( .A1(n4810), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4803)
         );
  OAI22_X1 U5998 ( .A1(n4811), .A2(n6265), .B1(n6294), .B2(n6149), .ZN(n4801)
         );
  AOI21_X1 U5999 ( .B1(n4813), .B2(n6261), .A(n4801), .ZN(n4802) );
  OAI211_X1 U6000 ( .C1(n4816), .C2(n6193), .A(n4803), .B(n4802), .ZN(U3103)
         );
  NAND2_X1 U6001 ( .A1(n4810), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4806)
         );
  OAI22_X1 U6002 ( .A1(n4811), .A2(n6259), .B1(n6294), .B2(n4925), .ZN(n4804)
         );
  AOI21_X1 U6003 ( .B1(n4813), .B2(n6255), .A(n4804), .ZN(n4805) );
  OAI211_X1 U6004 ( .C1(n4816), .C2(n6189), .A(n4806), .B(n4805), .ZN(U3102)
         );
  NAND2_X1 U6005 ( .A1(n4810), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4809)
         );
  OAI22_X1 U6006 ( .A1(n4811), .A2(n6285), .B1(n6294), .B2(n6158), .ZN(n4807)
         );
  AOI21_X1 U6007 ( .B1(n4813), .B2(n6281), .A(n4807), .ZN(n4808) );
  OAI211_X1 U6008 ( .C1(n4816), .C2(n6203), .A(n4809), .B(n4808), .ZN(U3106)
         );
  NAND2_X1 U6009 ( .A1(n4810), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4815)
         );
  OAI22_X1 U6010 ( .A1(n4811), .A2(n6228), .B1(n6294), .B2(n6279), .ZN(n4812)
         );
  AOI21_X1 U6011 ( .B1(n4813), .B2(n6274), .A(n4812), .ZN(n4814) );
  OAI211_X1 U6012 ( .C1(n4816), .C2(n6199), .A(n4815), .B(n4814), .ZN(U3105)
         );
  AOI22_X1 U6013 ( .A1(n4833), .A2(n6186), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4832), .ZN(n4817) );
  OAI21_X1 U6014 ( .B1(n4925), .B2(n4835), .A(n4817), .ZN(n4818) );
  AOI21_X1 U6015 ( .B1(n6255), .B2(n4837), .A(n4818), .ZN(n4819) );
  OAI21_X1 U6016 ( .B1(n6189), .B2(n4839), .A(n4819), .ZN(U3126) );
  AOI22_X1 U6017 ( .A1(n4833), .A2(n6272), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4832), .ZN(n4820) );
  OAI21_X1 U6018 ( .B1(n6279), .B2(n4835), .A(n4820), .ZN(n4821) );
  AOI21_X1 U6019 ( .B1(n6274), .B2(n4837), .A(n4821), .ZN(n4822) );
  OAI21_X1 U6020 ( .B1(n6199), .B2(n4839), .A(n4822), .ZN(U3129) );
  AOI22_X1 U6021 ( .A1(n4833), .A2(n6205), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4832), .ZN(n4823) );
  OAI21_X1 U6022 ( .B1(n6165), .B2(n4835), .A(n4823), .ZN(n4824) );
  AOI21_X1 U6023 ( .B1(n6288), .B2(n4837), .A(n4824), .ZN(n4825) );
  OAI21_X1 U6024 ( .B1(n6211), .B2(n4839), .A(n4825), .ZN(U3131) );
  AOI22_X1 U6025 ( .A1(n4833), .A2(n6200), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4832), .ZN(n4826) );
  OAI21_X1 U6026 ( .B1(n6158), .B2(n4835), .A(n4826), .ZN(n4827) );
  AOI21_X1 U6027 ( .B1(n6281), .B2(n4837), .A(n4827), .ZN(n4828) );
  OAI21_X1 U6028 ( .B1(n6203), .B2(n4839), .A(n4828), .ZN(U3130) );
  AOI22_X1 U6029 ( .A1(n4833), .A2(n6178), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4832), .ZN(n4829) );
  OAI21_X1 U6030 ( .B1(n4918), .B2(n4835), .A(n4829), .ZN(n4830) );
  AOI21_X1 U6031 ( .B1(n2958), .B2(n4837), .A(n4830), .ZN(n4831) );
  OAI21_X1 U6032 ( .B1(n6181), .B2(n4839), .A(n4831), .ZN(U3124) );
  AOI22_X1 U6033 ( .A1(n4833), .A2(n6266), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4832), .ZN(n4834) );
  OAI21_X1 U6034 ( .B1(n6271), .B2(n4835), .A(n4834), .ZN(n4836) );
  AOI21_X1 U6035 ( .B1(n6267), .B2(n4837), .A(n4836), .ZN(n4838) );
  OAI21_X1 U6036 ( .B1(n6196), .B2(n4839), .A(n4838), .ZN(U3128) );
  OAI222_X1 U6037 ( .A1(n4840), .A2(n5858), .B1(n4841), .B2(n5925), .C1(n5109), 
        .C2(n3722), .ZN(U2889) );
  INV_X1 U6038 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6517) );
  OAI222_X1 U6039 ( .A1(n5996), .A2(n5858), .B1(n4841), .B2(n5931), .C1(n5109), 
        .C2(n6517), .ZN(U2885) );
  NAND3_X1 U6040 ( .A1(n4842), .A2(n6233), .A3(n5812), .ZN(n4845) );
  NAND2_X1 U6041 ( .A1(n5490), .A2(n4843), .ZN(n4844) );
  AND2_X1 U6042 ( .A1(n4845), .A2(n4844), .ZN(n6213) );
  NOR2_X1 U6043 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4846), .ZN(n6220)
         );
  INV_X1 U6044 ( .A(n5479), .ZN(n4848) );
  OAI211_X1 U6045 ( .C1(n4193), .C2(n6220), .A(n4848), .B(n4847), .ZN(n4849)
         );
  INV_X1 U6046 ( .A(n4849), .ZN(n4854) );
  OAI21_X1 U6047 ( .B1(n6222), .B2(n6207), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4851) );
  OAI211_X1 U6048 ( .C1(n5481), .C2(n4852), .A(n4851), .B(n6233), .ZN(n4853)
         );
  NAND2_X1 U6049 ( .A1(n6224), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4857) );
  INV_X1 U6050 ( .A(n6222), .ZN(n4867) );
  OAI22_X1 U6051 ( .A1(n4867), .A2(n6253), .B1(n6144), .B2(n6227), .ZN(n4855)
         );
  AOI21_X1 U6052 ( .B1(n6249), .B2(n6220), .A(n4855), .ZN(n4856) );
  OAI211_X1 U6053 ( .C1(n6213), .C2(n6185), .A(n4857), .B(n4856), .ZN(U3085)
         );
  NAND2_X1 U6054 ( .A1(n6224), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4860) );
  OAI22_X1 U6055 ( .A1(n4867), .A2(n6158), .B1(n6285), .B2(n6227), .ZN(n4858)
         );
  AOI21_X1 U6056 ( .B1(n6281), .B2(n6220), .A(n4858), .ZN(n4859) );
  OAI211_X1 U6057 ( .C1(n6213), .C2(n6203), .A(n4860), .B(n4859), .ZN(U3090)
         );
  NAND2_X1 U6058 ( .A1(n6224), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4863) );
  OAI22_X1 U6059 ( .A1(n4867), .A2(n6149), .B1(n6265), .B2(n6227), .ZN(n4861)
         );
  AOI21_X1 U6060 ( .B1(n6261), .B2(n6220), .A(n4861), .ZN(n4862) );
  OAI211_X1 U6061 ( .C1(n6213), .C2(n6193), .A(n4863), .B(n4862), .ZN(U3087)
         );
  NAND2_X1 U6062 ( .A1(n6224), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4866) );
  OAI22_X1 U6063 ( .A1(n4867), .A2(n6165), .B1(n6295), .B2(n6227), .ZN(n4864)
         );
  AOI21_X1 U6064 ( .B1(n6288), .B2(n6220), .A(n4864), .ZN(n4865) );
  OAI211_X1 U6065 ( .C1(n6213), .C2(n6211), .A(n4866), .B(n4865), .ZN(U3091)
         );
  NAND2_X1 U6066 ( .A1(n6224), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4870) );
  OAI22_X1 U6067 ( .A1(n4867), .A2(n4918), .B1(n6247), .B2(n6227), .ZN(n4868)
         );
  AOI21_X1 U6068 ( .B1(n2958), .B2(n6220), .A(n4868), .ZN(n4869) );
  OAI211_X1 U6069 ( .C1(n6213), .C2(n6181), .A(n4870), .B(n4869), .ZN(U3084)
         );
  AOI21_X1 U6070 ( .B1(n4609), .B2(n4872), .A(n4871), .ZN(n5739) );
  INV_X1 U6071 ( .A(n5739), .ZN(n4942) );
  AOI22_X1 U6072 ( .A1(n5042), .A2(DATAI_10_), .B1(n5861), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4873) );
  OAI21_X1 U6073 ( .B1(n4942), .B2(n5858), .A(n4873), .ZN(U2881) );
  OAI21_X1 U6074 ( .B1(n4871), .B2(n4875), .A(n4874), .ZN(n5961) );
  INV_X1 U6075 ( .A(n3015), .ZN(n4990) );
  AOI21_X1 U6076 ( .B1(n4876), .B2(n4894), .A(n4990), .ZN(n6036) );
  AOI22_X1 U6077 ( .A1(n5849), .A2(n6036), .B1(n5261), .B2(EBX_REG_11__SCAN_IN), .ZN(n4877) );
  OAI21_X1 U6078 ( .B1(n5961), .B2(n5264), .A(n4877), .ZN(U2848) );
  AOI22_X1 U6079 ( .A1(n5042), .A2(DATAI_11_), .B1(n5861), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4878) );
  OAI21_X1 U6080 ( .B1(n5961), .B2(n5858), .A(n4878), .ZN(U2880) );
  NAND2_X1 U6081 ( .A1(n5954), .A2(n4879), .ZN(n4882) );
  XOR2_X1 U6082 ( .A(n4882), .B(n4881), .Z(n4900) );
  NAND2_X1 U6083 ( .A1(n5739), .A2(n6030), .ZN(n4887) );
  INV_X1 U6084 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4883) );
  OAI22_X1 U6085 ( .A1(n5315), .A2(n4884), .B1(n6071), .B2(n4883), .ZN(n4885)
         );
  AOI21_X1 U6086 ( .B1(n6012), .B2(n5740), .A(n4885), .ZN(n4886) );
  OAI211_X1 U6087 ( .C1(n4900), .C2(n5675), .A(n4887), .B(n4886), .ZN(U2976)
         );
  OAI21_X1 U6088 ( .B1(n6080), .B2(n6112), .A(n4888), .ZN(n6065) );
  INV_X1 U6089 ( .A(n6065), .ZN(n6093) );
  NOR2_X1 U6090 ( .A1(n4890), .A2(n6064), .ZN(n6044) );
  OAI211_X1 U6091 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6044), .B(n4889), .ZN(n4899) );
  INV_X1 U6092 ( .A(n4890), .ZN(n6049) );
  AOI21_X1 U6093 ( .B1(n6107), .B2(n4891), .A(n6066), .ZN(n4892) );
  OAI21_X1 U6094 ( .B1(n6068), .B2(n4893), .A(n4892), .ZN(n6060) );
  INV_X1 U6095 ( .A(n6060), .ZN(n6058) );
  OAI21_X1 U6096 ( .B1(n6122), .B2(n6049), .A(n6058), .ZN(n6042) );
  OAI21_X1 U6097 ( .B1(n4896), .B2(n4895), .A(n4894), .ZN(n5737) );
  OAI22_X1 U6098 ( .A1(n6120), .A2(n5737), .B1(n4883), .B2(n6071), .ZN(n4897)
         );
  AOI21_X1 U6099 ( .B1(n6042), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4897), 
        .ZN(n4898) );
  OAI211_X1 U6100 ( .C1(n4900), .C2(n6083), .A(n4899), .B(n4898), .ZN(U3008)
         );
  NOR2_X1 U6101 ( .A1(n4902), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4996)
         );
  AOI22_X1 U6102 ( .A1(n6134), .A2(n6233), .B1(n5490), .B2(n4996), .ZN(n4941)
         );
  NAND3_X1 U6103 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6490), .A3(n6309), .ZN(n6137) );
  NOR2_X1 U6104 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6137), .ZN(n4938)
         );
  NOR2_X1 U6105 ( .A1(n4446), .A2(n4903), .ZN(n4904) );
  NAND2_X1 U6106 ( .A1(n4905), .A2(n4904), .ZN(n5484) );
  OAI21_X1 U6107 ( .B1(n4907), .B2(n6159), .A(n5001), .ZN(n4909) );
  INV_X1 U6108 ( .A(n6134), .ZN(n4908) );
  NAND2_X1 U6109 ( .A1(n4909), .A2(n4908), .ZN(n4911) );
  NAND2_X1 U6110 ( .A1(n4935), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U6111 ( .A1(n6295), .A2(n4936), .B1(n6155), .B2(n6165), .ZN(n4912)
         );
  AOI21_X1 U6112 ( .B1(n6288), .B2(n4938), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6113 ( .C1(n4941), .C2(n6211), .A(n4914), .B(n4913), .ZN(U3043)
         );
  NAND2_X1 U6114 ( .A1(n4935), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4917) );
  OAI22_X1 U6115 ( .A1(n6265), .A2(n4936), .B1(n6155), .B2(n6149), .ZN(n4915)
         );
  AOI21_X1 U6116 ( .B1(n6261), .B2(n4938), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6117 ( .C1(n4941), .C2(n6193), .A(n4917), .B(n4916), .ZN(U3039)
         );
  NAND2_X1 U6118 ( .A1(n4935), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4921) );
  OAI22_X1 U6119 ( .A1(n6247), .A2(n4936), .B1(n6155), .B2(n4918), .ZN(n4919)
         );
  AOI21_X1 U6120 ( .B1(n2958), .B2(n4938), .A(n4919), .ZN(n4920) );
  OAI211_X1 U6121 ( .C1(n4941), .C2(n6181), .A(n4921), .B(n4920), .ZN(U3036)
         );
  NAND2_X1 U6122 ( .A1(n4935), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4924) );
  OAI22_X1 U6123 ( .A1(n6219), .A2(n4936), .B1(n6155), .B2(n6271), .ZN(n4922)
         );
  AOI21_X1 U6124 ( .B1(n6267), .B2(n4938), .A(n4922), .ZN(n4923) );
  OAI211_X1 U6125 ( .C1(n4941), .C2(n6196), .A(n4924), .B(n4923), .ZN(U3040)
         );
  NAND2_X1 U6126 ( .A1(n4935), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4928) );
  OAI22_X1 U6127 ( .A1(n6259), .A2(n4936), .B1(n6155), .B2(n4925), .ZN(n4926)
         );
  AOI21_X1 U6128 ( .B1(n6255), .B2(n4938), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6129 ( .C1(n4941), .C2(n6189), .A(n4928), .B(n4927), .ZN(U3038)
         );
  NAND2_X1 U6130 ( .A1(n4935), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6131 ( .A1(n6144), .A2(n4936), .B1(n6155), .B2(n6253), .ZN(n4929)
         );
  AOI21_X1 U6132 ( .B1(n6249), .B2(n4938), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6133 ( .C1(n4941), .C2(n6185), .A(n4931), .B(n4930), .ZN(U3037)
         );
  NAND2_X1 U6134 ( .A1(n4935), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6135 ( .A1(n6285), .A2(n4936), .B1(n6155), .B2(n6158), .ZN(n4932)
         );
  AOI21_X1 U6136 ( .B1(n6281), .B2(n4938), .A(n4932), .ZN(n4933) );
  OAI211_X1 U6137 ( .C1(n4941), .C2(n6203), .A(n4934), .B(n4933), .ZN(U3042)
         );
  NAND2_X1 U6138 ( .A1(n4935), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4940) );
  OAI22_X1 U6139 ( .A1(n6228), .A2(n4936), .B1(n6155), .B2(n6279), .ZN(n4937)
         );
  AOI21_X1 U6140 ( .B1(n6274), .B2(n4938), .A(n4937), .ZN(n4939) );
  OAI211_X1 U6141 ( .C1(n4941), .C2(n6199), .A(n4940), .B(n4939), .ZN(U3041)
         );
  INV_X1 U6142 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5736) );
  OAI222_X1 U6143 ( .A1(n5737), .A2(n5267), .B1(n5852), .B2(n5736), .C1(n5264), 
        .C2(n4942), .ZN(U2849) );
  INV_X1 U6144 ( .A(n5123), .ZN(n4945) );
  OR2_X1 U6145 ( .A1(n4943), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U6146 ( .A1(n5780), .A2(n4944), .ZN(n5828) );
  INV_X1 U6147 ( .A(n5828), .ZN(n5844) );
  INV_X1 U6148 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4955) );
  INV_X1 U6149 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6438) );
  NOR2_X1 U6150 ( .A1(n5804), .A2(n6438), .ZN(n4954) );
  NOR2_X1 U6151 ( .A1(n4946), .A2(n4945), .ZN(n4947) );
  NAND2_X1 U6152 ( .A1(n4947), .A2(n3560), .ZN(n5838) );
  NOR2_X1 U6153 ( .A1(n4955), .A2(n5834), .ZN(n4948) );
  NOR2_X1 U6154 ( .A1(n5817), .A2(REIP_REG_1__SCAN_IN), .ZN(n5802) );
  AOI211_X1 U6155 ( .C1(n5821), .C2(EBX_REG_1__SCAN_IN), .A(n4948), .B(n5802), 
        .ZN(n4951) );
  NAND2_X1 U6156 ( .A1(n4949), .A2(n5831), .ZN(n4950) );
  OAI211_X1 U6157 ( .C1(n4952), .C2(n5838), .A(n4951), .B(n4950), .ZN(n4953)
         );
  AOI211_X1 U6158 ( .C1(n5799), .C2(n4955), .A(n4954), .B(n4953), .ZN(n4956)
         );
  OAI21_X1 U6159 ( .B1(n5844), .B2(n4957), .A(n4956), .ZN(U2826) );
  AOI21_X1 U6160 ( .B1(n4874), .B2(n4959), .A(n4958), .ZN(n5723) );
  INV_X1 U6161 ( .A(n5723), .ZN(n4962) );
  AOI22_X1 U6162 ( .A1(n5042), .A2(DATAI_12_), .B1(n5861), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4960) );
  OAI21_X1 U6163 ( .B1(n4962), .B2(n5858), .A(n4960), .ZN(U2879) );
  XNOR2_X1 U6164 ( .A(n4990), .B(n4989), .ZN(n4969) );
  INV_X1 U6165 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4961) );
  OAI222_X1 U6166 ( .A1(n4962), .A2(n5264), .B1(n5267), .B2(n4969), .C1(n4961), 
        .C2(n5852), .ZN(U2847) );
  INV_X1 U6167 ( .A(n4965), .ZN(n4966) );
  NOR2_X1 U6168 ( .A1(n4967), .A2(n4966), .ZN(n4968) );
  XNOR2_X1 U6169 ( .A(n4964), .B(n4968), .ZN(n4984) );
  INV_X1 U6170 ( .A(n4969), .ZN(n5720) );
  INV_X1 U6171 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6390) );
  NOR2_X1 U6172 ( .A1(n6112), .A2(n4970), .ZN(n5429) );
  NAND2_X1 U6173 ( .A1(n6107), .A2(n4971), .ZN(n5055) );
  INV_X1 U6174 ( .A(n5055), .ZN(n4972) );
  NAND3_X1 U6175 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n4975), .A3(n6037), .ZN(n4973) );
  OAI21_X1 U6176 ( .B1(n6071), .B2(n6390), .A(n4973), .ZN(n4978) );
  OAI22_X1 U6177 ( .A1(n6070), .A2(n6066), .B1(n4974), .B2(n6060), .ZN(n6041)
         );
  OAI21_X1 U6178 ( .B1(n6107), .B2(n5429), .A(n5955), .ZN(n4976) );
  AOI21_X1 U6179 ( .B1(n6041), .B2(n4976), .A(n4975), .ZN(n4977) );
  AOI211_X1 U6180 ( .C1(n6106), .C2(n5720), .A(n4978), .B(n4977), .ZN(n4979)
         );
  OAI21_X1 U6181 ( .B1(n4984), .B2(n6083), .A(n4979), .ZN(U3006) );
  NAND2_X1 U6182 ( .A1(n5723), .A2(n6030), .ZN(n4983) );
  OAI22_X1 U6183 ( .A1(n5315), .A2(n4980), .B1(n6071), .B2(n6390), .ZN(n4981)
         );
  AOI21_X1 U6184 ( .B1(n6012), .B2(n5724), .A(n4981), .ZN(n4982) );
  OAI211_X1 U6185 ( .C1(n4984), .C2(n5675), .A(n4983), .B(n4982), .ZN(U2974)
         );
  OAI21_X1 U6186 ( .B1(n4958), .B2(n4987), .A(n4986), .ZN(n5719) );
  AOI21_X1 U6187 ( .B1(n4990), .B2(n4989), .A(n4988), .ZN(n4991) );
  INV_X1 U6188 ( .A(n5065), .ZN(n5045) );
  NOR2_X1 U6189 ( .A1(n4991), .A2(n5045), .ZN(n5710) );
  AOI22_X1 U6190 ( .A1(n5849), .A2(n5710), .B1(n5261), .B2(EBX_REG_13__SCAN_IN), .ZN(n4992) );
  OAI21_X1 U6191 ( .B1(n5719), .B2(n5264), .A(n4992), .ZN(U2846) );
  AOI22_X1 U6192 ( .A1(n5042), .A2(DATAI_13_), .B1(n5861), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4993) );
  OAI21_X1 U6193 ( .B1(n5719), .B2(n5858), .A(n4993), .ZN(U2878) );
  INV_X1 U6194 ( .A(n6169), .ZN(n4994) );
  NOR3_X1 U6195 ( .A1(n4994), .A2(n6238), .A3(n5812), .ZN(n4995) );
  AOI21_X1 U6196 ( .B1(n5479), .B2(n4996), .A(n4995), .ZN(n5034) );
  NAND2_X1 U6197 ( .A1(n4997), .A2(n6177), .ZN(n5004) );
  INV_X1 U6198 ( .A(n5004), .ZN(n5032) );
  INV_X1 U6199 ( .A(n6204), .ZN(n5000) );
  NAND3_X1 U6200 ( .A1(n6233), .A2(n5030), .A3(n5000), .ZN(n5002) );
  AOI21_X1 U6201 ( .B1(n5002), .B2(n5001), .A(n6169), .ZN(n5003) );
  AOI21_X1 U6202 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5004), .A(n5003), .ZN(
        n5006) );
  NAND3_X1 U6203 ( .A1(n6490), .A2(n5006), .A3(n5005), .ZN(n5028) );
  AOI22_X1 U6204 ( .A1(n6204), .A2(n6260), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5028), .ZN(n5007) );
  OAI21_X1 U6205 ( .B1(n5030), .B2(n6265), .A(n5007), .ZN(n5008) );
  AOI21_X1 U6206 ( .B1(n6261), .B2(n5032), .A(n5008), .ZN(n5009) );
  OAI21_X1 U6207 ( .B1(n6193), .B2(n5034), .A(n5009), .ZN(U3071) );
  AOI22_X1 U6208 ( .A1(n6204), .A2(n6216), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5028), .ZN(n5010) );
  OAI21_X1 U6209 ( .B1(n5030), .B2(n6219), .A(n5010), .ZN(n5011) );
  AOI21_X1 U6210 ( .B1(n6267), .B2(n5032), .A(n5011), .ZN(n5012) );
  OAI21_X1 U6211 ( .B1(n6196), .B2(n5034), .A(n5012), .ZN(U3072) );
  AOI22_X1 U6212 ( .A1(n6204), .A2(n6182), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5028), .ZN(n5013) );
  OAI21_X1 U6213 ( .B1(n5030), .B2(n6144), .A(n5013), .ZN(n5014) );
  AOI21_X1 U6214 ( .B1(n6249), .B2(n5032), .A(n5014), .ZN(n5015) );
  OAI21_X1 U6215 ( .B1(n6185), .B2(n5034), .A(n5015), .ZN(U3069) );
  AOI22_X1 U6216 ( .A1(n6204), .A2(n6230), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5028), .ZN(n5016) );
  OAI21_X1 U6217 ( .B1(n5030), .B2(n6247), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6218 ( .B1(n2958), .B2(n5032), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6219 ( .B1(n6181), .B2(n5034), .A(n5018), .ZN(U3068) );
  AOI22_X1 U6220 ( .A1(n6204), .A2(n6223), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5028), .ZN(n5019) );
  OAI21_X1 U6221 ( .B1(n5030), .B2(n6228), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6222 ( .B1(n6274), .B2(n5032), .A(n5020), .ZN(n5021) );
  OAI21_X1 U6223 ( .B1(n6199), .B2(n5034), .A(n5021), .ZN(U3073) );
  AOI22_X1 U6224 ( .A1(n6204), .A2(n6287), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n5028), .ZN(n5022) );
  OAI21_X1 U6225 ( .B1(n5030), .B2(n6295), .A(n5022), .ZN(n5023) );
  AOI21_X1 U6226 ( .B1(n6288), .B2(n5032), .A(n5023), .ZN(n5024) );
  OAI21_X1 U6227 ( .B1(n6211), .B2(n5034), .A(n5024), .ZN(U3075) );
  AOI22_X1 U6228 ( .A1(n6204), .A2(n6280), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n5028), .ZN(n5025) );
  OAI21_X1 U6229 ( .B1(n5030), .B2(n6285), .A(n5025), .ZN(n5026) );
  AOI21_X1 U6230 ( .B1(n6281), .B2(n5032), .A(n5026), .ZN(n5027) );
  OAI21_X1 U6231 ( .B1(n6203), .B2(n5034), .A(n5027), .ZN(U3074) );
  AOI22_X1 U6232 ( .A1(n6204), .A2(n6254), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5028), .ZN(n5029) );
  OAI21_X1 U6233 ( .B1(n5030), .B2(n6259), .A(n5029), .ZN(n5031) );
  AOI21_X1 U6234 ( .B1(n6255), .B2(n5032), .A(n5031), .ZN(n5033) );
  OAI21_X1 U6235 ( .B1(n6189), .B2(n5034), .A(n5033), .ZN(U3070) );
  AOI21_X1 U6236 ( .B1(n4986), .B2(n5036), .A(n5035), .ZN(n5846) );
  INV_X1 U6237 ( .A(n5846), .ZN(n5038) );
  AOI22_X1 U6238 ( .A1(n5042), .A2(DATAI_14_), .B1(n5861), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U6239 ( .B1(n5038), .B2(n5858), .A(n5037), .ZN(U2877) );
  OAI21_X1 U6240 ( .B1(n5035), .B2(n5041), .A(n5040), .ZN(n5700) );
  AOI22_X1 U6241 ( .A1(n5042), .A2(DATAI_15_), .B1(n5861), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5043) );
  OAI21_X1 U6242 ( .B1(n5700), .B2(n5858), .A(n5043), .ZN(U2876) );
  AOI21_X1 U6243 ( .B1(n5045), .B2(n5064), .A(n5044), .ZN(n5046) );
  NOR2_X1 U6244 ( .A1(n5046), .A2(n5081), .ZN(n5696) );
  AOI22_X1 U6245 ( .A1(n5696), .A2(n5849), .B1(n5261), .B2(EBX_REG_15__SCAN_IN), .ZN(n5047) );
  OAI21_X1 U6246 ( .B1(n5700), .B2(n5264), .A(n5047), .ZN(U2844) );
  XNOR2_X1 U6247 ( .A(n3439), .B(n5465), .ZN(n5050) );
  XNOR2_X1 U6248 ( .A(n5049), .B(n5050), .ZN(n5070) );
  NAND2_X1 U6249 ( .A1(n6012), .A2(n5704), .ZN(n5051) );
  NAND2_X1 U6250 ( .A1(n6104), .A2(REIP_REG_14__SCAN_IN), .ZN(n5066) );
  OAI211_X1 U6251 ( .C1(n5315), .C2(n5052), .A(n5051), .B(n5066), .ZN(n5053)
         );
  AOI21_X1 U6252 ( .B1(n5846), .B2(n6030), .A(n5053), .ZN(n5054) );
  OAI21_X1 U6253 ( .B1(n5675), .B2(n5070), .A(n5054), .ZN(U2972) );
  NOR2_X1 U6255 ( .A1(n5663), .A2(n5466), .ZN(n5062) );
  NAND3_X1 U6256 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n3452), .ZN(n5662) );
  AOI21_X1 U6257 ( .B1(n5056), .B2(n5055), .A(n5662), .ZN(n5061) );
  NAND2_X1 U6258 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U6259 ( .A1(n5059), .A2(n5466), .B1(n5058), .B2(n5057), .ZN(n5060)
         );
  NAND2_X1 U6260 ( .A1(n5060), .A2(n6041), .ZN(n5658) );
  OAI33_X1 U6261 ( .A1(1'b0), .A2(n5062), .A3(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .B1(n5465), .B2(n5061), .B3(n5658), .ZN(n5069) );
  XNOR2_X1 U6262 ( .A(n5065), .B(n5064), .ZN(n5845) );
  INV_X1 U6263 ( .A(n5066), .ZN(n5067) );
  AOI21_X1 U6264 ( .B1(n6106), .B2(n5845), .A(n5067), .ZN(n5068) );
  OAI211_X1 U6265 ( .C1(n5070), .C2(n6083), .A(n5069), .B(n5068), .ZN(U3004)
         );
  AOI21_X1 U6266 ( .B1(n5072), .B2(n5040), .A(n5071), .ZN(n5866) );
  INV_X1 U6267 ( .A(n5866), .ZN(n5074) );
  XNOR2_X1 U6268 ( .A(n5081), .B(n5080), .ZN(n5464) );
  INV_X1 U6269 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5073) );
  OAI222_X1 U6270 ( .A1(n5074), .A2(n5264), .B1(n5267), .B2(n5464), .C1(n5073), 
        .C2(n5852), .ZN(U2843) );
  OAI21_X1 U6271 ( .B1(n5071), .B2(n5077), .A(n5076), .ZN(n5859) );
  AOI21_X1 U6272 ( .B1(n5081), .B2(n5080), .A(n5079), .ZN(n5082) );
  OR2_X1 U6273 ( .A1(n5078), .A2(n5082), .ZN(n5458) );
  INV_X1 U6274 ( .A(n5458), .ZN(n5083) );
  AOI22_X1 U6275 ( .A1(n5083), .A2(n5849), .B1(n5261), .B2(EBX_REG_17__SCAN_IN), .ZN(n5084) );
  OAI21_X1 U6276 ( .B1(n5859), .B2(n5264), .A(n5084), .ZN(U2842) );
  NOR2_X1 U6277 ( .A1(n5676), .A2(n6428), .ZN(n5085) );
  AOI21_X1 U6278 ( .B1(n6329), .B2(n6300), .A(n5085), .ZN(n5669) );
  INV_X1 U6279 ( .A(n5086), .ZN(n6429) );
  NAND2_X1 U6280 ( .A1(n5669), .A2(n6429), .ZN(n6432) );
  OAI21_X1 U6281 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6338), .A(n6432), 
        .ZN(n6433) );
  INV_X1 U6282 ( .A(n6433), .ZN(n5095) );
  INV_X1 U6283 ( .A(n6338), .ZN(n5097) );
  INV_X1 U6284 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U6285 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5088), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6507), .ZN(n5098) );
  NAND2_X1 U6286 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5099) );
  INV_X1 U6287 ( .A(n5099), .ZN(n5093) );
  NAND2_X1 U6288 ( .A1(n4455), .A2(n6297), .ZN(n5091) );
  OAI21_X1 U6289 ( .B1(n5089), .B2(n5087), .A(n3527), .ZN(n5090) );
  OAI211_X1 U6290 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n5092), .A(n5091), .B(n5090), .ZN(n6301) );
  AOI222_X1 U6291 ( .A1(n5097), .A2(n5087), .B1(n5098), .B2(n5093), .C1(n6301), 
        .C2(n5665), .ZN(n5094) );
  INV_X1 U6292 ( .A(n6432), .ZN(n5104) );
  OAI22_X1 U6293 ( .A1(n5095), .A2(n3471), .B1(n5094), .B2(n5104), .ZN(U3460)
         );
  INV_X1 U6294 ( .A(n5096), .ZN(n5100) );
  AOI21_X1 U6295 ( .B1(n5100), .B2(n5097), .A(n5104), .ZN(n5107) );
  NOR2_X1 U6296 ( .A1(n5099), .A2(n5098), .ZN(n5102) );
  NOR3_X1 U6297 ( .A1(n5100), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6338), 
        .ZN(n5101) );
  AOI211_X1 U6298 ( .C1(n5103), .C2(n5665), .A(n5102), .B(n5101), .ZN(n5105)
         );
  OAI22_X1 U6299 ( .A1(n5107), .A2(n5106), .B1(n5105), .B2(n5104), .ZN(U3459)
         );
  NAND2_X1 U6300 ( .A1(n5109), .A2(n5108), .ZN(n5111) );
  AOI22_X1 U6301 ( .A1(n5864), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5861), .ZN(n5110) );
  OAI21_X1 U6302 ( .B1(n5130), .B2(n5111), .A(n5110), .ZN(U2860) );
  NAND2_X1 U6303 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5112), .ZN(n5113) );
  NOR2_X1 U6304 ( .A1(n5113), .A2(REIP_REG_31__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6305 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n5820), .B1(
        REIP_REG_31__SCAN_IN), .B2(n5114), .ZN(n5115) );
  INV_X1 U6306 ( .A(n5115), .ZN(n5127) );
  NAND2_X1 U6307 ( .A1(n3580), .A2(n5214), .ZN(n5208) );
  NAND2_X1 U6308 ( .A1(n5213), .A2(n5117), .ZN(n5119) );
  NAND2_X1 U6309 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  OAI22_X1 U6310 ( .A1(n5120), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4156), .ZN(n5121) );
  NAND2_X1 U6311 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5123), .ZN(n5125) );
  OAI22_X1 U6312 ( .A1(n5341), .A2(n5824), .B1(n5125), .B2(n5124), .ZN(n5126)
         );
  NOR3_X1 U6313 ( .A1(n5128), .A2(n5127), .A3(n5126), .ZN(n5129) );
  OAI21_X1 U6314 ( .B1(n5130), .B2(n5780), .A(n5129), .ZN(U2796) );
  INV_X1 U6315 ( .A(n5131), .ZN(n5134) );
  INV_X1 U6316 ( .A(n5132), .ZN(n5133) );
  OAI21_X1 U6317 ( .B1(n5134), .B2(n5133), .A(n5232), .ZN(n5393) );
  OAI21_X1 U6318 ( .B1(n5137), .B2(n5136), .A(n5135), .ZN(n5626) );
  INV_X1 U6319 ( .A(n5626), .ZN(n5142) );
  AOI22_X1 U6320 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5821), .B1(n5622), .B2(n5799), .ZN(n5139) );
  INV_X1 U6321 ( .A(n5143), .ZN(n5560) );
  INV_X1 U6322 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6410) );
  NAND3_X1 U6323 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5560), .A3(n6410), .ZN(
        n5138) );
  OAI211_X1 U6324 ( .C1(n5834), .C2(n5140), .A(n5139), .B(n5138), .ZN(n5141)
         );
  AOI21_X1 U6325 ( .B1(n5142), .B2(n5770), .A(n5141), .ZN(n5145) );
  NOR2_X1 U6326 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5143), .ZN(n5149) );
  OAI21_X1 U6327 ( .B1(n5149), .B2(n5574), .A(REIP_REG_25__SCAN_IN), .ZN(n5144) );
  OAI211_X1 U6328 ( .C1(n5393), .C2(n5824), .A(n5145), .B(n5144), .ZN(U2802)
         );
  AOI22_X1 U6329 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5820), .ZN(n5148) );
  AOI22_X1 U6330 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5574), .B1(n5146), .B2(
        n5799), .ZN(n5147) );
  OAI211_X1 U6331 ( .C1(n5276), .C2(n5780), .A(n5148), .B(n5147), .ZN(n5150)
         );
  NOR2_X1 U6332 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  OAI21_X1 U6333 ( .B1(n5824), .B2(n5240), .A(n5151), .ZN(U2803) );
  NOR2_X1 U6334 ( .A1(n5152), .A2(n5153), .ZN(n5154) );
  NOR2_X1 U6335 ( .A1(n4190), .A2(n5154), .ZN(n5605) );
  INV_X1 U6336 ( .A(n5605), .ZN(n5244) );
  INV_X1 U6337 ( .A(n5593), .ZN(n5579) );
  NAND2_X1 U6338 ( .A1(n5155), .A2(n5160), .ZN(n5582) );
  INV_X1 U6339 ( .A(n5582), .ZN(n5156) );
  OAI21_X1 U6340 ( .B1(n5579), .B2(n5156), .A(REIP_REG_22__SCAN_IN), .ZN(n5164) );
  AND2_X1 U6341 ( .A1(n5247), .A2(n5157), .ZN(n5158) );
  NOR2_X1 U6342 ( .A1(n5159), .A2(n5158), .ZN(n5401) );
  INV_X1 U6343 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5245) );
  OAI22_X1 U6344 ( .A1(n5245), .A2(n5836), .B1(n3954), .B2(n5834), .ZN(n5162)
         );
  NAND2_X1 U6345 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5160), .ZN(n5572) );
  OAI22_X1 U6346 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5572), .B1(n5301), .B2(
        n5835), .ZN(n5161) );
  AOI211_X1 U6347 ( .C1(n5401), .C2(n5831), .A(n5162), .B(n5161), .ZN(n5163)
         );
  OAI211_X1 U6348 ( .C1(n5244), .C2(n5780), .A(n5164), .B(n5163), .ZN(U2805)
         );
  OR2_X1 U6349 ( .A1(n5166), .A2(n5165), .ZN(n5182) );
  NAND2_X1 U6350 ( .A1(n5078), .A2(n5182), .ZN(n5184) );
  XNOR2_X1 U6351 ( .A(n5184), .B(n5167), .ZN(n5262) );
  INV_X1 U6352 ( .A(n5262), .ZN(n5644) );
  INV_X1 U6353 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U6354 ( .A1(n5832), .A2(n5168), .ZN(n5191) );
  OAI21_X1 U6355 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5181), .A(n5191), .ZN(n5173) );
  AOI22_X1 U6356 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5821), .B1(n5317), .B2(n5799), .ZN(n5170) );
  NAND2_X1 U6357 ( .A1(n5804), .A2(n5169), .ZN(n5782) );
  OAI211_X1 U6358 ( .C1(n5834), .C2(n5171), .A(n5170), .B(n5782), .ZN(n5172)
         );
  AOI221_X1 U6359 ( .B1(n5174), .B2(n6402), .C1(n5173), .C2(
        REIP_REG_19__SCAN_IN), .A(n5172), .ZN(n5178) );
  XOR2_X1 U6360 ( .A(n5175), .B(n5176), .Z(n5613) );
  NAND2_X1 U6361 ( .A1(n5613), .A2(n5770), .ZN(n5177) );
  OAI211_X1 U6362 ( .C1(n5644), .C2(n5824), .A(n5178), .B(n5177), .ZN(U2808)
         );
  AOI21_X1 U6363 ( .B1(n5076), .B2(n5179), .A(n5175), .ZN(n5853) );
  INV_X1 U6364 ( .A(n5853), .ZN(n5266) );
  OAI22_X1 U6365 ( .A1(n5635), .A2(n5835), .B1(n5780), .B2(n5266), .ZN(n5188)
         );
  AOI21_X1 U6366 ( .B1(n5820), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5793), 
        .ZN(n5180) );
  OAI221_X1 U6367 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5181), .C1(n6399), .C2(
        n5191), .A(n5180), .ZN(n5187) );
  OR2_X1 U6368 ( .A1(n5078), .A2(n5182), .ZN(n5183) );
  NAND2_X1 U6369 ( .A1(n5184), .A2(n5183), .ZN(n5440) );
  INV_X1 U6370 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5185) );
  OAI22_X1 U6371 ( .A1(n5440), .A2(n5824), .B1(n5185), .B2(n5836), .ZN(n5186)
         );
  OR3_X1 U6372 ( .A1(n5188), .A2(n5187), .A3(n5186), .ZN(U2809) );
  NOR2_X1 U6373 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5189), .ZN(n5192) );
  OAI22_X1 U6374 ( .A1(n5192), .A2(n5191), .B1(n5190), .B2(n5834), .ZN(n5197)
         );
  INV_X1 U6375 ( .A(n5859), .ZN(n5193) );
  AOI22_X1 U6376 ( .A1(n5636), .A2(n5799), .B1(n5770), .B2(n5193), .ZN(n5195)
         );
  NAND2_X1 U6377 ( .A1(n5821), .A2(EBX_REG_17__SCAN_IN), .ZN(n5194) );
  OAI211_X1 U6378 ( .C1(n5458), .C2(n5824), .A(n5195), .B(n5194), .ZN(n5196)
         );
  OR3_X1 U6379 ( .A1(n5197), .A2(n5793), .A3(n5196), .ZN(U2810) );
  OAI21_X1 U6380 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5198), .ZN(n5202) );
  NOR2_X1 U6381 ( .A1(n5200), .A2(n5199), .ZN(n5701) );
  AOI22_X1 U6382 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5821), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5701), .ZN(n5201) );
  OAI21_X1 U6383 ( .B1(n5693), .B2(n5202), .A(n5201), .ZN(n5203) );
  AOI211_X1 U6384 ( .C1(n5820), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5793), 
        .B(n5203), .ZN(n5205) );
  AOI22_X1 U6385 ( .A1(n5326), .A2(n2956), .B1(n5770), .B2(n5866), .ZN(n5204)
         );
  OAI211_X1 U6386 ( .C1(n5464), .C2(n5824), .A(n5205), .B(n5204), .ZN(U2811)
         );
  OAI22_X1 U6387 ( .A1(n5341), .A2(n5267), .B1(n4182), .B2(n5852), .ZN(U2828)
         );
  AOI22_X1 U6388 ( .A1(n5349), .A2(n5849), .B1(EBX_REG_30__SCAN_IN), .B2(n5261), .ZN(n5206) );
  OAI21_X1 U6389 ( .B1(n4215), .B2(n5264), .A(n5206), .ZN(U2829) );
  INV_X1 U6390 ( .A(n5207), .ZN(n5539) );
  OAI21_X1 U6391 ( .B1(n5209), .B2(n3580), .A(n5208), .ZN(n5210) );
  INV_X1 U6392 ( .A(n5210), .ZN(n5211) );
  AND2_X1 U6393 ( .A1(n5220), .A2(n5211), .ZN(n5212) );
  OAI222_X1 U6394 ( .A1(n5539), .A2(n5264), .B1(n5852), .B2(n5214), .C1(n5267), 
        .C2(n5529), .ZN(U2830) );
  NAND2_X1 U6395 ( .A1(n2967), .A2(n5215), .ZN(n5216) );
  INV_X1 U6396 ( .A(n5594), .ZN(n5222) );
  INV_X1 U6397 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5221) );
  OR2_X1 U6398 ( .A1(n5227), .A2(n5218), .ZN(n5219) );
  NAND2_X1 U6399 ( .A1(n5220), .A2(n5219), .ZN(n5543) );
  OAI222_X1 U6400 ( .A1(n5222), .A2(n5264), .B1(n5852), .B2(n5221), .C1(n5267), 
        .C2(n5543), .ZN(U2831) );
  OAI21_X1 U6401 ( .B1(n5223), .B2(n5224), .A(n2967), .ZN(n5558) );
  INV_X1 U6402 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5228) );
  NOR2_X1 U6403 ( .A1(n5234), .A2(n5225), .ZN(n5226) );
  OR2_X1 U6404 ( .A1(n5227), .A2(n5226), .ZN(n5553) );
  OAI222_X1 U6405 ( .A1(n5558), .A2(n5264), .B1(n5852), .B2(n5228), .C1(n5553), 
        .C2(n5267), .ZN(U2832) );
  AND2_X1 U6406 ( .A1(n5135), .A2(n5229), .ZN(n5230) );
  OR2_X1 U6407 ( .A1(n5230), .A2(n5223), .ZN(n5617) );
  INV_X1 U6408 ( .A(n5617), .ZN(n5566) );
  NAND2_X1 U6409 ( .A1(n5566), .A2(n5850), .ZN(n5236) );
  AND2_X1 U6410 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NOR2_X1 U6411 ( .A1(n5234), .A2(n5233), .ZN(n5561) );
  NAND2_X1 U6412 ( .A1(n5561), .A2(n5849), .ZN(n5235) );
  OAI211_X1 U6413 ( .C1(n5237), .C2(n5852), .A(n5236), .B(n5235), .ZN(U2833)
         );
  INV_X1 U6414 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5238) );
  OAI222_X1 U6415 ( .A1(n5393), .A2(n5267), .B1(n5852), .B2(n5238), .C1(n5264), 
        .C2(n5626), .ZN(U2834) );
  INV_X1 U6416 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5239) );
  OAI222_X1 U6417 ( .A1(n5240), .A2(n5267), .B1(n5852), .B2(n5239), .C1(n5264), 
        .C2(n5276), .ZN(U2835) );
  OAI22_X1 U6418 ( .A1(n5241), .A2(n5267), .B1(n6485), .B2(n5852), .ZN(n5242)
         );
  INV_X1 U6419 ( .A(n5242), .ZN(n5243) );
  OAI21_X1 U6420 ( .B1(n5578), .B2(n5264), .A(n5243), .ZN(U2836) );
  INV_X1 U6421 ( .A(n5401), .ZN(n5246) );
  OAI222_X1 U6422 ( .A1(n5246), .A2(n5267), .B1(n5852), .B2(n5245), .C1(n5264), 
        .C2(n5244), .ZN(U2837) );
  INV_X1 U6423 ( .A(n5247), .ZN(n5248) );
  AOI21_X1 U6424 ( .B1(n5250), .B2(n5249), .A(n5248), .ZN(n5581) );
  INV_X1 U6425 ( .A(n5581), .ZN(n5254) );
  XOR2_X1 U6426 ( .A(n5251), .B(n5252), .Z(n5608) );
  AOI22_X1 U6427 ( .A1(n5850), .A2(n5608), .B1(EBX_REG_21__SCAN_IN), .B2(n5261), .ZN(n5253) );
  OAI21_X1 U6428 ( .B1(n5254), .B2(n5267), .A(n5253), .ZN(U2838) );
  AOI21_X1 U6429 ( .B1(n5256), .B2(n5255), .A(n5251), .ZN(n5628) );
  INV_X1 U6430 ( .A(n5628), .ZN(n5588) );
  MUX2_X1 U6431 ( .A(n2963), .B(n5258), .S(n5257), .Z(n5260) );
  XNOR2_X1 U6432 ( .A(n5260), .B(n5259), .ZN(n5587) );
  OAI222_X1 U6433 ( .A1(n5264), .A2(n5588), .B1(n5267), .B2(n5587), .C1(n5852), 
        .C2(n3639), .ZN(U2839) );
  INV_X1 U6434 ( .A(n5613), .ZN(n5265) );
  AOI22_X1 U6435 ( .A1(n5262), .A2(n5849), .B1(n5261), .B2(EBX_REG_19__SCAN_IN), .ZN(n5263) );
  OAI21_X1 U6436 ( .B1(n5265), .B2(n5264), .A(n5263), .ZN(U2840) );
  OAI222_X1 U6437 ( .A1(n5440), .A2(n5267), .B1(n5852), .B2(n5185), .C1(n5264), 
        .C2(n5266), .ZN(U2841) );
  INV_X1 U6438 ( .A(DATAI_29_), .ZN(n5269) );
  NAND2_X1 U6439 ( .A1(EAX_REG_29__SCAN_IN), .A2(n5861), .ZN(n5268) );
  OAI21_X1 U6440 ( .B1(n5857), .B2(n5269), .A(n5268), .ZN(n5270) );
  AOI21_X1 U6441 ( .B1(n5867), .B2(DATAI_13_), .A(n5270), .ZN(n5271) );
  OAI21_X1 U6442 ( .B1(n5539), .B2(n5858), .A(n5271), .ZN(U2862) );
  AOI22_X1 U6443 ( .A1(n5867), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5861), .ZN(n5273) );
  NAND2_X1 U6444 ( .A1(n5864), .A2(DATAI_27_), .ZN(n5272) );
  OAI211_X1 U6445 ( .C1(n5558), .C2(n5858), .A(n5273), .B(n5272), .ZN(U2864)
         );
  AOI22_X1 U6446 ( .A1(n5867), .A2(DATAI_8_), .B1(n5861), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6447 ( .A1(n5864), .A2(DATAI_24_), .ZN(n5274) );
  OAI211_X1 U6448 ( .C1(n5276), .C2(n5858), .A(n5275), .B(n5274), .ZN(U2867)
         );
  AOI22_X1 U6449 ( .A1(n5867), .A2(DATAI_7_), .B1(n5861), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6450 ( .A1(n5864), .A2(DATAI_23_), .ZN(n5277) );
  OAI211_X1 U6451 ( .C1(n5578), .C2(n5858), .A(n5278), .B(n5277), .ZN(U2868)
         );
  INV_X1 U6452 ( .A(n5279), .ZN(n5280) );
  NAND3_X1 U6453 ( .A1(n5280), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n2965), .ZN(n5283) );
  AND2_X1 U6454 ( .A1(n5381), .A2(n5386), .ZN(n5282) );
  NAND2_X1 U6455 ( .A1(n5392), .A2(n5282), .ZN(n5291) );
  AOI22_X1 U6456 ( .A1(n5283), .A2(n5291), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5385), .ZN(n5284) );
  XNOR2_X1 U6457 ( .A(n5284), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5370)
         );
  NOR2_X1 U6458 ( .A1(n6071), .A2(n5545), .ZN(n5366) );
  AOI21_X1 U6459 ( .B1(n6025), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5366), 
        .ZN(n5285) );
  OAI21_X1 U6460 ( .B1(n6035), .B2(n5540), .A(n5285), .ZN(n5286) );
  AOI21_X1 U6461 ( .B1(n5594), .B2(n6030), .A(n5286), .ZN(n5287) );
  OAI21_X1 U6462 ( .B1(n5675), .B2(n5370), .A(n5287), .ZN(U2958) );
  NOR2_X1 U6463 ( .A1(n6071), .A2(n6413), .ZN(n5372) );
  NOR2_X1 U6464 ( .A1(n5315), .A2(n5288), .ZN(n5289) );
  AOI211_X1 U6465 ( .C1(n6012), .C2(n5552), .A(n5372), .B(n5289), .ZN(n5295)
         );
  INV_X1 U6466 ( .A(n5291), .ZN(n5292) );
  NOR2_X1 U6467 ( .A1(n5290), .A2(n5292), .ZN(n5293) );
  XNOR2_X1 U6468 ( .A(n5293), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5377)
         );
  NAND2_X1 U6469 ( .A1(n5377), .A2(n6029), .ZN(n5294) );
  OAI211_X1 U6470 ( .C1(n5558), .C2(n4314), .A(n5295), .B(n5294), .ZN(U2959)
         );
  AOI21_X1 U6471 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2965), .A(n5297), 
        .ZN(n5298) );
  XNOR2_X1 U6472 ( .A(n5299), .B(n5298), .ZN(n5409) );
  NOR2_X1 U6473 ( .A1(n6071), .A2(n6598), .ZN(n5402) );
  AOI21_X1 U6474 ( .B1(n6025), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5402), 
        .ZN(n5300) );
  OAI21_X1 U6475 ( .B1(n6035), .B2(n5301), .A(n5300), .ZN(n5302) );
  AOI21_X1 U6476 ( .B1(n5605), .B2(n6030), .A(n5302), .ZN(n5303) );
  OAI21_X1 U6477 ( .B1(n5409), .B2(n5675), .A(n5303), .ZN(U2964) );
  AOI21_X1 U6478 ( .B1(n5306), .B2(n5305), .A(n5304), .ZN(n5416) );
  NOR2_X1 U6479 ( .A1(n6071), .A2(n5155), .ZN(n5410) );
  AOI21_X1 U6480 ( .B1(n6030), .B2(n5608), .A(n5410), .ZN(n5307) );
  OAI21_X1 U6481 ( .B1(n5315), .B2(n5308), .A(n5307), .ZN(n5309) );
  AOI21_X1 U6482 ( .B1(n6012), .B2(n5580), .A(n5309), .ZN(n5310) );
  OAI21_X1 U6483 ( .B1(n5416), .B2(n5675), .A(n5310), .ZN(U2965) );
  INV_X1 U6484 ( .A(n5312), .ZN(n5313) );
  AOI21_X1 U6485 ( .B1(n5311), .B2(n5314), .A(n5313), .ZN(n5645) );
  NAND2_X1 U6486 ( .A1(n5613), .A2(n6030), .ZN(n5319) );
  OAI22_X1 U6487 ( .A1(n5315), .A2(n5171), .B1(n6071), .B2(n6402), .ZN(n5316)
         );
  AOI21_X1 U6488 ( .B1(n6012), .B2(n5317), .A(n5316), .ZN(n5318) );
  OAI211_X1 U6489 ( .C1(n5645), .C2(n5675), .A(n5319), .B(n5318), .ZN(U2967)
         );
  NOR2_X1 U6490 ( .A1(n3439), .A2(n5467), .ZN(n5453) );
  INV_X1 U6491 ( .A(n5323), .ZN(n5324) );
  NOR2_X1 U6492 ( .A1(n5453), .A2(n5324), .ZN(n5325) );
  OAI22_X1 U6493 ( .A1(n5321), .A2(n5453), .B1(n5322), .B2(n5325), .ZN(n5472)
         );
  INV_X1 U6494 ( .A(n5326), .ZN(n5328) );
  AOI22_X1 U6495 ( .A1(n6025), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6104), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5327) );
  OAI21_X1 U6496 ( .B1(n6035), .B2(n5328), .A(n5327), .ZN(n5329) );
  AOI21_X1 U6497 ( .B1(n5866), .B2(n6030), .A(n5329), .ZN(n5330) );
  OAI21_X1 U6498 ( .B1(n5675), .B2(n5472), .A(n5330), .ZN(U2970) );
  NAND2_X1 U6499 ( .A1(n5331), .A2(n6126), .ZN(n5340) );
  NAND2_X1 U6500 ( .A1(n5332), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6501 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5361) );
  INV_X1 U6502 ( .A(n5363), .ZN(n5333) );
  NOR3_X1 U6503 ( .A1(n5371), .A2(n5333), .A3(n5354), .ZN(n5343) );
  NAND3_X1 U6504 ( .A1(n5343), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5088), .ZN(n5338) );
  OAI21_X1 U6505 ( .B1(n5361), .B2(n5333), .A(n6070), .ZN(n5334) );
  NAND2_X1 U6506 ( .A1(n5383), .A2(n5334), .ZN(n5353) );
  AOI21_X1 U6507 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6122), .ZN(n5335) );
  OAI21_X1 U6508 ( .B1(n5353), .B2(n5335), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n5336) );
  AND3_X1 U6509 ( .A1(n5338), .A2(n5337), .A3(n5336), .ZN(n5339) );
  OAI211_X1 U6510 ( .C1(n5341), .C2(n6120), .A(n5340), .B(n5339), .ZN(U2987)
         );
  INV_X1 U6511 ( .A(n5342), .ZN(n5351) );
  INV_X1 U6512 ( .A(n5343), .ZN(n5347) );
  NAND2_X1 U6513 ( .A1(n5383), .A2(n6122), .ZN(n5344) );
  OAI211_X1 U6514 ( .C1(n5353), .C2(n5354), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5344), .ZN(n5346) );
  OAI211_X1 U6515 ( .C1(n5347), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5346), .B(n5345), .ZN(n5348) );
  AOI21_X1 U6516 ( .B1(n5349), .B2(n6106), .A(n5348), .ZN(n5350) );
  OAI21_X1 U6517 ( .B1(n5351), .B2(n6083), .A(n5350), .ZN(U2988) );
  AOI21_X1 U6518 ( .B1(n5353), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5352), 
        .ZN(n5357) );
  INV_X1 U6519 ( .A(n5371), .ZN(n5355) );
  NAND3_X1 U6520 ( .A1(n5355), .A2(n5363), .A3(n5354), .ZN(n5356) );
  OAI211_X1 U6521 ( .C1(n5529), .C2(n6120), .A(n5357), .B(n5356), .ZN(n5358)
         );
  AOI21_X1 U6522 ( .B1(n5359), .B2(n6126), .A(n5358), .ZN(n5360) );
  INV_X1 U6523 ( .A(n5360), .ZN(U2989) );
  NAND2_X1 U6524 ( .A1(n6070), .A2(n5361), .ZN(n5362) );
  NAND2_X1 U6525 ( .A1(n5383), .A2(n5362), .ZN(n5373) );
  NOR3_X1 U6526 ( .A1(n5371), .A2(n5364), .A3(n5363), .ZN(n5365) );
  AOI211_X1 U6527 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5373), .A(n5366), .B(n5365), .ZN(n5369) );
  INV_X1 U6528 ( .A(n5543), .ZN(n5367) );
  NAND2_X1 U6529 ( .A1(n5367), .A2(n6106), .ZN(n5368) );
  OAI211_X1 U6530 ( .C1(n5370), .C2(n6083), .A(n5369), .B(n5368), .ZN(U2990)
         );
  NOR2_X1 U6531 ( .A1(n5371), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5376)
         );
  AOI21_X1 U6532 ( .B1(n5373), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5372), 
        .ZN(n5374) );
  OAI21_X1 U6533 ( .B1(n5553), .B2(n6120), .A(n5374), .ZN(n5375) );
  AOI211_X1 U6534 ( .C1(n5377), .C2(n6126), .A(n5376), .B(n5375), .ZN(n5378)
         );
  INV_X1 U6535 ( .A(n5378), .ZN(U2991) );
  INV_X1 U6536 ( .A(n5379), .ZN(n5380) );
  NOR2_X1 U6537 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  XNOR2_X1 U6538 ( .A(n5279), .B(n5382), .ZN(n5616) );
  OAI22_X1 U6539 ( .A1(n5383), .A2(n5385), .B1(n6071), .B2(n6519), .ZN(n5384)
         );
  AOI21_X1 U6540 ( .B1(n5561), .B2(n6106), .A(n5384), .ZN(n5390) );
  AOI22_X1 U6541 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .B1(n5386), .B2(n5385), .ZN(n5387)
         );
  INV_X1 U6542 ( .A(n5387), .ZN(n5388) );
  OR2_X1 U6543 ( .A1(n5398), .A2(n5388), .ZN(n5389) );
  OAI211_X1 U6544 ( .C1(n5616), .C2(n6083), .A(n5390), .B(n5389), .ZN(U2992)
         );
  OAI21_X1 U6545 ( .B1(n5392), .B2(n5391), .A(n4271), .ZN(n5623) );
  NAND2_X1 U6546 ( .A1(n5623), .A2(n6126), .ZN(n5397) );
  OAI22_X1 U6547 ( .A1(n5393), .A2(n6120), .B1(n6071), .B2(n6410), .ZN(n5394)
         );
  AOI21_X1 U6548 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5395), .A(n5394), 
        .ZN(n5396) );
  OAI211_X1 U6549 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5398), .A(n5397), .B(n5396), .ZN(U2993) );
  NOR2_X1 U6550 ( .A1(n5400), .A2(n5399), .ZN(n5407) );
  INV_X1 U6551 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6552 ( .A1(n5401), .A2(n6106), .ZN(n5404) );
  INV_X1 U6553 ( .A(n5402), .ZN(n5403) );
  OAI211_X1 U6554 ( .C1(n5412), .C2(n5405), .A(n5404), .B(n5403), .ZN(n5406)
         );
  AOI21_X1 U6555 ( .B1(n5414), .B2(n5407), .A(n5406), .ZN(n5408) );
  OAI21_X1 U6556 ( .B1(n5409), .B2(n6083), .A(n5408), .ZN(U2996) );
  AOI21_X1 U6557 ( .B1(n5581), .B2(n6106), .A(n5410), .ZN(n5411) );
  OAI21_X1 U6558 ( .B1(n5412), .B2(n4220), .A(n5411), .ZN(n5413) );
  AOI21_X1 U6559 ( .B1(n5414), .B2(n4220), .A(n5413), .ZN(n5415) );
  OAI21_X1 U6560 ( .B1(n5416), .B2(n6083), .A(n5415), .ZN(U2997) );
  XNOR2_X1 U6561 ( .A(n3439), .B(n5418), .ZN(n5419) );
  XNOR2_X1 U6562 ( .A(n5417), .B(n5419), .ZN(n5627) );
  INV_X1 U6563 ( .A(n5627), .ZN(n5432) );
  NAND3_X1 U6564 ( .A1(n5420), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6037), .ZN(n5650) );
  NOR2_X1 U6565 ( .A1(n5421), .A2(n5650), .ZN(n5425) );
  INV_X1 U6566 ( .A(n5422), .ZN(n5424) );
  OAI22_X1 U6567 ( .A1(n5587), .A2(n6120), .B1(n6071), .B2(n6404), .ZN(n5423)
         );
  AOI21_X1 U6568 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(n5431) );
  NOR2_X1 U6569 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5426), .ZN(n5460)
         );
  OAI21_X1 U6570 ( .B1(n6068), .B2(n5428), .A(n5427), .ZN(n5456) );
  AOI21_X1 U6571 ( .B1(n5429), .B2(n5460), .A(n5456), .ZN(n5443) );
  OAI21_X1 U6572 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6122), .A(n5443), 
        .ZN(n5648) );
  NAND2_X1 U6573 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5430) );
  OAI211_X1 U6574 ( .C1(n5432), .C2(n6083), .A(n5431), .B(n5430), .ZN(U2998)
         );
  INV_X1 U6575 ( .A(n5433), .ZN(n5434) );
  NOR2_X1 U6576 ( .A1(n3439), .A2(n5434), .ZN(n5435) );
  INV_X1 U6577 ( .A(n5435), .ZN(n5437) );
  INV_X1 U6578 ( .A(n5322), .ZN(n5436) );
  AOI22_X1 U6579 ( .A1(n5436), .A2(n5435), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n2965), .ZN(n5455) );
  AOI21_X1 U6580 ( .B1(n5321), .B2(n5437), .A(n5455), .ZN(n5439) );
  XNOR2_X1 U6581 ( .A(n5439), .B(n5438), .ZN(n5632) );
  INV_X1 U6582 ( .A(n5632), .ZN(n5448) );
  INV_X1 U6583 ( .A(n5440), .ZN(n5446) );
  INV_X1 U6584 ( .A(n5441), .ZN(n5444) );
  NAND2_X1 U6585 ( .A1(n6104), .A2(REIP_REG_18__SCAN_IN), .ZN(n5442) );
  OAI221_X1 U6586 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5444), .C1(
        n5438), .C2(n5443), .A(n5442), .ZN(n5445) );
  AOI21_X1 U6587 ( .B1(n5446), .B2(n6106), .A(n5445), .ZN(n5447) );
  OAI21_X1 U6588 ( .B1(n5448), .B2(n6083), .A(n5447), .ZN(U3000) );
  MUX2_X1 U6589 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n5451), .S(n3439), 
        .Z(n5452) );
  OAI21_X1 U6590 ( .B1(n5450), .B2(n5453), .A(n5452), .ZN(n5454) );
  OAI21_X1 U6591 ( .B1(n5455), .B2(n5450), .A(n5454), .ZN(n5637) );
  INV_X1 U6592 ( .A(n5637), .ZN(n5462) );
  AOI22_X1 U6593 ( .A1(n6104), .A2(REIP_REG_17__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5456), .ZN(n5457) );
  OAI21_X1 U6594 ( .B1(n6120), .B2(n5458), .A(n5457), .ZN(n5459) );
  AOI21_X1 U6595 ( .B1(n6037), .B2(n5460), .A(n5459), .ZN(n5461) );
  OAI21_X1 U6596 ( .B1(n5462), .B2(n6083), .A(n5461), .ZN(U3001) );
  OAI21_X1 U6597 ( .B1(n6122), .B2(n5463), .A(n6041), .ZN(n5651) );
  INV_X1 U6598 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6397) );
  OAI22_X1 U6599 ( .A1(n6120), .A2(n5464), .B1(n6397), .B2(n6071), .ZN(n5470)
         );
  INV_X1 U6600 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5467) );
  NOR3_X1 U6601 ( .A1(n5663), .A2(n5466), .A3(n5465), .ZN(n5652) );
  OAI221_X1 U6602 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5656), .C2(n5467), .A(n5652), 
        .ZN(n5468) );
  INV_X1 U6603 ( .A(n5468), .ZN(n5469) );
  AOI211_X1 U6604 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5651), .A(n5470), .B(n5469), .ZN(n5471) );
  OAI21_X1 U6605 ( .B1(n5472), .B2(n6083), .A(n5471), .ZN(U3002) );
  XNOR2_X1 U6606 ( .A(n6232), .B(n4446), .ZN(n5474) );
  OAI22_X1 U6607 ( .A1(n5474), .A2(n6238), .B1(n4416), .B2(n5473), .ZN(n5475)
         );
  MUX2_X1 U6608 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5475), .S(n6130), 
        .Z(U3463) );
  INV_X1 U6609 ( .A(n5665), .ZN(n6436) );
  OAI22_X1 U6610 ( .A1(n5477), .A2(n6436), .B1(n5476), .B2(n6338), .ZN(n5478)
         );
  MUX2_X1 U6611 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5478), .S(n6432), 
        .Z(U3456) );
  AOI22_X1 U6612 ( .A1(n5482), .A2(n5481), .B1(n5480), .B2(n5479), .ZN(n5519)
         );
  NOR2_X1 U6613 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5483), .ZN(n5517)
         );
  OAI21_X1 U6614 ( .B1(n5514), .B2(n6152), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5486) );
  AND3_X1 U6615 ( .A1(n6233), .A2(n5487), .A3(n5486), .ZN(n5489) );
  NOR3_X1 U6616 ( .A1(n5490), .A2(n5489), .A3(n5488), .ZN(n5491) );
  AOI22_X1 U6617 ( .A1(n5514), .A2(n6230), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5513), .ZN(n5492) );
  OAI21_X1 U6618 ( .B1(n6247), .B2(n6164), .A(n5492), .ZN(n5493) );
  AOI21_X1 U6619 ( .B1(n2958), .B2(n5517), .A(n5493), .ZN(n5494) );
  OAI21_X1 U6620 ( .B1(n5519), .B2(n6181), .A(n5494), .ZN(U3052) );
  AOI22_X1 U6621 ( .A1(n5514), .A2(n6182), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5513), .ZN(n5495) );
  OAI21_X1 U6622 ( .B1(n6144), .B2(n6164), .A(n5495), .ZN(n5496) );
  AOI21_X1 U6623 ( .B1(n6249), .B2(n5517), .A(n5496), .ZN(n5497) );
  OAI21_X1 U6624 ( .B1(n5519), .B2(n6185), .A(n5497), .ZN(U3053) );
  AOI22_X1 U6625 ( .A1(n5514), .A2(n6254), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5513), .ZN(n5498) );
  OAI21_X1 U6626 ( .B1(n6259), .B2(n6164), .A(n5498), .ZN(n5499) );
  AOI21_X1 U6627 ( .B1(n6255), .B2(n5517), .A(n5499), .ZN(n5500) );
  OAI21_X1 U6628 ( .B1(n5519), .B2(n6189), .A(n5500), .ZN(U3054) );
  AOI22_X1 U6629 ( .A1(n5514), .A2(n6260), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5513), .ZN(n5501) );
  OAI21_X1 U6630 ( .B1(n6265), .B2(n6164), .A(n5501), .ZN(n5502) );
  AOI21_X1 U6631 ( .B1(n6261), .B2(n5517), .A(n5502), .ZN(n5503) );
  OAI21_X1 U6632 ( .B1(n5519), .B2(n6193), .A(n5503), .ZN(U3055) );
  AOI22_X1 U6633 ( .A1(n5514), .A2(n6216), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5513), .ZN(n5504) );
  OAI21_X1 U6634 ( .B1(n6219), .B2(n6164), .A(n5504), .ZN(n5505) );
  AOI21_X1 U6635 ( .B1(n6267), .B2(n5517), .A(n5505), .ZN(n5506) );
  OAI21_X1 U6636 ( .B1(n5519), .B2(n6196), .A(n5506), .ZN(U3056) );
  AOI22_X1 U6637 ( .A1(n5514), .A2(n6223), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5513), .ZN(n5507) );
  OAI21_X1 U6638 ( .B1(n6228), .B2(n6164), .A(n5507), .ZN(n5508) );
  AOI21_X1 U6639 ( .B1(n6274), .B2(n5517), .A(n5508), .ZN(n5509) );
  OAI21_X1 U6640 ( .B1(n5519), .B2(n6199), .A(n5509), .ZN(U3057) );
  AOI22_X1 U6641 ( .A1(n5514), .A2(n6280), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5513), .ZN(n5510) );
  OAI21_X1 U6642 ( .B1(n6285), .B2(n6164), .A(n5510), .ZN(n5511) );
  AOI21_X1 U6643 ( .B1(n6281), .B2(n5517), .A(n5511), .ZN(n5512) );
  OAI21_X1 U6644 ( .B1(n5519), .B2(n6203), .A(n5512), .ZN(U3058) );
  AOI22_X1 U6645 ( .A1(n5514), .A2(n6287), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5513), .ZN(n5515) );
  OAI21_X1 U6646 ( .B1(n6295), .B2(n6164), .A(n5515), .ZN(n5516) );
  AOI21_X1 U6647 ( .B1(n6288), .B2(n5517), .A(n5516), .ZN(n5518) );
  OAI21_X1 U6648 ( .B1(n5519), .B2(n6211), .A(n5518), .ZN(U3059) );
  AOI22_X1 U6649 ( .A1(n6104), .A2(REIP_REG_15__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6650 ( .A1(n2978), .A2(n5522), .ZN(n5523) );
  XNOR2_X1 U6651 ( .A(n5521), .B(n5523), .ZN(n5653) );
  AOI22_X1 U6652 ( .A1(n5653), .A2(n6029), .B1(n6012), .B2(n5697), .ZN(n5524)
         );
  OAI211_X1 U6653 ( .C1(n4314), .C2(n5700), .A(n5525), .B(n5524), .ZN(U2971)
         );
  INV_X1 U6654 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6521) );
  NOR2_X1 U6655 ( .A1(n6521), .A2(n5888), .ZN(U2892) );
  AOI21_X1 U6656 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5527), .A(n5526), .ZN(
        n5528) );
  INV_X1 U6657 ( .A(n5528), .ZN(U2788) );
  INV_X1 U6658 ( .A(n5529), .ZN(n5537) );
  AOI22_X1 U6659 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5821), .B1(n5530), .B2(n5799), .ZN(n5531) );
  OAI21_X1 U6660 ( .B1(n5532), .B2(n5834), .A(n5531), .ZN(n5536) );
  AOI21_X1 U6661 ( .B1(n6571), .B2(n5534), .A(n5533), .ZN(n5535) );
  AOI211_X1 U6662 ( .C1(n5537), .C2(n5831), .A(n5536), .B(n5535), .ZN(n5538)
         );
  OAI21_X1 U6663 ( .B1(n5539), .B2(n5780), .A(n5538), .ZN(U2798) );
  AOI22_X1 U6664 ( .A1(EBX_REG_28__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5820), .ZN(n5549) );
  INV_X1 U6665 ( .A(n5540), .ZN(n5542) );
  AOI22_X1 U6666 ( .A1(n5542), .A2(n2956), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5541), .ZN(n5548) );
  NOR2_X1 U6667 ( .A1(n5543), .A2(n5824), .ZN(n5544) );
  AOI21_X1 U6668 ( .B1(n5594), .B2(n5770), .A(n5544), .ZN(n5547) );
  NAND3_X1 U6669 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5555), .A3(n5545), .ZN(
        n5546) );
  NAND4_X1 U6670 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(U2799)
         );
  AOI22_X1 U6671 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5820), .ZN(n5550) );
  OAI21_X1 U6672 ( .B1(n5563), .B2(n6413), .A(n5550), .ZN(n5551) );
  AOI21_X1 U6673 ( .B1(n5552), .B2(n2956), .A(n5551), .ZN(n5557) );
  INV_X1 U6674 ( .A(n5553), .ZN(n5554) );
  AOI22_X1 U6675 ( .A1(n5555), .A2(n6413), .B1(n5831), .B2(n5554), .ZN(n5556)
         );
  OAI211_X1 U6676 ( .C1(n5558), .C2(n5780), .A(n5557), .B(n5556), .ZN(U2800)
         );
  AOI22_X1 U6677 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5820), .ZN(n5568) );
  NOR2_X1 U6678 ( .A1(n4230), .A2(n6410), .ZN(n5559) );
  AOI21_X1 U6679 ( .B1(n5560), .B2(n5559), .A(REIP_REG_26__SCAN_IN), .ZN(n5564) );
  INV_X1 U6680 ( .A(n5561), .ZN(n5562) );
  OAI22_X1 U6681 ( .A1(n5564), .A2(n5563), .B1(n5824), .B2(n5562), .ZN(n5565)
         );
  AOI21_X1 U6682 ( .B1(n5566), .B2(n5770), .A(n5565), .ZN(n5567) );
  OAI211_X1 U6683 ( .C1(n5621), .C2(n5835), .A(n5568), .B(n5567), .ZN(U2801)
         );
  OAI22_X1 U6684 ( .A1(n6485), .A2(n5836), .B1(n5569), .B2(n5834), .ZN(n5570)
         );
  AOI21_X1 U6685 ( .B1(n5571), .B2(n2956), .A(n5570), .ZN(n5577) );
  OAI21_X1 U6686 ( .B1(n6598), .B2(n5572), .A(n3652), .ZN(n5575) );
  AOI22_X1 U6687 ( .A1(n5575), .A2(n5574), .B1(n5831), .B2(n5573), .ZN(n5576)
         );
  OAI211_X1 U6688 ( .C1(n5578), .C2(n5780), .A(n5577), .B(n5576), .ZN(U2804)
         );
  AOI22_X1 U6689 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5820), .ZN(n5585) );
  AOI22_X1 U6690 ( .A1(n5580), .A2(n2956), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5579), .ZN(n5584) );
  AOI22_X1 U6691 ( .A1(n5831), .A2(n5581), .B1(n5770), .B2(n5608), .ZN(n5583)
         );
  NAND4_X1 U6692 ( .A1(n5585), .A2(n5584), .A3(n5583), .A4(n5582), .ZN(U2806)
         );
  INV_X1 U6693 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5586) );
  OAI22_X1 U6694 ( .A1(n5586), .A2(n5834), .B1(n5631), .B2(n5835), .ZN(n5590)
         );
  OAI22_X1 U6695 ( .A1(n5780), .A2(n5588), .B1(n5587), .B2(n5824), .ZN(n5589)
         );
  AOI211_X1 U6696 ( .C1(EBX_REG_20__SCAN_IN), .C2(n5821), .A(n5590), .B(n5589), 
        .ZN(n5591) );
  OAI221_X1 U6697 ( .B1(n5593), .B2(n6404), .C1(n5593), .C2(n5592), .A(n5591), 
        .ZN(U2807) );
  AOI22_X1 U6698 ( .A1(n5594), .A2(n5865), .B1(n5864), .B2(DATAI_28_), .ZN(
        n5596) );
  AOI22_X1 U6699 ( .A1(n5867), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5861), .ZN(n5595) );
  NAND2_X1 U6700 ( .A1(n5596), .A2(n5595), .ZN(U2863) );
  INV_X1 U6701 ( .A(DATAI_26_), .ZN(n5597) );
  OAI22_X1 U6702 ( .A1(n5617), .A2(n5858), .B1(n5857), .B2(n5597), .ZN(n5598)
         );
  INV_X1 U6703 ( .A(n5598), .ZN(n5600) );
  AOI22_X1 U6704 ( .A1(n5867), .A2(DATAI_10_), .B1(n5861), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6705 ( .A1(n5600), .A2(n5599), .ZN(U2865) );
  OAI22_X1 U6706 ( .A1(n5626), .A2(n5858), .B1(n5857), .B2(n5601), .ZN(n5602)
         );
  INV_X1 U6707 ( .A(n5602), .ZN(n5604) );
  AOI22_X1 U6708 ( .A1(n5867), .A2(DATAI_9_), .B1(n5861), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6709 ( .A1(n5604), .A2(n5603), .ZN(U2866) );
  AOI22_X1 U6710 ( .A1(n5605), .A2(n5865), .B1(n5864), .B2(DATAI_22_), .ZN(
        n5607) );
  AOI22_X1 U6711 ( .A1(n5867), .A2(DATAI_6_), .B1(n5861), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6712 ( .A1(n5607), .A2(n5606), .ZN(U2869) );
  AOI22_X1 U6713 ( .A1(n5864), .A2(DATAI_21_), .B1(n5865), .B2(n5608), .ZN(
        n5610) );
  AOI22_X1 U6714 ( .A1(n5867), .A2(DATAI_5_), .B1(n5861), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6715 ( .A1(n5610), .A2(n5609), .ZN(U2870) );
  AOI22_X1 U6716 ( .A1(n5628), .A2(n5865), .B1(n5864), .B2(DATAI_20_), .ZN(
        n5612) );
  AOI22_X1 U6717 ( .A1(n5867), .A2(DATAI_4_), .B1(n5861), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6718 ( .A1(n5612), .A2(n5611), .ZN(U2871) );
  AOI22_X1 U6719 ( .A1(n5613), .A2(n5865), .B1(n5864), .B2(DATAI_19_), .ZN(
        n5615) );
  AOI22_X1 U6720 ( .A1(n5867), .A2(DATAI_3_), .B1(n5861), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6721 ( .A1(n5615), .A2(n5614), .ZN(U2872) );
  AOI22_X1 U6722 ( .A1(n6104), .A2(REIP_REG_26__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5620) );
  OAI22_X1 U6723 ( .A1(n5617), .A2(n4314), .B1(n5616), .B2(n5675), .ZN(n5618)
         );
  INV_X1 U6724 ( .A(n5618), .ZN(n5619) );
  OAI211_X1 U6725 ( .C1(n6035), .C2(n5621), .A(n5620), .B(n5619), .ZN(U2960)
         );
  AOI22_X1 U6726 ( .A1(n6104), .A2(REIP_REG_25__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5625) );
  AOI22_X1 U6727 ( .A1(n5623), .A2(n6029), .B1(n6012), .B2(n5622), .ZN(n5624)
         );
  OAI211_X1 U6728 ( .C1(n4314), .C2(n5626), .A(n5625), .B(n5624), .ZN(U2961)
         );
  AOI22_X1 U6729 ( .A1(n6104), .A2(REIP_REG_20__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5630) );
  AOI22_X1 U6730 ( .A1(n5628), .A2(n6030), .B1(n6029), .B2(n5627), .ZN(n5629)
         );
  OAI211_X1 U6731 ( .C1(n6035), .C2(n5631), .A(n5630), .B(n5629), .ZN(U2966)
         );
  AOI22_X1 U6732 ( .A1(n6104), .A2(REIP_REG_18__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5634) );
  AOI22_X1 U6733 ( .A1(n6029), .A2(n5632), .B1(n6030), .B2(n5853), .ZN(n5633)
         );
  OAI211_X1 U6734 ( .C1(n6035), .C2(n5635), .A(n5634), .B(n5633), .ZN(U2968)
         );
  AOI22_X1 U6735 ( .A1(n6104), .A2(REIP_REG_17__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5639) );
  AOI22_X1 U6736 ( .A1(n5637), .A2(n6029), .B1(n6012), .B2(n5636), .ZN(n5638)
         );
  OAI211_X1 U6737 ( .C1(n4314), .C2(n5859), .A(n5639), .B(n5638), .ZN(U2969)
         );
  AOI22_X1 U6738 ( .A1(n6104), .A2(REIP_REG_13__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5643) );
  XNOR2_X1 U6739 ( .A(n5640), .B(n5641), .ZN(n5659) );
  AOI22_X1 U6740 ( .A1(n5659), .A2(n6029), .B1(n6012), .B2(n5715), .ZN(n5642)
         );
  OAI211_X1 U6741 ( .C1(n4314), .C2(n5719), .A(n5643), .B(n5642), .ZN(U2973)
         );
  NOR2_X1 U6742 ( .A1(n6071), .A2(n6402), .ZN(n5647) );
  OAI22_X1 U6743 ( .A1(n5645), .A2(n6083), .B1(n5644), .B2(n6120), .ZN(n5646)
         );
  AOI211_X1 U6744 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5649) );
  OAI21_X1 U6745 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5650), .A(n5649), 
        .ZN(U2999) );
  INV_X1 U6746 ( .A(n5651), .ZN(n5657) );
  AOI22_X1 U6747 ( .A1(n6106), .A2(n5696), .B1(n6104), .B2(
        REIP_REG_15__SCAN_IN), .ZN(n5655) );
  AOI22_X1 U6748 ( .A1(n5653), .A2(n6126), .B1(n5652), .B2(n5656), .ZN(n5654)
         );
  OAI211_X1 U6749 ( .C1(n5657), .C2(n5656), .A(n5655), .B(n5654), .ZN(U3003)
         );
  AOI22_X1 U6750 ( .A1(n6106), .A2(n5710), .B1(n6104), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5661) );
  AOI22_X1 U6751 ( .A1(n5659), .A2(n6126), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5658), .ZN(n5660) );
  OAI211_X1 U6752 ( .C1(n5663), .C2(n5662), .A(n5661), .B(n5660), .ZN(U3005)
         );
  INV_X1 U6753 ( .A(n5796), .ZN(n5667) );
  INV_X1 U6754 ( .A(n5664), .ZN(n5666) );
  NAND3_X1 U6755 ( .A1(n5667), .A2(n5666), .A3(n5665), .ZN(n5668) );
  OAI22_X1 U6756 ( .A1(n5669), .A2(n5668), .B1(n4432), .B2(n6432), .ZN(U3455)
         );
  INV_X1 U6757 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6500) );
  AOI221_X2 U6758 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6363), .C2(STATE_REG_0__SCAN_IN), .A(n6458), .ZN(n6427) );
  INV_X1 U6759 ( .A(n6427), .ZN(n6424) );
  OAI21_X1 U6760 ( .B1(n6458), .B2(n6500), .A(n6424), .ZN(U2789) );
  NAND2_X1 U6761 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6453), .ZN(n5672) );
  OAI21_X1 U6762 ( .B1(n5670), .B2(n6347), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5671) );
  OAI21_X1 U6763 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5672), .A(n5671), .ZN(
        U2790) );
  NAND2_X1 U6764 ( .A1(n6514), .A2(n6577), .ZN(n6467) );
  INV_X1 U6765 ( .A(n6467), .ZN(n5674) );
  OAI21_X1 U6766 ( .B1(n5674), .B2(D_C_N_REG_SCAN_IN), .A(n6418), .ZN(n5673)
         );
  OAI21_X1 U6767 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6447), .A(n5673), .ZN(
        U2791) );
  OAI21_X1 U6768 ( .B1(n5674), .B2(BS16_N), .A(n6427), .ZN(n6425) );
  OAI21_X1 U6769 ( .B1(n6427), .B2(n4534), .A(n6425), .ZN(U2792) );
  OAI21_X1 U6770 ( .B1(n5677), .B2(n5676), .A(n5675), .ZN(U2793) );
  NOR4_X1 U6771 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5681) );
  NOR4_X1 U6772 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5680) );
  NOR4_X1 U6773 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U6774 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U6775 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5687)
         );
  NOR4_X1 U6776 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5685) );
  AOI211_X1 U6777 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_28__SCAN_IN), .B(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n5684) );
  NOR4_X1 U6778 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n5683) );
  NOR4_X1 U6779 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5682) );
  NAND4_X1 U6780 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n5686)
         );
  NOR2_X1 U6781 ( .A1(n5687), .A2(n5686), .ZN(n6442) );
  INV_X1 U6782 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5689) );
  NOR3_X1 U6783 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5690) );
  OAI21_X1 U6784 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5690), .A(n6442), .ZN(n5688)
         );
  OAI21_X1 U6785 ( .B1(n6442), .B2(n5689), .A(n5688), .ZN(U2794) );
  INV_X1 U6786 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6426) );
  AOI21_X1 U6787 ( .B1(n6438), .B2(n6426), .A(n5690), .ZN(n5692) );
  INV_X1 U6788 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5691) );
  INV_X1 U6789 ( .A(n6442), .ZN(n6445) );
  AOI22_X1 U6790 ( .A1(n6442), .A2(n5692), .B1(n5691), .B2(n6445), .ZN(U2795)
         );
  OAI21_X1 U6791 ( .B1(n5834), .B2(n6536), .A(n5782), .ZN(n5695) );
  OAI22_X1 U6792 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5693), .B1(n6547), .B2(
        n5836), .ZN(n5694) );
  AOI211_X1 U6793 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5701), .A(n5695), .B(n5694), .ZN(n5699) );
  AOI22_X1 U6794 ( .A1(n2956), .A2(n5697), .B1(n5831), .B2(n5696), .ZN(n5698)
         );
  OAI211_X1 U6795 ( .C1(n5780), .C2(n5700), .A(n5699), .B(n5698), .ZN(U2812)
         );
  AOI22_X1 U6796 ( .A1(n5701), .A2(REIP_REG_14__SCAN_IN), .B1(n5831), .B2(
        n5845), .ZN(n5708) );
  AOI22_X1 U6797 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5821), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n5820), .ZN(n5707) );
  NOR2_X1 U6798 ( .A1(n5817), .A2(REIP_REG_14__SCAN_IN), .ZN(n5702) );
  AOI21_X1 U6799 ( .B1(n5703), .B2(n5702), .A(n5793), .ZN(n5706) );
  AOI22_X1 U6800 ( .A1(n5704), .A2(n5799), .B1(n5770), .B2(n5846), .ZN(n5705)
         );
  NAND4_X1 U6801 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(U2813)
         );
  NOR3_X1 U6802 ( .A1(n5817), .A2(REIP_REG_13__SCAN_IN), .A3(n5709), .ZN(n5714) );
  AOI22_X1 U6803 ( .A1(n5710), .A2(n5831), .B1(n5821), .B2(EBX_REG_13__SCAN_IN), .ZN(n5711) );
  OAI211_X1 U6804 ( .C1(n5834), .C2(n5712), .A(n5711), .B(n5782), .ZN(n5713)
         );
  AOI211_X1 U6805 ( .C1(n5799), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5718)
         );
  INV_X1 U6806 ( .A(n5817), .ZN(n5744) );
  AND3_X1 U6807 ( .A1(n5744), .A2(n6390), .A3(n5716), .ZN(n5722) );
  OAI21_X1 U6808 ( .B1(n5716), .B2(n5817), .A(n5804), .ZN(n5733) );
  OAI21_X1 U6809 ( .B1(n5722), .B2(n5733), .A(REIP_REG_13__SCAN_IN), .ZN(n5717) );
  OAI211_X1 U6810 ( .C1(n5719), .C2(n5780), .A(n5718), .B(n5717), .ZN(U2814)
         );
  AOI22_X1 U6811 ( .A1(n5720), .A2(n5831), .B1(PHYADDRPOINTER_REG_12__SCAN_IN), 
        .B2(n5820), .ZN(n5727) );
  AND2_X1 U6812 ( .A1(n5733), .A2(REIP_REG_12__SCAN_IN), .ZN(n5721) );
  AOI211_X1 U6813 ( .C1(n5821), .C2(EBX_REG_12__SCAN_IN), .A(n5722), .B(n5721), 
        .ZN(n5726) );
  AOI22_X1 U6814 ( .A1(n5724), .A2(n5799), .B1(n5770), .B2(n5723), .ZN(n5725)
         );
  NAND4_X1 U6815 ( .A1(n5727), .A2(n5726), .A3(n5725), .A4(n5782), .ZN(U2815)
         );
  INV_X1 U6816 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5729) );
  OAI22_X1 U6817 ( .A1(n5836), .A2(n5729), .B1(n5834), .B2(n5728), .ZN(n5730)
         );
  AOI211_X1 U6818 ( .C1(n6036), .C2(n5831), .A(n5730), .B(n5793), .ZN(n5735)
         );
  OAI21_X1 U6819 ( .B1(n5817), .B2(n5731), .A(n6388), .ZN(n5732) );
  AOI22_X1 U6820 ( .A1(n5958), .A2(n2956), .B1(n5733), .B2(n5732), .ZN(n5734)
         );
  OAI211_X1 U6821 ( .C1(n5780), .C2(n5961), .A(n5735), .B(n5734), .ZN(U2816)
         );
  OAI22_X1 U6822 ( .A1(n5737), .A2(n5824), .B1(n5736), .B2(n5836), .ZN(n5738)
         );
  AOI211_X1 U6823 ( .C1(n5820), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5793), 
        .B(n5738), .ZN(n5748) );
  AOI22_X1 U6824 ( .A1(n5740), .A2(n2956), .B1(n5770), .B2(n5739), .ZN(n5747)
         );
  INV_X1 U6825 ( .A(n5742), .ZN(n5741) );
  OAI21_X1 U6826 ( .B1(n5741), .B2(n5817), .A(n5804), .ZN(n5760) );
  NOR3_X1 U6827 ( .A1(n5817), .A2(REIP_REG_9__SCAN_IN), .A3(n5742), .ZN(n5749)
         );
  OAI21_X1 U6828 ( .B1(n5760), .B2(n5749), .A(REIP_REG_10__SCAN_IN), .ZN(n5746) );
  NAND3_X1 U6829 ( .A1(n5744), .A2(n4883), .A3(n5743), .ZN(n5745) );
  NAND4_X1 U6830 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(U2817)
         );
  AOI21_X1 U6831 ( .B1(n5760), .B2(REIP_REG_9__SCAN_IN), .A(n5749), .ZN(n5753)
         );
  AOI22_X1 U6832 ( .A1(n6043), .A2(n5831), .B1(n5820), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5750) );
  OAI211_X1 U6833 ( .C1(n5780), .C2(n5971), .A(n5750), .B(n5782), .ZN(n5751)
         );
  AOI21_X1 U6834 ( .B1(n5968), .B2(n2956), .A(n5751), .ZN(n5752) );
  OAI211_X1 U6835 ( .C1(n5754), .C2(n5836), .A(n5753), .B(n5752), .ZN(U2818)
         );
  INV_X1 U6836 ( .A(n5755), .ZN(n6052) );
  OAI22_X1 U6837 ( .A1(n6052), .A2(n5824), .B1(n5756), .B2(n5836), .ZN(n5757)
         );
  AOI211_X1 U6838 ( .C1(n5820), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5793), 
        .B(n5757), .ZN(n5762) );
  NAND2_X1 U6839 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5765) );
  NOR2_X1 U6840 ( .A1(n5817), .A2(n5758), .ZN(n5787) );
  NAND2_X1 U6841 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5787), .ZN(n5777) );
  INV_X1 U6842 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U6843 ( .B1(n5765), .B2(n5777), .A(n6599), .ZN(n5759) );
  AOI22_X1 U6844 ( .A1(n5975), .A2(n2956), .B1(n5760), .B2(n5759), .ZN(n5761)
         );
  OAI211_X1 U6845 ( .C1(n5780), .C2(n5979), .A(n5762), .B(n5761), .ZN(U2819)
         );
  OR2_X1 U6846 ( .A1(n5817), .A2(n5763), .ZN(n5764) );
  AND2_X1 U6847 ( .A1(n5804), .A2(n5764), .ZN(n5776) );
  INV_X1 U6848 ( .A(n5776), .ZN(n5786) );
  INV_X1 U6849 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6516) );
  INV_X1 U6850 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6381) );
  AOI21_X1 U6851 ( .B1(n6516), .B2(n6381), .A(n5777), .ZN(n5766) );
  AOI22_X1 U6852 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5786), .B1(n5766), .B2(n5765), .ZN(n5772) );
  INV_X1 U6853 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5768) );
  AOI22_X1 U6854 ( .A1(n6059), .A2(n5831), .B1(n5821), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5767) );
  OAI211_X1 U6855 ( .C1(n5834), .C2(n5768), .A(n5767), .B(n5782), .ZN(n5769)
         );
  AOI21_X1 U6856 ( .B1(n5770), .B2(n5984), .A(n5769), .ZN(n5771) );
  OAI211_X1 U6857 ( .C1(n5987), .C2(n5835), .A(n5772), .B(n5771), .ZN(U2820)
         );
  OAI22_X1 U6858 ( .A1(n6072), .A2(n5824), .B1(n5773), .B2(n5836), .ZN(n5774)
         );
  AOI211_X1 U6859 ( .C1(n5820), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5793), 
        .B(n5774), .ZN(n5775) );
  OAI221_X1 U6860 ( .B1(REIP_REG_6__SCAN_IN), .B2(n5777), .C1(n6381), .C2(
        n5776), .A(n5775), .ZN(n5778) );
  AOI21_X1 U6861 ( .B1(n5993), .B2(n2956), .A(n5778), .ZN(n5779) );
  OAI21_X1 U6862 ( .B1(n5780), .B2(n5996), .A(n5779), .ZN(U2821) );
  INV_X1 U6863 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5784) );
  INV_X1 U6864 ( .A(n5781), .ZN(n6079) );
  AOI22_X1 U6865 ( .A1(n6079), .A2(n5831), .B1(n5821), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5783) );
  OAI211_X1 U6866 ( .C1(n5834), .C2(n5784), .A(n5783), .B(n5782), .ZN(n5785)
         );
  AOI21_X1 U6867 ( .B1(n6002), .B2(n5828), .A(n5785), .ZN(n5789) );
  OAI21_X1 U6868 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5787), .A(n5786), .ZN(n5788)
         );
  OAI211_X1 U6869 ( .C1(n5835), .C2(n6005), .A(n5789), .B(n5788), .ZN(U2822)
         );
  OAI21_X1 U6870 ( .B1(n5790), .B2(n5794), .A(n5832), .ZN(n5816) );
  OAI22_X1 U6871 ( .A1(n5816), .A2(n6377), .B1(n5791), .B2(n5834), .ZN(n5792)
         );
  AOI211_X1 U6872 ( .C1(n5821), .C2(EBX_REG_4__SCAN_IN), .A(n5793), .B(n5792), 
        .ZN(n5801) );
  NOR3_X1 U6873 ( .A1(n5817), .A2(n5794), .A3(REIP_REG_4__SCAN_IN), .ZN(n5798)
         );
  OAI22_X1 U6874 ( .A1(n5796), .A2(n5838), .B1(n5824), .B2(n5795), .ZN(n5797)
         );
  AOI211_X1 U6875 ( .C1(n5799), .C2(n6011), .A(n5798), .B(n5797), .ZN(n5800)
         );
  OAI211_X1 U6876 ( .C1(n5844), .C2(n6015), .A(n5801), .B(n5800), .ZN(U2823)
         );
  INV_X1 U6877 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6375) );
  INV_X1 U6878 ( .A(n5802), .ZN(n5803) );
  NAND3_X1 U6879 ( .A1(n5804), .A2(REIP_REG_2__SCAN_IN), .A3(n5803), .ZN(n5819) );
  INV_X1 U6880 ( .A(n5838), .ZN(n5811) );
  OR2_X1 U6881 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U6882 ( .A1(n5808), .A2(n5807), .ZN(n5848) );
  AOI22_X1 U6883 ( .A1(n5821), .A2(EBX_REG_3__SCAN_IN), .B1(n5820), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5809) );
  OAI21_X1 U6884 ( .B1(n5848), .B2(n5824), .A(n5809), .ZN(n5810) );
  AOI21_X1 U6885 ( .B1(n5812), .B2(n5811), .A(n5810), .ZN(n5813) );
  OAI21_X1 U6886 ( .B1(n5835), .B2(n6024), .A(n5813), .ZN(n5814) );
  AOI21_X1 U6887 ( .B1(n6021), .B2(n5828), .A(n5814), .ZN(n5815) );
  OAI221_X1 U6888 ( .B1(n5816), .B2(n6375), .C1(n5816), .C2(n5819), .A(n5815), 
        .ZN(U2824) );
  NOR2_X1 U6889 ( .A1(n4416), .A2(n5838), .ZN(n5827) );
  INV_X1 U6890 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6373) );
  OAI21_X1 U6891 ( .B1(n6438), .B2(n5817), .A(n6373), .ZN(n5818) );
  AOI22_X1 U6892 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n5820), .B1(n5819), 
        .B2(n5818), .ZN(n5823) );
  NAND2_X1 U6893 ( .A1(n5821), .A2(EBX_REG_2__SCAN_IN), .ZN(n5822) );
  OAI211_X1 U6894 ( .C1(n5825), .C2(n5824), .A(n5823), .B(n5822), .ZN(n5826)
         );
  AOI211_X1 U6895 ( .C1(n5828), .C2(n6031), .A(n5827), .B(n5826), .ZN(n5829)
         );
  OAI21_X1 U6896 ( .B1(n6034), .B2(n5835), .A(n5829), .ZN(U2825) );
  AOI22_X1 U6897 ( .A1(n5832), .A2(REIP_REG_0__SCAN_IN), .B1(n5831), .B2(n5830), .ZN(n5842) );
  AOI21_X1 U6898 ( .B1(n5835), .B2(n5834), .A(n5833), .ZN(n5840) );
  OAI22_X1 U6899 ( .A1(n3712), .A2(n5838), .B1(n5837), .B2(n5836), .ZN(n5839)
         );
  NOR2_X1 U6900 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  OAI211_X1 U6901 ( .C1(n5844), .C2(n5843), .A(n5842), .B(n5841), .ZN(U2827)
         );
  INV_X1 U6902 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6481) );
  AOI22_X1 U6903 ( .A1(n5846), .A2(n5850), .B1(n5849), .B2(n5845), .ZN(n5847)
         );
  OAI21_X1 U6904 ( .B1(n6481), .B2(n5852), .A(n5847), .ZN(U2845) );
  INV_X1 U6905 ( .A(n5848), .ZN(n6097) );
  AOI22_X1 U6906 ( .A1(n6021), .A2(n5850), .B1(n5849), .B2(n6097), .ZN(n5851)
         );
  OAI21_X1 U6907 ( .B1(n6482), .B2(n5852), .A(n5851), .ZN(U2856) );
  AOI22_X1 U6908 ( .A1(n5853), .A2(n5865), .B1(n5864), .B2(DATAI_18_), .ZN(
        n5855) );
  AOI22_X1 U6909 ( .A1(n5867), .A2(DATAI_2_), .B1(n5861), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6910 ( .A1(n5855), .A2(n5854), .ZN(U2873) );
  INV_X1 U6911 ( .A(DATAI_17_), .ZN(n5856) );
  OAI22_X1 U6912 ( .A1(n5859), .A2(n5858), .B1(n5857), .B2(n5856), .ZN(n5860)
         );
  INV_X1 U6913 ( .A(n5860), .ZN(n5863) );
  AOI22_X1 U6914 ( .A1(n5867), .A2(DATAI_1_), .B1(n5861), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6915 ( .A1(n5863), .A2(n5862), .ZN(U2874) );
  AOI22_X1 U6916 ( .A1(n5866), .A2(n5865), .B1(n5864), .B2(DATAI_16_), .ZN(
        n5869) );
  AOI22_X1 U6917 ( .A1(n5867), .A2(DATAI_0_), .B1(n5861), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6918 ( .A1(n5869), .A2(n5868), .ZN(U2875) );
  INV_X1 U6919 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6584) );
  INV_X1 U6920 ( .A(n5870), .ZN(n5872) );
  AOI22_X1 U6921 ( .A1(n5872), .A2(EAX_REG_23__SCAN_IN), .B1(n6450), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5871) );
  OAI21_X1 U6922 ( .B1(n6584), .B2(n5888), .A(n5871), .ZN(U2900) );
  AOI22_X1 U6923 ( .A1(n5895), .A2(DATAO_REG_16__SCAN_IN), .B1(n5872), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U6924 ( .B1(n5892), .B2(n6553), .A(n5873), .ZN(U2907) );
  INV_X1 U6925 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5952) );
  AOI22_X1 U6926 ( .A1(n5883), .A2(LWORD_REG_15__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5874) );
  OAI21_X1 U6927 ( .B1(n5952), .B2(n5897), .A(n5874), .ZN(U2908) );
  INV_X1 U6928 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5948) );
  AOI22_X1 U6929 ( .A1(n6450), .A2(LWORD_REG_14__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5875) );
  OAI21_X1 U6930 ( .B1(n5948), .B2(n5897), .A(n5875), .ZN(U2909) );
  INV_X1 U6931 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U6932 ( .A1(EAX_REG_13__SCAN_IN), .A2(n5890), .B1(n5895), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5876) );
  OAI21_X1 U6933 ( .B1(n5892), .B2(n6535), .A(n5876), .ZN(U2910) );
  INV_X1 U6934 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5943) );
  AOI22_X1 U6935 ( .A1(n6450), .A2(LWORD_REG_12__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5877) );
  OAI21_X1 U6936 ( .B1(n5943), .B2(n5897), .A(n5877), .ZN(U2911) );
  AOI22_X1 U6937 ( .A1(EAX_REG_11__SCAN_IN), .A2(n5890), .B1(n5895), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6938 ( .B1(n5892), .B2(n6506), .A(n5878), .ZN(U2912) );
  INV_X1 U6939 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5940) );
  AOI22_X1 U6940 ( .A1(n6450), .A2(LWORD_REG_10__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5879) );
  OAI21_X1 U6941 ( .B1(n5940), .B2(n5897), .A(n5879), .ZN(U2913) );
  INV_X1 U6942 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5881) );
  AOI22_X1 U6943 ( .A1(n6450), .A2(LWORD_REG_9__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5880) );
  OAI21_X1 U6944 ( .B1(n5881), .B2(n5897), .A(n5880), .ZN(U2914) );
  INV_X1 U6945 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5936) );
  AOI22_X1 U6946 ( .A1(n6450), .A2(LWORD_REG_8__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5882) );
  OAI21_X1 U6947 ( .B1(n5936), .B2(n5897), .A(n5882), .ZN(U2915) );
  INV_X1 U6948 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5885) );
  AOI22_X1 U6949 ( .A1(n5883), .A2(LWORD_REG_7__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U6950 ( .B1(n5885), .B2(n5897), .A(n5884), .ZN(U2916) );
  AOI22_X1 U6951 ( .A1(n6450), .A2(LWORD_REG_6__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5886) );
  OAI21_X1 U6952 ( .B1(n6517), .B2(n5897), .A(n5886), .ZN(U2917) );
  INV_X1 U6953 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6484) );
  INV_X1 U6954 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n5887) );
  OAI222_X1 U6955 ( .A1(n5888), .A2(n6484), .B1(n5897), .B2(n3735), .C1(n5892), 
        .C2(n5887), .ZN(U2918) );
  AOI22_X1 U6956 ( .A1(n6450), .A2(LWORD_REG_4__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5889) );
  OAI21_X1 U6957 ( .B1(n6555), .B2(n5897), .A(n5889), .ZN(U2919) );
  INV_X1 U6958 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U6959 ( .A1(EAX_REG_3__SCAN_IN), .A2(n5890), .B1(n5895), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U6960 ( .B1(n5892), .B2(n6587), .A(n5891), .ZN(U2920) );
  AOI22_X1 U6961 ( .A1(n6450), .A2(LWORD_REG_2__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U6962 ( .B1(n3722), .B2(n5897), .A(n5893), .ZN(U2921) );
  AOI22_X1 U6963 ( .A1(n6450), .A2(LWORD_REG_1__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5894) );
  OAI21_X1 U6964 ( .B1(n3703), .B2(n5897), .A(n5894), .ZN(U2922) );
  AOI22_X1 U6965 ( .A1(n6450), .A2(LWORD_REG_0__SCAN_IN), .B1(n5895), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5896) );
  OAI21_X1 U6966 ( .B1(n3714), .B2(n5897), .A(n5896), .ZN(U2923) );
  AOI22_X1 U6967 ( .A1(n6614), .A2(UWORD_REG_1__SCAN_IN), .B1(n5949), .B2(
        DATAI_1_), .ZN(n5898) );
  OAI21_X1 U6968 ( .B1(n5899), .B2(n5951), .A(n5898), .ZN(U2925) );
  AOI22_X1 U6969 ( .A1(n6614), .A2(UWORD_REG_2__SCAN_IN), .B1(n5949), .B2(
        DATAI_2_), .ZN(n5901) );
  OAI21_X1 U6970 ( .B1(n6488), .B2(n5951), .A(n5901), .ZN(U2926) );
  AOI22_X1 U6971 ( .A1(n4297), .A2(UWORD_REG_3__SCAN_IN), .B1(n5949), .B2(
        DATAI_3_), .ZN(n5902) );
  OAI21_X1 U6972 ( .B1(n6503), .B2(n5951), .A(n5902), .ZN(U2927) );
  AOI22_X1 U6973 ( .A1(n4297), .A2(UWORD_REG_4__SCAN_IN), .B1(n5949), .B2(
        DATAI_4_), .ZN(n5903) );
  OAI21_X1 U6974 ( .B1(n5904), .B2(n5951), .A(n5903), .ZN(U2928) );
  AOI22_X1 U6975 ( .A1(n4297), .A2(UWORD_REG_6__SCAN_IN), .B1(n5949), .B2(
        DATAI_6_), .ZN(n5905) );
  OAI21_X1 U6976 ( .B1(n5906), .B2(n5951), .A(n5905), .ZN(U2930) );
  AOI22_X1 U6977 ( .A1(n4297), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6613), .ZN(n5907) );
  OAI21_X1 U6978 ( .B1(n5945), .B2(n5933), .A(n5907), .ZN(U2931) );
  INV_X1 U6979 ( .A(DATAI_8_), .ZN(n5908) );
  NOR2_X1 U6980 ( .A1(n5945), .A2(n5908), .ZN(n5934) );
  AOI21_X1 U6981 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n4297), .A(n5934), .ZN(n5909) );
  OAI21_X1 U6982 ( .B1(n5910), .B2(n5951), .A(n5909), .ZN(U2932) );
  INV_X1 U6983 ( .A(DATAI_10_), .ZN(n5911) );
  NOR2_X1 U6984 ( .A1(n5945), .A2(n5911), .ZN(n5938) );
  AOI21_X1 U6985 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n4297), .A(n5938), .ZN(
        n5912) );
  OAI21_X1 U6986 ( .B1(n5913), .B2(n5951), .A(n5912), .ZN(U2934) );
  AOI21_X1 U6987 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6614), .A(n5914), .ZN(
        n5915) );
  OAI21_X1 U6988 ( .B1(n4048), .B2(n5951), .A(n5915), .ZN(U2935) );
  INV_X1 U6989 ( .A(DATAI_13_), .ZN(n6578) );
  AOI22_X1 U6990 ( .A1(n4297), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6613), .ZN(n5916) );
  OAI21_X1 U6991 ( .B1(n5945), .B2(n6578), .A(n5916), .ZN(U2937) );
  INV_X1 U6992 ( .A(DATAI_14_), .ZN(n5917) );
  NOR2_X1 U6993 ( .A1(n5945), .A2(n5917), .ZN(n5946) );
  AOI21_X1 U6994 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6614), .A(n5946), .ZN(
        n5918) );
  OAI21_X1 U6995 ( .B1(n5919), .B2(n5951), .A(n5918), .ZN(U2938) );
  AOI22_X1 U6996 ( .A1(n4297), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6613), .ZN(n5920) );
  OAI21_X1 U6997 ( .B1(n5945), .B2(n5921), .A(n5920), .ZN(U2939) );
  AOI22_X1 U6998 ( .A1(n4297), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6613), .ZN(n5922) );
  OAI21_X1 U6999 ( .B1(n5945), .B2(n5923), .A(n5922), .ZN(U2940) );
  AOI22_X1 U7000 ( .A1(n6614), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6613), .ZN(n5924) );
  OAI21_X1 U7001 ( .B1(n5945), .B2(n5925), .A(n5924), .ZN(U2941) );
  AOI22_X1 U7002 ( .A1(n6614), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6613), .ZN(n5926) );
  OAI21_X1 U7003 ( .B1(n5945), .B2(n4477), .A(n5926), .ZN(U2942) );
  AOI22_X1 U7004 ( .A1(n6614), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6613), .ZN(n5927) );
  OAI21_X1 U7005 ( .B1(n5945), .B2(n5928), .A(n5927), .ZN(U2943) );
  AOI22_X1 U7006 ( .A1(n6614), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6613), .ZN(n5929) );
  OAI21_X1 U7007 ( .B1(n5945), .B2(n4298), .A(n5929), .ZN(U2944) );
  AOI22_X1 U7008 ( .A1(n6614), .A2(LWORD_REG_6__SCAN_IN), .B1(n6613), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n5930) );
  OAI21_X1 U7009 ( .B1(n5945), .B2(n5931), .A(n5930), .ZN(U2945) );
  AOI22_X1 U7010 ( .A1(n6614), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6613), .ZN(n5932) );
  OAI21_X1 U7011 ( .B1(n5945), .B2(n5933), .A(n5932), .ZN(U2946) );
  AOI21_X1 U7012 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6614), .A(n5934), .ZN(n5935) );
  OAI21_X1 U7013 ( .B1(n5936), .B2(n5951), .A(n5935), .ZN(U2947) );
  AOI22_X1 U7014 ( .A1(n6614), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6613), .ZN(n5937) );
  NAND2_X1 U7015 ( .A1(n5949), .A2(DATAI_9_), .ZN(n6615) );
  NAND2_X1 U7016 ( .A1(n5937), .A2(n6615), .ZN(U2948) );
  AOI21_X1 U7017 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6614), .A(n5938), .ZN(
        n5939) );
  OAI21_X1 U7018 ( .B1(n5940), .B2(n5951), .A(n5939), .ZN(U2949) );
  AOI21_X1 U7019 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6614), .A(n5941), .ZN(
        n5942) );
  OAI21_X1 U7020 ( .B1(n5943), .B2(n5951), .A(n5942), .ZN(U2951) );
  AOI22_X1 U7021 ( .A1(n6614), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6613), .ZN(n5944) );
  OAI21_X1 U7022 ( .B1(n5945), .B2(n6578), .A(n5944), .ZN(U2952) );
  AOI21_X1 U7023 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6614), .A(n5946), .ZN(
        n5947) );
  OAI21_X1 U7024 ( .B1(n5948), .B2(n5951), .A(n5947), .ZN(U2953) );
  AOI22_X1 U7025 ( .A1(n4297), .A2(LWORD_REG_15__SCAN_IN), .B1(n5949), .B2(
        DATAI_15_), .ZN(n5950) );
  OAI21_X1 U7026 ( .B1(n5952), .B2(n5951), .A(n5950), .ZN(U2954) );
  AOI22_X1 U7027 ( .A1(n6104), .A2(REIP_REG_11__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7028 ( .A1(n5953), .A2(n5954), .ZN(n5957) );
  XNOR2_X1 U7029 ( .A(n2965), .B(n5955), .ZN(n5956) );
  XNOR2_X1 U7030 ( .A(n5957), .B(n5956), .ZN(n6038) );
  AOI22_X1 U7031 ( .A1(n6029), .A2(n6038), .B1(n6012), .B2(n5958), .ZN(n5959)
         );
  OAI211_X1 U7032 ( .C1(n4314), .C2(n5961), .A(n5960), .B(n5959), .ZN(U2975)
         );
  AOI22_X1 U7033 ( .A1(n6104), .A2(REIP_REG_9__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7034 ( .A1(n5963), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7035 ( .A1(n5974), .A2(n5964), .ZN(n5967) );
  XNOR2_X1 U7036 ( .A(n2965), .B(n5965), .ZN(n5966) );
  XNOR2_X1 U7037 ( .A(n5967), .B(n5966), .ZN(n6045) );
  AOI22_X1 U7038 ( .A1(n6045), .A2(n6029), .B1(n6012), .B2(n5968), .ZN(n5969)
         );
  OAI211_X1 U7039 ( .C1(n4314), .C2(n5971), .A(n5970), .B(n5969), .ZN(U2977)
         );
  AOI22_X1 U7040 ( .A1(n6104), .A2(REIP_REG_8__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7041 ( .A1(n5963), .A2(n5972), .ZN(n5973) );
  NAND2_X1 U7042 ( .A1(n5974), .A2(n5973), .ZN(n6051) );
  INV_X1 U7043 ( .A(n6051), .ZN(n5976) );
  AOI22_X1 U7044 ( .A1(n5976), .A2(n6029), .B1(n6012), .B2(n5975), .ZN(n5977)
         );
  OAI211_X1 U7045 ( .C1(n4314), .C2(n5979), .A(n5978), .B(n5977), .ZN(U2978)
         );
  AOI22_X1 U7046 ( .A1(n6104), .A2(REIP_REG_7__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5986) );
  OR2_X1 U7047 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  AND2_X1 U7048 ( .A1(n5983), .A2(n5982), .ZN(n6061) );
  AOI22_X1 U7049 ( .A1(n5984), .A2(n6030), .B1(n6029), .B2(n6061), .ZN(n5985)
         );
  OAI211_X1 U7050 ( .C1(n6035), .C2(n5987), .A(n5986), .B(n5985), .ZN(U2979)
         );
  AOI22_X1 U7051 ( .A1(n6104), .A2(REIP_REG_6__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5995) );
  OAI21_X1 U7052 ( .B1(n5989), .B2(n5991), .A(n5990), .ZN(n5992) );
  INV_X1 U7053 ( .A(n5992), .ZN(n6074) );
  AOI22_X1 U7054 ( .A1(n6074), .A2(n6029), .B1(n6012), .B2(n5993), .ZN(n5994)
         );
  OAI211_X1 U7055 ( .C1(n4314), .C2(n5996), .A(n5995), .B(n5994), .ZN(U2980)
         );
  AOI22_X1 U7056 ( .A1(n6104), .A2(REIP_REG_5__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7057 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7058 ( .A1(n5997), .A2(n6000), .ZN(n6084) );
  INV_X1 U7059 ( .A(n6084), .ZN(n6001) );
  AOI22_X1 U7060 ( .A1(n6002), .A2(n6030), .B1(n6029), .B2(n6001), .ZN(n6003)
         );
  OAI211_X1 U7061 ( .C1(n6035), .C2(n6005), .A(n6004), .B(n6003), .ZN(U2981)
         );
  AOI22_X1 U7062 ( .A1(n6104), .A2(REIP_REG_4__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7063 ( .B1(n6006), .B2(n6009), .A(n6008), .ZN(n6010) );
  INV_X1 U7064 ( .A(n6010), .ZN(n6091) );
  AOI22_X1 U7065 ( .A1(n6091), .A2(n6029), .B1(n6012), .B2(n6011), .ZN(n6013)
         );
  OAI211_X1 U7066 ( .C1(n4314), .C2(n6015), .A(n6014), .B(n6013), .ZN(U2982)
         );
  AOI22_X1 U7067 ( .A1(n6104), .A2(REIP_REG_3__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7068 ( .B1(n6019), .B2(n6017), .A(n6018), .ZN(n6020) );
  INV_X1 U7069 ( .A(n6020), .ZN(n6098) );
  AOI22_X1 U7070 ( .A1(n6098), .A2(n6029), .B1(n6021), .B2(n6030), .ZN(n6022)
         );
  OAI211_X1 U7071 ( .C1(n6035), .C2(n6024), .A(n6023), .B(n6022), .ZN(U2983)
         );
  AOI22_X1 U7072 ( .A1(n6104), .A2(REIP_REG_2__SCAN_IN), .B1(n6025), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7073 ( .A(n6027), .B(n3312), .ZN(n6028) );
  XNOR2_X1 U7074 ( .A(n6026), .B(n6028), .ZN(n6110) );
  AOI22_X1 U7075 ( .A1(n6031), .A2(n6030), .B1(n6110), .B2(n6029), .ZN(n6032)
         );
  OAI211_X1 U7076 ( .C1(n6035), .C2(n6034), .A(n6033), .B(n6032), .ZN(U2984)
         );
  AOI22_X1 U7077 ( .A1(n6106), .A2(n6036), .B1(n6104), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6040) );
  AOI22_X1 U7078 ( .A1(n6126), .A2(n6038), .B1(n5955), .B2(n6037), .ZN(n6039)
         );
  OAI211_X1 U7079 ( .C1(n5955), .C2(n6041), .A(n6040), .B(n6039), .ZN(U3007)
         );
  INV_X1 U7080 ( .A(n6042), .ZN(n6048) );
  AOI22_X1 U7081 ( .A1(n6106), .A2(n6043), .B1(n6104), .B2(REIP_REG_9__SCAN_IN), .ZN(n6047) );
  AOI22_X1 U7082 ( .A1(n6045), .A2(n6126), .B1(n6044), .B2(n5965), .ZN(n6046)
         );
  OAI211_X1 U7083 ( .C1(n6048), .C2(n5965), .A(n6047), .B(n6046), .ZN(U3009)
         );
  AOI211_X1 U7084 ( .C1(n6050), .C2(n6057), .A(n6049), .B(n6064), .ZN(n6055)
         );
  NOR2_X1 U7085 ( .A1(n6051), .A2(n6083), .ZN(n6054) );
  OAI22_X1 U7086 ( .A1(n6120), .A2(n6052), .B1(n6599), .B2(n6071), .ZN(n6053)
         );
  NOR3_X1 U7087 ( .A1(n6055), .A2(n6054), .A3(n6053), .ZN(n6056) );
  OAI21_X1 U7088 ( .B1(n6058), .B2(n6057), .A(n6056), .ZN(U3010) );
  AOI22_X1 U7089 ( .A1(n6106), .A2(n6059), .B1(n6104), .B2(REIP_REG_7__SCAN_IN), .ZN(n6063) );
  AOI22_X1 U7090 ( .A1(n6061), .A2(n6126), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6060), .ZN(n6062) );
  OAI211_X1 U7091 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6064), .A(n6063), 
        .B(n6062), .ZN(U3011) );
  NAND3_X1 U7092 ( .A1(n6078), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6065), 
        .ZN(n6077) );
  NAND2_X1 U7093 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6078), .ZN(n6069)
         );
  INV_X1 U7094 ( .A(n6080), .ZN(n6108) );
  INV_X1 U7095 ( .A(n6066), .ZN(n6067) );
  OAI21_X1 U7096 ( .B1(n6068), .B2(n6108), .A(n6067), .ZN(n6111) );
  AOI21_X1 U7097 ( .B1(n6070), .B2(n6069), .A(n6111), .ZN(n6090) );
  OAI22_X1 U7098 ( .A1(n6120), .A2(n6072), .B1(n6381), .B2(n6071), .ZN(n6073)
         );
  AOI21_X1 U7099 ( .B1(n6074), .B2(n6126), .A(n6073), .ZN(n6075) );
  OAI221_X1 U7100 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6077), .C1(n6076), .C2(n6090), .A(n6075), .ZN(U3012) );
  AOI21_X1 U7101 ( .B1(n6107), .B2(n6078), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6089) );
  AOI22_X1 U7102 ( .A1(n6106), .A2(n6079), .B1(n6104), .B2(REIP_REG_5__SCAN_IN), .ZN(n6088) );
  NOR2_X1 U7103 ( .A1(n6080), .A2(n6094), .ZN(n6081) );
  NAND2_X1 U7104 ( .A1(n6082), .A2(n6081), .ZN(n6085) );
  OAI22_X1 U7105 ( .A1(n6112), .A2(n6085), .B1(n6084), .B2(n6083), .ZN(n6086)
         );
  INV_X1 U7106 ( .A(n6086), .ZN(n6087) );
  OAI211_X1 U7107 ( .C1(n6090), .C2(n6089), .A(n6088), .B(n6087), .ZN(U3013)
         );
  AOI21_X1 U7108 ( .B1(n6107), .B2(n6109), .A(n6111), .ZN(n6103) );
  AOI222_X1 U7109 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6104), .B1(n6106), .B2(
        n6092), .C1(n6126), .C2(n6091), .ZN(n6096) );
  NOR2_X1 U7110 ( .A1(n6109), .A2(n6093), .ZN(n6099) );
  OAI211_X1 U7111 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6099), .B(n6094), .ZN(n6095) );
  OAI211_X1 U7112 ( .C1(n6103), .C2(n6522), .A(n6096), .B(n6095), .ZN(U3014)
         );
  AOI22_X1 U7113 ( .A1(n6106), .A2(n6097), .B1(n6104), .B2(REIP_REG_3__SCAN_IN), .ZN(n6101) );
  AOI22_X1 U7114 ( .A1(n6099), .A2(n6102), .B1(n6098), .B2(n6126), .ZN(n6100)
         );
  OAI211_X1 U7115 ( .C1(n6103), .C2(n6102), .A(n6101), .B(n6100), .ZN(U3015)
         );
  AOI22_X1 U7116 ( .A1(n6106), .A2(n6105), .B1(n6104), .B2(REIP_REG_2__SCAN_IN), .ZN(n6117) );
  OAI221_X1 U7117 ( .B1(n6109), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6109), .C2(n6108), .A(n6107), .ZN(n6116) );
  AOI22_X1 U7118 ( .A1(n6111), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6126), 
        .B2(n6110), .ZN(n6115) );
  INV_X1 U7119 ( .A(n6112), .ZN(n6113) );
  NAND3_X1 U7120 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6113), .A3(n3312), 
        .ZN(n6114) );
  NAND4_X1 U7121 ( .A1(n6117), .A2(n6116), .A3(n6115), .A4(n6114), .ZN(U3016)
         );
  OAI21_X1 U7122 ( .B1(n6120), .B2(n6119), .A(n6118), .ZN(n6124) );
  NOR3_X1 U7123 ( .A1(n6122), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6121), 
        .ZN(n6123) );
  AOI211_X1 U7124 ( .C1(n6126), .C2(n6125), .A(n6124), .B(n6123), .ZN(n6127)
         );
  OAI221_X1 U7125 ( .B1(n6507), .B2(n6129), .C1(n6507), .C2(n6128), .A(n6127), 
        .ZN(U3017) );
  NOR2_X1 U7126 ( .A1(n6314), .A2(n6130), .ZN(U3019) );
  AOI22_X1 U7127 ( .A1(n2958), .A2(n3014), .B1(n6230), .B2(n6152), .ZN(n6141)
         );
  NAND3_X1 U7128 ( .A1(n6132), .A2(n6232), .A3(n6131), .ZN(n6133) );
  NAND2_X1 U7129 ( .A1(n6133), .A2(n6233), .ZN(n6139) );
  AOI21_X1 U7130 ( .B1(n6134), .B2(n6298), .A(n3014), .ZN(n6138) );
  INV_X1 U7131 ( .A(n6138), .ZN(n6136) );
  AOI21_X1 U7132 ( .B1(n6238), .B2(n6137), .A(n6237), .ZN(n6135) );
  OAI22_X1 U7133 ( .A1(n6139), .A2(n6138), .B1(n6137), .B2(n6326), .ZN(n6160)
         );
  AOI22_X1 U7134 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6161), .B1(n6244), 
        .B2(n6160), .ZN(n6140) );
  OAI211_X1 U7135 ( .C1(n6247), .C2(n6155), .A(n6141), .B(n6140), .ZN(U3044)
         );
  AOI22_X1 U7136 ( .A1(n6249), .A2(n3014), .B1(n6182), .B2(n6152), .ZN(n6143)
         );
  AOI22_X1 U7137 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6161), .B1(n6250), 
        .B2(n6160), .ZN(n6142) );
  OAI211_X1 U7138 ( .C1(n6155), .C2(n6144), .A(n6143), .B(n6142), .ZN(U3045)
         );
  AOI22_X1 U7139 ( .A1(n6255), .A2(n3014), .B1(n6254), .B2(n6152), .ZN(n6146)
         );
  AOI22_X1 U7140 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6161), .B1(n6256), 
        .B2(n6160), .ZN(n6145) );
  OAI211_X1 U7141 ( .C1(n6155), .C2(n6259), .A(n6146), .B(n6145), .ZN(U3046)
         );
  AOI22_X1 U7142 ( .A1(n6261), .A2(n3014), .B1(n6190), .B2(n6159), .ZN(n6148)
         );
  AOI22_X1 U7143 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6161), .B1(n6262), 
        .B2(n6160), .ZN(n6147) );
  OAI211_X1 U7144 ( .C1(n6149), .C2(n6164), .A(n6148), .B(n6147), .ZN(U3047)
         );
  AOI22_X1 U7145 ( .A1(n6267), .A2(n3014), .B1(n6216), .B2(n6152), .ZN(n6151)
         );
  AOI22_X1 U7146 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6161), .B1(n6268), 
        .B2(n6160), .ZN(n6150) );
  OAI211_X1 U7147 ( .C1(n6155), .C2(n6219), .A(n6151), .B(n6150), .ZN(U3048)
         );
  AOI22_X1 U7148 ( .A1(n6274), .A2(n3014), .B1(n6223), .B2(n6152), .ZN(n6154)
         );
  AOI22_X1 U7149 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6161), .B1(n6275), 
        .B2(n6160), .ZN(n6153) );
  OAI211_X1 U7150 ( .C1(n6155), .C2(n6228), .A(n6154), .B(n6153), .ZN(U3049)
         );
  AOI22_X1 U7151 ( .A1(n6281), .A2(n3014), .B1(n6200), .B2(n6159), .ZN(n6157)
         );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6161), .B1(n6282), 
        .B2(n6160), .ZN(n6156) );
  OAI211_X1 U7153 ( .C1(n6158), .C2(n6164), .A(n6157), .B(n6156), .ZN(U3050)
         );
  AOI22_X1 U7154 ( .A1(n6288), .A2(n3014), .B1(n6205), .B2(n6159), .ZN(n6163)
         );
  AOI22_X1 U7155 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6161), .B1(n6290), 
        .B2(n6160), .ZN(n6162) );
  OAI211_X1 U7156 ( .C1(n6165), .C2(n6164), .A(n6163), .B(n6162), .ZN(U3051)
         );
  NOR2_X1 U7157 ( .A1(n3712), .A2(n6167), .ZN(n6168) );
  NAND2_X1 U7158 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7159 ( .A1(n6170), .A2(n6171), .ZN(n6172) );
  AOI22_X1 U7160 ( .A1(n6174), .A2(n6172), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6177), .ZN(n6212) );
  INV_X1 U7161 ( .A(n6171), .ZN(n6206) );
  AOI22_X1 U7162 ( .A1(n2958), .A2(n6206), .B1(n6230), .B2(n6207), .ZN(n6180)
         );
  INV_X1 U7163 ( .A(n6172), .ZN(n6173) );
  NAND2_X1 U7164 ( .A1(n6174), .A2(n6173), .ZN(n6176) );
  OAI211_X1 U7165 ( .C1(n6233), .C2(n6177), .A(n6176), .B(n6175), .ZN(n6208)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6208), .B1(n6178), 
        .B2(n6204), .ZN(n6179) );
  OAI211_X1 U7167 ( .C1(n6212), .C2(n6181), .A(n6180), .B(n6179), .ZN(U3076)
         );
  AOI22_X1 U7168 ( .A1(n6249), .A2(n6206), .B1(n6182), .B2(n6207), .ZN(n6184)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6208), .B1(n6248), 
        .B2(n6204), .ZN(n6183) );
  OAI211_X1 U7170 ( .C1(n6212), .C2(n6185), .A(n6184), .B(n6183), .ZN(U3077)
         );
  AOI22_X1 U7171 ( .A1(n6255), .A2(n6206), .B1(n6186), .B2(n6204), .ZN(n6188)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6208), .B1(n6254), 
        .B2(n6207), .ZN(n6187) );
  OAI211_X1 U7173 ( .C1(n6212), .C2(n6189), .A(n6188), .B(n6187), .ZN(U3078)
         );
  AOI22_X1 U7174 ( .A1(n6261), .A2(n6206), .B1(n6260), .B2(n6207), .ZN(n6192)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6208), .B1(n6190), 
        .B2(n6204), .ZN(n6191) );
  OAI211_X1 U7176 ( .C1(n6212), .C2(n6193), .A(n6192), .B(n6191), .ZN(U3079)
         );
  AOI22_X1 U7177 ( .A1(n6267), .A2(n6206), .B1(n6216), .B2(n6207), .ZN(n6195)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6208), .B1(n6266), 
        .B2(n6204), .ZN(n6194) );
  OAI211_X1 U7179 ( .C1(n6212), .C2(n6196), .A(n6195), .B(n6194), .ZN(U3080)
         );
  AOI22_X1 U7180 ( .A1(n6274), .A2(n6206), .B1(n6272), .B2(n6204), .ZN(n6198)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6208), .B1(n6223), 
        .B2(n6207), .ZN(n6197) );
  OAI211_X1 U7182 ( .C1(n6212), .C2(n6199), .A(n6198), .B(n6197), .ZN(U3081)
         );
  AOI22_X1 U7183 ( .A1(n6281), .A2(n6206), .B1(n6200), .B2(n6204), .ZN(n6202)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6208), .B1(n6280), 
        .B2(n6207), .ZN(n6201) );
  OAI211_X1 U7185 ( .C1(n6212), .C2(n6203), .A(n6202), .B(n6201), .ZN(U3082)
         );
  AOI22_X1 U7186 ( .A1(n6288), .A2(n6206), .B1(n6205), .B2(n6204), .ZN(n6210)
         );
  AOI22_X1 U7187 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6208), .B1(n6287), 
        .B2(n6207), .ZN(n6209) );
  OAI211_X1 U7188 ( .C1(n6212), .C2(n6211), .A(n6210), .B(n6209), .ZN(U3083)
         );
  INV_X1 U7189 ( .A(n6213), .ZN(n6221) );
  AOI22_X1 U7190 ( .A1(n6256), .A2(n6221), .B1(n6255), .B2(n6220), .ZN(n6215)
         );
  AOI22_X1 U7191 ( .A1(n6224), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6254), 
        .B2(n6222), .ZN(n6214) );
  OAI211_X1 U7192 ( .C1(n6259), .C2(n6227), .A(n6215), .B(n6214), .ZN(U3086)
         );
  AOI22_X1 U7193 ( .A1(n6268), .A2(n6221), .B1(n6267), .B2(n6220), .ZN(n6218)
         );
  AOI22_X1 U7194 ( .A1(n6224), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6216), 
        .B2(n6222), .ZN(n6217) );
  OAI211_X1 U7195 ( .C1(n6219), .C2(n6227), .A(n6218), .B(n6217), .ZN(U3088)
         );
  AOI22_X1 U7196 ( .A1(n6275), .A2(n6221), .B1(n6274), .B2(n6220), .ZN(n6226)
         );
  AOI22_X1 U7197 ( .A1(n6224), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6223), 
        .B2(n6222), .ZN(n6225) );
  OAI211_X1 U7198 ( .C1(n6228), .C2(n6227), .A(n6226), .B(n6225), .ZN(U3089)
         );
  AOI22_X1 U7199 ( .A1(n2958), .A2(n3012), .B1(n6230), .B2(n6286), .ZN(n6246)
         );
  INV_X1 U7200 ( .A(n6232), .ZN(n6234) );
  OAI21_X1 U7201 ( .B1(n6235), .B2(n6234), .A(n6233), .ZN(n6243) );
  AOI21_X1 U7202 ( .B1(n6236), .B2(n6298), .A(n3012), .ZN(n6242) );
  INV_X1 U7203 ( .A(n6242), .ZN(n6240) );
  AOI21_X1 U7204 ( .B1(n6238), .B2(n6241), .A(n6237), .ZN(n6239) );
  OAI21_X1 U7205 ( .B1(n6243), .B2(n6240), .A(n6239), .ZN(n6291) );
  OAI22_X1 U7206 ( .A1(n6243), .A2(n6242), .B1(n6241), .B2(n6326), .ZN(n6289)
         );
  AOI22_X1 U7207 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6291), .B1(n6244), 
        .B2(n6289), .ZN(n6245) );
  OAI211_X1 U7208 ( .C1(n6247), .C2(n6294), .A(n6246), .B(n6245), .ZN(U3108)
         );
  INV_X1 U7209 ( .A(n6294), .ZN(n6273) );
  AOI22_X1 U7210 ( .A1(n6249), .A2(n3012), .B1(n6273), .B2(n6248), .ZN(n6252)
         );
  AOI22_X1 U7211 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6291), .B1(n6250), 
        .B2(n6289), .ZN(n6251) );
  OAI211_X1 U7212 ( .C1(n6253), .C2(n6278), .A(n6252), .B(n6251), .ZN(U3109)
         );
  AOI22_X1 U7213 ( .A1(n6255), .A2(n3012), .B1(n6254), .B2(n6286), .ZN(n6258)
         );
  AOI22_X1 U7214 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6291), .B1(n6256), 
        .B2(n6289), .ZN(n6257) );
  OAI211_X1 U7215 ( .C1(n6259), .C2(n6294), .A(n6258), .B(n6257), .ZN(U3110)
         );
  AOI22_X1 U7216 ( .A1(n6261), .A2(n3012), .B1(n6260), .B2(n6286), .ZN(n6264)
         );
  AOI22_X1 U7217 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6291), .B1(n6262), 
        .B2(n6289), .ZN(n6263) );
  OAI211_X1 U7218 ( .C1(n6265), .C2(n6294), .A(n6264), .B(n6263), .ZN(U3111)
         );
  AOI22_X1 U7219 ( .A1(n6267), .A2(n3012), .B1(n6273), .B2(n6266), .ZN(n6270)
         );
  AOI22_X1 U7220 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6291), .B1(n6268), 
        .B2(n6289), .ZN(n6269) );
  OAI211_X1 U7221 ( .C1(n6271), .C2(n6278), .A(n6270), .B(n6269), .ZN(U3112)
         );
  AOI22_X1 U7222 ( .A1(n6274), .A2(n3012), .B1(n6273), .B2(n6272), .ZN(n6277)
         );
  AOI22_X1 U7223 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6291), .B1(n6275), 
        .B2(n6289), .ZN(n6276) );
  OAI211_X1 U7224 ( .C1(n6279), .C2(n6278), .A(n6277), .B(n6276), .ZN(U3113)
         );
  AOI22_X1 U7225 ( .A1(n6281), .A2(n3012), .B1(n6280), .B2(n6286), .ZN(n6284)
         );
  AOI22_X1 U7226 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6291), .B1(n6282), 
        .B2(n6289), .ZN(n6283) );
  OAI211_X1 U7227 ( .C1(n6285), .C2(n6294), .A(n6284), .B(n6283), .ZN(U3114)
         );
  AOI22_X1 U7228 ( .A1(n6288), .A2(n3012), .B1(n6287), .B2(n6286), .ZN(n6293)
         );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6291), .B1(n6290), 
        .B2(n6289), .ZN(n6292) );
  OAI211_X1 U7230 ( .C1(n6295), .C2(n6294), .A(n6293), .B(n6292), .ZN(U3115)
         );
  AOI22_X1 U7231 ( .A1(n6298), .A2(n6297), .B1(n3527), .B2(n6296), .ZN(n6431)
         );
  NAND2_X1 U7232 ( .A1(n6299), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6437) );
  NAND3_X1 U7233 ( .A1(n6431), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6437), .ZN(n6302) );
  OAI211_X1 U7234 ( .C1(n6303), .C2(n6302), .A(n6301), .B(n6300), .ZN(n6305)
         );
  NAND2_X1 U7235 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  NAND2_X1 U7236 ( .A1(n6305), .A2(n6304), .ZN(n6310) );
  NAND2_X1 U7237 ( .A1(n6309), .A2(n6310), .ZN(n6306) );
  NAND2_X1 U7238 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  OAI21_X1 U7239 ( .B1(n6310), .B2(n6309), .A(n6308), .ZN(n6311) );
  OAI21_X1 U7240 ( .B1(n6312), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6311), 
        .ZN(n6315) );
  NAND2_X1 U7241 ( .A1(n6312), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6313) );
  NAND3_X1 U7242 ( .A1(n6315), .A2(n6314), .A3(n6313), .ZN(n6325) );
  NOR2_X1 U7243 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6319) );
  NOR2_X1 U7244 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  OAI21_X1 U7245 ( .B1(n6320), .B2(n6319), .A(n6318), .ZN(n6321) );
  NOR2_X1 U7246 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  NAND2_X1 U7247 ( .A1(READY_N), .A2(n6326), .ZN(n6354) );
  OAI211_X1 U7248 ( .C1(n6330), .C2(n6328), .A(n6327), .B(n6354), .ZN(n6337)
         );
  NAND2_X1 U7249 ( .A1(n6330), .A2(n6329), .ZN(n6332) );
  NAND2_X1 U7250 ( .A1(READY_N), .A2(n6450), .ZN(n6331) );
  NAND2_X1 U7251 ( .A1(n6332), .A2(n6331), .ZN(n6336) );
  OR2_X1 U7252 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  NOR2_X1 U7253 ( .A1(n6337), .A2(n6345), .ZN(n6341) );
  OAI21_X1 U7254 ( .B1(n6339), .B2(n6338), .A(n6530), .ZN(n6340) );
  OAI22_X1 U7255 ( .A1(n6530), .A2(n6341), .B1(n6345), .B2(n6340), .ZN(n6342)
         );
  OR2_X1 U7256 ( .A1(n6343), .A2(n6342), .ZN(U3148) );
  INV_X1 U7257 ( .A(n6345), .ZN(n6430) );
  INV_X1 U7258 ( .A(n6354), .ZN(n6350) );
  NOR2_X1 U7259 ( .A1(n6344), .A2(n6453), .ZN(n6353) );
  AOI221_X1 U7260 ( .B1(READY_N), .B2(n6347), .C1(n6346), .C2(n6347), .A(n6345), .ZN(n6348) );
  AOI211_X1 U7261 ( .C1(n6350), .C2(n6353), .A(n6349), .B(n6348), .ZN(n6351)
         );
  OAI21_X1 U7262 ( .B1(n6352), .B2(n6430), .A(n6351), .ZN(U3149) );
  NAND3_X1 U7263 ( .A1(n6354), .A2(n6353), .A3(n6428), .ZN(n6356) );
  NAND2_X1 U7264 ( .A1(n6356), .A2(n6355), .ZN(U3150) );
  AND2_X1 U7265 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6424), .ZN(U3151) );
  AND2_X1 U7266 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6424), .ZN(U3152) );
  AND2_X1 U7267 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6424), .ZN(U3153) );
  INV_X1 U7268 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6491) );
  NOR2_X1 U7269 ( .A1(n6427), .A2(n6491), .ZN(U3154) );
  AND2_X1 U7270 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6424), .ZN(U3155) );
  AND2_X1 U7271 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6424), .ZN(U3156) );
  AND2_X1 U7272 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6424), .ZN(U3157) );
  INV_X1 U7273 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6566) );
  NOR2_X1 U7274 ( .A1(n6427), .A2(n6566), .ZN(U3158) );
  AND2_X1 U7275 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6424), .ZN(U3159) );
  AND2_X1 U7276 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6424), .ZN(U3160) );
  AND2_X1 U7277 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6424), .ZN(U3161) );
  AND2_X1 U7278 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6424), .ZN(U3162) );
  AND2_X1 U7279 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6424), .ZN(U3163) );
  AND2_X1 U7280 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6424), .ZN(U3164) );
  AND2_X1 U7281 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6424), .ZN(U3165) );
  AND2_X1 U7282 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6424), .ZN(U3166) );
  AND2_X1 U7283 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6424), .ZN(U3167) );
  INV_X1 U7284 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6498) );
  NOR2_X1 U7285 ( .A1(n6427), .A2(n6498), .ZN(U3168) );
  AND2_X1 U7286 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6424), .ZN(U3169) );
  AND2_X1 U7287 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6424), .ZN(U3170) );
  INV_X1 U7288 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6583) );
  NOR2_X1 U7289 ( .A1(n6427), .A2(n6583), .ZN(U3171) );
  AND2_X1 U7290 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6424), .ZN(U3172) );
  AND2_X1 U7291 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6424), .ZN(U3173) );
  AND2_X1 U7292 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6424), .ZN(U3174) );
  AND2_X1 U7293 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6424), .ZN(U3175) );
  AND2_X1 U7294 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6424), .ZN(U3176) );
  AND2_X1 U7295 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6424), .ZN(U3177) );
  AND2_X1 U7296 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6424), .ZN(U3178) );
  AND2_X1 U7297 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6424), .ZN(U3179) );
  AND2_X1 U7298 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6424), .ZN(U3180) );
  AOI22_X1 U7299 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6369) );
  AND2_X1 U7300 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6360) );
  INV_X1 U7301 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6358) );
  INV_X1 U7302 ( .A(NA_N), .ZN(n6366) );
  AOI211_X1 U7303 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6366), .A(
        STATE_REG_0__SCAN_IN), .B(n6365), .ZN(n6371) );
  AOI221_X1 U7304 ( .B1(n6360), .B2(n6418), .C1(n6358), .C2(n6418), .A(n6371), 
        .ZN(n6357) );
  OAI21_X1 U7305 ( .B1(n6365), .B2(n6369), .A(n6357), .ZN(U3181) );
  NOR2_X1 U7306 ( .A1(n6514), .A2(n6358), .ZN(n6367) );
  NAND2_X1 U7307 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6359) );
  OAI21_X1 U7308 ( .B1(n6367), .B2(n6360), .A(n6359), .ZN(n6361) );
  OAI211_X1 U7309 ( .C1(n6363), .C2(n4295), .A(n6362), .B(n6361), .ZN(U3182)
         );
  AOI221_X1 U7310 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4295), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6364) );
  AOI221_X1 U7311 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6364), .C2(HOLD), .A(n6514), .ZN(n6370) );
  AOI21_X1 U7312 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6368) );
  OAI22_X1 U7313 ( .A1(n6371), .A2(n6370), .B1(n6369), .B2(n6368), .ZN(U3183)
         );
  AND2_X1 U7314 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6458), .ZN(n6414) );
  INV_X1 U7315 ( .A(n6414), .ZN(n6421) );
  AOI22_X1 U7316 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6447), .ZN(n6372) );
  OAI21_X1 U7317 ( .B1(n6438), .B2(n6421), .A(n6372), .ZN(U3184) );
  INV_X1 U7318 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6602) );
  OAI222_X1 U7319 ( .A1(n6421), .A2(n6373), .B1(n6602), .B2(n6458), .C1(n6375), 
        .C2(n6416), .ZN(U3185) );
  AOI22_X1 U7320 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6447), .ZN(n6374) );
  OAI21_X1 U7321 ( .B1(n6375), .B2(n6421), .A(n6374), .ZN(U3186) );
  AOI22_X1 U7322 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6447), .ZN(n6376) );
  OAI21_X1 U7323 ( .B1(n6377), .B2(n6421), .A(n6376), .ZN(U3187) );
  AOI22_X1 U7324 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6447), .ZN(n6378) );
  OAI21_X1 U7325 ( .B1(n6379), .B2(n6421), .A(n6378), .ZN(U3188) );
  AOI22_X1 U7326 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6447), .ZN(n6380) );
  OAI21_X1 U7327 ( .B1(n6381), .B2(n6421), .A(n6380), .ZN(U3189) );
  AOI22_X1 U7328 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6447), .ZN(n6382) );
  OAI21_X1 U7329 ( .B1(n6516), .B2(n6421), .A(n6382), .ZN(U3190) );
  AOI22_X1 U7330 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6447), .ZN(n6383) );
  OAI21_X1 U7331 ( .B1(n6599), .B2(n6421), .A(n6383), .ZN(U3191) );
  AOI22_X1 U7332 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6447), .ZN(n6384) );
  OAI21_X1 U7333 ( .B1(n6385), .B2(n6421), .A(n6384), .ZN(U3192) );
  AOI22_X1 U7334 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6447), .ZN(n6386) );
  OAI21_X1 U7335 ( .B1(n4883), .B2(n6421), .A(n6386), .ZN(U3193) );
  AOI22_X1 U7336 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6447), .ZN(n6387) );
  OAI21_X1 U7337 ( .B1(n6388), .B2(n6421), .A(n6387), .ZN(U3194) );
  AOI22_X1 U7338 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6447), .ZN(n6389) );
  OAI21_X1 U7339 ( .B1(n6390), .B2(n6421), .A(n6389), .ZN(U3195) );
  AOI22_X1 U7340 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6447), .ZN(n6391) );
  OAI21_X1 U7341 ( .B1(n6392), .B2(n6421), .A(n6391), .ZN(U3196) );
  INV_X1 U7342 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6394) );
  AOI22_X1 U7343 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6418), .ZN(n6393) );
  OAI21_X1 U7344 ( .B1(n6394), .B2(n6421), .A(n6393), .ZN(U3197) );
  AOI22_X1 U7345 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6447), .ZN(n6395) );
  OAI21_X1 U7346 ( .B1(n6397), .B2(n6416), .A(n6395), .ZN(U3198) );
  AOI22_X1 U7347 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6418), .ZN(n6396) );
  OAI21_X1 U7348 ( .B1(n6397), .B2(n6421), .A(n6396), .ZN(U3199) );
  AOI22_X1 U7349 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6447), .ZN(n6398) );
  OAI21_X1 U7350 ( .B1(n6399), .B2(n6416), .A(n6398), .ZN(U3200) );
  AOI22_X1 U7351 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6447), .ZN(n6400) );
  OAI21_X1 U7352 ( .B1(n6402), .B2(n6416), .A(n6400), .ZN(U3201) );
  AOI22_X1 U7353 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6447), .ZN(n6401) );
  OAI21_X1 U7354 ( .B1(n6402), .B2(n6421), .A(n6401), .ZN(U3202) );
  AOI22_X1 U7355 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6447), .ZN(n6403) );
  OAI21_X1 U7356 ( .B1(n6404), .B2(n6421), .A(n6403), .ZN(U3203) );
  AOI22_X1 U7357 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6418), .ZN(n6405) );
  OAI21_X1 U7358 ( .B1(n6598), .B2(n6416), .A(n6405), .ZN(U3204) );
  AOI22_X1 U7359 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6418), .ZN(n6406) );
  OAI21_X1 U7360 ( .B1(n3652), .B2(n6416), .A(n6406), .ZN(U3205) );
  AOI22_X1 U7361 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6418), .ZN(n6407) );
  OAI21_X1 U7362 ( .B1(n3652), .B2(n6421), .A(n6407), .ZN(U3206) );
  AOI22_X1 U7363 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6418), .ZN(n6408) );
  OAI21_X1 U7364 ( .B1(n4230), .B2(n6421), .A(n6408), .ZN(U3207) );
  AOI22_X1 U7365 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6418), .ZN(n6409) );
  OAI21_X1 U7366 ( .B1(n6410), .B2(n6421), .A(n6409), .ZN(U3208) );
  INV_X1 U7367 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6519) );
  AOI22_X1 U7368 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6418), .ZN(n6411) );
  OAI21_X1 U7369 ( .B1(n6519), .B2(n6421), .A(n6411), .ZN(U3209) );
  AOI22_X1 U7370 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6418), .ZN(n6412) );
  OAI21_X1 U7371 ( .B1(n6413), .B2(n6421), .A(n6412), .ZN(U3210) );
  AOI22_X1 U7372 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6414), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6418), .ZN(n6415) );
  OAI21_X1 U7373 ( .B1(n6571), .B2(n6416), .A(n6415), .ZN(U3211) );
  AOI22_X1 U7374 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6418), .ZN(n6417) );
  OAI21_X1 U7375 ( .B1(n6571), .B2(n6421), .A(n6417), .ZN(U3212) );
  AOI22_X1 U7376 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6419), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6418), .ZN(n6420) );
  OAI21_X1 U7377 ( .B1(n6422), .B2(n6421), .A(n6420), .ZN(U3213) );
  MUX2_X1 U7378 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6458), .Z(U3445) );
  MUX2_X1 U7379 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6458), .Z(U3446) );
  MUX2_X1 U7380 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6458), .Z(U3447) );
  MUX2_X1 U7381 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6458), .Z(U3448) );
  INV_X1 U7382 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6586) );
  INV_X1 U7383 ( .A(n6425), .ZN(n6423) );
  AOI21_X1 U7384 ( .B1(n6586), .B2(n6424), .A(n6423), .ZN(U3451) );
  OAI21_X1 U7385 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(U3452) );
  OAI211_X1 U7386 ( .C1(n4193), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3453)
         );
  OAI22_X1 U7387 ( .A1(n6431), .A2(n6436), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6513), .ZN(n6434) );
  OAI22_X1 U7388 ( .A1(n6434), .A2(n6433), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6432), .ZN(n6435) );
  OAI21_X1 U7389 ( .B1(n6437), .B2(n6436), .A(n6435), .ZN(U3461) );
  AOI21_X1 U7390 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6439) );
  AOI22_X1 U7391 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6439), .B2(n6438), .ZN(n6441) );
  INV_X1 U7392 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6440) );
  AOI22_X1 U7393 ( .A1(n6442), .A2(n6441), .B1(n6440), .B2(n6445), .ZN(U3468)
         );
  INV_X1 U7394 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6594) );
  NOR2_X1 U7395 ( .A1(n6445), .A2(REIP_REG_1__SCAN_IN), .ZN(n6443) );
  AOI22_X1 U7396 ( .A1(n6594), .A2(n6445), .B1(n6444), .B2(n6443), .ZN(U3469)
         );
  NAND2_X1 U7397 ( .A1(n6447), .A2(W_R_N_REG_SCAN_IN), .ZN(n6446) );
  OAI21_X1 U7398 ( .B1(n6447), .B2(READREQUEST_REG_SCAN_IN), .A(n6446), .ZN(
        U3470) );
  AOI211_X1 U7399 ( .C1(n6450), .C2(n4295), .A(n6449), .B(n6448), .ZN(n6457)
         );
  OAI211_X1 U7400 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6452), .A(n6451), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6454) );
  AOI21_X1 U7401 ( .B1(n6454), .B2(STATE2_REG_0__SCAN_IN), .A(n6453), .ZN(
        n6456) );
  NAND2_X1 U7402 ( .A1(n6457), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6455) );
  OAI21_X1 U7403 ( .B1(n6457), .B2(n6456), .A(n6455), .ZN(U3472) );
  MUX2_X1 U7404 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6458), .Z(U3473) );
  INV_X1 U7405 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6487) );
  NOR4_X1 U7406 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        INSTQUEUE_REG_8__3__SCAN_IN), .A3(n6504), .A4(n6487), .ZN(n6462) );
  NOR4_X1 U7407 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(
        INSTQUEUE_REG_7__3__SCAN_IN), .A3(n6565), .A4(n6581), .ZN(n6461) );
  NOR4_X1 U7408 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(LWORD_REG_11__SCAN_IN), 
        .A3(UWORD_REG_0__SCAN_IN), .A4(ADS_N_REG_SCAN_IN), .ZN(n6460) );
  NOR4_X1 U7409 ( .A1(EAX_REG_4__SCAN_IN), .A2(BYTEENABLE_REG_0__SCAN_IN), 
        .A3(LWORD_REG_3__SCAN_IN), .A4(LWORD_REG_13__SCAN_IN), .ZN(n6459) );
  NAND4_X1 U7410 ( .A1(n6462), .A2(n6461), .A3(n6460), .A4(n6459), .ZN(n6479)
         );
  NAND4_X1 U7411 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6478) );
  NOR4_X1 U7412 ( .A1(EBX_REG_23__SCAN_IN), .A2(EBX_REG_14__SCAN_IN), .A3(
        UWORD_REG_5__SCAN_IN), .A4(DATAO_REG_28__SCAN_IN), .ZN(n6465) );
  NOR4_X1 U7413 ( .A1(EAX_REG_19__SCAN_IN), .A2(EAX_REG_27__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6464) );
  NOR3_X1 U7414 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        REIP_REG_29__SCAN_IN), .A3(REIP_REG_26__SCAN_IN), .ZN(n6463) );
  NAND4_X1 U7415 ( .A1(n6465), .A2(n6464), .A3(ADDRESS_REG_1__SCAN_IN), .A4(
        n6463), .ZN(n6477) );
  INV_X1 U7416 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6593) );
  NOR4_X1 U7417 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        INSTQUEUE_REG_10__1__SCAN_IN), .A3(n6593), .A4(n6490), .ZN(n6475) );
  INV_X1 U7418 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6497) );
  INV_X1 U7419 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6532) );
  NOR4_X1 U7420 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6497), .A3(n6513), 
        .A4(n6532), .ZN(n6474) );
  INV_X1 U7421 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6533) );
  INV_X1 U7422 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6570) );
  NAND4_X1 U7423 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), .A3(INSTQUEUE_REG_7__4__SCAN_IN), .A4(n6570), .ZN(n6466) );
  NOR4_X1 U7424 ( .A1(n3201), .A2(n6533), .A3(n6467), .A4(n6466), .ZN(n6473)
         );
  NAND4_X1 U7425 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(EAX_REG_1__SCAN_IN), .A3(EAX_REG_6__SCAN_IN), .A4(DATAO_REG_21__SCAN_IN), .ZN(n6471) );
  NAND4_X1 U7426 ( .A1(EAX_REG_18__SCAN_IN), .A2(DATAO_REG_5__SCAN_IN), .A3(
        UWORD_REG_12__SCAN_IN), .A4(DATAO_REG_23__SCAN_IN), .ZN(n6470) );
  NAND4_X1 U7427 ( .A1(EBX_REG_3__SCAN_IN), .A2(EBX_REG_15__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .A4(DATAI_13_), .ZN(n6469) );
  NAND4_X1 U7428 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        REIP_REG_22__SCAN_IN), .A3(DATAI_25_), .A4(DATAO_REG_31__SCAN_IN), 
        .ZN(n6468) );
  NOR4_X1 U7429 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6472)
         );
  NAND4_X1 U7430 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n6476)
         );
  NOR4_X1 U7431 ( .A1(n6479), .A2(n6478), .A3(n6477), .A4(n6476), .ZN(n6620)
         );
  AOI22_X1 U7432 ( .A1(n6482), .A2(keyinput9), .B1(keyinput59), .B2(n6481), 
        .ZN(n6480) );
  OAI221_X1 U7433 ( .B1(n6482), .B2(keyinput9), .C1(n6481), .C2(keyinput59), 
        .A(n6480), .ZN(n6495) );
  AOI22_X1 U7434 ( .A1(n6485), .A2(keyinput26), .B1(keyinput52), .B2(n6484), 
        .ZN(n6483) );
  OAI221_X1 U7435 ( .B1(n6485), .B2(keyinput26), .C1(n6484), .C2(keyinput52), 
        .A(n6483), .ZN(n6494) );
  AOI22_X1 U7436 ( .A1(n6488), .A2(keyinput4), .B1(n6487), .B2(keyinput50), 
        .ZN(n6486) );
  OAI221_X1 U7437 ( .B1(n6488), .B2(keyinput4), .C1(n6487), .C2(keyinput50), 
        .A(n6486), .ZN(n6493) );
  AOI22_X1 U7438 ( .A1(n6491), .A2(keyinput22), .B1(n6490), .B2(keyinput47), 
        .ZN(n6489) );
  OAI221_X1 U7439 ( .B1(n6491), .B2(keyinput22), .C1(n6490), .C2(keyinput47), 
        .A(n6489), .ZN(n6492) );
  NOR4_X1 U7440 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6544)
         );
  AOI22_X1 U7441 ( .A1(n6498), .A2(keyinput25), .B1(n6497), .B2(keyinput39), 
        .ZN(n6496) );
  OAI221_X1 U7442 ( .B1(n6498), .B2(keyinput25), .C1(n6497), .C2(keyinput39), 
        .A(n6496), .ZN(n6511) );
  AOI22_X1 U7443 ( .A1(n6501), .A2(keyinput19), .B1(n6500), .B2(keyinput27), 
        .ZN(n6499) );
  OAI221_X1 U7444 ( .B1(n6501), .B2(keyinput19), .C1(n6500), .C2(keyinput27), 
        .A(n6499), .ZN(n6510) );
  AOI22_X1 U7445 ( .A1(n6504), .A2(keyinput63), .B1(keyinput21), .B2(n6503), 
        .ZN(n6502) );
  OAI221_X1 U7446 ( .B1(n6504), .B2(keyinput63), .C1(n6503), .C2(keyinput21), 
        .A(n6502), .ZN(n6509) );
  AOI22_X1 U7447 ( .A1(n6507), .A2(keyinput31), .B1(keyinput12), .B2(n6506), 
        .ZN(n6505) );
  OAI221_X1 U7448 ( .B1(n6507), .B2(keyinput31), .C1(n6506), .C2(keyinput12), 
        .A(n6505), .ZN(n6508) );
  NOR4_X1 U7449 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(n6543)
         );
  AOI22_X1 U7450 ( .A1(n6514), .A2(keyinput49), .B1(n6513), .B2(keyinput43), 
        .ZN(n6512) );
  OAI221_X1 U7451 ( .B1(n6514), .B2(keyinput49), .C1(n6513), .C2(keyinput43), 
        .A(n6512), .ZN(n6526) );
  AOI22_X1 U7452 ( .A1(n6517), .A2(keyinput32), .B1(keyinput60), .B2(n6516), 
        .ZN(n6515) );
  OAI221_X1 U7453 ( .B1(n6517), .B2(keyinput32), .C1(n6516), .C2(keyinput60), 
        .A(n6515), .ZN(n6525) );
  AOI22_X1 U7454 ( .A1(n6519), .A2(keyinput57), .B1(n3703), .B2(keyinput42), 
        .ZN(n6518) );
  OAI221_X1 U7455 ( .B1(n6519), .B2(keyinput57), .C1(n3703), .C2(keyinput42), 
        .A(n6518), .ZN(n6524) );
  AOI22_X1 U7456 ( .A1(n6522), .A2(keyinput17), .B1(keyinput29), .B2(n6521), 
        .ZN(n6520) );
  OAI221_X1 U7457 ( .B1(n6522), .B2(keyinput17), .C1(n6521), .C2(keyinput29), 
        .A(n6520), .ZN(n6523) );
  NOR4_X1 U7458 ( .A1(n6526), .A2(n6525), .A3(n6524), .A4(n6523), .ZN(n6542)
         );
  INV_X1 U7459 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7460 ( .A1(n6528), .A2(keyinput7), .B1(keyinput56), .B2(n4067), 
        .ZN(n6527) );
  OAI221_X1 U7461 ( .B1(n6528), .B2(keyinput7), .C1(n4067), .C2(keyinput56), 
        .A(n6527), .ZN(n6540) );
  AOI22_X1 U7462 ( .A1(n4048), .A2(keyinput40), .B1(n6530), .B2(keyinput44), 
        .ZN(n6529) );
  OAI221_X1 U7463 ( .B1(n4048), .B2(keyinput40), .C1(n6530), .C2(keyinput44), 
        .A(n6529), .ZN(n6539) );
  AOI22_X1 U7464 ( .A1(n6533), .A2(keyinput54), .B1(n6532), .B2(keyinput2), 
        .ZN(n6531) );
  OAI221_X1 U7465 ( .B1(n6533), .B2(keyinput54), .C1(n6532), .C2(keyinput2), 
        .A(n6531), .ZN(n6538) );
  NOR4_X1 U7466 ( .A1(n6540), .A2(n6539), .A3(n6538), .A4(n6537), .ZN(n6541)
         );
  NAND4_X1 U7467 ( .A1(n6544), .A2(n6543), .A3(n6542), .A4(n6541), .ZN(n6612)
         );
  AOI22_X1 U7468 ( .A1(n6547), .A2(keyinput15), .B1(keyinput33), .B2(n6546), 
        .ZN(n6545) );
  OAI221_X1 U7469 ( .B1(n6547), .B2(keyinput15), .C1(n6546), .C2(keyinput33), 
        .A(n6545), .ZN(n6560) );
  AOI22_X1 U7470 ( .A1(n6550), .A2(keyinput62), .B1(n6549), .B2(keyinput41), 
        .ZN(n6548) );
  OAI221_X1 U7471 ( .B1(n6550), .B2(keyinput62), .C1(n6549), .C2(keyinput41), 
        .A(n6548), .ZN(n6559) );
  INV_X1 U7472 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6552) );
  AOI22_X1 U7473 ( .A1(n6553), .A2(keyinput13), .B1(n6552), .B2(keyinput46), 
        .ZN(n6551) );
  OAI221_X1 U7474 ( .B1(n6553), .B2(keyinput13), .C1(n6552), .C2(keyinput46), 
        .A(n6551), .ZN(n6558) );
  INV_X1 U7475 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6556) );
  AOI22_X1 U7476 ( .A1(n6556), .A2(keyinput20), .B1(keyinput11), .B2(n6555), 
        .ZN(n6554) );
  OAI221_X1 U7477 ( .B1(n6556), .B2(keyinput20), .C1(n6555), .C2(keyinput11), 
        .A(n6554), .ZN(n6557) );
  NOR4_X1 U7478 ( .A1(n6560), .A2(n6559), .A3(n6558), .A4(n6557), .ZN(n6610)
         );
  INV_X1 U7479 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6563) );
  INV_X1 U7480 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U7481 ( .A1(n6563), .A2(keyinput30), .B1(n6562), .B2(keyinput35), 
        .ZN(n6561) );
  OAI221_X1 U7482 ( .B1(n6563), .B2(keyinput30), .C1(n6562), .C2(keyinput35), 
        .A(n6561), .ZN(n6575) );
  AOI22_X1 U7483 ( .A1(n6566), .A2(keyinput45), .B1(n6565), .B2(keyinput53), 
        .ZN(n6564) );
  OAI221_X1 U7484 ( .B1(n6566), .B2(keyinput45), .C1(n6565), .C2(keyinput53), 
        .A(n6564), .ZN(n6574) );
  INV_X1 U7485 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6568) );
  AOI22_X1 U7486 ( .A1(n5601), .A2(keyinput0), .B1(n6568), .B2(keyinput38), 
        .ZN(n6567) );
  OAI221_X1 U7487 ( .B1(n5601), .B2(keyinput0), .C1(n6568), .C2(keyinput38), 
        .A(n6567), .ZN(n6573) );
  AOI22_X1 U7488 ( .A1(n6571), .A2(keyinput55), .B1(n6570), .B2(keyinput5), 
        .ZN(n6569) );
  OAI221_X1 U7489 ( .B1(n6571), .B2(keyinput55), .C1(n6570), .C2(keyinput5), 
        .A(n6569), .ZN(n6572) );
  NOR4_X1 U7490 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(n6609)
         );
  AOI22_X1 U7491 ( .A1(n6578), .A2(keyinput34), .B1(n6577), .B2(keyinput24), 
        .ZN(n6576) );
  OAI221_X1 U7492 ( .B1(n6578), .B2(keyinput34), .C1(n6577), .C2(keyinput24), 
        .A(n6576), .ZN(n6591) );
  INV_X1 U7493 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6580) );
  AOI22_X1 U7494 ( .A1(n6581), .A2(keyinput58), .B1(n6580), .B2(keyinput51), 
        .ZN(n6579) );
  OAI221_X1 U7495 ( .B1(n6581), .B2(keyinput58), .C1(n6580), .C2(keyinput51), 
        .A(n6579), .ZN(n6590) );
  AOI22_X1 U7496 ( .A1(n6584), .A2(keyinput8), .B1(n6583), .B2(keyinput18), 
        .ZN(n6582) );
  OAI221_X1 U7497 ( .B1(n6584), .B2(keyinput8), .C1(n6583), .C2(keyinput18), 
        .A(n6582), .ZN(n6589) );
  AOI22_X1 U7498 ( .A1(n6587), .A2(keyinput37), .B1(keyinput6), .B2(n6586), 
        .ZN(n6585) );
  OAI221_X1 U7499 ( .B1(n6587), .B2(keyinput37), .C1(n6586), .C2(keyinput6), 
        .A(n6585), .ZN(n6588) );
  NOR4_X1 U7500 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6608)
         );
  AOI22_X1 U7501 ( .A1(n6594), .A2(keyinput23), .B1(n6593), .B2(keyinput10), 
        .ZN(n6592) );
  OAI221_X1 U7502 ( .B1(n6594), .B2(keyinput23), .C1(n6593), .C2(keyinput10), 
        .A(n6592), .ZN(n6606) );
  AOI22_X1 U7503 ( .A1(n3201), .A2(keyinput1), .B1(n6596), .B2(keyinput28), 
        .ZN(n6595) );
  OAI221_X1 U7504 ( .B1(n3201), .B2(keyinput1), .C1(n6596), .C2(keyinput28), 
        .A(n6595), .ZN(n6605) );
  AOI22_X1 U7505 ( .A1(n6599), .A2(keyinput36), .B1(n6598), .B2(keyinput61), 
        .ZN(n6597) );
  OAI221_X1 U7506 ( .B1(n6599), .B2(keyinput36), .C1(n6598), .C2(keyinput61), 
        .A(n6597), .ZN(n6604) );
  INV_X1 U7507 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7508 ( .A1(n6602), .A2(keyinput48), .B1(n6601), .B2(keyinput14), 
        .ZN(n6600) );
  OAI221_X1 U7509 ( .B1(n6602), .B2(keyinput48), .C1(n6601), .C2(keyinput14), 
        .A(n6600), .ZN(n6603) );
  NOR4_X1 U7510 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6607)
         );
  NAND4_X1 U7511 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n6611)
         );
  NOR2_X1 U7512 ( .A1(n6612), .A2(n6611), .ZN(n6618) );
  AOI22_X1 U7513 ( .A1(n6614), .A2(UWORD_REG_9__SCAN_IN), .B1(n6613), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U7514 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  XNOR2_X1 U7515 ( .A(n6618), .B(n6617), .ZN(n6619) );
  XNOR2_X1 U7516 ( .A(n6620), .B(n6619), .ZN(U2933) );
  AND2_X2 U34650 ( .A1(n3018), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U4209 ( .A(n3294), .B(n3298), .ZN(n3242) );
  BUF_X2 U3837 ( .A(n3702), .Z(n4447) );
  CLKBUF_X1 U3407 ( .A(n3184), .Z(n3325) );
  AND2_X2 U3438 ( .A1(n5087), .A2(n4394), .ZN(n3331) );
  CLKBUF_X1 U34560 ( .A(n3138), .Z(n3557) );
  INV_X1 U34720 ( .A(n3439), .ZN(n4219) );
  CLKBUF_X1 U3766 ( .A(n5296), .Z(n5299) );
  OR2_X1 U4042 ( .A1(n4520), .A2(n2961), .ZN(n6621) );
endmodule

