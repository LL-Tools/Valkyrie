

module b22_C_SARLock_k_64_9 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6430, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15177;

  OAI21_X1 U7179 ( .B1(n13282), .B2(n12952), .A(n11727), .ZN(n13087) );
  XNOR2_X1 U7180 ( .A(n8265), .B(n8264), .ZN(n13367) );
  AND2_X1 U7181 ( .A1(n6749), .A2(n6463), .ZN(n9019) );
  NAND2_X1 U7182 ( .A1(n10652), .A2(n10540), .ZN(n10529) );
  INV_X1 U7183 ( .A(n13535), .ZN(n13485) );
  NAND2_X2 U7184 ( .A1(n7988), .A2(n7989), .ZN(n11644) );
  CLKBUF_X1 U7185 ( .A(n7488), .Z(n7886) );
  CLKBUF_X2 U7186 ( .A(n7458), .Z(n7906) );
  CLKBUF_X2 U7187 ( .A(n7816), .Z(n7801) );
  CLKBUF_X2 U7188 ( .A(n7509), .Z(n7912) );
  CLKBUF_X2 U7189 ( .A(n7411), .Z(n6622) );
  BUF_X2 U7190 ( .A(n9953), .Z(n6435) );
  INV_X2 U7191 ( .A(n9198), .ZN(n11741) );
  OR2_X1 U7192 ( .A1(n8258), .A2(n8251), .ZN(n6957) );
  AND2_X2 U7193 ( .A1(n13365), .A2(n11773), .ZN(n9138) );
  XNOR2_X1 U7194 ( .A(n9087), .B(P2_IR_REG_22__SCAN_IN), .ZN(n11777) );
  INV_X1 U7195 ( .A(n9088), .ZN(n9089) );
  INV_X1 U7196 ( .A(n14231), .ZN(n6430) );
  INV_X2 U7197 ( .A(n6430), .ZN(P3_U3151) );
  INV_X1 U7198 ( .A(P3_STATE_REG_SCAN_IN), .ZN(n14231) );
  INV_X2 U7200 ( .A(n15177), .ZN(n6433) );
  NOR2_X1 U7201 ( .A1(n13911), .A2(n13914), .ZN(n6805) );
  AND3_X1 U7202 ( .A1(n8248), .A2(n8247), .A3(n8922), .ZN(n8928) );
  INV_X1 U7203 ( .A(n10529), .ZN(n10619) );
  NAND2_X1 U7204 ( .A1(n11757), .A2(n11756), .ZN(n13136) );
  NAND2_X1 U7206 ( .A1(n9086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U7207 ( .A1(n14375), .A2(n14371), .ZN(n14372) );
  INV_X1 U7208 ( .A(n8694), .ZN(n8641) );
  OAI21_X1 U7209 ( .B1(n14822), .B2(n7568), .A(n8000), .ZN(n11652) );
  INV_X1 U7210 ( .A(n9236), .ZN(n9198) );
  NAND2_X1 U7211 ( .A1(n7065), .A2(n7064), .ZN(n11146) );
  INV_X1 U7212 ( .A(n8691), .ZN(n8697) );
  AND2_X1 U7213 ( .A1(n8512), .A2(n8511), .ZN(n8735) );
  AND3_X1 U7214 ( .A1(n7485), .A2(n7484), .A3(n7483), .ZN(n14864) );
  NAND2_X1 U7215 ( .A1(n9290), .A2(n9289), .ZN(n11847) );
  NAND2_X1 U7216 ( .A1(n9235), .A2(n9234), .ZN(n14755) );
  XNOR2_X1 U7217 ( .A(n9089), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9573) );
  OR2_X1 U7218 ( .A1(n14006), .A2(n14125), .ZN(n13979) );
  INV_X1 U7219 ( .A(n14840), .ZN(n12254) );
  INV_X1 U7221 ( .A(n8269), .ZN(n8261) );
  AOI21_X2 U7222 ( .B1(n11231), .B2(n6469), .A(n7075), .ZN(n11579) );
  NOR2_X2 U7223 ( .A1(n9377), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n9379) );
  OAI21_X2 U7224 ( .B1(n14018), .B2(n7216), .A(n7214), .ZN(n13981) );
  OAI22_X2 U7225 ( .A1(n12546), .A2(n12438), .B1(n12553), .B2(n12558), .ZN(
        n12533) );
  XNOR2_X2 U7226 ( .A(n8225), .B(SI_24_), .ZN(n8656) );
  AND2_X4 U7227 ( .A1(n8260), .A2(n8261), .ZN(n8539) );
  NAND2_X2 U7229 ( .A1(n7621), .A2(n8012), .ZN(n14278) );
  OAI21_X2 U7230 ( .B1(n7824), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7825), .ZN(
        n7836) );
  OAI21_X2 U7231 ( .B1(n11233), .B2(n11232), .A(n11235), .ZN(n11396) );
  AOI21_X2 U7232 ( .B1(n6976), .B2(n6980), .A(n6519), .ZN(n6975) );
  AND2_X2 U7233 ( .A1(n7293), .A2(n6597), .ZN(n9481) );
  NOR2_X2 U7234 ( .A1(n9377), .A2(n9076), .ZN(n9077) );
  AND2_X2 U7235 ( .A1(n9379), .A2(n9079), .ZN(n7401) );
  OAI22_X2 U7237 ( .A1(n14271), .A2(n12414), .B1(n12668), .B2(n12413), .ZN(
        n12665) );
  NAND2_X2 U7238 ( .A1(n12412), .A2(n12411), .ZN(n14271) );
  AOI211_X2 U7239 ( .C1(n14799), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n12377), .B(
        n12376), .ZN(n12378) );
  INV_X1 U7240 ( .A(n10123), .ZN(n11278) );
  INV_X1 U7241 ( .A(n10123), .ZN(n13536) );
  NAND2_X1 U7242 ( .A1(n10424), .A2(n9737), .ZN(n6434) );
  NAND2_X2 U7243 ( .A1(n7518), .A2(n7517), .ZN(n7530) );
  OAI21_X2 U7244 ( .B1(n12665), .B2(n7340), .A(n7338), .ZN(n12598) );
  NAND2_X2 U7245 ( .A1(n7550), .A2(n7994), .ZN(n14822) );
  XNOR2_X2 U7246 ( .A(n9019), .B(n7116), .ZN(n14225) );
  XNOR2_X2 U7247 ( .A(n8219), .B(SI_22_), .ZN(n9454) );
  NOR4_X2 U7249 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  OR2_X1 U7250 ( .A1(n12479), .A2(n12485), .ZN(n8079) );
  NAND2_X1 U7251 ( .A1(n13583), .A2(n13582), .ZN(n13581) );
  NAND2_X1 U7252 ( .A1(n6783), .A2(n8289), .ZN(n14093) );
  OR2_X1 U7253 ( .A1(n7754), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7755) );
  AND2_X1 U7254 ( .A1(n14836), .A2(n11648), .ZN(n14824) );
  NAND2_X1 U7255 ( .A1(n9366), .A2(n9365), .ZN(n14332) );
  NOR2_X1 U7256 ( .A1(n14233), .A2(n14654), .ZN(n14232) );
  OAI21_X1 U7257 ( .B1(n10971), .B2(n10973), .A(n10970), .ZN(n10771) );
  NOR2_X1 U7258 ( .A1(n11163), .A2(n7028), .ZN(n7027) );
  AND2_X1 U7259 ( .A1(n7638), .A2(n7625), .ZN(n7637) );
  INV_X1 U7260 ( .A(n11644), .ZN(n11313) );
  AND4_X1 U7261 ( .A1(n7528), .A2(n7527), .A3(n7526), .A4(n7525), .ZN(n14840)
         );
  INV_X4 U7262 ( .A(n13536), .ZN(n13481) );
  NAND2_X1 U7263 ( .A1(n14891), .A2(n11298), .ZN(n7973) );
  INV_X1 U7264 ( .A(n12257), .ZN(n14918) );
  INV_X4 U7265 ( .A(n13206), .ZN(n13221) );
  INV_X1 U7266 ( .A(n11793), .ZN(n10060) );
  CLKBUF_X2 U7267 ( .A(n9191), .Z(n11959) );
  AND2_X2 U7268 ( .A1(n7422), .A2(n7420), .ZN(n7509) );
  INV_X1 U7269 ( .A(n12040), .ZN(n12031) );
  CLKBUF_X2 U7270 ( .A(n8116), .Z(n8117) );
  INV_X1 U7271 ( .A(n6646), .ZN(n10557) );
  NAND2_X1 U7272 ( .A1(n6875), .A2(n8079), .ZN(n6874) );
  MUX2_X1 U7273 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13344), .S(n14754), .Z(
        P2_U3496) );
  NAND2_X1 U7274 ( .A1(n12863), .A2(n9522), .ZN(n12929) );
  AND2_X1 U7275 ( .A1(n6675), .A2(n9678), .ZN(n12164) );
  NOR2_X1 U7276 ( .A1(n14091), .A2(n6598), .ZN(n14094) );
  NAND2_X1 U7277 ( .A1(n7877), .A2(n7876), .ZN(n12479) );
  NAND2_X1 U7278 ( .A1(n13815), .A2(n13814), .ZN(n13875) );
  NAND2_X1 U7279 ( .A1(n11976), .A2(n11975), .ZN(n13059) );
  NAND2_X1 U7280 ( .A1(n13846), .A2(n13845), .ZN(n14078) );
  NAND2_X1 U7281 ( .A1(n6600), .A2(n6599), .ZN(n6598) );
  NAND2_X1 U7282 ( .A1(n14093), .A2(n14588), .ZN(n6599) );
  AND2_X1 U7283 ( .A1(n9528), .A2(n9527), .ZN(n13092) );
  OAI21_X1 U7284 ( .B1(n13807), .B2(n6947), .A(n6447), .ZN(n13985) );
  OR2_X1 U7285 ( .A1(n14033), .A2(n13805), .ZN(n13807) );
  XNOR2_X1 U7286 ( .A(n12322), .B(n6851), .ZN(n12323) );
  NAND2_X1 U7287 ( .A1(n7732), .A2(n12602), .ZN(n12605) );
  AND2_X1 U7288 ( .A1(n13290), .A2(n13145), .ZN(n13126) );
  AOI21_X1 U7289 ( .B1(n6683), .B2(n6681), .A(n6518), .ZN(n6680) );
  NAND3_X1 U7290 ( .A1(n7171), .A2(n7787), .A3(n7169), .ZN(n7799) );
  NAND2_X1 U7291 ( .A1(n7274), .A2(n7271), .ZN(n8300) );
  NAND2_X1 U7292 ( .A1(n8658), .A2(n8657), .ZN(n14106) );
  NAND2_X1 U7293 ( .A1(n8656), .A2(n6786), .ZN(n7274) );
  NOR2_X2 U7294 ( .A1(n13222), .A2(n13321), .ZN(n13209) );
  OR2_X1 U7295 ( .A1(n12624), .A2(n12617), .ZN(n12423) );
  AND2_X1 U7296 ( .A1(n8226), .A2(n7275), .ZN(n6786) );
  OR2_X1 U7297 ( .A1(n12421), .A2(n12420), .ZN(n12617) );
  NAND2_X1 U7298 ( .A1(n7769), .A2(n7755), .ZN(n7756) );
  NAND2_X1 U7299 ( .A1(n7754), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7769) );
  AND2_X1 U7300 ( .A1(n6751), .A2(n14450), .ZN(n9026) );
  OAI21_X1 U7301 ( .B1(n14451), .B2(n14452), .A(n6752), .ZN(n6751) );
  NAND2_X1 U7302 ( .A1(n7092), .A2(n14234), .ZN(n14451) );
  NAND2_X1 U7303 ( .A1(n10916), .A2(n10851), .ZN(n10852) );
  NAND2_X1 U7304 ( .A1(n6507), .A2(n7018), .ZN(n11283) );
  OAI21_X1 U7305 ( .B1(n14235), .B2(n14236), .A(n7093), .ZN(n7092) );
  OAI21_X1 U7306 ( .B1(n11108), .B2(n7228), .A(n7226), .ZN(n11215) );
  NOR2_X1 U7307 ( .A1(n14232), .A2(n9024), .ZN(n14235) );
  XNOR2_X1 U7308 ( .A(n8211), .B(SI_20_), .ZN(n8335) );
  AOI21_X1 U7309 ( .B1(n7027), .B2(n10770), .A(n6581), .ZN(n7026) );
  OR2_X1 U7310 ( .A1(n7624), .A2(n10055), .ZN(n7625) );
  NAND2_X1 U7311 ( .A1(n8472), .A2(n8471), .ZN(n11193) );
  INV_X2 U7312 ( .A(n14927), .ZN(n14865) );
  AOI21_X1 U7313 ( .B1(n11313), .B2(n6883), .A(n6882), .ZN(n6881) );
  CLKBUF_X1 U7314 ( .A(n12911), .Z(n12943) );
  NOR2_X1 U7315 ( .A1(n10048), .A2(n10301), .ZN(n14379) );
  NAND2_X2 U7316 ( .A1(n10827), .A2(n14716), .ZN(n14714) );
  NAND2_X1 U7317 ( .A1(n9576), .A2(n9571), .ZN(n12928) );
  INV_X4 U7318 ( .A(n12045), .ZN(n9682) );
  NAND2_X1 U7319 ( .A1(n8574), .A2(n8573), .ZN(n14557) );
  INV_X2 U7320 ( .A(n14776), .ZN(n6436) );
  NAND2_X1 U7321 ( .A1(n15162), .A2(n15161), .ZN(n15160) );
  INV_X1 U7322 ( .A(n10890), .ZN(n14890) );
  NAND2_X2 U7323 ( .A1(n10037), .A2(n10346), .ZN(n13535) );
  NAND2_X1 U7324 ( .A1(n10350), .A2(n8527), .ZN(n10353) );
  XNOR2_X1 U7325 ( .A(n9006), .B(n7094), .ZN(n15162) );
  AND4_X1 U7326 ( .A1(n7474), .A2(n7473), .A3(n7472), .A4(n7471), .ZN(n10890)
         );
  NAND2_X1 U7327 ( .A1(n9166), .A2(n9165), .ZN(n11806) );
  NAND4_X1 U7328 ( .A1(n7450), .A2(n7449), .A3(n7448), .A4(n7447), .ZN(n12257)
         );
  NAND2_X2 U7329 ( .A1(n9151), .A2(n9150), .ZN(n14730) );
  CLKBUF_X1 U7330 ( .A(n10034), .Z(n10038) );
  BUF_X2 U7331 ( .A(n7671), .Z(n7911) );
  NAND2_X1 U7332 ( .A1(n8935), .A2(n8934), .ZN(n10034) );
  CLKBUF_X1 U7333 ( .A(n10321), .Z(n14548) );
  OR2_X1 U7334 ( .A1(n13627), .A2(n14532), .ZN(n10311) );
  AOI21_X1 U7335 ( .B1(n6437), .B2(n6803), .A(n7260), .ZN(n6798) );
  NAND2_X1 U7336 ( .A1(n6517), .A2(n6927), .ZN(n13627) );
  NAND4_X1 U7337 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(n13628)
         );
  NAND2_X1 U7338 ( .A1(n8889), .A2(n10602), .ZN(n10033) );
  CLKBUF_X1 U7339 ( .A(n8676), .Z(n8698) );
  XNOR2_X1 U7340 ( .A(n8933), .B(n8932), .ZN(n9793) );
  OR2_X2 U7341 ( .A1(n10323), .A2(n9908), .ZN(n14576) );
  NAND2_X1 U7342 ( .A1(n7419), .A2(n12810), .ZN(n7420) );
  NAND2_X1 U7343 ( .A1(n8142), .A2(n8141), .ZN(n8508) );
  BUF_X2 U7344 ( .A(n11777), .Z(n12040) );
  OAI21_X1 U7345 ( .B1(n8931), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8933) );
  NOR2_X1 U7346 ( .A1(n8435), .A2(n7263), .ZN(n7262) );
  INV_X1 U7348 ( .A(n9908), .ZN(n10602) );
  NAND2_X1 U7349 ( .A1(n8713), .A2(n8712), .ZN(n10738) );
  MUX2_X1 U7350 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7417), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7419) );
  NAND2_X1 U7351 ( .A1(n7418), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7416) );
  CLKBUF_X1 U7352 ( .A(n7418), .Z(n12810) );
  MUX2_X1 U7353 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8710), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8713) );
  NAND2_X4 U7354 ( .A1(n8937), .A2(n14191), .ZN(n8326) );
  INV_X1 U7355 ( .A(n8230), .ZN(n7272) );
  OR2_X1 U7356 ( .A1(n6622), .A2(n6856), .ZN(n6855) );
  INV_X2 U7357 ( .A(n13366), .ZN(n13373) );
  OR2_X1 U7358 ( .A1(n9553), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9541) );
  NOR2_X1 U7359 ( .A1(n15170), .A2(n8995), .ZN(n8999) );
  NAND2_X1 U7360 ( .A1(n6861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6860) );
  NAND2_X2 U7361 ( .A1(n9771), .A2(P2_U3088), .ZN(n13377) );
  XNOR2_X1 U7362 ( .A(n8144), .B(SI_3_), .ZN(n8507) );
  INV_X2 U7363 ( .A(n14184), .ZN(n14198) );
  NAND2_X2 U7364 ( .A1(n6781), .A2(n6778), .ZN(n8178) );
  NAND4_X1 U7365 ( .A1(n7432), .A2(n13787), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6782), .ZN(n6781) );
  NAND4_X1 U7366 ( .A1(n8130), .A2(n8520), .A3(n7207), .A4(n7206), .ZN(n8358)
         );
  AND3_X1 U7367 ( .A1(n9055), .A2(n9056), .A3(n9080), .ZN(n9075) );
  NAND4_X1 U7368 ( .A1(n6780), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n6779), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U7369 ( .A1(n8993), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8992) );
  AND3_X1 U7370 ( .A1(n9053), .A2(n9054), .A3(n9052), .ZN(n9074) );
  AND4_X2 U7371 ( .A1(n6896), .A2(n6895), .A3(n6894), .A4(n7701), .ZN(n6478)
         );
  INV_X1 U7372 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9047) );
  INV_X1 U7373 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6906) );
  INV_X1 U7374 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8102) );
  INV_X1 U7375 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8130) );
  INV_X1 U7376 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7207) );
  INV_X1 U7377 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8109) );
  INV_X4 U7378 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7379 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n9051) );
  NOR2_X1 U7380 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n9054) );
  NOR2_X1 U7381 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n9052) );
  INV_X1 U7382 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9080) );
  NOR2_X1 U7383 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8123) );
  INV_X1 U7384 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13787) );
  INV_X1 U7385 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7432) );
  INV_X4 U7386 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7387 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8421) );
  INV_X1 U7388 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9163) );
  OAI21_X1 U7389 ( .B1(n11958), .B2(n6494), .A(n6610), .ZN(n6609) );
  OAI21_X2 U7390 ( .B1(n11693), .B2(n7306), .A(n7305), .ZN(n12870) );
  OAI22_X4 U7391 ( .A1(n11658), .A2(n9376), .B1(n12936), .B2(n12932), .ZN(
        n11693) );
  NOR2_X2 U7392 ( .A1(n11236), .A2(n11867), .ZN(n11388) );
  XNOR2_X2 U7393 ( .A(n9481), .B(n9479), .ZN(n12823) );
  XNOR2_X2 U7394 ( .A(n10060), .B(n10187), .ZN(n10185) );
  AOI21_X2 U7395 ( .B1(n11770), .B2(n11974), .A(n11729), .ZN(n13260) );
  INV_X1 U7396 ( .A(n12075), .ZN(n6984) );
  NAND2_X1 U7397 ( .A1(n9610), .A2(n9609), .ZN(n9619) );
  AOI21_X1 U7398 ( .B1(n6975), .B2(n6977), .A(n6684), .ZN(n6683) );
  INV_X1 U7399 ( .A(n12158), .ZN(n6684) );
  NAND2_X1 U7400 ( .A1(n12428), .A2(n7341), .ZN(n7340) );
  INV_X1 U7401 ( .A(n7934), .ZN(n7411) );
  INV_X1 U7402 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9050) );
  INV_X1 U7403 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9049) );
  INV_X1 U7404 ( .A(n7026), .ZN(n7024) );
  NOR2_X1 U7405 ( .A1(n14428), .A2(n14406), .ZN(n6864) );
  NOR2_X1 U7406 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8247) );
  NAND2_X1 U7407 ( .A1(n6799), .A2(n6801), .ZN(n8167) );
  OR2_X1 U7408 ( .A1(n8450), .A2(n6803), .ZN(n6799) );
  NAND2_X1 U7409 ( .A1(n6960), .A2(n9618), .ZN(n6958) );
  INV_X1 U7410 ( .A(n7911), .ZN(n7891) );
  NAND2_X1 U7411 ( .A1(n6925), .A2(n6465), .ZN(n13141) );
  INV_X1 U7412 ( .A(n9148), .ZN(n9953) );
  NAND2_X2 U7413 ( .A1(n9969), .A2(n9967), .ZN(n9148) );
  XNOR2_X1 U7414 ( .A(n9010), .B(n9009), .ZN(n14219) );
  AOI21_X1 U7415 ( .B1(n8822), .B2(n6441), .A(n8821), .ZN(n7137) );
  AOI21_X1 U7416 ( .B1(n7137), .B2(n7138), .A(n7136), .ZN(n7135) );
  INV_X1 U7417 ( .A(n6521), .ZN(n7136) );
  INV_X1 U7418 ( .A(n8822), .ZN(n7138) );
  OR2_X1 U7419 ( .A1(n13059), .A2(n13057), .ZN(n11982) );
  NOR2_X1 U7420 ( .A1(n13307), .A2(n13195), .ZN(n6771) );
  NAND2_X1 U7421 ( .A1(n8735), .A2(n13625), .ZN(n8732) );
  INV_X1 U7422 ( .A(n8166), .ZN(n7263) );
  OR2_X1 U7423 ( .A1(n10433), .A2(n10448), .ZN(n6639) );
  OR2_X1 U7424 ( .A1(n14783), .A2(n6566), .ZN(n6653) );
  NOR2_X1 U7425 ( .A1(n12307), .A2(n6852), .ZN(n12329) );
  NOR2_X1 U7426 ( .A1(n6853), .A2(n7650), .ZN(n6852) );
  INV_X1 U7427 ( .A(n12308), .ZN(n6853) );
  NAND2_X1 U7428 ( .A1(n12476), .A2(n7871), .ZN(n12451) );
  OR2_X1 U7429 ( .A1(n12453), .A2(n12502), .ZN(n7871) );
  OR2_X1 U7430 ( .A1(n12782), .A2(n12574), .ZN(n8041) );
  OR2_X1 U7431 ( .A1(n12609), .A2(n12622), .ZN(n8034) );
  AOI21_X1 U7432 ( .B1(n6881), .B2(n11644), .A(n14837), .ZN(n6880) );
  NOR2_X1 U7433 ( .A1(n7407), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n6986) );
  INV_X1 U7434 ( .A(n7479), .ZN(n6985) );
  NAND2_X1 U7435 ( .A1(n7753), .A2(n7752), .ZN(n7754) );
  INV_X1 U7436 ( .A(n7179), .ZN(n7178) );
  OAI21_X1 U7437 ( .B1(n7714), .B2(n7180), .A(n7733), .ZN(n7179) );
  INV_X1 U7438 ( .A(n7185), .ZN(n7184) );
  OAI21_X1 U7439 ( .B1(n7641), .B2(n7186), .A(n7676), .ZN(n7185) );
  INV_X1 U7440 ( .A(n13365), .ZN(n9100) );
  INV_X1 U7441 ( .A(n13019), .ZN(n6718) );
  NAND2_X1 U7442 ( .A1(n13036), .A2(n13035), .ZN(n13037) );
  INV_X1 U7443 ( .A(n7072), .ZN(n7071) );
  OAI21_X1 U7444 ( .B1(n13122), .B2(n7073), .A(n11759), .ZN(n7072) );
  NOR2_X1 U7445 ( .A1(n6774), .A2(n12876), .ZN(n6773) );
  INV_X1 U7446 ( .A(n6775), .ZN(n6774) );
  NAND2_X1 U7447 ( .A1(n12004), .A2(n6470), .ZN(n6908) );
  AND2_X1 U7448 ( .A1(n13126), .A2(n13282), .ZN(n13104) );
  AND3_X2 U7449 ( .A1(n6905), .A2(n6906), .A3(n9047), .ZN(n7322) );
  AOI21_X1 U7450 ( .B1(n14068), .B2(n8884), .A(n8883), .ZN(n8901) );
  NOR2_X1 U7451 ( .A1(n13876), .A2(n7246), .ZN(n7245) );
  INV_X1 U7452 ( .A(n7249), .ZN(n7246) );
  OR2_X1 U7453 ( .A1(n13412), .A2(n11604), .ZN(n11598) );
  OR2_X1 U7454 ( .A1(n14557), .A2(n13623), .ZN(n10390) );
  OR2_X1 U7455 ( .A1(n13625), .A2(n8735), .ZN(n10375) );
  NAND2_X1 U7456 ( .A1(n8212), .A2(SI_20_), .ZN(n8213) );
  NAND2_X1 U7457 ( .A1(n8418), .A2(n7396), .ZN(n8420) );
  NAND2_X1 U7458 ( .A1(n8167), .A2(n7262), .ZN(n8438) );
  NAND2_X1 U7459 ( .A1(n7256), .A2(n7257), .ZN(n8450) );
  INV_X1 U7460 ( .A(n7258), .ZN(n7257) );
  OAI21_X1 U7461 ( .B1(n8157), .B2(n8464), .A(n8160), .ZN(n7258) );
  XNOR2_X1 U7462 ( .A(n8945), .B(n7122), .ZN(n8991) );
  INV_X1 U7463 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7122) );
  OAI21_X1 U7464 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n8961), .A(n8960), .ZN(
        n8986) );
  NAND2_X1 U7465 ( .A1(n6979), .A2(n9645), .ZN(n6978) );
  AOI21_X1 U7466 ( .B1(n12164), .B2(n12547), .A(n6973), .ZN(n6972) );
  INV_X1 U7467 ( .A(n12165), .ZN(n6973) );
  NAND2_X1 U7468 ( .A1(n6692), .A2(n6489), .ZN(n12173) );
  NOR2_X1 U7469 ( .A1(n8092), .A2(n7187), .ZN(n7957) );
  NAND2_X1 U7470 ( .A1(n8090), .A2(n6484), .ZN(n7187) );
  AND2_X1 U7471 ( .A1(n12062), .A2(n7421), .ZN(n7671) );
  NAND2_X1 U7472 ( .A1(n10577), .A2(n6812), .ZN(n6811) );
  NAND2_X1 U7473 ( .A1(n6815), .A2(n6810), .ZN(n6809) );
  AND2_X1 U7474 ( .A1(n6644), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6641) );
  XNOR2_X1 U7475 ( .A(n12329), .B(n6851), .ZN(n12311) );
  OR2_X1 U7476 ( .A1(n12311), .A2(n12310), .ZN(n6850) );
  AND2_X1 U7477 ( .A1(n7851), .A2(n7850), .ZN(n12486) );
  INV_X1 U7478 ( .A(n12451), .ZN(n12492) );
  OR2_X1 U7479 ( .A1(n7819), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7829) );
  OAI21_X1 U7480 ( .B1(n12541), .B2(n6888), .A(n6885), .ZN(n12515) );
  AOI21_X1 U7481 ( .B1(n6887), .B2(n12439), .A(n6886), .ZN(n6885) );
  INV_X1 U7482 ( .A(n8062), .ZN(n6886) );
  NOR2_X1 U7483 ( .A1(n6485), .A2(n7331), .ZN(n7330) );
  OAI21_X1 U7484 ( .B1(n12593), .B2(n6889), .A(n8041), .ZN(n12569) );
  INV_X1 U7485 ( .A(n8042), .ZN(n6889) );
  INV_X1 U7486 ( .A(n7339), .ZN(n7338) );
  OAI21_X1 U7487 ( .B1(n7340), .B2(n12422), .A(n12431), .ZN(n7339) );
  INV_X1 U7488 ( .A(n10592), .ZN(n10540) );
  AND2_X1 U7489 ( .A1(n9734), .A2(n12805), .ZN(n10660) );
  INV_X1 U7490 ( .A(n14892), .ZN(n14917) );
  NAND2_X1 U7491 ( .A1(n10424), .A2(n9737), .ZN(n7816) );
  INV_X1 U7492 ( .A(n7758), .ZN(n7923) );
  NAND2_X1 U7493 ( .A1(n7430), .A2(n7429), .ZN(n8118) );
  MUX2_X1 U7494 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7427), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7430) );
  OAI21_X1 U7495 ( .B1(n7932), .B2(n6460), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7427) );
  NAND2_X1 U7496 ( .A1(n7855), .A2(n7854), .ZN(n7857) );
  OR2_X1 U7497 ( .A1(n6858), .A2(n6856), .ZN(n6854) );
  NOR2_X1 U7498 ( .A1(n8113), .A2(n6467), .ZN(n9605) );
  OR2_X1 U7499 ( .A1(n7613), .A2(n7612), .ZN(n7199) );
  BUF_X4 U7500 ( .A(n9137), .Z(n12840) );
  AND2_X1 U7501 ( .A1(n10336), .A2(n9171), .ZN(n7282) );
  NAND2_X1 U7502 ( .A1(n9433), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11703) );
  AND2_X1 U7503 ( .A1(n13077), .A2(n13094), .ZN(n13079) );
  AOI22_X1 U7504 ( .A1(n13087), .A2(n13098), .B1(n11934), .B2(n13272), .ZN(
        n13071) );
  NAND2_X1 U7505 ( .A1(n9433), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9527) );
  AND2_X1 U7506 ( .A1(n13209), .A2(n6767), .ZN(n13145) );
  NOR2_X1 U7507 ( .A1(n6768), .A2(n13296), .ZN(n6767) );
  INV_X1 U7508 ( .A(n6769), .ZN(n6768) );
  NAND2_X1 U7509 ( .A1(n13156), .A2(n11721), .ZN(n6925) );
  AOI21_X1 U7510 ( .B1(n7082), .B2(n7081), .A(n6503), .ZN(n7080) );
  INV_X1 U7511 ( .A(n11752), .ZN(n7081) );
  AOI21_X1 U7512 ( .B1(n6456), .B2(n11713), .A(n6915), .ZN(n6914) );
  INV_X1 U7513 ( .A(n11716), .ZN(n6915) );
  NOR2_X1 U7514 ( .A1(n13247), .A2(n7087), .ZN(n7086) );
  INV_X1 U7515 ( .A(n11879), .ZN(n7087) );
  INV_X1 U7516 ( .A(n6920), .ZN(n6919) );
  NAND2_X1 U7517 ( .A1(n9435), .A2(n9434), .ZN(n13326) );
  NOR2_X1 U7518 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n9060) );
  OR2_X1 U7519 ( .A1(n13406), .A2(n13405), .ZN(n7402) );
  AND2_X1 U7520 ( .A1(n11362), .A2(n11359), .ZN(n11360) );
  INV_X1 U7521 ( .A(n11191), .ZN(n7020) );
  XNOR2_X1 U7522 ( .A(n6994), .B(n10689), .ZN(n10128) );
  OAI22_X1 U7523 ( .A1(n11278), .A2(n10125), .B1(n10124), .B2(n14532), .ZN(
        n6994) );
  OAI21_X1 U7524 ( .B1(n13822), .B2(n7212), .A(n7209), .ZN(n14034) );
  INV_X1 U7525 ( .A(n13824), .ZN(n7212) );
  AND2_X1 U7526 ( .A1(n6521), .A2(n7210), .ZN(n7209) );
  NAND2_X1 U7527 ( .A1(n7211), .A2(n13824), .ZN(n7210) );
  NAND2_X1 U7528 ( .A1(n13822), .A2(n7213), .ZN(n14049) );
  NOR2_X1 U7529 ( .A1(n6863), .A2(n14149), .ZN(n6862) );
  INV_X1 U7530 ( .A(n6864), .ZN(n6863) );
  NOR2_X1 U7531 ( .A1(n6488), .A2(n7233), .ZN(n7232) );
  NOR2_X1 U7532 ( .A1(n14575), .A2(n13621), .ZN(n7233) );
  INV_X1 U7533 ( .A(n8326), .ZN(n9815) );
  NAND2_X1 U7534 ( .A1(n9919), .A2(n10738), .ZN(n10323) );
  AND2_X1 U7535 ( .A1(n7390), .A2(n7241), .ZN(n7238) );
  NOR2_X1 U7536 ( .A1(n14211), .A2(n9000), .ZN(n9001) );
  NAND2_X1 U7537 ( .A1(n15160), .A2(n9008), .ZN(n9010) );
  INV_X1 U7538 ( .A(n6732), .ZN(n14204) );
  NAND2_X1 U7539 ( .A1(n12259), .A2(n9612), .ZN(n11294) );
  NAND2_X1 U7540 ( .A1(n9617), .A2(n9614), .ZN(n10642) );
  NAND2_X1 U7541 ( .A1(n9433), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U7542 ( .A1(n14682), .A2(n11438), .ZN(n11442) );
  AND2_X1 U7543 ( .A1(n7049), .A2(n7055), .ZN(n7048) );
  NAND2_X1 U7544 ( .A1(n14776), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7055) );
  OR2_X1 U7545 ( .A1(n7054), .A2(n14776), .ZN(n7049) );
  NAND2_X1 U7546 ( .A1(n6746), .A2(n6744), .ZN(n6749) );
  INV_X1 U7547 ( .A(n15166), .ZN(n6745) );
  INV_X1 U7548 ( .A(n9020), .ZN(n7116) );
  NAND2_X1 U7549 ( .A1(n14225), .A2(n14224), .ZN(n14223) );
  NOR2_X1 U7550 ( .A1(n11780), .A2(n12028), .ZN(n7347) );
  OR2_X1 U7551 ( .A1(n11807), .A2(n11809), .ZN(n7373) );
  NAND2_X1 U7552 ( .A1(n11856), .A2(n11858), .ZN(n7356) );
  INV_X1 U7553 ( .A(n11874), .ZN(n7354) );
  AOI21_X1 U7554 ( .B1(n7131), .B2(n7134), .A(n7130), .ZN(n7129) );
  INV_X1 U7555 ( .A(n7135), .ZN(n7134) );
  NAND2_X1 U7556 ( .A1(n8835), .A2(n8836), .ZN(n8834) );
  NAND2_X1 U7557 ( .A1(n11904), .A2(n11902), .ZN(n7371) );
  NAND2_X1 U7558 ( .A1(n7369), .A2(n11913), .ZN(n7368) );
  INV_X1 U7559 ( .A(n8201), .ZN(n7255) );
  AOI22_X1 U7560 ( .A1(n11928), .A2(n11927), .B1(n11926), .B2(n11925), .ZN(
        n11932) );
  NAND2_X1 U7561 ( .A1(n11953), .A2(n11952), .ZN(n11946) );
  INV_X1 U7562 ( .A(n11947), .ZN(n11936) );
  NOR2_X1 U7563 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  AND2_X1 U7564 ( .A1(n11999), .A2(n11998), .ZN(n7059) );
  INV_X1 U7565 ( .A(n10823), .ZN(n7062) );
  OAI21_X1 U7566 ( .B1(n10786), .B2(n13622), .A(n10390), .ZN(n6942) );
  NOR2_X1 U7567 ( .A1(n10389), .A2(n6940), .ZN(n6937) );
  NOR2_X1 U7568 ( .A1(n14561), .A2(n10776), .ZN(n6940) );
  INV_X1 U7569 ( .A(n8312), .ZN(n7275) );
  OAI21_X1 U7570 ( .B1(n8196), .B2(n6794), .A(n6792), .ZN(n8211) );
  AOI21_X1 U7571 ( .B1(n6795), .B2(n6793), .A(n6524), .ZN(n6792) );
  INV_X1 U7572 ( .A(n6795), .ZN(n6794) );
  INV_X1 U7573 ( .A(n8195), .ZN(n6793) );
  NAND2_X1 U7574 ( .A1(n8405), .A2(n7392), .ZN(n8196) );
  AND2_X1 U7575 ( .A1(n8185), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U7576 ( .A1(n7269), .A2(n8183), .ZN(n7268) );
  INV_X1 U7577 ( .A(n7396), .ZN(n7269) );
  NAND2_X1 U7578 ( .A1(n7267), .A2(n7270), .ZN(n7266) );
  INV_X1 U7579 ( .A(n8183), .ZN(n7270) );
  INV_X1 U7580 ( .A(n6802), .ZN(n6801) );
  OAI21_X1 U7581 ( .B1(n8161), .B2(n6803), .A(n8164), .ZN(n6802) );
  OAI21_X1 U7582 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(n8944), .A(n8943), .ZN(
        n8945) );
  INV_X1 U7583 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n8944) );
  INV_X1 U7584 ( .A(n10429), .ZN(n6668) );
  OR2_X1 U7585 ( .A1(n6671), .A2(n14904), .ZN(n6665) );
  NAND2_X1 U7586 ( .A1(n10453), .A2(n10452), .ZN(n10487) );
  NAND2_X1 U7587 ( .A1(n10487), .A2(n6755), .ZN(n11047) );
  OR2_X1 U7588 ( .A1(n10488), .A2(n10414), .ZN(n6755) );
  INV_X1 U7589 ( .A(n11461), .ZN(n6847) );
  INV_X1 U7590 ( .A(n6837), .ZN(n6834) );
  INV_X1 U7591 ( .A(n11539), .ZN(n6835) );
  NAND2_X1 U7592 ( .A1(n12343), .A2(n6753), .ZN(n12370) );
  AOI21_X1 U7593 ( .B1(n12366), .B2(n14210), .A(n12365), .ZN(n12386) );
  OR2_X1 U7594 ( .A1(n12465), .A2(n12473), .ZN(n8086) );
  OR2_X1 U7595 ( .A1(n12507), .A2(n12486), .ZN(n8071) );
  NAND2_X1 U7596 ( .A1(n8066), .A2(n8067), .ZN(n12446) );
  OR2_X1 U7597 ( .A1(n12714), .A2(n12558), .ZN(n8054) );
  INV_X1 U7598 ( .A(n7988), .ZN(n6882) );
  INV_X1 U7599 ( .A(n7987), .ZN(n6883) );
  INV_X1 U7600 ( .A(n10652), .ZN(n12685) );
  AND2_X1 U7601 ( .A1(n6622), .A2(n6991), .ZN(n8103) );
  AND2_X1 U7602 ( .A1(n6442), .A2(n6992), .ZN(n6991) );
  INV_X1 U7603 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n6992) );
  INV_X1 U7604 ( .A(n7716), .ZN(n7180) );
  INV_X1 U7605 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7405) );
  INV_X1 U7606 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7404) );
  INV_X1 U7607 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7403) );
  INV_X1 U7608 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7333) );
  INV_X1 U7609 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U7610 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n6896) );
  NOR2_X1 U7611 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n6895) );
  NOR2_X1 U7612 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n6894) );
  INV_X1 U7613 ( .A(n7659), .ZN(n7186) );
  AND2_X1 U7614 ( .A1(n9820), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7612) );
  INV_X1 U7615 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7408) );
  AND2_X1 U7616 ( .A1(n7194), .A2(n7546), .ZN(n7193) );
  INV_X1 U7617 ( .A(n7531), .ZN(n7191) );
  NOR2_X1 U7618 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7465) );
  INV_X1 U7619 ( .A(n7294), .ZN(n7291) );
  XNOR2_X1 U7620 ( .A(n12840), .B(n11793), .ZN(n9144) );
  INV_X1 U7621 ( .A(n12840), .ZN(n9529) );
  INV_X1 U7622 ( .A(n11773), .ZN(n9099) );
  INV_X1 U7623 ( .A(n9998), .ZN(n6713) );
  INV_X1 U7624 ( .A(n14635), .ZN(n6712) );
  AND2_X1 U7625 ( .A1(n6713), .A2(n10084), .ZN(n6706) );
  INV_X1 U7626 ( .A(n11758), .ZN(n7073) );
  INV_X1 U7627 ( .A(n11718), .ZN(n6913) );
  INV_X1 U7628 ( .A(n11634), .ZN(n6921) );
  NAND2_X1 U7629 ( .A1(n12013), .A2(n7077), .ZN(n7076) );
  INV_X1 U7630 ( .A(n11382), .ZN(n7077) );
  NOR2_X1 U7631 ( .A1(n6924), .A2(n6923), .ZN(n6922) );
  INV_X1 U7632 ( .A(n11570), .ZN(n6924) );
  INV_X1 U7633 ( .A(n7067), .ZN(n7066) );
  OAI21_X1 U7634 ( .B1(n10863), .B2(n7068), .A(n11073), .ZN(n7067) );
  INV_X1 U7635 ( .A(n10999), .ZN(n7068) );
  NOR2_X1 U7636 ( .A1(n9274), .A2(n15122), .ZN(n9273) );
  INV_X1 U7637 ( .A(n10832), .ZN(n6902) );
  OR2_X1 U7638 ( .A1(n13236), .A2(n13326), .ZN(n13222) );
  INV_X1 U7639 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U7640 ( .A1(n9540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9545) );
  OR2_X1 U7641 ( .A1(n9541), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9540) );
  INV_X1 U7642 ( .A(n10124), .ZN(n10037) );
  INV_X1 U7643 ( .A(n10738), .ZN(n8889) );
  INV_X1 U7644 ( .A(n13403), .ZN(n7034) );
  NAND2_X1 U7645 ( .A1(n7253), .A2(n7244), .ZN(n7247) );
  INV_X1 U7646 ( .A(n13966), .ZN(n13833) );
  NAND2_X1 U7647 ( .A1(n14020), .A2(n14019), .ZN(n14018) );
  NAND2_X1 U7648 ( .A1(n6945), .A2(n6946), .ZN(n6944) );
  OR2_X1 U7649 ( .A1(n14141), .A2(n13568), .ZN(n13825) );
  AND2_X1 U7650 ( .A1(n14050), .A2(n13821), .ZN(n7213) );
  INV_X1 U7651 ( .A(n11109), .ZN(n7228) );
  OR2_X1 U7652 ( .A1(n7229), .A2(n7228), .ZN(n7227) );
  AND2_X1 U7653 ( .A1(n11137), .A2(n11107), .ZN(n7229) );
  NOR2_X1 U7654 ( .A1(n11358), .A2(n6869), .ZN(n6868) );
  INV_X1 U7655 ( .A(n14573), .ZN(n6867) );
  NAND2_X1 U7656 ( .A1(n11293), .A2(n6866), .ZN(n6869) );
  INV_X1 U7657 ( .A(n11193), .ZN(n6866) );
  NAND2_X1 U7658 ( .A1(n8525), .A2(n8526), .ZN(n10350) );
  NOR2_X2 U7659 ( .A1(n14093), .A2(n13897), .ZN(n13887) );
  AND2_X1 U7660 ( .A1(n14034), .A2(n13825), .ZN(n14020) );
  INV_X1 U7661 ( .A(n10033), .ZN(n10031) );
  INV_X1 U7662 ( .A(n10967), .ZN(n10693) );
  NAND2_X1 U7663 ( .A1(n10384), .A2(n10383), .ZN(n10605) );
  AND2_X1 U7664 ( .A1(n9796), .A2(n9795), .ZN(n10024) );
  INV_X1 U7665 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U7666 ( .A1(n8420), .A2(n8183), .ZN(n8375) );
  NAND2_X1 U7667 ( .A1(n6788), .A2(n6787), .ZN(n8479) );
  AOI21_X1 U7668 ( .B1(n6790), .B2(n6791), .A(n6515), .ZN(n6787) );
  INV_X1 U7669 ( .A(n8153), .ZN(n6791) );
  NAND2_X1 U7670 ( .A1(n8146), .A2(n8145), .ZN(n8493) );
  INV_X1 U7671 ( .A(n8507), .ZN(n8143) );
  NAND2_X1 U7672 ( .A1(n8949), .A2(n8950), .ZN(n8951) );
  XNOR2_X1 U7673 ( .A(n8951), .B(n7095), .ZN(n9005) );
  INV_X1 U7674 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7095) );
  OR2_X1 U7675 ( .A1(n8955), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n8954) );
  OAI21_X1 U7676 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n13729), .A(n8965), .ZN(
        n8980) );
  AOI21_X1 U7677 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n8967), .A(n8966), .ZN(
        n9028) );
  NOR2_X1 U7678 ( .A1(n8981), .A2(n8980), .ZN(n8966) );
  OAI21_X1 U7679 ( .B1(n12216), .B2(n6963), .A(n6497), .ZN(n12063) );
  OR2_X1 U7680 ( .A1(n12215), .A2(n6963), .ZN(n6962) );
  INV_X1 U7681 ( .A(n9628), .ZN(n6963) );
  AOI21_X1 U7682 ( .B1(n6680), .B2(n6682), .A(n6678), .ZN(n6677) );
  INV_X1 U7683 ( .A(n12207), .ZN(n6678) );
  NOR2_X1 U7684 ( .A1(n10893), .A2(n6691), .ZN(n6690) );
  INV_X1 U7685 ( .A(n6961), .ZN(n6691) );
  NAND2_X1 U7686 ( .A1(n12091), .A2(n9635), .ZN(n12117) );
  AOI22_X1 U7687 ( .A1(n12150), .A2(n12149), .B1(n9625), .B2(n14873), .ZN(
        n12216) );
  NAND2_X1 U7688 ( .A1(n12216), .A2(n12215), .ZN(n12214) );
  OR2_X1 U7689 ( .A1(n12804), .A2(n9711), .ZN(n10655) );
  NAND2_X1 U7690 ( .A1(n6756), .A2(n10442), .ZN(n10509) );
  OR2_X1 U7691 ( .A1(n10441), .A2(n10502), .ZN(n6756) );
  OR2_X1 U7692 ( .A1(n8117), .A2(n10503), .ZN(n6827) );
  NAND2_X1 U7693 ( .A1(n8117), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6826) );
  AND2_X1 U7694 ( .A1(n10429), .A2(n10586), .ZN(n6671) );
  NAND2_X1 U7695 ( .A1(n6639), .A2(n10432), .ZN(n10742) );
  OR2_X1 U7696 ( .A1(n10742), .A2(n14862), .ZN(n7114) );
  NOR2_X1 U7697 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  INV_X1 U7698 ( .A(n6459), .ZN(n6814) );
  NAND2_X1 U7699 ( .A1(n6816), .A2(n6821), .ZN(n6815) );
  INV_X1 U7700 ( .A(n6817), .ZN(n6816) );
  AOI21_X1 U7701 ( .B1(n10576), .B2(n6459), .A(n6818), .ZN(n6817) );
  XNOR2_X1 U7702 ( .A(n11047), .B(n10489), .ZN(n10490) );
  NOR2_X1 U7703 ( .A1(n10489), .A2(n7112), .ZN(n6634) );
  NAND2_X1 U7704 ( .A1(n6440), .A2(n11046), .ZN(n6630) );
  NAND2_X1 U7705 ( .A1(n10434), .A2(n6635), .ZN(n6631) );
  NOR2_X1 U7706 ( .A1(n10435), .A2(n10489), .ZN(n6635) );
  NAND2_X1 U7707 ( .A1(n6633), .A2(n6639), .ZN(n7111) );
  AND2_X1 U7708 ( .A1(n10432), .A2(n6440), .ZN(n6633) );
  NAND2_X1 U7709 ( .A1(n6651), .A2(n6653), .ZN(n6657) );
  AND2_X1 U7710 ( .A1(n6654), .A2(n6452), .ZN(n6651) );
  NAND2_X1 U7711 ( .A1(n6844), .A2(n6847), .ZN(n6843) );
  INV_X1 U7712 ( .A(n14779), .ZN(n6844) );
  NAND2_X1 U7713 ( .A1(n6845), .A2(n6847), .ZN(n6842) );
  NAND2_X1 U7714 ( .A1(n6846), .A2(n11462), .ZN(n6845) );
  INV_X1 U7715 ( .A(n6848), .ZN(n6846) );
  AND3_X1 U7716 ( .A1(n7101), .A2(n11520), .A3(P3_REG2_REG_11__SCAN_IN), .ZN(
        n11521) );
  NAND2_X1 U7717 ( .A1(n7103), .A2(n11526), .ZN(n7101) );
  INV_X1 U7718 ( .A(n11478), .ZN(n7103) );
  NOR2_X1 U7719 ( .A1(n6838), .A2(n12267), .ZN(n6837) );
  INV_X1 U7720 ( .A(n12264), .ZN(n6838) );
  NAND2_X1 U7721 ( .A1(n6836), .A2(n6835), .ZN(n6832) );
  INV_X1 U7722 ( .A(n11538), .ZN(n6836) );
  INV_X1 U7723 ( .A(n6832), .ZN(n12262) );
  AND2_X1 U7724 ( .A1(n6850), .A2(n6849), .ZN(n12334) );
  NAND2_X1 U7725 ( .A1(n12331), .A2(n12332), .ZN(n6849) );
  NAND2_X1 U7726 ( .A1(n12318), .A2(n7105), .ZN(n7104) );
  NAND2_X1 U7727 ( .A1(n6658), .A2(n6454), .ZN(n6662) );
  INV_X1 U7728 ( .A(n12301), .ZN(n6658) );
  XNOR2_X1 U7729 ( .A(n12370), .B(n12359), .ZN(n12345) );
  NOR2_X1 U7730 ( .A1(n12344), .A2(n12320), .ZN(n6664) );
  NAND2_X1 U7731 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n12345), .ZN(n12372) );
  NAND2_X1 U7732 ( .A1(n12388), .A2(n7380), .ZN(n6859) );
  AND2_X1 U7733 ( .A1(n8086), .A2(n8081), .ZN(n12457) );
  AOI22_X1 U7734 ( .A1(n12462), .A2(n12461), .B1(n12460), .B2(n14892), .ZN(
        n12463) );
  NAND2_X1 U7735 ( .A1(n12493), .A2(n12492), .ZN(n12491) );
  INV_X1 U7736 ( .A(n12446), .ZN(n12514) );
  AND3_X1 U7737 ( .A1(n7833), .A2(n7832), .A3(n7831), .ZN(n12526) );
  INV_X1 U7738 ( .A(n12569), .ZN(n7767) );
  NAND2_X1 U7739 ( .A1(n12432), .A2(n12608), .ZN(n12599) );
  OR2_X1 U7740 ( .A1(n7605), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U7741 ( .A1(n14285), .A2(n14284), .ZN(n6890) );
  AND2_X1 U7742 ( .A1(n7570), .A2(n7569), .ZN(n7590) );
  AOI21_X1 U7743 ( .B1(n7327), .B2(n7329), .A(n6516), .ZN(n7326) );
  NOR2_X1 U7744 ( .A1(n7538), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7570) );
  AOI21_X1 U7745 ( .B1(n11645), .B2(n11644), .A(n11643), .ZN(n14838) );
  NAND3_X1 U7746 ( .A1(n7469), .A2(n7468), .A3(n7467), .ZN(n11298) );
  AND4_X1 U7747 ( .A1(n7426), .A2(n7425), .A3(n7424), .A4(n7423), .ZN(n14916)
         );
  INV_X1 U7748 ( .A(n14915), .ZN(n14889) );
  NAND2_X1 U7749 ( .A1(n6693), .A2(SI_1_), .ZN(n7456) );
  INV_X1 U7750 ( .A(n9740), .ZN(n6884) );
  INV_X1 U7751 ( .A(n7816), .ZN(n6693) );
  INV_X1 U7752 ( .A(n12686), .ZN(n6893) );
  INV_X1 U7753 ( .A(n12463), .ZN(n6892) );
  OR2_X1 U7754 ( .A1(n7801), .A2(n11518), .ZN(n7860) );
  AND2_X1 U7755 ( .A1(n14924), .A2(n14955), .ZN(n14305) );
  INV_X1 U7756 ( .A(n14305), .ZN(n14972) );
  NAND2_X1 U7757 ( .A1(n10521), .A2(n10619), .ZN(n14915) );
  INV_X1 U7758 ( .A(n7202), .ZN(n7201) );
  OAI22_X1 U7759 ( .A1(n7204), .A2(n7203), .B1(n11701), .B2(
        P1_DATAO_REG_28__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U7760 ( .A1(n6586), .A2(n7874), .ZN(n7203) );
  NAND2_X1 U7761 ( .A1(n7838), .A2(n7837), .ZN(n7853) );
  NAND2_X1 U7762 ( .A1(n8103), .A2(n8102), .ZN(n8108) );
  NAND2_X1 U7763 ( .A1(n7172), .A2(n7173), .ZN(n7171) );
  INV_X1 U7764 ( .A(n8103), .ZN(n8099) );
  OR2_X1 U7765 ( .A1(n7756), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7770) );
  NOR2_X1 U7766 ( .A1(n6457), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n6987) );
  AND2_X1 U7767 ( .A1(n7735), .A2(n7717), .ZN(n7733) );
  INV_X1 U7768 ( .A(n6457), .ZN(n6988) );
  NAND2_X1 U7769 ( .A1(n7698), .A2(n7697), .ZN(n7715) );
  AND2_X1 U7770 ( .A1(n7716), .A2(n7699), .ZN(n7714) );
  AND2_X1 U7771 ( .A1(n7678), .A2(n7661), .ZN(n7676) );
  AND2_X1 U7772 ( .A1(n7659), .A2(n7640), .ZN(n7641) );
  NAND2_X1 U7773 ( .A1(n7642), .A2(n7641), .ZN(n7660) );
  INV_X1 U7774 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7647) );
  INV_X1 U7775 ( .A(n7616), .ZN(n7198) );
  NAND2_X1 U7776 ( .A1(n7599), .A2(n7598), .ZN(n7613) );
  NAND2_X1 U7777 ( .A1(n7558), .A2(n7557), .ZN(n7577) );
  XNOR2_X1 U7778 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7515) );
  OR2_X1 U7779 ( .A1(n7504), .A2(n7503), .ZN(n10448) );
  XNOR2_X1 U7780 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7496) );
  NOR2_X1 U7781 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7334) );
  NAND2_X1 U7782 ( .A1(n9465), .A2(n9464), .ZN(n6597) );
  NOR2_X1 U7783 ( .A1(n7317), .A2(n12838), .ZN(n7316) );
  INV_X1 U7784 ( .A(n9522), .ZN(n7317) );
  INV_X1 U7785 ( .A(n11694), .ZN(n7307) );
  XNOR2_X1 U7786 ( .A(n12840), .B(n11806), .ZN(n10467) );
  NOR2_X1 U7787 ( .A1(n10370), .A2(n7284), .ZN(n7283) );
  INV_X1 U7788 ( .A(n9147), .ZN(n7284) );
  NAND2_X1 U7789 ( .A1(n9108), .A2(n12031), .ZN(n9477) );
  NAND2_X1 U7790 ( .A1(n9464), .A2(n7291), .ZN(n7290) );
  OR2_X1 U7791 ( .A1(n12849), .A2(n7292), .ZN(n7288) );
  INV_X1 U7792 ( .A(n9464), .ZN(n7292) );
  NAND2_X1 U7793 ( .A1(n12849), .A2(n7289), .ZN(n7285) );
  NOR2_X1 U7794 ( .A1(n9464), .A2(n7291), .ZN(n7289) );
  AND2_X1 U7795 ( .A1(n9211), .A2(n9190), .ZN(n7312) );
  NOR2_X1 U7796 ( .A1(n10826), .A2(n9569), .ZN(n9576) );
  NAND2_X1 U7797 ( .A1(n6609), .A2(n11989), .ZN(n11988) );
  AND4_X1 U7798 ( .A1(n9535), .A2(n9534), .A3(n9533), .A4(n9532), .ZN(n11934)
         );
  AND4_X1 U7799 ( .A1(n9503), .A2(n9502), .A3(n9501), .A4(n9500), .ZN(n12918)
         );
  NAND2_X1 U7800 ( .A1(n6713), .A2(n6708), .ZN(n6707) );
  INV_X1 U7801 ( .A(n6710), .ZN(n6708) );
  AOI21_X1 U7802 ( .B1(n10084), .B2(n10085), .A(n6711), .ZN(n6710) );
  INV_X1 U7803 ( .A(n9999), .ZN(n6711) );
  INV_X1 U7804 ( .A(n10163), .ZN(n6721) );
  OR2_X1 U7805 ( .A1(n6723), .A2(n6724), .ZN(n6720) );
  NAND2_X1 U7806 ( .A1(n9250), .A2(n9074), .ZN(n9377) );
  INV_X1 U7807 ( .A(n6727), .ZN(n13040) );
  AND2_X1 U7808 ( .A1(n13104), .A2(n13092), .ZN(n13094) );
  XNOR2_X1 U7809 ( .A(n13272), .B(n12951), .ZN(n13098) );
  AOI21_X1 U7810 ( .B1(n13136), .B2(n13139), .A(n7400), .ZN(n13123) );
  NAND2_X1 U7811 ( .A1(n13123), .A2(n13122), .ZN(n13125) );
  INV_X1 U7812 ( .A(n13203), .ZN(n6916) );
  OR2_X1 U7813 ( .A1(n13326), .A2(n11712), .ZN(n6917) );
  OR2_X1 U7814 ( .A1(n13218), .A2(n11713), .ZN(n6918) );
  NAND2_X1 U7815 ( .A1(n6455), .A2(n6922), .ZN(n11635) );
  NOR2_X1 U7816 ( .A1(n11380), .A2(n7079), .ZN(n7078) );
  INV_X1 U7817 ( .A(n11230), .ZN(n7079) );
  NAND2_X1 U7818 ( .A1(n11149), .A2(n11148), .ZN(n11233) );
  NOR2_X1 U7819 ( .A1(n11078), .A2(n14345), .ZN(n11150) );
  AOI21_X1 U7820 ( .B1(n6909), .B2(n10863), .A(n6496), .ZN(n6907) );
  NAND2_X1 U7821 ( .A1(n10852), .A2(n10863), .ZN(n11000) );
  OAI21_X1 U7822 ( .B1(n11990), .B2(n10296), .A(n10061), .ZN(n10186) );
  NAND2_X1 U7823 ( .A1(n11990), .A2(n10276), .ZN(n10059) );
  INV_X1 U7824 ( .A(n11784), .ZN(n10931) );
  NAND2_X1 U7825 ( .A1(n11969), .A2(n11777), .ZN(n7303) );
  XNOR2_X1 U7826 ( .A(n11736), .B(n12019), .ZN(n7057) );
  NAND2_X1 U7827 ( .A1(n11779), .A2(n12031), .ZN(n14761) );
  NAND2_X1 U7828 ( .A1(n9933), .A2(n12030), .ZN(n14753) );
  INV_X1 U7829 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13357) );
  NOR2_X1 U7830 ( .A1(n9162), .A2(n7345), .ZN(n9248) );
  AND2_X1 U7831 ( .A1(n9792), .A2(n9803), .ZN(n8935) );
  INV_X1 U7832 ( .A(n10769), .ZN(n7028) );
  INV_X1 U7833 ( .A(n7402), .ZN(n7036) );
  AND2_X1 U7834 ( .A1(n7041), .A2(n7040), .ZN(n13515) );
  NAND2_X1 U7835 ( .A1(n10686), .A2(n10687), .ZN(n7040) );
  AND2_X1 U7836 ( .A1(n13575), .A2(n6999), .ZN(n6998) );
  OR2_X1 U7837 ( .A1(n13507), .A2(n7000), .ZN(n6999) );
  INV_X1 U7838 ( .A(n13474), .ZN(n7000) );
  AOI21_X1 U7839 ( .B1(n13513), .B2(n10695), .A(n10696), .ZN(n10971) );
  NAND2_X1 U7840 ( .A1(n14372), .A2(n13403), .ZN(n14398) );
  OR2_X1 U7841 ( .A1(n8909), .A2(n8915), .ZN(n7385) );
  NAND2_X1 U7842 ( .A1(n8881), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U7843 ( .A1(n8255), .A2(n8254), .ZN(n13790) );
  INV_X1 U7844 ( .A(n14071), .ZN(n13789) );
  INV_X1 U7845 ( .A(n14085), .ZN(n13869) );
  OAI21_X1 U7846 ( .B1(n13875), .B2(n13816), .A(n13818), .ZN(n13859) );
  AOI21_X1 U7847 ( .B1(n7245), .B2(n7243), .A(n7248), .ZN(n7242) );
  NAND2_X1 U7848 ( .A1(n7245), .A2(n6805), .ZN(n6804) );
  AND2_X1 U7849 ( .A1(n14093), .A2(n13840), .ZN(n7248) );
  XNOR2_X1 U7850 ( .A(n14093), .B(n13840), .ZN(n13876) );
  OR2_X1 U7851 ( .A1(n13911), .A2(n13914), .ZN(n7253) );
  NAND2_X1 U7852 ( .A1(n13788), .A2(n13908), .ZN(n13909) );
  NAND2_X1 U7853 ( .A1(n13833), .A2(n13832), .ZN(n13964) );
  INV_X1 U7854 ( .A(n7215), .ZN(n7214) );
  OAI21_X1 U7855 ( .B1(n7217), .B2(n7216), .A(n13982), .ZN(n7215) );
  INV_X1 U7856 ( .A(n13829), .ZN(n7216) );
  NAND2_X1 U7857 ( .A1(n13999), .A2(n13829), .ZN(n13983) );
  OR2_X1 U7858 ( .A1(n14134), .A2(n14001), .ZN(n6949) );
  NAND2_X1 U7859 ( .A1(n6948), .A2(n6946), .ZN(n14012) );
  NAND2_X1 U7860 ( .A1(n14018), .A2(n7217), .ZN(n13999) );
  NAND2_X1 U7861 ( .A1(n11600), .A2(n11599), .ZN(n13822) );
  AND2_X1 U7862 ( .A1(n11598), .A2(n8805), .ZN(n11625) );
  NAND2_X1 U7863 ( .A1(n11420), .A2(n11419), .ZN(n11608) );
  NAND2_X1 U7864 ( .A1(n11595), .A2(n11596), .ZN(n11419) );
  NAND2_X1 U7865 ( .A1(n10807), .A2(n10806), .ZN(n11108) );
  NAND2_X1 U7866 ( .A1(n11108), .A2(n7229), .ZN(n11136) );
  AOI21_X1 U7867 ( .B1(n6931), .B2(n6933), .A(n6501), .ZN(n6929) );
  OAI21_X1 U7868 ( .B1(n7236), .B2(n10389), .A(n6471), .ZN(n7230) );
  NAND2_X1 U7869 ( .A1(n10376), .A2(n10375), .ZN(n10603) );
  INV_X1 U7870 ( .A(n13949), .ZN(n14252) );
  NAND2_X1 U7871 ( .A1(n10311), .A2(n10313), .ZN(n10308) );
  AND2_X1 U7872 ( .A1(n14199), .A2(n8326), .ZN(n14120) );
  OR2_X1 U7873 ( .A1(n8694), .A2(n9752), .ZN(n6926) );
  OR2_X1 U7874 ( .A1(n10323), .A2(n10030), .ZN(n14592) );
  INV_X1 U7875 ( .A(n14578), .ZN(n14597) );
  NAND2_X1 U7876 ( .A1(n8241), .A2(n8240), .ZN(n8684) );
  XNOR2_X1 U7877 ( .A(n8684), .B(n8683), .ZN(n13363) );
  XNOR2_X1 U7878 ( .A(n8288), .B(n8287), .ZN(n11775) );
  INV_X1 U7879 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6780) );
  INV_X1 U7880 ( .A(n8178), .ZN(n8324) );
  AOI22_X1 U7881 ( .A1(n8711), .A2(n7127), .B1(n7125), .B2(n7124), .ZN(n7123)
         );
  AND2_X1 U7882 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7127) );
  XNOR2_X1 U7883 ( .A(n8714), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9908) );
  XNOR2_X1 U7884 ( .A(n8640), .B(n8639), .ZN(n10595) );
  NAND2_X1 U7885 ( .A1(n8438), .A2(n8172), .ZN(n8587) );
  INV_X2 U7886 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U7887 ( .A1(n9123), .A2(n8550), .ZN(n8531) );
  INV_X1 U7888 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n8993) );
  XNOR2_X1 U7889 ( .A(n9005), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U7890 ( .A1(n15157), .A2(n9004), .ZN(n9006) );
  AOI21_X1 U7891 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n13712), .A(n8962), .ZN(
        n8984) );
  NOR2_X1 U7892 ( .A1(n8987), .A2(n8986), .ZN(n8962) );
  NAND2_X1 U7893 ( .A1(n14456), .A2(n14454), .ZN(n9029) );
  OR2_X1 U7894 ( .A1(n11328), .A2(n8115), .ZN(n9734) );
  NOR2_X1 U7895 ( .A1(n12237), .A2(n9691), .ZN(n6970) );
  AND2_X1 U7896 ( .A1(n9691), .A2(n12229), .ZN(n6969) );
  NAND2_X1 U7897 ( .A1(n12164), .A2(n6673), .ZN(n12083) );
  NAND2_X1 U7898 ( .A1(n12191), .A2(n6674), .ZN(n6673) );
  NAND2_X1 U7899 ( .A1(n7773), .A2(n7772), .ZN(n12562) );
  OR2_X1 U7900 ( .A1(n7801), .A2(n10590), .ZN(n7772) );
  AOI21_X1 U7901 ( .B1(n9616), .B2(n9615), .A(n10642), .ZN(n10640) );
  AND4_X1 U7902 ( .A1(n7713), .A2(n7712), .A3(n7711), .A4(n7710), .ZN(n12637)
         );
  NAND2_X1 U7903 ( .A1(n7724), .A2(n7723), .ZN(n12609) );
  AND2_X1 U7904 ( .A1(n9727), .A2(n9726), .ZN(n12242) );
  OAI211_X1 U7905 ( .C1(n8098), .C2(n10518), .A(n7168), .B(n7167), .ZN(n7166)
         );
  INV_X1 U7906 ( .A(n12486), .ZN(n12512) );
  OAI211_X1 U7907 ( .C1(n7891), .C2(n12705), .A(n7822), .B(n7821), .ZN(n12536)
         );
  NAND2_X1 U7908 ( .A1(n7488), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7448) );
  OAI22_X1 U7909 ( .A1(n10717), .A2(n10501), .B1(n6825), .B2(n10502), .ZN(
        n10544) );
  NAND2_X1 U7910 ( .A1(n6827), .A2(n6826), .ZN(n6825) );
  NAND2_X1 U7911 ( .A1(n6643), .A2(n6574), .ZN(n6642) );
  INV_X1 U7912 ( .A(n12260), .ZN(n6643) );
  NAND2_X1 U7913 ( .A1(n12260), .A2(n14216), .ZN(n6640) );
  NAND2_X1 U7914 ( .A1(n6662), .A2(n7104), .ZN(n12340) );
  INV_X1 U7915 ( .A(n12393), .ZN(n14801) );
  INV_X1 U7916 ( .A(n14810), .ZN(n14781) );
  OAI21_X1 U7917 ( .B1(n12490), .B2(n14877), .A(n12489), .ZN(n12693) );
  NOR2_X1 U7918 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  NAND2_X1 U7919 ( .A1(n12541), .A2(n12540), .ZN(n12707) );
  NAND2_X1 U7920 ( .A1(n7803), .A2(n7802), .ZN(n12709) );
  OR2_X1 U7921 ( .A1(n7801), .A2(n10886), .ZN(n7802) );
  INV_X1 U7922 ( .A(n12453), .ZN(n12762) );
  NOR2_X1 U7923 ( .A1(n9538), .A2(n7319), .ZN(n7318) );
  INV_X1 U7924 ( .A(n9526), .ZN(n7319) );
  NAND2_X1 U7925 ( .A1(n9433), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U7926 ( .A1(n10291), .A2(n9147), .ZN(n10371) );
  INV_X1 U7927 ( .A(n9492), .ZN(n6595) );
  OR2_X1 U7928 ( .A1(n9374), .A2(n9375), .ZN(n9373) );
  NAND2_X1 U7929 ( .A1(n9382), .A2(n9381), .ZN(n14321) );
  NAND2_X1 U7930 ( .A1(n9397), .A2(n9396), .ZN(n12876) );
  NAND2_X1 U7931 ( .A1(n9264), .A2(n11015), .ZN(n11022) );
  NAND2_X1 U7932 ( .A1(n9331), .A2(n9330), .ZN(n14339) );
  INV_X1 U7933 ( .A(n12929), .ZN(n6592) );
  INV_X1 U7934 ( .A(n11934), .ZN(n12951) );
  NAND2_X1 U7935 ( .A1(n11442), .A2(n6694), .ZN(n11584) );
  NOR2_X1 U7936 ( .A1(n6580), .A2(n6695), .ZN(n6694) );
  NOR2_X1 U7937 ( .A1(n11444), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6695) );
  AND2_X1 U7938 ( .A1(n9981), .A2(n12039), .ZN(n14696) );
  CLKBUF_X1 U7939 ( .A(n9573), .Z(n12027) );
  AND2_X1 U7940 ( .A1(n9511), .A2(n9510), .ZN(n13282) );
  NAND2_X1 U7941 ( .A1(n9433), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9510) );
  OR3_X1 U7942 ( .A1(n13127), .A2(n13126), .A3(n13221), .ZN(n13289) );
  NAND2_X1 U7943 ( .A1(n9433), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U7944 ( .A1(n7057), .A2(n7051), .ZN(n7050) );
  NOR2_X1 U7945 ( .A1(n14776), .A2(n7052), .ZN(n7051) );
  AND2_X1 U7946 ( .A1(n13263), .A2(n6450), .ZN(n7054) );
  NAND2_X1 U7947 ( .A1(n7057), .A2(n14753), .ZN(n7056) );
  NOR2_X1 U7948 ( .A1(n9162), .A2(n7365), .ZN(n7364) );
  NAND2_X1 U7949 ( .A1(n9070), .A2(n9098), .ZN(n7365) );
  NAND2_X1 U7950 ( .A1(n8621), .A2(n8620), .ZN(n14428) );
  NAND2_X1 U7951 ( .A1(n8670), .A2(n8669), .ZN(n14112) );
  NOR2_X1 U7952 ( .A1(n10129), .A2(n10130), .ZN(n10146) );
  NAND2_X1 U7953 ( .A1(n7002), .A2(n7001), .ZN(n14375) );
  AOI21_X1 U7954 ( .B1(n7003), .B2(n7006), .A(n6502), .ZN(n7001) );
  AND4_X1 U7955 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n10712)
         );
  NAND2_X1 U7956 ( .A1(n8398), .A2(n8397), .ZN(n14146) );
  INV_X1 U7957 ( .A(n13627), .ZN(n10125) );
  NOR2_X1 U7958 ( .A1(n6466), .A2(n8515), .ZN(n8516) );
  NOR2_X1 U7959 ( .A1(n8513), .A2(n7391), .ZN(n8517) );
  NAND2_X1 U7960 ( .A1(n8315), .A2(n8314), .ZN(n13924) );
  NAND2_X1 U7961 ( .A1(n8411), .A2(n8410), .ZN(n14149) );
  INV_X1 U7962 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14179) );
  AND2_X1 U7963 ( .A1(n7390), .A2(n7240), .ZN(n7239) );
  AND2_X1 U7964 ( .A1(n7241), .A2(n8259), .ZN(n7240) );
  INV_X1 U7965 ( .A(n9002), .ZN(n6750) );
  NAND2_X1 U7966 ( .A1(n6748), .A2(n6747), .ZN(n6746) );
  NAND2_X1 U7967 ( .A1(n6737), .A2(n6735), .ZN(n14233) );
  AOI22_X1 U7968 ( .A1(n14225), .A2(n6448), .B1(n9022), .B2(n6736), .ZN(n6735)
         );
  NAND2_X1 U7969 ( .A1(n14457), .A2(n14458), .ZN(n14454) );
  INV_X1 U7970 ( .A(n14455), .ZN(n14456) );
  XNOR2_X1 U7971 ( .A(n9029), .B(n7096), .ZN(n14461) );
  INV_X1 U7972 ( .A(n9030), .ZN(n7096) );
  NAND2_X1 U7973 ( .A1(n14461), .A2(n14460), .ZN(n14459) );
  NAND2_X1 U7974 ( .A1(n6734), .A2(n6733), .ZN(n6732) );
  NAND2_X1 U7975 ( .A1(n9036), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6733) );
  OAI21_X1 U7976 ( .B1(n14204), .B2(n14205), .A(n14706), .ZN(n7110) );
  NAND2_X1 U7977 ( .A1(n14204), .A2(n14205), .ZN(n14203) );
  NOR2_X1 U7978 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  OAI211_X1 U7979 ( .C1(n11796), .C2(n11794), .A(n11792), .B(n11791), .ZN(
        n7349) );
  INV_X1 U7980 ( .A(n11794), .ZN(n7351) );
  OR2_X1 U7981 ( .A1(n7375), .A2(n11808), .ZN(n7374) );
  INV_X1 U7982 ( .A(n11807), .ZN(n7375) );
  INV_X1 U7983 ( .A(n11820), .ZN(n7360) );
  INV_X1 U7984 ( .A(n11831), .ZN(n7358) );
  AND3_X1 U7985 ( .A1(n8742), .A2(n8741), .A3(n8740), .ZN(n8752) );
  INV_X1 U7986 ( .A(n11844), .ZN(n7362) );
  OR2_X1 U7987 ( .A1(n7160), .A2(n8762), .ZN(n7159) );
  INV_X1 U7988 ( .A(n8761), .ZN(n7160) );
  NAND2_X1 U7989 ( .A1(n8773), .A2(n7151), .ZN(n7150) );
  NAND2_X1 U7990 ( .A1(n8783), .A2(n8785), .ZN(n7143) );
  AOI21_X1 U7991 ( .B1(n7353), .B2(n11874), .A(n6923), .ZN(n7352) );
  INV_X1 U7992 ( .A(n11875), .ZN(n7353) );
  INV_X1 U7993 ( .A(n8794), .ZN(n7144) );
  NOR2_X1 U7994 ( .A1(n8797), .A2(n8794), .ZN(n7145) );
  AOI21_X1 U7995 ( .B1(n7135), .B2(n7133), .A(n7132), .ZN(n7131) );
  INV_X1 U7996 ( .A(n8824), .ZN(n7132) );
  INV_X1 U7997 ( .A(n7137), .ZN(n7133) );
  OAI22_X1 U7998 ( .A1(n8830), .A2(n7140), .B1(n8831), .B2(n7139), .ZN(n8835)
         );
  NOR2_X1 U7999 ( .A1(n8832), .A2(n8829), .ZN(n7140) );
  INV_X1 U8000 ( .A(n8829), .ZN(n7139) );
  NAND2_X1 U8001 ( .A1(n7157), .A2(n8841), .ZN(n7156) );
  NAND2_X1 U8002 ( .A1(n8859), .A2(n7154), .ZN(n7153) );
  NAND2_X1 U8003 ( .A1(n12950), .A2(n11967), .ZN(n7280) );
  NAND2_X1 U8004 ( .A1(n13266), .A2(n11985), .ZN(n7281) );
  NAND2_X1 U8005 ( .A1(n7279), .A2(n7277), .ZN(n11952) );
  NAND2_X1 U8006 ( .A1(n11933), .A2(n7278), .ZN(n7277) );
  NAND2_X1 U8007 ( .A1(n13077), .A2(n11967), .ZN(n7279) );
  INV_X1 U8008 ( .A(n11967), .ZN(n7278) );
  CLKBUF_X1 U8009 ( .A(n8726), .Z(n8764) );
  NOR2_X1 U8010 ( .A1(n8203), .A2(n6796), .ZN(n6795) );
  INV_X1 U8011 ( .A(n8394), .ZN(n6796) );
  NAND2_X1 U8012 ( .A1(n8204), .A2(n7255), .ZN(n7254) );
  OR2_X1 U8013 ( .A1(n10562), .A2(n10431), .ZN(n10433) );
  AND2_X1 U8014 ( .A1(n7938), .A2(n12476), .ZN(n8077) );
  NAND2_X1 U8015 ( .A1(n7344), .A2(n7414), .ZN(n7343) );
  INV_X1 U8016 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7414) );
  INV_X1 U8017 ( .A(n7413), .ZN(n7344) );
  NAND2_X1 U8018 ( .A1(n7163), .A2(n8869), .ZN(n7162) );
  NOR2_X1 U8019 ( .A1(n6446), .A2(n7252), .ZN(n7244) );
  INV_X1 U8020 ( .A(n6950), .ZN(n6945) );
  NOR2_X1 U8021 ( .A1(n8312), .A2(n8655), .ZN(n7273) );
  NAND2_X1 U8022 ( .A1(n8198), .A2(n8197), .ZN(n8201) );
  NAND2_X1 U8023 ( .A1(n8192), .A2(n8191), .ZN(n8195) );
  AOI21_X1 U8024 ( .B1(n8567), .B2(n8153), .A(n8555), .ZN(n6790) );
  NAND2_X1 U8025 ( .A1(n7121), .A2(n8946), .ZN(n8947) );
  NAND2_X1 U8026 ( .A1(n8991), .A2(n13659), .ZN(n7121) );
  INV_X1 U8027 ( .A(SI_13_), .ZN(n8179) );
  NOR2_X1 U8028 ( .A1(n7956), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U8029 ( .A1(n12477), .A2(n7955), .ZN(n7189) );
  NAND2_X1 U8030 ( .A1(n14298), .A2(n7954), .ZN(n8089) );
  NOR2_X1 U8031 ( .A1(n12754), .A2(n12251), .ZN(n8092) );
  NAND2_X1 U8032 ( .A1(n10743), .A2(n10450), .ZN(n10453) );
  NAND2_X1 U8033 ( .A1(n7111), .A2(n7112), .ZN(n6637) );
  NAND2_X1 U8034 ( .A1(n6556), .A2(n11474), .ZN(n6655) );
  NAND2_X1 U8035 ( .A1(n14786), .A2(n6754), .ZN(n11467) );
  OR2_X1 U8036 ( .A1(n14789), .A2(n14986), .ZN(n6754) );
  NAND2_X1 U8037 ( .A1(n12266), .A2(n6765), .ZN(n12281) );
  OR2_X1 U8038 ( .A1(n12267), .A2(n11528), .ZN(n6765) );
  AND2_X1 U8039 ( .A1(n6612), .A2(n6611), .ZN(n12322) );
  NAND2_X1 U8040 ( .A1(n12309), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8041 ( .A1(n12303), .A2(n12302), .ZN(n6612) );
  INV_X1 U8042 ( .A(n12321), .ZN(n7105) );
  OR2_X1 U8043 ( .A1(n12387), .A2(n14230), .ZN(n7380) );
  AOI21_X1 U8044 ( .B1(n12492), .B2(n6878), .A(n6877), .ZN(n6876) );
  INV_X1 U8045 ( .A(n8072), .ZN(n6878) );
  INV_X1 U8046 ( .A(n8077), .ZN(n6877) );
  INV_X1 U8047 ( .A(n12435), .ZN(n7331) );
  INV_X1 U8048 ( .A(n7328), .ZN(n7327) );
  OAI21_X1 U8049 ( .B1(n11649), .B2(n7329), .A(n11669), .ZN(n7328) );
  INV_X1 U8050 ( .A(n11650), .ZN(n7329) );
  AND2_X1 U8051 ( .A1(n8002), .A2(n8000), .ZN(n14821) );
  NAND2_X1 U8052 ( .A1(n11307), .A2(n11306), .ZN(n14852) );
  INV_X1 U8053 ( .A(SI_16_), .ZN(n8191) );
  NAND2_X1 U8054 ( .A1(n9611), .A2(n14899), .ZN(n14869) );
  OR2_X1 U8055 ( .A1(n9694), .A2(n9707), .ZN(n10524) );
  NAND2_X1 U8056 ( .A1(n9604), .A2(n6964), .ZN(n6965) );
  AND2_X1 U8057 ( .A1(n9605), .A2(n6966), .ZN(n6964) );
  NAND2_X1 U8058 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), 
        .ZN(n6856) );
  NOR2_X1 U8059 ( .A1(n7343), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U8060 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  OR2_X1 U8061 ( .A1(n7814), .A2(n11559), .ZN(n7825) );
  AOI21_X1 U8062 ( .B1(n7769), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n7785), .ZN(
        n7173) );
  NAND2_X1 U8063 ( .A1(n7197), .A2(n7195), .ZN(n7624) );
  AOI21_X1 U8064 ( .B1(n6555), .B2(n7612), .A(n7196), .ZN(n7195) );
  INV_X1 U8065 ( .A(n7622), .ZN(n7196) );
  OR2_X1 U8066 ( .A1(n7626), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7644) );
  INV_X1 U8067 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n15124) );
  CLKBUF_X1 U8068 ( .A(n7479), .Z(n7480) );
  NAND2_X1 U8069 ( .A1(n9451), .A2(n7295), .ZN(n7294) );
  INV_X1 U8070 ( .A(n9452), .ZN(n7295) );
  AND2_X1 U8071 ( .A1(n9292), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9311) );
  AND2_X1 U8072 ( .A1(n9273), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9292) );
  INV_X1 U8073 ( .A(n11978), .ZN(n6610) );
  OR2_X1 U8074 ( .A1(n13039), .A2(n14693), .ZN(n6727) );
  NOR2_X1 U8075 ( .A1(n13159), .A2(n6770), .ZN(n6769) );
  INV_X1 U8076 ( .A(n6771), .ZN(n6770) );
  NAND2_X1 U8077 ( .A1(n11751), .A2(n11752), .ZN(n7084) );
  OAI21_X1 U8078 ( .B1(n6922), .B2(n6921), .A(n11705), .ZN(n6920) );
  NOR2_X1 U8079 ( .A1(n14332), .A2(n14321), .ZN(n6775) );
  NAND2_X1 U8080 ( .A1(n9311), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9350) );
  AOI21_X1 U8081 ( .B1(n11999), .B2(n7062), .A(n6500), .ZN(n7061) );
  INV_X1 U8082 ( .A(n11777), .ZN(n7304) );
  INV_X1 U8083 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9554) );
  NOR2_X1 U8084 ( .A1(n9078), .A2(n9247), .ZN(n6594) );
  INV_X1 U8085 ( .A(n9086), .ZN(n6605) );
  AND2_X1 U8086 ( .A1(n9048), .A2(n9058), .ZN(n7321) );
  INV_X1 U8087 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6905) );
  AND2_X1 U8088 ( .A1(n7010), .A2(n13601), .ZN(n7009) );
  NAND2_X1 U8089 ( .A1(n7011), .A2(n7017), .ZN(n7010) );
  INV_X1 U8090 ( .A(n7012), .ZN(n7011) );
  INV_X1 U8091 ( .A(n7244), .ZN(n7243) );
  NAND2_X1 U8092 ( .A1(n7250), .A2(n13839), .ZN(n7249) );
  OAI21_X1 U8093 ( .B1(n13960), .B2(n6953), .A(n6952), .ZN(n13915) );
  NAND2_X1 U8094 ( .A1(n13811), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8095 ( .A1(n6955), .A2(n13811), .ZN(n6952) );
  INV_X1 U8096 ( .A(n13961), .ZN(n6954) );
  NAND2_X1 U8097 ( .A1(n13915), .A2(n13914), .ZN(n13913) );
  NAND2_X1 U8098 ( .A1(n13929), .A2(n6956), .ZN(n6955) );
  INV_X1 U8099 ( .A(n7399), .ZN(n6956) );
  OR2_X1 U8100 ( .A1(n7223), .A2(n13836), .ZN(n7221) );
  AND2_X1 U8101 ( .A1(n13961), .A2(n6530), .ZN(n7223) );
  NAND2_X1 U8102 ( .A1(n7225), .A2(n13834), .ZN(n7222) );
  NOR2_X1 U8103 ( .A1(n13947), .A2(n14106), .ZN(n13908) );
  NOR2_X1 U8104 ( .A1(n13979), .A2(n14120), .ZN(n6872) );
  NOR2_X1 U8105 ( .A1(n14019), .A2(n6951), .ZN(n6950) );
  INV_X1 U8106 ( .A(n13806), .ZN(n6951) );
  NOR2_X1 U8107 ( .A1(n14013), .A2(n7218), .ZN(n7217) );
  INV_X1 U8108 ( .A(n13827), .ZN(n7218) );
  INV_X1 U8109 ( .A(n7213), .ZN(n7211) );
  AND2_X1 U8110 ( .A1(n7379), .A2(n11100), .ZN(n6936) );
  INV_X1 U8111 ( .A(n6932), .ZN(n6931) );
  OAI21_X1 U8112 ( .B1(n10810), .B2(n6933), .A(n11098), .ZN(n6932) );
  INV_X1 U8113 ( .A(n10812), .ZN(n6933) );
  NAND2_X1 U8114 ( .A1(n6939), .A2(n6938), .ZN(n14566) );
  OR2_X1 U8115 ( .A1(n6941), .A2(n6940), .ZN(n6938) );
  INV_X1 U8116 ( .A(n6942), .ZN(n6941) );
  NAND2_X1 U8117 ( .A1(n13887), .A2(n13869), .ZN(n13868) );
  NOR2_X1 U8118 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8127) );
  NOR2_X1 U8119 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n8128) );
  NOR2_X1 U8120 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8126) );
  NAND2_X1 U8121 ( .A1(n6785), .A2(n6784), .ZN(n8226) );
  AOI21_X1 U8122 ( .B1(n8224), .B2(n10886), .A(n11269), .ZN(n6784) );
  INV_X1 U8123 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6782) );
  INV_X1 U8124 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8125 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n8251), .ZN(n7124) );
  NAND2_X1 U8126 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7126), .ZN(n7125) );
  NAND2_X1 U8127 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n7126) );
  NAND2_X1 U8128 ( .A1(n8709), .A2(n8707), .ZN(n7045) );
  INV_X1 U8129 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U8130 ( .A1(n8202), .A2(n8201), .ZN(n8634) );
  NAND2_X1 U8131 ( .A1(n8395), .A2(n8394), .ZN(n8202) );
  NAND2_X1 U8132 ( .A1(n8196), .A2(n8195), .ZN(n8395) );
  AND2_X1 U8133 ( .A1(n7266), .A2(n8190), .ZN(n7265) );
  OR2_X1 U8134 ( .A1(n8439), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8588) );
  OAI21_X1 U8135 ( .B1(n8178), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n8133), .ZN(
        n8135) );
  OAI22_X1 U8136 ( .A1(n7117), .A2(n8992), .B1(P1_ADDR_REG_1__SCAN_IN), .B2(
        n7118), .ZN(n8997) );
  AND2_X1 U8137 ( .A1(n7118), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7117) );
  INV_X1 U8138 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7118) );
  XNOR2_X1 U8139 ( .A(n8947), .B(n7120), .ZN(n8988) );
  INV_X1 U8140 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8141 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  INV_X1 U8142 ( .A(n11684), .ZN(n6983) );
  NAND2_X1 U8143 ( .A1(n11545), .A2(n6989), .ZN(n12091) );
  NOR2_X1 U8144 ( .A1(n12094), .A2(n6990), .ZN(n6989) );
  INV_X1 U8145 ( .A(n9633), .ZN(n6990) );
  AND3_X1 U8146 ( .A1(n7587), .A2(n7586), .A3(n7585), .ZN(n11671) );
  NAND2_X1 U8147 ( .A1(n9620), .A2(n11299), .ZN(n6961) );
  AND3_X1 U8148 ( .A1(n7440), .A2(n7439), .A3(n7438), .ZN(n11302) );
  NAND2_X1 U8149 ( .A1(n12063), .A2(n9629), .ZN(n11342) );
  NOR2_X1 U8150 ( .A1(n7708), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7726) );
  OR2_X1 U8151 ( .A1(n7686), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7708) );
  AND2_X1 U8152 ( .A1(n12129), .A2(n9681), .ZN(n12165) );
  OR2_X1 U8153 ( .A1(n11547), .A2(n11548), .ZN(n11545) );
  AND2_X1 U8154 ( .A1(n12259), .A2(n10668), .ZN(n7962) );
  INV_X1 U8155 ( .A(n6683), .ZN(n6682) );
  INV_X1 U8156 ( .A(n6975), .ZN(n6681) );
  NAND2_X1 U8157 ( .A1(n6981), .A2(n6979), .ZN(n12236) );
  NAND2_X1 U8158 ( .A1(n7669), .A2(n7668), .ZN(n7686) );
  NAND2_X1 U8159 ( .A1(n6614), .A2(n6613), .ZN(n10551) );
  OR2_X1 U8160 ( .A1(n10557), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U8161 ( .A1(n10557), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U8162 ( .A1(n10550), .A2(n10551), .ZN(n10549) );
  INV_X1 U8163 ( .A(n7119), .ZN(n10564) );
  OAI211_X1 U8164 ( .C1(n6669), .C2(n10545), .A(n6665), .B(n6667), .ZN(n7119)
         );
  NAND2_X1 U8165 ( .A1(n6668), .A2(n10444), .ZN(n6667) );
  NAND2_X1 U8166 ( .A1(n7111), .A2(n7113), .ZN(n10477) );
  INV_X1 U8167 ( .A(n6809), .ZN(n6806) );
  NAND2_X1 U8168 ( .A1(n11048), .A2(n11049), .ZN(n14787) );
  NAND2_X1 U8169 ( .A1(n14787), .A2(n14788), .ZN(n14786) );
  XNOR2_X1 U8170 ( .A(n11467), .B(n11057), .ZN(n11050) );
  AND2_X1 U8171 ( .A1(n11041), .A2(n14789), .ZN(n6848) );
  NOR2_X1 U8172 ( .A1(n14780), .A2(n14779), .ZN(n14778) );
  AND2_X1 U8173 ( .A1(n6657), .A2(n6656), .ZN(n14814) );
  AOI21_X1 U8174 ( .B1(n6843), .B2(n6842), .A(n6840), .ZN(n6839) );
  INV_X1 U8175 ( .A(n14803), .ZN(n6840) );
  NAND2_X1 U8176 ( .A1(n11525), .A2(n6473), .ZN(n11530) );
  NAND2_X1 U8177 ( .A1(n11530), .A2(n11529), .ZN(n12266) );
  NOR2_X1 U8178 ( .A1(n11523), .A2(n14295), .ZN(n7100) );
  XNOR2_X1 U8179 ( .A(n12281), .B(n12278), .ZN(n12268) );
  NAND2_X1 U8180 ( .A1(n6828), .A2(n6830), .ZN(n12290) );
  INV_X1 U8181 ( .A(n6831), .ZN(n6830) );
  OAI21_X1 U8182 ( .B1(n6833), .B2(n6835), .A(n6563), .ZN(n6831) );
  NAND2_X1 U8183 ( .A1(n6664), .A2(n14210), .ZN(n6663) );
  INV_X1 U8184 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U8185 ( .A1(n12369), .A2(n12368), .ZN(n12388) );
  OR2_X1 U8186 ( .A1(n7878), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12407) );
  NOR2_X1 U8187 ( .A1(n12477), .A2(n7337), .ZN(n7336) );
  INV_X1 U8188 ( .A(n12454), .ZN(n7337) );
  OR2_X1 U8189 ( .A1(n7829), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7845) );
  INV_X1 U8190 ( .A(n7806), .ZN(n7805) );
  NAND2_X1 U8191 ( .A1(n7775), .A2(n7774), .ZN(n7791) );
  INV_X1 U8192 ( .A(n7776), .ZN(n7775) );
  OR2_X1 U8193 ( .A1(n7791), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7806) );
  AND2_X1 U8194 ( .A1(n8054), .A2(n8055), .ZN(n12549) );
  NAND2_X1 U8195 ( .A1(n12573), .A2(n12568), .ZN(n7332) );
  AND2_X1 U8196 ( .A1(n8041), .A2(n8042), .ZN(n12584) );
  NAND2_X1 U8197 ( .A1(n12599), .A2(n12433), .ZN(n12585) );
  NAND2_X1 U8198 ( .A1(n12599), .A2(n7342), .ZN(n12587) );
  AND2_X1 U8199 ( .A1(n12592), .A2(n12433), .ZN(n7342) );
  AND2_X1 U8200 ( .A1(n7726), .A2(n7725), .ZN(n7746) );
  NOR2_X1 U8201 ( .A1(n7382), .A2(n7692), .ZN(n7693) );
  AND4_X1 U8202 ( .A1(n7658), .A2(n7657), .A3(n7656), .A4(n7655), .ZN(n12652)
         );
  AND2_X1 U8203 ( .A1(n12655), .A2(n8020), .ZN(n12664) );
  NOR2_X1 U8204 ( .A1(n7654), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7669) );
  OR2_X1 U8205 ( .A1(n7631), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7654) );
  AND4_X1 U8206 ( .A1(n7610), .A2(n7609), .A3(n7608), .A4(n7607), .ZN(n14289)
         );
  AND4_X1 U8207 ( .A1(n7575), .A2(n7574), .A3(n7573), .A4(n7572), .ZN(n14290)
         );
  NAND2_X1 U8208 ( .A1(n14824), .A2(n11649), .ZN(n14823) );
  NAND2_X1 U8209 ( .A1(n11399), .A2(n7987), .ZN(n11314) );
  AND4_X1 U8210 ( .A1(n7543), .A2(n7542), .A3(n7541), .A4(n7540), .ZN(n11647)
         );
  NAND2_X1 U8211 ( .A1(n14852), .A2(n7335), .ZN(n11402) );
  AND2_X1 U8212 ( .A1(n11310), .A2(n11309), .ZN(n7335) );
  AND2_X1 U8213 ( .A1(n7987), .A2(n7985), .ZN(n11401) );
  NOR2_X1 U8214 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7490) );
  INV_X1 U8215 ( .A(n14920), .ZN(n14877) );
  AND2_X1 U8216 ( .A1(n14869), .A2(n7976), .ZN(n14893) );
  AND2_X1 U8217 ( .A1(n10539), .A2(n10538), .ZN(n14924) );
  NAND2_X1 U8218 ( .A1(n7973), .A2(n14885), .ZN(n14914) );
  CLKBUF_X1 U8219 ( .A(n11295), .Z(n7941) );
  NAND2_X1 U8220 ( .A1(n10519), .A2(n10518), .ZN(n14920) );
  CLKBUF_X1 U8221 ( .A(n7940), .Z(n10638) );
  NAND2_X1 U8222 ( .A1(n7905), .A2(n7904), .ZN(n7925) );
  NAND2_X1 U8223 ( .A1(n7828), .A2(n7827), .ZN(n12699) );
  OR2_X1 U8224 ( .A1(n7801), .A2(n11327), .ZN(n7827) );
  NAND2_X1 U8225 ( .A1(n7818), .A2(n7817), .ZN(n12443) );
  OR2_X1 U8226 ( .A1(n7801), .A2(n11269), .ZN(n7817) );
  AND2_X1 U8227 ( .A1(n7653), .A2(n7652), .ZN(n12415) );
  NAND2_X1 U8228 ( .A1(n7899), .A2(n7898), .ZN(n7919) );
  OR2_X1 U8229 ( .A1(n7897), .A2(n7896), .ZN(n7899) );
  OR2_X1 U8230 ( .A1(n7919), .A2(n7918), .ZN(n7921) );
  NOR2_X1 U8231 ( .A1(n7205), .A2(n7872), .ZN(n7204) );
  INV_X1 U8232 ( .A(n7856), .ZN(n7205) );
  XNOR2_X1 U8233 ( .A(n8100), .B(n8102), .ZN(n10422) );
  NAND2_X1 U8234 ( .A1(n8099), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8100) );
  XNOR2_X1 U8235 ( .A(n7936), .B(P3_IR_REG_20__SCAN_IN), .ZN(n10618) );
  CLKBUF_X1 U8236 ( .A(n7934), .Z(n7935) );
  AOI21_X1 U8237 ( .B1(n7178), .B2(n7180), .A(n7176), .ZN(n7175) );
  INV_X1 U8238 ( .A(n7735), .ZN(n7176) );
  AND2_X1 U8239 ( .A1(n7752), .A2(n7736), .ZN(n7737) );
  AND2_X1 U8240 ( .A1(n7697), .A2(n7679), .ZN(n7695) );
  AOI21_X1 U8241 ( .B1(n7184), .B2(n7186), .A(n7183), .ZN(n7182) );
  INV_X1 U8242 ( .A(n7678), .ZN(n7183) );
  NAND2_X1 U8243 ( .A1(n7579), .A2(n7578), .ZN(n7597) );
  AOI21_X1 U8244 ( .B1(n7193), .B2(n7191), .A(n6520), .ZN(n7190) );
  INV_X1 U8245 ( .A(n7193), .ZN(n7192) );
  XNOR2_X1 U8246 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7555) );
  AND2_X1 U8247 ( .A1(n9786), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7529) );
  XNOR2_X1 U8248 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7546) );
  OR2_X1 U8249 ( .A1(n7533), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7544) );
  XNOR2_X1 U8250 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7475) );
  OR2_X1 U8251 ( .A1(n7466), .A2(n6647), .ZN(n6646) );
  NAND2_X1 U8252 ( .A1(n6650), .A2(n6648), .ZN(n6647) );
  NAND2_X1 U8253 ( .A1(n8112), .A2(n6649), .ZN(n6648) );
  AND2_X1 U8254 ( .A1(n12916), .A2(n9521), .ZN(n9522) );
  NOR2_X1 U8255 ( .A1(n11560), .A2(n7311), .ZN(n7310) );
  INV_X1 U8256 ( .A(n9327), .ZN(n7311) );
  NAND2_X1 U8257 ( .A1(n7299), .A2(n12879), .ZN(n6596) );
  NOR2_X1 U8258 ( .A1(n7300), .A2(n7298), .ZN(n7297) );
  INV_X1 U8259 ( .A(n9478), .ZN(n7298) );
  NAND2_X1 U8260 ( .A1(n9932), .A2(n11992), .ZN(n12028) );
  OR2_X1 U8261 ( .A1(n11741), .A2(n9962), .ZN(n9169) );
  AND3_X1 U8262 ( .A1(n9113), .A2(n9114), .A3(n9115), .ZN(n7046) );
  OR2_X1 U8263 ( .A1(n11731), .A2(n10292), .ZN(n9117) );
  NAND2_X1 U8264 ( .A1(n6704), .A2(n6712), .ZN(n6702) );
  NAND2_X1 U8265 ( .A1(n14620), .A2(n6706), .ZN(n6705) );
  OR2_X1 U8266 ( .A1(n10170), .A2(n10169), .ZN(n10213) );
  AOI21_X1 U8267 ( .B1(n6716), .B2(n6720), .A(n6715), .ZN(n6714) );
  INV_X1 U8268 ( .A(n13020), .ZN(n6715) );
  NAND2_X1 U8269 ( .A1(n6727), .A2(n6726), .ZN(n14692) );
  NAND2_X1 U8270 ( .A1(n13039), .A2(n14693), .ZN(n6726) );
  NOR2_X1 U8271 ( .A1(n14692), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14691) );
  NAND2_X1 U8272 ( .A1(n11961), .A2(n11960), .ZN(n13055) );
  NAND2_X1 U8273 ( .A1(n9433), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11960) );
  NOR2_X1 U8274 ( .A1(n13055), .A2(n13062), .ZN(n13063) );
  NOR2_X1 U8275 ( .A1(n9134), .A2(n11772), .ZN(n11729) );
  OAI21_X1 U8276 ( .B1(n11934), .B2(n13092), .A(n13274), .ZN(n13076) );
  AOI21_X1 U8277 ( .B1(n7071), .B2(n7073), .A(n6495), .ZN(n7069) );
  INV_X1 U8278 ( .A(n13290), .ZN(n13131) );
  NAND2_X1 U8279 ( .A1(n13209), .A2(n6769), .ZN(n13157) );
  OR2_X1 U8280 ( .A1(n13172), .A2(n13173), .ZN(n13174) );
  OAI21_X1 U8281 ( .B1(n6914), .B2(n6913), .A(n6510), .ZN(n6912) );
  NAND2_X1 U8282 ( .A1(n13209), .A2(n13314), .ZN(n13189) );
  NAND2_X1 U8283 ( .A1(n11750), .A2(n11749), .ZN(n13201) );
  AND2_X1 U8284 ( .A1(n6480), .A2(n11748), .ZN(n7085) );
  AND2_X1 U8285 ( .A1(n13243), .A2(n6773), .ZN(n6772) );
  NAND2_X1 U8286 ( .A1(n11388), .A2(n6775), .ZN(n11636) );
  NAND2_X1 U8287 ( .A1(n11388), .A2(n11387), .ZN(n11572) );
  NAND2_X1 U8288 ( .A1(n7076), .A2(n6482), .ZN(n7075) );
  AOI21_X1 U8289 ( .B1(n7066), .B2(n7068), .A(n6490), .ZN(n7064) );
  NAND2_X1 U8290 ( .A1(n11069), .A2(n11068), .ZN(n11149) );
  NAND2_X1 U8291 ( .A1(n10921), .A2(n14765), .ZN(n11007) );
  OR2_X1 U8292 ( .A1(n11007), .A2(n11847), .ZN(n11078) );
  OR2_X1 U8293 ( .A1(n9257), .A2(n9090), .ZN(n9274) );
  NOR2_X1 U8294 ( .A1(n11029), .A2(n14755), .ZN(n10920) );
  AND2_X1 U8295 ( .A1(n10920), .A2(n10925), .ZN(n10921) );
  INV_X1 U8296 ( .A(n6901), .ZN(n6900) );
  AOI21_X1 U8297 ( .B1(n6901), .B2(n11998), .A(n6514), .ZN(n6899) );
  NOR2_X1 U8298 ( .A1(n10833), .A2(n6902), .ZN(n6901) );
  OR2_X1 U8299 ( .A1(n11028), .A2(n14746), .ZN(n11029) );
  NAND2_X1 U8300 ( .A1(n10246), .A2(n10941), .ZN(n11028) );
  AND2_X1 U8301 ( .A1(n10906), .A2(n10950), .ZN(n10246) );
  NOR2_X1 U8302 ( .A1(n10957), .A2(n11806), .ZN(n10906) );
  OR2_X1 U8303 ( .A1(n10959), .A2(n14730), .ZN(n10957) );
  XNOR2_X1 U8304 ( .A(n13260), .B(n12949), .ZN(n12019) );
  OR3_X1 U8305 ( .A1(n13094), .A2(n13093), .A3(n13221), .ZN(n13275) );
  OR3_X1 U8306 ( .A1(n13104), .A2(n13103), .A3(n13221), .ZN(n13281) );
  NAND2_X1 U8307 ( .A1(n9433), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U8308 ( .A1(n9096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9071) );
  XNOR2_X1 U8309 ( .A(n9547), .B(P2_IR_REG_26__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U8310 ( .A1(n6606), .A2(n6603), .ZN(n9107) );
  NOR2_X1 U8311 ( .A1(n6605), .A2(n6604), .ZN(n6603) );
  NAND2_X1 U8312 ( .A1(n9083), .A2(n6594), .ZN(n6606) );
  NOR2_X1 U8313 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6604) );
  AND2_X1 U8314 ( .A1(n9080), .A2(n9081), .ZN(n6617) );
  INV_X1 U8315 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9079) );
  CLKBUF_X1 U8316 ( .A(n9250), .Z(n9287) );
  AND2_X1 U8317 ( .A1(n9233), .A2(n9232), .ZN(n10166) );
  OR2_X1 U8318 ( .A1(n9213), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U8319 ( .A1(n6906), .A2(n6905), .ZN(n6904) );
  INV_X1 U8320 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8485) );
  AOI21_X1 U8321 ( .B1(n7023), .B2(n7022), .A(n6523), .ZN(n7021) );
  INV_X1 U8322 ( .A(n7027), .ZN(n7022) );
  INV_X1 U8323 ( .A(n11180), .ZN(n7029) );
  NAND2_X1 U8324 ( .A1(n7019), .A2(n7023), .ZN(n7018) );
  NAND2_X1 U8325 ( .A1(n13581), .A2(n7030), .ZN(n13549) );
  AND2_X1 U8326 ( .A1(n13456), .A2(n13454), .ZN(n7030) );
  NAND2_X1 U8327 ( .A1(n7016), .A2(n6458), .ZN(n7015) );
  INV_X1 U8328 ( .A(n14384), .ZN(n7016) );
  NAND2_X1 U8329 ( .A1(n11284), .A2(n11285), .ZN(n11361) );
  NOR2_X1 U8330 ( .A1(n13536), .A2(n10669), .ZN(n10039) );
  AND2_X1 U8331 ( .A1(n10036), .A2(n10035), .ZN(n10121) );
  NAND2_X1 U8332 ( .A1(n10037), .A2(n10307), .ZN(n10035) );
  NOR2_X1 U8333 ( .A1(n10038), .A2(n8543), .ZN(n10032) );
  NOR2_X1 U8334 ( .A1(n8594), .A2(n8428), .ZN(n8622) );
  NOR2_X1 U8335 ( .A1(n8608), .A2(n9882), .ZN(n8607) );
  AND2_X1 U8336 ( .A1(n11496), .A2(n7004), .ZN(n7003) );
  NAND2_X1 U8337 ( .A1(n11360), .A2(n7005), .ZN(n7004) );
  INV_X1 U8338 ( .A(n11285), .ZN(n7005) );
  INV_X1 U8339 ( .A(n11360), .ZN(n7006) );
  INV_X1 U8340 ( .A(n10148), .ZN(n7037) );
  NOR2_X1 U8341 ( .A1(n13567), .A2(n7013), .ZN(n7012) );
  INV_X1 U8342 ( .A(n7015), .ZN(n7013) );
  INV_X1 U8343 ( .A(n7033), .ZN(n7031) );
  AOI21_X1 U8344 ( .B1(n7035), .B2(n7034), .A(n6493), .ZN(n7033) );
  AND2_X1 U8345 ( .A1(n10038), .A2(n8936), .ZN(n10707) );
  INV_X1 U8346 ( .A(n8542), .ZN(n8687) );
  AND2_X1 U8347 ( .A1(n8625), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8513) );
  INV_X1 U8348 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n13712) );
  OR2_X1 U8349 ( .A1(n8406), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U8350 ( .A1(n8696), .A2(n8695), .ZN(n13844) );
  OR2_X1 U8351 ( .A1(n13909), .A2(n14098), .ZN(n13897) );
  OR2_X1 U8352 ( .A1(n13959), .A2(n6955), .ZN(n13927) );
  NOR2_X1 U8353 ( .A1(n13959), .A2(n7399), .ZN(n13928) );
  INV_X1 U8354 ( .A(n13908), .ZN(n13942) );
  NOR2_X1 U8355 ( .A1(n13960), .A2(n13961), .ZN(n13959) );
  NAND2_X1 U8356 ( .A1(n6872), .A2(n6871), .ZN(n13947) );
  INV_X1 U8357 ( .A(n14112), .ZN(n6871) );
  INV_X1 U8358 ( .A(n6872), .ZN(n13967) );
  NAND2_X1 U8359 ( .A1(n13807), .A2(n6950), .ZN(n6948) );
  NAND2_X1 U8360 ( .A1(n14005), .A2(n14011), .ZN(n14006) );
  OR2_X1 U8361 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  NAND2_X1 U8362 ( .A1(n10321), .A2(n13782), .ZN(n10346) );
  NOR2_X1 U8363 ( .A1(n8415), .A2(n8399), .ZN(n8400) );
  NOR2_X1 U8364 ( .A1(n14054), .A2(n14146), .ZN(n14057) );
  INV_X1 U8365 ( .A(n13823), .ZN(n14050) );
  AOI21_X1 U8366 ( .B1(n6602), .B2(n11595), .A(n6601), .ZN(n11626) );
  INV_X1 U8367 ( .A(n11596), .ZN(n6601) );
  INV_X1 U8368 ( .A(n11597), .ZN(n6602) );
  AND2_X1 U8369 ( .A1(n8622), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U8370 ( .A1(n8624), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U8371 ( .A1(n14245), .A2(n14434), .ZN(n14244) );
  INV_X1 U8372 ( .A(n11418), .ZN(n14249) );
  AND2_X1 U8373 ( .A1(n7227), .A2(n11212), .ZN(n7226) );
  NAND2_X1 U8374 ( .A1(n6935), .A2(n6934), .ZN(n11417) );
  AND2_X1 U8375 ( .A1(n11217), .A2(n6483), .ZN(n6934) );
  NAND2_X1 U8376 ( .A1(n6867), .A2(n6444), .ZN(n11211) );
  NAND2_X1 U8377 ( .A1(n6867), .A2(n6868), .ZN(n11134) );
  OR2_X1 U8378 ( .A1(n8562), .A2(n8485), .ZN(n8487) );
  NAND2_X1 U8379 ( .A1(n6930), .A2(n10812), .ZN(n11099) );
  NAND2_X1 U8380 ( .A1(n10811), .A2(n10810), .ZN(n6930) );
  NOR2_X1 U8381 ( .A1(n14573), .A2(n11193), .ZN(n10816) );
  OR2_X1 U8382 ( .A1(n7231), .A2(n10728), .ZN(n7236) );
  INV_X1 U8383 ( .A(n10380), .ZN(n7231) );
  NAND2_X1 U8384 ( .A1(n10793), .A2(n10389), .ZN(n7237) );
  AND2_X1 U8385 ( .A1(n8498), .A2(n8497), .ZN(n10967) );
  AND2_X1 U8386 ( .A1(n10671), .A2(n10355), .ZN(n10348) );
  OR2_X1 U8387 ( .A1(n13628), .A2(n10669), .ZN(n10312) );
  NOR2_X1 U8388 ( .A1(n14576), .A2(n13782), .ZN(n10305) );
  INV_X1 U8389 ( .A(n14092), .ZN(n6600) );
  NAND2_X1 U8390 ( .A1(n8337), .A2(n8336), .ZN(n14130) );
  AOI222_X1 U8391 ( .A1(n14554), .A2(n14023), .B1(n14022), .B2(n14254), .C1(
        n14021), .C2(n14252), .ZN(n14137) );
  NAND2_X1 U8392 ( .A1(n13807), .A2(n13806), .ZN(n14028) );
  NAND2_X1 U8393 ( .A1(n8456), .A2(n8455), .ZN(n14587) );
  INV_X1 U8394 ( .A(n10024), .ZN(n9912) );
  NOR2_X1 U8395 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7241) );
  XNOR2_X1 U8396 ( .A(n8693), .B(n8692), .ZN(n11770) );
  NAND2_X1 U8397 ( .A1(n8931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8927) );
  OR2_X1 U8398 ( .A1(n8708), .A2(n7045), .ZN(n8711) );
  NOR2_X1 U8399 ( .A1(n8708), .A2(n7042), .ZN(n8921) );
  NAND2_X1 U8400 ( .A1(n7044), .A2(n7043), .ZN(n7042) );
  INV_X1 U8401 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7043) );
  INV_X1 U8402 ( .A(n7045), .ZN(n7044) );
  INV_X1 U8403 ( .A(n8250), .ZN(n8708) );
  XNOR2_X1 U8404 ( .A(n8381), .B(n8380), .ZN(n10259) );
  NAND2_X1 U8405 ( .A1(n8167), .A2(n8166), .ZN(n8436) );
  NAND2_X1 U8406 ( .A1(n6800), .A2(n8163), .ZN(n8601) );
  NAND2_X1 U8407 ( .A1(n8450), .A2(n8161), .ZN(n6800) );
  NOR2_X1 U8408 ( .A1(n8468), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8602) );
  OR2_X1 U8409 ( .A1(n8480), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8466) );
  OR2_X1 U8410 ( .A1(n8466), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U8411 ( .A1(n7259), .A2(n8157), .ZN(n8465) );
  AND2_X1 U8412 ( .A1(n8569), .A2(n8359), .ZN(n8571) );
  NOR2_X1 U8413 ( .A1(n8358), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U8414 ( .A1(n8178), .A2(n6506), .ZN(n8550) );
  XNOR2_X1 U8415 ( .A(n6461), .B(n8992), .ZN(n8994) );
  NAND2_X1 U8416 ( .A1(n8953), .A2(n8952), .ZN(n9011) );
  INV_X1 U8417 ( .A(n9022), .ZN(n6738) );
  INV_X1 U8418 ( .A(n9021), .ZN(n6736) );
  AOI21_X1 U8419 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n8964), .A(n8963), .ZN(
        n8983) );
  OR2_X1 U8420 ( .A1(n14466), .A2(n7090), .ZN(n7089) );
  INV_X1 U8421 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7091) );
  NAND2_X1 U8422 ( .A1(n12214), .A2(n9628), .ZN(n12065) );
  NAND2_X1 U8423 ( .A1(n6981), .A2(n6464), .ZN(n12074) );
  INV_X1 U8424 ( .A(n12083), .ZN(n6974) );
  NAND2_X1 U8425 ( .A1(n11545), .A2(n9633), .ZN(n12093) );
  NAND2_X1 U8426 ( .A1(n6686), .A2(n6476), .ZN(n12057) );
  AND3_X1 U8427 ( .A1(n7507), .A2(n7506), .A3(n7505), .ZN(n14859) );
  OR2_X1 U8428 ( .A1(n7816), .A2(SI_4_), .ZN(n7485) );
  AND2_X1 U8429 ( .A1(n6692), .A2(n6449), .ZN(n12174) );
  AND3_X1 U8430 ( .A1(n7566), .A2(n7565), .A3(n7564), .ZN(n14830) );
  NAND2_X1 U8431 ( .A1(n7790), .A2(n7789), .ZN(n12714) );
  AND3_X1 U8432 ( .A1(n7604), .A2(n7603), .A3(n7602), .ZN(n12201) );
  INV_X1 U8433 ( .A(n12244), .ZN(n12220) );
  INV_X1 U8434 ( .A(n12245), .ZN(n12219) );
  AND2_X1 U8435 ( .A1(n7870), .A2(n7869), .ZN(n12502) );
  AND4_X1 U8436 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n12651)
         );
  AND2_X1 U8437 ( .A1(n7917), .A2(n7893), .ZN(n12473) );
  NAND4_X1 U8438 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n12575)
         );
  INV_X1 U8439 ( .A(n12637), .ZN(n12429) );
  INV_X1 U8440 ( .A(n12651), .ZN(n12416) );
  INV_X1 U8441 ( .A(n12652), .ZN(n14273) );
  NAND4_X1 U8442 ( .A1(n7636), .A2(n7635), .A3(n7634), .A4(n7633), .ZN(n12668)
         );
  INV_X1 U8443 ( .A(n14289), .ZN(n14272) );
  NAND4_X1 U8444 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .ZN(n12252)
         );
  INV_X1 U8445 ( .A(n14290), .ZN(n14825) );
  INV_X1 U8446 ( .A(n14916), .ZN(n9611) );
  OAI211_X1 U8447 ( .C1(n6824), .C2(n6826), .A(n6823), .B(n6822), .ZN(n10501)
         );
  NAND2_X1 U8448 ( .A1(n6670), .A2(n6672), .ZN(n10578) );
  INV_X1 U8449 ( .A(n7114), .ZN(n10741) );
  NAND2_X1 U8450 ( .A1(n6815), .A2(n6811), .ZN(n10749) );
  NAND2_X1 U8451 ( .A1(n6819), .A2(n10418), .ZN(n10485) );
  OAI21_X1 U8452 ( .B1(n6809), .B2(n10577), .A(n6807), .ZN(n6819) );
  AOI21_X1 U8453 ( .B1(n6815), .B2(n6808), .A(n10750), .ZN(n6807) );
  NOR2_X1 U8454 ( .A1(n6812), .A2(n10751), .ZN(n6808) );
  NAND2_X1 U8455 ( .A1(n6632), .A2(n6627), .ZN(n10478) );
  AND2_X1 U8456 ( .A1(n6631), .A2(n6628), .ZN(n6627) );
  NOR2_X1 U8457 ( .A1(n14778), .A2(n6848), .ZN(n11463) );
  NAND2_X1 U8458 ( .A1(n7101), .A2(n11520), .ZN(n11479) );
  INV_X1 U8459 ( .A(n11521), .ZN(n7099) );
  NAND2_X1 U8460 ( .A1(n6568), .A2(n14216), .ZN(n6644) );
  NAND2_X1 U8461 ( .A1(n6832), .A2(n6829), .ZN(n12288) );
  AND2_X1 U8462 ( .A1(n6645), .A2(n6474), .ZN(n12280) );
  NAND2_X1 U8463 ( .A1(n7106), .A2(n12317), .ZN(n12301) );
  NAND2_X1 U8464 ( .A1(n7107), .A2(n6851), .ZN(n7106) );
  INV_X1 U8465 ( .A(n6850), .ZN(n12330) );
  NOR2_X1 U8466 ( .A1(n12301), .A2(n15036), .ZN(n12319) );
  OAI211_X1 U8467 ( .C1(n12359), .C2(n6662), .A(n6660), .B(n6659), .ZN(n12341)
         );
  INV_X1 U8468 ( .A(n6661), .ZN(n6660) );
  NAND3_X1 U8469 ( .A1(n6662), .A2(n7104), .A3(n6573), .ZN(n6659) );
  OAI21_X1 U8470 ( .B1(n7104), .B2(n12359), .A(n6663), .ZN(n6661) );
  NOR2_X1 U8471 ( .A1(n12341), .A2(n12342), .ZN(n12358) );
  NOR2_X1 U8472 ( .A1(n12340), .A2(n6664), .ZN(n12360) );
  AOI21_X1 U8473 ( .B1(n12363), .B2(n12362), .A(n12361), .ZN(n12385) );
  XNOR2_X1 U8474 ( .A(n6763), .B(n12396), .ZN(n6762) );
  OR2_X1 U8475 ( .A1(n12394), .A2(n6764), .ZN(n6763) );
  AND2_X1 U8476 ( .A1(n14230), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U8477 ( .A1(n6761), .A2(n6572), .ZN(n6759) );
  NAND2_X1 U8478 ( .A1(n12401), .A2(n14810), .ZN(n6761) );
  NAND2_X1 U8479 ( .A1(n12398), .A2(n12397), .ZN(n6760) );
  INV_X1 U8480 ( .A(n7953), .ZN(n14298) );
  NAND2_X1 U8481 ( .A1(n7842), .A2(n7841), .ZN(n12507) );
  CLKBUF_X1 U8482 ( .A(n12521), .Z(n12522) );
  NAND2_X1 U8483 ( .A1(n12707), .A2(n6887), .ZN(n12527) );
  NAND2_X1 U8484 ( .A1(n7760), .A2(n7759), .ZN(n12721) );
  OR2_X1 U8485 ( .A1(n7801), .A2(n10344), .ZN(n7759) );
  CLKBUF_X1 U8486 ( .A(n12598), .Z(n12601) );
  AND3_X1 U8487 ( .A1(n7537), .A2(n7536), .A3(n7535), .ZN(n12067) );
  INV_X1 U8488 ( .A(n12466), .ZN(n14902) );
  NOR2_X1 U8489 ( .A1(n14954), .A2(n11298), .ZN(n14933) );
  NAND2_X1 U8490 ( .A1(n10660), .A2(n10534), .ZN(n14910) );
  INV_X1 U8491 ( .A(n12583), .ZN(n14281) );
  NAND2_X1 U8492 ( .A1(n10424), .A2(n6481), .ZN(n7445) );
  NAND2_X1 U8493 ( .A1(n6693), .A2(SI_0_), .ZN(n7446) );
  INV_X1 U8494 ( .A(n12677), .ZN(n14268) );
  INV_X1 U8495 ( .A(n14910), .ZN(n14901) );
  INV_X1 U8496 ( .A(n6624), .ZN(n6623) );
  OAI21_X1 U8497 ( .B1(n12687), .B2(n14305), .A(n6891), .ZN(n6624) );
  NOR2_X1 U8498 ( .A1(n6893), .A2(n6892), .ZN(n6891) );
  NOR2_X1 U8499 ( .A1(n12693), .A2(n7383), .ZN(n12759) );
  OR2_X1 U8500 ( .A1(n12713), .A2(n12712), .ZN(n12772) );
  NAND2_X1 U8501 ( .A1(n7744), .A2(n7743), .ZN(n12782) );
  AND2_X1 U8502 ( .A1(n12748), .A2(n12747), .ZN(n12799) );
  AND2_X1 U8503 ( .A1(n9696), .A2(n9695), .ZN(n12804) );
  INV_X1 U8504 ( .A(n12805), .ZN(n12803) );
  AND2_X1 U8505 ( .A1(n10422), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12805) );
  INV_X1 U8506 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12807) );
  NAND2_X1 U8507 ( .A1(n7200), .A2(n7874), .ZN(n7883) );
  CLKBUF_X1 U8508 ( .A(n8118), .Z(n8119) );
  NAND2_X1 U8509 ( .A1(n8108), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8110) );
  AND2_X1 U8510 ( .A1(n7959), .A2(n8099), .ZN(n10652) );
  NAND2_X1 U8511 ( .A1(n7933), .A2(n6525), .ZN(n10592) );
  NAND2_X1 U8512 ( .A1(n7769), .A2(n7770), .ZN(n7786) );
  INV_X1 U8513 ( .A(n10618), .ZN(n10345) );
  XNOR2_X1 U8514 ( .A(n7741), .B(n7740), .ZN(n12392) );
  NAND2_X1 U8515 ( .A1(n7177), .A2(n7716), .ZN(n7734) );
  NAND2_X1 U8516 ( .A1(n7715), .A2(n7714), .ZN(n7177) );
  INV_X1 U8517 ( .A(SI_15_), .ZN(n9928) );
  NAND2_X1 U8518 ( .A1(n7660), .A2(n7659), .ZN(n7677) );
  INV_X1 U8519 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7663) );
  INV_X1 U8520 ( .A(SI_12_), .ZN(n15112) );
  NAND2_X1 U8521 ( .A1(n7199), .A2(n6555), .ZN(n7623) );
  NAND2_X1 U8522 ( .A1(n7199), .A2(n7614), .ZN(n7617) );
  OR2_X1 U8523 ( .A1(n7584), .A2(n7583), .ZN(n11475) );
  INV_X1 U8524 ( .A(n14789), .ZN(n11056) );
  AOI22_X1 U8525 ( .A1(n6522), .A2(P3_IR_REG_0__SCAN_IN), .B1(n6758), .B2(
        n8112), .ZN(n6757) );
  NAND2_X1 U8526 ( .A1(n7309), .A2(n9344), .ZN(n11659) );
  NAND2_X1 U8527 ( .A1(n11022), .A2(n9268), .ZN(n11202) );
  AND2_X1 U8528 ( .A1(n10273), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12898) );
  NAND2_X1 U8529 ( .A1(n7315), .A2(n12837), .ZN(n7314) );
  INV_X1 U8530 ( .A(n7318), .ZN(n7315) );
  OR2_X1 U8531 ( .A1(n9134), .A2(n9777), .ZN(n9109) );
  OAI21_X1 U8532 ( .B1(n9111), .B2(n9776), .A(n9110), .ZN(n6589) );
  NOR2_X1 U8533 ( .A1(n11693), .A2(n11694), .ZN(n11692) );
  NAND2_X1 U8534 ( .A1(n9186), .A2(n10468), .ZN(n10474) );
  NAND2_X1 U8535 ( .A1(n7308), .A2(n9393), .ZN(n7305) );
  NAND2_X1 U8536 ( .A1(n7308), .A2(n7307), .ZN(n7306) );
  INV_X1 U8537 ( .A(n12871), .ZN(n7308) );
  NAND2_X1 U8538 ( .A1(n12880), .A2(n12879), .ZN(n12861) );
  NAND2_X1 U8539 ( .A1(n12822), .A2(n7387), .ZN(n12880) );
  XNOR2_X1 U8540 ( .A(n10467), .B(n9172), .ZN(n10336) );
  NAND2_X1 U8541 ( .A1(n11119), .A2(n9243), .ZN(n11129) );
  NAND2_X1 U8542 ( .A1(n11507), .A2(n9327), .ZN(n11561) );
  NOR2_X1 U8543 ( .A1(n7287), .A2(n7381), .ZN(n7286) );
  INV_X1 U8544 ( .A(n7290), .ZN(n7287) );
  NAND2_X1 U8545 ( .A1(n9456), .A2(n9455), .ZN(n13307) );
  NAND2_X1 U8546 ( .A1(n9433), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U8547 ( .A1(n11203), .A2(n9285), .ZN(n11331) );
  NAND2_X1 U8548 ( .A1(n9143), .A2(n10284), .ZN(n10291) );
  NAND2_X1 U8549 ( .A1(n10474), .A2(n9190), .ZN(n10986) );
  NAND2_X1 U8550 ( .A1(n9576), .A2(n9575), .ZN(n12908) );
  OAI21_X1 U8551 ( .B1(n9574), .B2(n10840), .A(n14716), .ZN(n12911) );
  INV_X1 U8552 ( .A(n11933), .ZN(n12950) );
  NAND2_X1 U8553 ( .A1(n6709), .A2(n10084), .ZN(n10087) );
  OR2_X1 U8554 ( .A1(n14620), .A2(n10085), .ZN(n6709) );
  AND2_X1 U8555 ( .A1(n6722), .A2(n6721), .ZN(n10207) );
  INV_X1 U8556 ( .A(n10164), .ZN(n6722) );
  INV_X1 U8557 ( .A(n10207), .ZN(n6719) );
  NOR2_X1 U8558 ( .A1(n10207), .A2(n6720), .ZN(n13021) );
  AND2_X1 U8559 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  NAND2_X1 U8560 ( .A1(n11584), .A2(n6582), .ZN(n13036) );
  OAI21_X1 U8561 ( .B1(n13049), .B2(n14700), .A(n13048), .ZN(n6700) );
  OAI22_X1 U8562 ( .A1(n13052), .A2(n14700), .B1(n13051), .B2(n13050), .ZN(
        n6698) );
  INV_X1 U8563 ( .A(n13055), .ZN(n13258) );
  OR3_X1 U8564 ( .A1(n13079), .A2(n13078), .A3(n13221), .ZN(n13264) );
  AND2_X1 U8565 ( .A1(n13073), .A2(n13072), .ZN(n13268) );
  INV_X1 U8566 ( .A(n13092), .ZN(n13272) );
  NAND2_X1 U8567 ( .A1(n13125), .A2(n11758), .ZN(n13111) );
  NAND2_X1 U8568 ( .A1(n6925), .A2(n11722), .ZN(n13138) );
  NAND2_X1 U8569 ( .A1(n6911), .A2(n6914), .ZN(n13188) );
  NAND2_X1 U8570 ( .A1(n13218), .A2(n6456), .ZN(n6911) );
  NAND2_X1 U8571 ( .A1(n9441), .A2(n9440), .ZN(n13321) );
  NAND2_X1 U8572 ( .A1(n9433), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U8573 ( .A1(n6918), .A2(n6917), .ZN(n13202) );
  NAND2_X1 U8574 ( .A1(n13244), .A2(n11748), .ZN(n13216) );
  NAND2_X1 U8575 ( .A1(n11746), .A2(n11879), .ZN(n13246) );
  NAND2_X1 U8576 ( .A1(n11635), .A2(n11634), .ZN(n11706) );
  NAND2_X1 U8577 ( .A1(n7074), .A2(n11382), .ZN(n11578) );
  NAND2_X1 U8578 ( .A1(n11231), .A2(n7078), .ZN(n7074) );
  NAND2_X1 U8579 ( .A1(n11231), .A2(n11230), .ZN(n11381) );
  NAND2_X1 U8580 ( .A1(n9349), .A2(n9348), .ZN(n11867) );
  NAND2_X1 U8581 ( .A1(n9310), .A2(n9309), .ZN(n14345) );
  NAND2_X1 U8582 ( .A1(n6910), .A2(n6909), .ZN(n11066) );
  AND2_X1 U8583 ( .A1(n6910), .A2(n6470), .ZN(n7376) );
  NAND2_X1 U8584 ( .A1(n11001), .A2(n12002), .ZN(n6910) );
  NAND2_X1 U8585 ( .A1(n11000), .A2(n10999), .ZN(n11074) );
  NAND2_X1 U8586 ( .A1(n7063), .A2(n10823), .ZN(n11026) );
  NAND2_X1 U8587 ( .A1(n10822), .A2(n11998), .ZN(n7063) );
  NAND2_X1 U8588 ( .A1(n6903), .A2(n10832), .ZN(n11027) );
  NAND2_X1 U8589 ( .A1(n10830), .A2(n10829), .ZN(n6903) );
  NAND2_X1 U8590 ( .A1(n14714), .A2(n10841), .ZN(n13242) );
  INV_X1 U8591 ( .A(n13242), .ZN(n13194) );
  INV_X1 U8592 ( .A(n13197), .ZN(n13251) );
  AND2_X1 U8593 ( .A1(n14714), .A2(n10873), .ZN(n13183) );
  OR3_X1 U8594 ( .A1(n13293), .A2(n13292), .A3(n13291), .ZN(n13348) );
  NAND2_X1 U8595 ( .A1(n13360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U8596 ( .A1(n6898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6897) );
  CLKBUF_X1 U8597 ( .A(n9969), .Z(n12039) );
  INV_X1 U8598 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10239) );
  INV_X1 U8599 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10161) );
  INV_X1 U8600 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10237) );
  INV_X1 U8601 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10057) );
  INV_X1 U8602 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9950) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9786) );
  INV_X1 U8604 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9775) );
  INV_X1 U8605 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9781) );
  INV_X1 U8606 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9773) );
  INV_X1 U8607 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9779) );
  INV_X1 U8608 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9777) );
  XNOR2_X1 U8609 ( .A(n6728), .B(P2_IR_REG_1__SCAN_IN), .ZN(n12985) );
  NOR2_X1 U8610 ( .A1(n9976), .A2(n9247), .ZN(n6728) );
  NAND2_X1 U8611 ( .A1(n7025), .A2(n7026), .ZN(n11182) );
  NAND2_X1 U8612 ( .A1(n10771), .A2(n7027), .ZN(n7025) );
  NAND2_X1 U8613 ( .A1(n14398), .A2(n7402), .ZN(n14359) );
  NAND2_X1 U8614 ( .A1(n11361), .A2(n11360), .ZN(n11499) );
  AND2_X1 U8615 ( .A1(n14379), .A2(n14254), .ZN(n14415) );
  NAND2_X1 U8616 ( .A1(n7018), .A2(n7021), .ZN(n11192) );
  NAND2_X1 U8617 ( .A1(n13581), .A2(n13454), .ZN(n13551) );
  AOI21_X1 U8618 ( .B1(n6998), .B2(n7000), .A(n6499), .ZN(n6996) );
  NAND2_X1 U8619 ( .A1(n7014), .A2(n7015), .ZN(n13566) );
  NAND2_X1 U8620 ( .A1(n13506), .A2(n13507), .ZN(n6997) );
  NOR2_X1 U8621 ( .A1(n10146), .A2(n10145), .ZN(n10149) );
  NAND2_X1 U8622 ( .A1(n7008), .A2(n7017), .ZN(n13600) );
  NAND2_X1 U8623 ( .A1(n7014), .A2(n7012), .ZN(n7008) );
  NAND2_X1 U8624 ( .A1(n8365), .A2(n8364), .ZN(n14141) );
  OAI21_X1 U8625 ( .B1(n10771), .B2(n10770), .A(n10769), .ZN(n11164) );
  NAND2_X1 U8626 ( .A1(n10047), .A2(n10046), .ZN(n14401) );
  INV_X1 U8627 ( .A(n14401), .ZN(n14421) );
  OR2_X1 U8628 ( .A1(n8715), .A2(n8887), .ZN(n7386) );
  INV_X1 U8629 ( .A(n10712), .ZN(n13624) );
  NAND4_X1 U8630 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n13625)
         );
  OR2_X1 U8631 ( .A1(n8542), .A2(n10363), .ZN(n8505) );
  NAND2_X1 U8632 ( .A1(n8697), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6927) );
  AND2_X1 U8633 ( .A1(n8686), .A2(n8685), .ZN(n14071) );
  INV_X1 U8634 ( .A(n14078), .ZN(n14072) );
  NAND2_X1 U8635 ( .A1(n8267), .A2(n8266), .ZN(n14085) );
  NAND2_X1 U8636 ( .A1(n11775), .A2(n8534), .ZN(n6783) );
  NAND2_X1 U8637 ( .A1(n13884), .A2(n13883), .ZN(n14091) );
  NAND2_X1 U8638 ( .A1(n7253), .A2(n7251), .ZN(n13895) );
  NAND2_X1 U8639 ( .A1(n13964), .A2(n13834), .ZN(n13946) );
  NAND2_X1 U8640 ( .A1(n8347), .A2(n8346), .ZN(n14125) );
  AND3_X1 U8641 ( .A1(n13992), .A2(n13991), .A3(n13990), .ZN(n14127) );
  NAND2_X1 U8642 ( .A1(n8643), .A2(n8642), .ZN(n14134) );
  NAND2_X1 U8643 ( .A1(n14049), .A2(n13824), .ZN(n14035) );
  OR2_X1 U8644 ( .A1(n13412), .A2(n6865), .ZN(n11616) );
  NAND2_X1 U8645 ( .A1(n11608), .A2(n11607), .ZN(n11622) );
  NAND2_X1 U8646 ( .A1(n8591), .A2(n8590), .ZN(n14238) );
  NAND2_X1 U8647 ( .A1(n11101), .A2(n11100), .ZN(n11216) );
  NAND2_X1 U8648 ( .A1(n11136), .A2(n11109), .ZN(n11213) );
  NAND2_X1 U8649 ( .A1(n15146), .A2(n14597), .ZN(n14065) );
  AOI211_X1 U8650 ( .C1(n14554), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n14541) );
  NAND2_X1 U8651 ( .A1(n15146), .A2(n10324), .ZN(n14260) );
  INV_X1 U8652 ( .A(n14065), .ZN(n14248) );
  INV_X2 U8653 ( .A(n14613), .ZN(n14615) );
  OR2_X1 U8654 ( .A1(n14105), .A2(n14104), .ZN(n14168) );
  INV_X2 U8655 ( .A(n14599), .ZN(n14601) );
  AND2_X1 U8656 ( .A1(n10706), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9797) );
  XNOR2_X1 U8657 ( .A(n8246), .B(n8245), .ZN(n14185) );
  OAI22_X1 U8658 ( .A1(n8684), .A2(n8243), .B1(n8242), .B2(n12060), .ZN(n8246)
         );
  NAND2_X1 U8659 ( .A1(n14182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U8660 ( .A1(n8250), .A2(n7390), .ZN(n6943) );
  INV_X1 U8661 ( .A(n9919), .ZN(n14200) );
  INV_X1 U8662 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n15099) );
  INV_X1 U8663 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10240) );
  INV_X1 U8664 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10261) );
  INV_X1 U8665 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10206) );
  INV_X1 U8666 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10055) );
  INV_X1 U8667 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9951) );
  INV_X1 U8668 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9820) );
  INV_X1 U8669 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9807) );
  INV_X1 U8670 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9801) );
  INV_X1 U8671 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9788) );
  INV_X1 U8672 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U8673 ( .A1(n7208), .A2(n8520), .ZN(n8509) );
  XNOR2_X1 U8674 ( .A(n8994), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U8675 ( .A1(n15167), .A2(n9003), .ZN(n15158) );
  INV_X1 U8676 ( .A(n9007), .ZN(n7094) );
  NAND2_X1 U8677 ( .A1(n14223), .A2(n9021), .ZN(n9023) );
  NAND2_X1 U8678 ( .A1(n14235), .A2(n14236), .ZN(n14234) );
  NAND2_X1 U8679 ( .A1(n14451), .A2(n14452), .ZN(n14450) );
  NOR2_X1 U8680 ( .A1(n9026), .A2(n9025), .ZN(n14455) );
  NAND2_X1 U8681 ( .A1(n14459), .A2(n9031), .ZN(n14463) );
  NAND2_X1 U8682 ( .A1(n14463), .A2(n14464), .ZN(n14462) );
  NAND2_X1 U8683 ( .A1(n6739), .A2(n14462), .ZN(n14467) );
  OAI21_X1 U8684 ( .B1(n14463), .B2(n14464), .A(n6740), .ZN(n6739) );
  INV_X1 U8685 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8686 ( .A1(n7089), .A2(n7088), .ZN(n14473) );
  INV_X1 U8687 ( .A(n9035), .ZN(n7088) );
  AOI21_X1 U8688 ( .B1(n9692), .B2(n6969), .A(n9731), .ZN(n6967) );
  NOR2_X1 U8689 ( .A1(n10640), .A2(n9618), .ZN(n10632) );
  OAI21_X1 U8690 ( .B1(n10577), .B2(n10576), .A(n6459), .ZN(n10560) );
  OAI21_X1 U8691 ( .B1(n6625), .B2(n14815), .A(n12402), .ZN(P3_U3201) );
  XNOR2_X1 U8692 ( .A(n6626), .B(n12389), .ZN(n6625) );
  AOI21_X1 U8693 ( .B1(n6762), .B2(n14809), .A(n6759), .ZN(n12402) );
  OR2_X1 U8694 ( .A1(n12385), .A2(n12384), .ZN(n6626) );
  INV_X1 U8695 ( .A(n6619), .ZN(n6618) );
  OAI22_X1 U8696 ( .A1(n12758), .A2(n12751), .B1(n14993), .B2(n12691), .ZN(
        n6619) );
  NAND2_X1 U8697 ( .A1(n7324), .A2(n7323), .ZN(P3_U3456) );
  NAND2_X1 U8698 ( .A1(n14973), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U8699 ( .A1(n12755), .A2(n14975), .ZN(n7324) );
  INV_X1 U8700 ( .A(n6621), .ZN(n6620) );
  OAI22_X1 U8701 ( .A1(n12758), .A2(n12802), .B1(n14975), .B2(n12757), .ZN(
        n6621) );
  NAND2_X1 U8702 ( .A1(n6593), .A2(n6590), .ZN(P2_U3212) );
  AOI21_X1 U8703 ( .B1(n6592), .B2(n6591), .A(n12925), .ZN(n6590) );
  NAND2_X1 U8704 ( .A1(n6699), .A2(n6696), .ZN(P2_U3233) );
  AOI21_X1 U8705 ( .B1(n6698), .B2(n13053), .A(n6697), .ZN(n6696) );
  NAND2_X1 U8706 ( .A1(n6700), .A2(n12027), .ZN(n6699) );
  OAI21_X1 U8707 ( .B1(n14705), .B2(n7432), .A(n13054), .ZN(n6697) );
  NOR2_X1 U8708 ( .A1(n14776), .A2(n14749), .ZN(n7053) );
  AND2_X1 U8709 ( .A1(n7058), .A2(n7056), .ZN(n6777) );
  NAND2_X1 U8710 ( .A1(n6746), .A2(n6743), .ZN(n15165) );
  INV_X1 U8711 ( .A(n6749), .ZN(n15164) );
  OAI21_X1 U8712 ( .B1(n14217), .B2(n9013), .A(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n6743) );
  NAND2_X1 U8713 ( .A1(n14203), .A2(n6730), .ZN(n6729) );
  NAND2_X1 U8714 ( .A1(n6732), .A2(n6731), .ZN(n6730) );
  XNOR2_X1 U8715 ( .A(n7109), .B(n7108), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8716 ( .A(n9046), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U8717 ( .A1(n14203), .A2(n7110), .ZN(n7109) );
  CLKBUF_X3 U8718 ( .A(n11797), .Z(n11967) );
  AND2_X1 U8719 ( .A1(n6801), .A2(n8172), .ZN(n6437) );
  INV_X2 U8720 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8112) );
  AND2_X1 U8721 ( .A1(n6974), .A2(n12525), .ZN(n6438) );
  OR2_X1 U8722 ( .A1(n15148), .A2(n11165), .ZN(n6439) );
  AND2_X1 U8723 ( .A1(n7115), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6440) );
  INV_X1 U8724 ( .A(n8178), .ZN(n9737) );
  NAND2_X1 U8725 ( .A1(n8302), .A2(n8301), .ZN(n14098) );
  INV_X1 U8726 ( .A(n14098), .ZN(n7250) );
  XNOR2_X1 U8727 ( .A(n8110), .B(n8109), .ZN(n9602) );
  AND2_X1 U8728 ( .A1(n8806), .A2(n8892), .ZN(n6441) );
  AND2_X1 U8729 ( .A1(n7410), .A2(n6993), .ZN(n6442) );
  OR2_X1 U8730 ( .A1(n14783), .A2(n6556), .ZN(n6443) );
  AND2_X1 U8731 ( .A1(n6870), .A2(n6868), .ZN(n6444) );
  AND2_X1 U8732 ( .A1(n13416), .A2(n6458), .ZN(n6445) );
  INV_X1 U8733 ( .A(n6980), .ZN(n6979) );
  NAND2_X1 U8734 ( .A1(n6984), .A2(n6464), .ZN(n6980) );
  NOR2_X1 U8735 ( .A1(n7250), .A2(n13839), .ZN(n6446) );
  INV_X1 U8736 ( .A(n8163), .ZN(n6803) );
  AND2_X1 U8737 ( .A1(n13808), .A2(n6944), .ZN(n6447) );
  NOR2_X1 U8738 ( .A1(n6738), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8739 ( .A1(n9622), .A2(n9611), .ZN(n6449) );
  AND2_X1 U8740 ( .A1(n13262), .A2(n6557), .ZN(n6450) );
  AND2_X1 U8741 ( .A1(n7056), .A2(n6557), .ZN(n6451) );
  INV_X1 U8742 ( .A(n14019), .ZN(n7130) );
  AND2_X1 U8743 ( .A1(n6655), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6452) );
  INV_X1 U8744 ( .A(n12359), .ZN(n14210) );
  NAND2_X1 U8745 ( .A1(n9946), .A2(n9945), .ZN(n14776) );
  NAND2_X1 U8746 ( .A1(n10794), .A2(n10390), .ZN(n10725) );
  INV_X1 U8747 ( .A(n11523), .ZN(n7102) );
  NAND2_X1 U8748 ( .A1(n6719), .A2(n6725), .ZN(n6453) );
  AND2_X1 U8749 ( .A1(n7105), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6454) );
  INV_X4 U8750 ( .A(n8324), .ZN(n8231) );
  OR2_X1 U8751 ( .A1(n11568), .A2(n11567), .ZN(n6455) );
  AND2_X1 U8752 ( .A1(n6916), .A2(n6917), .ZN(n6456) );
  NAND2_X1 U8753 ( .A1(n7408), .A2(n7409), .ZN(n6457) );
  NAND2_X1 U8754 ( .A1(n13422), .A2(n13421), .ZN(n6458) );
  OR2_X1 U8755 ( .A1(n10410), .A2(n10444), .ZN(n6459) );
  INV_X1 U8756 ( .A(n12008), .ZN(n6923) );
  INV_X1 U8757 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U8758 ( .A1(n7560), .A2(n6988), .ZN(n7582) );
  OR2_X1 U8759 ( .A1(n7343), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n6460) );
  XOR2_X1 U8760 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), .Z(
        n6461) );
  NAND2_X1 U8761 ( .A1(n7334), .A2(n6649), .ZN(n7436) );
  INV_X1 U8762 ( .A(n7322), .ZN(n9132) );
  OR2_X1 U8763 ( .A1(n12665), .A2(n12664), .ZN(n6462) );
  OR2_X1 U8764 ( .A1(n9015), .A2(n9016), .ZN(n6463) );
  OR2_X1 U8765 ( .A1(n9643), .A2(n9644), .ZN(n6464) );
  INV_X1 U8766 ( .A(n6977), .ZN(n6976) );
  NAND2_X1 U8767 ( .A1(n9648), .A2(n6978), .ZN(n6977) );
  AND2_X1 U8768 ( .A1(n11724), .A2(n11722), .ZN(n6465) );
  INV_X1 U8769 ( .A(n12602), .ZN(n12608) );
  AND2_X1 U8770 ( .A1(n8034), .A2(n8037), .ZN(n12602) );
  NOR2_X1 U8771 ( .A1(n8542), .A2(n8514), .ZN(n6466) );
  NAND2_X1 U8772 ( .A1(n8605), .A2(n8604), .ZN(n11358) );
  AND2_X1 U8773 ( .A1(n6622), .A2(n6858), .ZN(n6467) );
  OR2_X1 U8774 ( .A1(n8326), .A2(n13631), .ZN(n6468) );
  AND2_X1 U8775 ( .A1(n7560), .A2(n7408), .ZN(n7562) );
  NOR2_X1 U8776 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7208) );
  NAND2_X1 U8777 ( .A1(n7332), .A2(n12435), .ZN(n12556) );
  NAND2_X1 U8778 ( .A1(n6997), .A2(n13474), .ZN(n13574) );
  AND2_X1 U8779 ( .A1(n12013), .A2(n7078), .ZN(n6469) );
  OR2_X1 U8780 ( .A1(n11843), .A2(n11002), .ZN(n6470) );
  NAND2_X1 U8781 ( .A1(n8387), .A2(n8386), .ZN(n13412) );
  OR2_X1 U8782 ( .A1(n10786), .A2(n10776), .ZN(n6471) );
  OR3_X1 U8783 ( .A1(n8711), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n6472) );
  OR2_X1 U8784 ( .A1(n11527), .A2(n11526), .ZN(n6473) );
  NAND2_X1 U8785 ( .A1(n8427), .A2(n8426), .ZN(n14406) );
  INV_X2 U8786 ( .A(n9619), .ZN(n12045) );
  INV_X1 U8787 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8259) );
  INV_X1 U8788 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9098) );
  OR2_X1 U8789 ( .A1(n12278), .A2(n12277), .ZN(n6474) );
  AND2_X1 U8790 ( .A1(n7242), .A2(n6804), .ZN(n6475) );
  INV_X1 U8791 ( .A(n12439), .ZN(n12540) );
  INV_X1 U8792 ( .A(n12879), .ZN(n7300) );
  AND2_X1 U8793 ( .A1(n9691), .A2(n6685), .ZN(n6476) );
  NAND2_X1 U8794 ( .A1(n9073), .A2(n9072), .ZN(n13195) );
  INV_X1 U8795 ( .A(n13839), .ZN(n13881) );
  INV_X1 U8796 ( .A(n10786), .ZN(n14561) );
  XOR2_X1 U8797 ( .A(n12709), .B(n9682), .Z(n6477) );
  NAND2_X1 U8798 ( .A1(n8517), .A2(n8516), .ZN(n13626) );
  INV_X1 U8799 ( .A(n13626), .ZN(n8526) );
  XOR2_X1 U8800 ( .A(n12022), .B(n12027), .Z(n6479) );
  INV_X1 U8801 ( .A(n10435), .ZN(n7115) );
  INV_X1 U8802 ( .A(n8860), .ZN(n7154) );
  OR2_X1 U8803 ( .A1(n13326), .A2(n12959), .ZN(n6480) );
  INV_X1 U8804 ( .A(n8774), .ZN(n7151) );
  INV_X1 U8805 ( .A(n8882), .ZN(n7148) );
  AND2_X1 U8806 ( .A1(n9771), .A2(n6884), .ZN(n6481) );
  OR2_X1 U8807 ( .A1(n14332), .A2(n12963), .ZN(n6482) );
  NAND2_X1 U8808 ( .A1(n11492), .A2(n13617), .ZN(n6483) );
  NOR2_X1 U8809 ( .A1(n14360), .A2(n7036), .ZN(n7035) );
  AND3_X1 U8810 ( .A1(n8085), .A2(n7188), .A3(n8089), .ZN(n6484) );
  AND2_X1 U8811 ( .A1(n12562), .A2(n12575), .ZN(n6485) );
  AND3_X1 U8812 ( .A1(n7288), .A2(n7290), .A3(n7285), .ZN(n6486) );
  NOR2_X1 U8813 ( .A1(n12535), .A2(n6477), .ZN(n6487) );
  NAND2_X1 U8814 ( .A1(n9467), .A2(n9466), .ZN(n13159) );
  AND3_X1 U8815 ( .A1(n6471), .A2(n7236), .A3(n6439), .ZN(n6488) );
  AND4_X1 U8816 ( .A1(n7513), .A2(n7512), .A3(n7511), .A4(n7510), .ZN(n11315)
         );
  INV_X1 U8817 ( .A(n11315), .ZN(n14855) );
  AND2_X1 U8818 ( .A1(n6449), .A2(n12175), .ZN(n6489) );
  AND2_X1 U8819 ( .A1(n11847), .A2(n12967), .ZN(n6490) );
  NOR2_X1 U8820 ( .A1(n12319), .A2(n12318), .ZN(n6491) );
  NOR2_X1 U8821 ( .A1(n14406), .A2(n14361), .ZN(n6492) );
  INV_X1 U8822 ( .A(n8172), .ZN(n7261) );
  AND2_X1 U8823 ( .A1(n13408), .A2(n13407), .ZN(n6493) );
  INV_X1 U8824 ( .A(n9645), .ZN(n6982) );
  INV_X1 U8825 ( .A(n10751), .ZN(n6810) );
  INV_X1 U8826 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8251) );
  INV_X1 U8827 ( .A(n10489), .ZN(n11046) );
  INV_X1 U8828 ( .A(n13834), .ZN(n7224) );
  OR2_X1 U8829 ( .A1(n11957), .A2(n11956), .ZN(n6494) );
  NOR2_X1 U8830 ( .A1(n11181), .A2(n7024), .ZN(n7023) );
  INV_X1 U8831 ( .A(n8842), .ZN(n7157) );
  INV_X1 U8832 ( .A(n8870), .ZN(n7163) );
  AND2_X1 U8833 ( .A1(n13282), .A2(n11929), .ZN(n6495) );
  INV_X1 U8834 ( .A(n11914), .ZN(n7369) );
  AND2_X1 U8835 ( .A1(n11847), .A2(n11065), .ZN(n6496) );
  AND2_X1 U8836 ( .A1(n6962), .A2(n12064), .ZN(n6497) );
  AND2_X1 U8837 ( .A1(n7050), .A2(n7048), .ZN(n6498) );
  AND2_X1 U8838 ( .A1(n13480), .A2(n13479), .ZN(n6499) );
  INV_X1 U8839 ( .A(n7252), .ZN(n7251) );
  NOR2_X1 U8840 ( .A1(n13788), .A2(n13933), .ZN(n7252) );
  NAND2_X1 U8841 ( .A1(n10412), .A2(n10573), .ZN(n6821) );
  INV_X1 U8842 ( .A(n6821), .ZN(n6813) );
  NOR2_X1 U8843 ( .A1(n14746), .A2(n12972), .ZN(n6500) );
  NOR2_X1 U8844 ( .A1(n14587), .A2(n13619), .ZN(n6501) );
  NOR2_X1 U8845 ( .A1(n13386), .A2(n13385), .ZN(n6502) );
  NOR2_X1 U8846 ( .A1(n13195), .A2(n12957), .ZN(n6503) );
  AND2_X1 U8847 ( .A1(n6918), .A2(n6456), .ZN(n6504) );
  AND2_X1 U8848 ( .A1(n7247), .A2(n7245), .ZN(n6505) );
  INV_X1 U8849 ( .A(n9107), .ZN(n9932) );
  AND2_X1 U8850 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n6506) );
  AND2_X1 U8851 ( .A1(n7021), .A2(n7020), .ZN(n6507) );
  AND2_X1 U8852 ( .A1(n11299), .A2(n7467), .ZN(n6508) );
  INV_X1 U8853 ( .A(n13812), .ZN(n13914) );
  INV_X1 U8854 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8256) );
  OR2_X1 U8855 ( .A1(n10849), .A2(n10856), .ZN(n6509) );
  NAND2_X1 U8856 ( .A1(n13195), .A2(n11717), .ZN(n6510) );
  NAND3_X1 U8857 ( .A1(n6987), .A2(n6478), .A3(n7560), .ZN(n6511) );
  OR2_X1 U8858 ( .A1(n8708), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6512) );
  AND4_X1 U8859 ( .A1(n8129), .A2(n8126), .A3(n8128), .A4(n8127), .ZN(n6513)
         );
  INV_X1 U8860 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7431) );
  NOR2_X1 U8861 ( .A1(n14746), .A2(n11120), .ZN(n6514) );
  AND2_X1 U8862 ( .A1(n8154), .A2(SI_6_), .ZN(n6515) );
  INV_X1 U8863 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7410) );
  AND2_X1 U8864 ( .A1(n14825), .A2(n11671), .ZN(n6516) );
  INV_X1 U8865 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7740) );
  INV_X1 U8866 ( .A(n6947), .ZN(n6946) );
  NAND2_X1 U8867 ( .A1(n14013), .A2(n6949), .ZN(n6947) );
  INV_X1 U8868 ( .A(n6888), .ZN(n6887) );
  NAND2_X1 U8869 ( .A1(n7823), .A2(n8059), .ZN(n6888) );
  AND3_X1 U8870 ( .A1(n8528), .A2(n8529), .A3(n8530), .ZN(n6517) );
  AND2_X1 U8871 ( .A1(n9655), .A2(n12429), .ZN(n6518) );
  OR2_X1 U8872 ( .A1(n7388), .A2(n7377), .ZN(n6519) );
  AND2_X1 U8873 ( .A1(n9788), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6520) );
  AND2_X1 U8874 ( .A1(n13825), .A2(n8823), .ZN(n6521) );
  OAI21_X1 U8875 ( .B1(n7262), .B2(n7261), .A(n7393), .ZN(n7260) );
  AND2_X1 U8876 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n6522) );
  AND2_X1 U8877 ( .A1(n11179), .A2(n7029), .ZN(n6523) );
  NAND2_X1 U8878 ( .A1(n8209), .A2(n7254), .ZN(n6524) );
  INV_X1 U8879 ( .A(n6704), .ZN(n6703) );
  NAND2_X1 U8880 ( .A1(n6707), .A2(n6564), .ZN(n6704) );
  INV_X1 U8881 ( .A(n9162), .ZN(n6766) );
  NAND2_X1 U8882 ( .A1(n6622), .A2(n6442), .ZN(n6525) );
  AND2_X1 U8883 ( .A1(n9021), .A2(n6738), .ZN(n6526) );
  AND2_X1 U8884 ( .A1(n8270), .A2(n8269), .ZN(n8625) );
  INV_X2 U8885 ( .A(n8625), .ZN(n8676) );
  AND2_X1 U8886 ( .A1(n6456), .A2(n11718), .ZN(n6527) );
  AND2_X1 U8887 ( .A1(n12707), .A2(n8059), .ZN(n6528) );
  AND2_X1 U8888 ( .A1(n11609), .A2(n11607), .ZN(n6529) );
  OR2_X1 U8889 ( .A1(n13832), .A2(n7224), .ZN(n6530) );
  AND2_X1 U8890 ( .A1(n8155), .A2(n8158), .ZN(n6531) );
  AND2_X1 U8891 ( .A1(n9280), .A2(n9268), .ZN(n6532) );
  AND2_X1 U8892 ( .A1(n9362), .A2(n9344), .ZN(n6533) );
  XNOR2_X1 U8893 ( .A(n11298), .B(n12045), .ZN(n9620) );
  AND2_X1 U8894 ( .A1(n12929), .A2(n7318), .ZN(n6534) );
  OR2_X1 U8895 ( .A1(n7163), .A2(n8869), .ZN(n6535) );
  OR2_X1 U8896 ( .A1(n7157), .A2(n8841), .ZN(n6536) );
  OR2_X1 U8897 ( .A1(n11904), .A2(n11902), .ZN(n6537) );
  AND2_X1 U8898 ( .A1(n14018), .A2(n13827), .ZN(n6538) );
  OR2_X1 U8899 ( .A1(n8785), .A2(n8783), .ZN(n6539) );
  OR2_X1 U8900 ( .A1(n8763), .A2(n8761), .ZN(n6540) );
  OR2_X1 U8901 ( .A1(n11822), .A2(n11820), .ZN(n6541) );
  OR2_X1 U8902 ( .A1(n11858), .A2(n11856), .ZN(n6542) );
  AND2_X1 U8903 ( .A1(n6706), .A2(n6712), .ZN(n6543) );
  OR2_X1 U8904 ( .A1(n7358), .A2(n11832), .ZN(n6544) );
  OR2_X1 U8905 ( .A1(n7360), .A2(n11821), .ZN(n6545) );
  OR2_X1 U8906 ( .A1(n7362), .A2(n11845), .ZN(n6546) );
  OR2_X1 U8907 ( .A1(n11913), .A2(n7369), .ZN(n6547) );
  OR2_X1 U8908 ( .A1(n7154), .A2(n8859), .ZN(n6548) );
  OR2_X1 U8909 ( .A1(n7148), .A2(n8881), .ZN(n6549) );
  OR2_X1 U8910 ( .A1(n7151), .A2(n8773), .ZN(n6550) );
  OR2_X1 U8911 ( .A1(n11831), .A2(n11833), .ZN(n6551) );
  OR2_X1 U8912 ( .A1(n11844), .A2(n11846), .ZN(n6552) );
  NAND2_X1 U8913 ( .A1(n9412), .A2(n9411), .ZN(n13330) );
  INV_X1 U8914 ( .A(n13836), .ZN(n7225) );
  NAND2_X1 U8915 ( .A1(n7354), .A2(n11875), .ZN(n6553) );
  INV_X1 U8916 ( .A(n7083), .ZN(n7082) );
  OR2_X1 U8917 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6554) );
  INV_X1 U8918 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6758) );
  OR2_X1 U8919 ( .A1(n13428), .A2(n13427), .ZN(n7017) );
  INV_X1 U8920 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8252) );
  INV_X1 U8921 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8922 ( .A1(n6445), .A2(n14411), .ZN(n7014) );
  XNOR2_X1 U8923 ( .A(n8927), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U8924 ( .A1(n11746), .A2(n7086), .ZN(n13244) );
  AND2_X1 U8925 ( .A1(n7198), .A2(n7614), .ZN(n6555) );
  INV_X1 U8926 ( .A(n12535), .ZN(n12558) );
  AND2_X1 U8927 ( .A1(n11056), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6556) );
  AND2_X1 U8928 ( .A1(n11743), .A2(n11742), .ZN(n6557) );
  NAND2_X1 U8929 ( .A1(n13209), .A2(n6771), .ZN(n6558) );
  NAND2_X1 U8930 ( .A1(n14823), .A2(n11650), .ZN(n11670) );
  OAI21_X1 U8931 ( .B1(n11684), .B2(n6682), .A(n6680), .ZN(n12206) );
  OAI21_X1 U8932 ( .B1(n11684), .B2(n6977), .A(n6975), .ZN(n12157) );
  NAND2_X1 U8933 ( .A1(n14245), .A2(n6864), .ZN(n6865) );
  NOR2_X1 U8934 ( .A1(n7479), .A2(n7407), .ZN(n7560) );
  INV_X1 U8935 ( .A(n14839), .ZN(n12253) );
  AND4_X1 U8936 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n14839)
         );
  NOR2_X1 U8937 ( .A1(n11692), .A2(n9393), .ZN(n6559) );
  NAND2_X1 U8938 ( .A1(n12252), .A2(n12201), .ZN(n6560) );
  NAND2_X1 U8939 ( .A1(n11388), .A2(n6773), .ZN(n6776) );
  AND2_X1 U8940 ( .A1(n6948), .A2(n6949), .ZN(n6561) );
  AND2_X1 U8941 ( .A1(n14398), .A2(n7035), .ZN(n6562) );
  NOR2_X1 U8942 ( .A1(n14039), .A2(n14134), .ZN(n14005) );
  OR2_X1 U8943 ( .A1(n12289), .A2(n14216), .ZN(n6563) );
  NAND2_X1 U8944 ( .A1(n9991), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6564) );
  INV_X1 U8945 ( .A(n10476), .ZN(n7112) );
  AND2_X1 U8946 ( .A1(n6455), .A2(n11570), .ZN(n6565) );
  OR2_X1 U8947 ( .A1(n6556), .A2(n11474), .ZN(n6566) );
  AND2_X1 U8948 ( .A1(n13822), .A2(n13821), .ZN(n6567) );
  INV_X1 U8949 ( .A(n6717), .ZN(n6716) );
  OAI21_X1 U8950 ( .B1(n6720), .B2(n6721), .A(n6718), .ZN(n6717) );
  INV_X1 U8951 ( .A(n12928), .ZN(n6591) );
  INV_X1 U8952 ( .A(n12332), .ZN(n6851) );
  NAND2_X1 U8953 ( .A1(n6965), .A2(n9606), .ZN(n9693) );
  NAND2_X1 U8954 ( .A1(n8442), .A2(n8441), .ZN(n11492) );
  INV_X1 U8955 ( .A(n11492), .ZN(n6870) );
  AND2_X1 U8956 ( .A1(n12263), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6568) );
  AND2_X1 U8957 ( .A1(n6806), .A2(n6811), .ZN(n6569) );
  INV_X1 U8958 ( .A(n6908), .ZN(n6909) );
  AND2_X1 U8959 ( .A1(n7237), .A2(n10380), .ZN(n6570) );
  INV_X1 U8960 ( .A(n12267), .ZN(n12263) );
  NAND2_X1 U8961 ( .A1(n6890), .A2(n8007), .ZN(n11668) );
  AND2_X1 U8962 ( .A1(n10666), .A2(n10665), .ZN(n14973) );
  INV_X1 U8963 ( .A(n12344), .ZN(n14222) );
  INV_X1 U8964 ( .A(n7230), .ZN(n7235) );
  NOR2_X1 U8965 ( .A1(n12262), .A2(n6837), .ZN(n6571) );
  NOR2_X1 U8966 ( .A1(n12400), .A2(n6760), .ZN(n6572) );
  NAND2_X1 U8967 ( .A1(n11478), .A2(n11536), .ZN(n11520) );
  NOR2_X1 U8968 ( .A1(n6664), .A2(n14210), .ZN(n6573) );
  NOR2_X1 U8969 ( .A1(n6568), .A2(n14216), .ZN(n6574) );
  AND2_X1 U8970 ( .A1(n7099), .A2(n11520), .ZN(n6575) );
  INV_X1 U8971 ( .A(n8655), .ZN(n7276) );
  AND2_X1 U8972 ( .A1(n6935), .A2(n6483), .ZN(n6576) );
  AND2_X1 U8973 ( .A1(n11108), .A2(n11107), .ZN(n6577) );
  AND2_X1 U8974 ( .A1(n14852), .A2(n11309), .ZN(n6578) );
  INV_X1 U8975 ( .A(n14753), .ZN(n7052) );
  INV_X2 U8976 ( .A(n14973), .ZN(n14975) );
  NOR2_X1 U8977 ( .A1(n10348), .A2(n10322), .ZN(n6579) );
  INV_X1 U8978 ( .A(n13951), .ZN(n14254) );
  AND2_X2 U8979 ( .A1(n10626), .A2(n10625), .ZN(n14993) );
  INV_X1 U8980 ( .A(n14954), .ZN(n14907) );
  AND2_X1 U8981 ( .A1(n9715), .A2(n10660), .ZN(n12229) );
  AND2_X1 U8982 ( .A1(n11444), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6580) );
  AND2_X1 U8983 ( .A1(n10779), .A2(n10778), .ZN(n6581) );
  INV_X1 U8984 ( .A(n10750), .ZN(n6820) );
  NAND2_X1 U8985 ( .A1(n12265), .A2(n6834), .ZN(n6833) );
  INV_X1 U8986 ( .A(n6833), .ZN(n6829) );
  OR2_X1 U8987 ( .A1(n11588), .A2(n11439), .ZN(n6582) );
  AND2_X1 U8988 ( .A1(n6705), .A2(n6703), .ZN(n6583) );
  AND2_X1 U8989 ( .A1(n7114), .A2(n10432), .ZN(n6584) );
  AND2_X1 U8990 ( .A1(n6705), .A2(n6707), .ZN(n6585) );
  OR2_X1 U8991 ( .A1(n13370), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U8992 ( .A1(n8937), .A2(n13639), .ZN(n6587) );
  INV_X1 U8993 ( .A(n10209), .ZN(n6723) );
  INV_X1 U8994 ( .A(n6725), .ZN(n6724) );
  NAND2_X1 U8995 ( .A1(n10210), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8996 ( .A1(n6757), .A2(n7454), .ZN(n10502) );
  INV_X1 U8997 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6752) );
  INV_X1 U8998 ( .A(n14571), .ZN(n13878) );
  NAND2_X1 U8999 ( .A1(n6472), .A2(n7123), .ZN(n9919) );
  AOI21_X1 U9000 ( .B1(n14080), .B2(n14554), .A(n14079), .ZN(n14081) );
  AND2_X1 U9001 ( .A1(n15146), .A2(n14554), .ZN(n13863) );
  NAND2_X1 U9002 ( .A1(n10474), .A2(n7312), .ZN(n10984) );
  NAND2_X1 U9003 ( .A1(n11022), .A2(n6532), .ZN(n11203) );
  NAND2_X2 U9004 ( .A1(n9148), .A2(n9771), .ZN(n9134) );
  NAND2_X1 U9005 ( .A1(n11507), .A2(n7310), .ZN(n7309) );
  OAI21_X2 U9006 ( .B1(n12891), .B2(n12887), .A(n12888), .ZN(n12851) );
  XNOR2_X1 U9007 ( .A(n10282), .B(n9128), .ZN(n10277) );
  NAND2_X1 U9008 ( .A1(n10330), .A2(n9174), .ZN(n9186) );
  NAND2_X2 U9009 ( .A1(n9109), .A2(n6588), .ZN(n11784) );
  INV_X1 U9010 ( .A(n6589), .ZN(n6588) );
  NAND2_X1 U9011 ( .A1(n12927), .A2(n12926), .ZN(n6593) );
  NAND3_X1 U9012 ( .A1(n6596), .A2(n7296), .A3(n6595), .ZN(n9509) );
  NAND2_X1 U9013 ( .A1(n12831), .A2(n12830), .ZN(n12829) );
  NAND2_X1 U9014 ( .A1(n13141), .A2(n11725), .ZN(n13118) );
  OAI21_X2 U9015 ( .B1(n13231), .B2(n11711), .A(n11710), .ZN(n13218) );
  OAI21_X1 U9016 ( .B1(n10830), .B2(n6900), .A(n6899), .ZN(n10857) );
  NAND3_X1 U9017 ( .A1(n9062), .A2(n6766), .A3(n7366), .ZN(n9096) );
  NAND2_X1 U9018 ( .A1(n13116), .A2(n7397), .ZN(n13102) );
  NAND2_X1 U9019 ( .A1(n10194), .A2(n10193), .ZN(n10249) );
  NAND2_X1 U9020 ( .A1(n10189), .A2(n10188), .ZN(n10960) );
  OAI21_X1 U9021 ( .B1(n6455), .B2(n6921), .A(n6919), .ZN(n11709) );
  NOR2_X2 U9022 ( .A1(n7345), .A2(n9061), .ZN(n7366) );
  AOI21_X1 U9023 ( .B1(n7221), .B2(n7222), .A(n13929), .ZN(n7219) );
  NAND2_X1 U9024 ( .A1(n8177), .A2(n8176), .ZN(n8418) );
  NAND2_X1 U9025 ( .A1(n7247), .A2(n7249), .ZN(n13877) );
  NAND2_X1 U9026 ( .A1(n8568), .A2(n6790), .ZN(n6788) );
  AOI22_X1 U9027 ( .A1(n12905), .A2(n12904), .B1(n9424), .B2(n9423), .ZN(
        n12831) );
  INV_X1 U9028 ( .A(n12931), .ZN(n11658) );
  INV_X1 U9029 ( .A(n7387), .ZN(n7299) );
  NAND2_X2 U9030 ( .A1(n6607), .A2(n13053), .ZN(n10917) );
  NAND3_X1 U9031 ( .A1(n7302), .A2(n7301), .A3(n7303), .ZN(n6607) );
  NAND2_X2 U9032 ( .A1(n12851), .A2(n12850), .ZN(n12849) );
  OAI21_X1 U9033 ( .B1(n9601), .B2(n6534), .A(n9600), .ZN(P2_U3186) );
  NAND2_X1 U9034 ( .A1(n12823), .A2(n9478), .ZN(n12822) );
  NAND2_X1 U9035 ( .A1(n6608), .A2(n7352), .ZN(n11881) );
  NAND3_X1 U9036 ( .A1(n6616), .A2(n6553), .A3(n6615), .ZN(n6608) );
  OR2_X2 U9037 ( .A1(n11229), .A2(n11228), .ZN(n11231) );
  NAND2_X1 U9038 ( .A1(n7070), .A2(n7069), .ZN(n13097) );
  XNOR2_X1 U9039 ( .A(n11762), .B(n11761), .ZN(n13259) );
  NAND2_X1 U9040 ( .A1(n10579), .A2(n10446), .ZN(n10566) );
  NAND2_X1 U9041 ( .A1(n10580), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10579) );
  NAND2_X1 U9042 ( .A1(n11873), .A2(n11872), .ZN(n6615) );
  NAND2_X1 U9043 ( .A1(n11869), .A2(n11868), .ZN(n6616) );
  NOR3_X4 U9044 ( .A1(n7932), .A2(n6460), .A3(P3_IR_REG_28__SCAN_IN), .ZN(
        n7428) );
  NAND3_X1 U9045 ( .A1(n7401), .A2(n9083), .A3(n6617), .ZN(n9085) );
  OAI21_X2 U9046 ( .B1(n12500), .B2(n12501), .A(n12450), .ZN(n12484) );
  NAND2_X1 U9047 ( .A1(n7321), .A2(n7322), .ZN(n7320) );
  NAND2_X1 U9048 ( .A1(n12464), .A2(n6623), .ZN(n12755) );
  AOI21_X1 U9049 ( .B1(n11673), .B2(n6560), .A(n7395), .ZN(n11675) );
  INV_X1 U9050 ( .A(n13139), .ZN(n11724) );
  NAND2_X1 U9051 ( .A1(n7054), .A2(n6777), .ZN(n13344) );
  NAND2_X1 U9052 ( .A1(n14918), .A2(n10517), .ZN(n7966) );
  XNOR2_X2 U9053 ( .A(n7416), .B(n12807), .ZN(n12062) );
  OAI21_X1 U9054 ( .B1(n12756), .B2(n14990), .A(n6618), .ZN(P3_U3487) );
  OAI21_X1 U9055 ( .B1(n12756), .B2(n14973), .A(n6620), .ZN(P3_U3455) );
  NAND2_X1 U9056 ( .A1(n9160), .A2(n9171), .ZN(n10370) );
  NAND2_X1 U9057 ( .A1(n7283), .A2(n10291), .ZN(n10329) );
  NAND2_X1 U9058 ( .A1(n12023), .A2(n11777), .ZN(n7302) );
  NAND3_X1 U9059 ( .A1(n7288), .A2(n7285), .A3(n7286), .ZN(n7293) );
  NAND2_X1 U9060 ( .A1(n12929), .A2(n9526), .ZN(n9539) );
  NAND2_X1 U9061 ( .A1(n9572), .A2(n6591), .ZN(n9601) );
  NAND4_X2 U9062 ( .A1(n9051), .A2(n9050), .A3(n9163), .A4(n9049), .ZN(n7345)
         );
  INV_X1 U9063 ( .A(n11067), .ZN(n11069) );
  NAND2_X1 U9064 ( .A1(n8568), .A2(n8151), .ZN(n6789) );
  NAND2_X1 U9065 ( .A1(n6789), .A2(n8153), .ZN(n8556) );
  NAND2_X1 U9066 ( .A1(n7738), .A2(n7737), .ZN(n7753) );
  NAND2_X1 U9067 ( .A1(n6876), .A2(n12451), .ZN(n6875) );
  NAND2_X1 U9068 ( .A1(n7478), .A2(n7477), .ZN(n7497) );
  NAND2_X1 U9069 ( .A1(n7499), .A2(n7498), .ZN(n7516) );
  NAND2_X1 U9070 ( .A1(n7696), .A2(n7695), .ZN(n7698) );
  AOI21_X1 U9071 ( .B1(n7929), .B2(n7928), .A(n7927), .ZN(n7930) );
  AOI21_X1 U9072 ( .B1(n7852), .B2(n6876), .A(n6874), .ZN(n6873) );
  NAND2_X1 U9073 ( .A1(n7556), .A2(n7555), .ZN(n7558) );
  OAI21_X2 U9074 ( .B1(n7799), .B2(n7798), .A(n7800), .ZN(n7811) );
  NAND2_X1 U9075 ( .A1(n12472), .A2(n12456), .ZN(n12458) );
  AOI21_X1 U9076 ( .B1(n6629), .B2(n6639), .A(n6634), .ZN(n6628) );
  NOR2_X1 U9077 ( .A1(n10434), .A2(n6630), .ZN(n6629) );
  NAND3_X1 U9078 ( .A1(n7113), .A2(n6638), .A3(n7111), .ZN(n6632) );
  NAND2_X1 U9079 ( .A1(n10434), .A2(n7115), .ZN(n7113) );
  OAI21_X1 U9080 ( .B1(n6637), .B2(n6636), .A(n11046), .ZN(n11053) );
  INV_X1 U9081 ( .A(n7113), .ZN(n6636) );
  NOR2_X1 U9082 ( .A1(n10476), .A2(n11046), .ZN(n6638) );
  NOR2_X1 U9083 ( .A1(n12260), .A2(n6568), .ZN(n12277) );
  NAND3_X1 U9084 ( .A1(n6642), .A2(n6644), .A3(n6640), .ZN(n12261) );
  NAND3_X1 U9085 ( .A1(n6642), .A2(n6641), .A3(n6640), .ZN(n6645) );
  INV_X1 U9086 ( .A(n6645), .ZN(n12279) );
  MUX2_X1 U9087 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n15096), .S(n6646), .Z(n10547) );
  INV_X2 U9088 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6649) );
  NAND3_X1 U9089 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7454), .A3(
        P3_IR_REG_2__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U9090 ( .A1(n6443), .A2(n11474), .ZN(n6656) );
  NAND2_X1 U9091 ( .A1(n6654), .A2(n6652), .ZN(n11058) );
  AND2_X1 U9092 ( .A1(n6653), .A2(n6655), .ZN(n6652) );
  NAND2_X1 U9093 ( .A1(n14783), .A2(n11474), .ZN(n6654) );
  INV_X1 U9094 ( .A(n6657), .ZN(n11473) );
  NAND2_X1 U9095 ( .A1(n10545), .A2(n6671), .ZN(n6672) );
  NAND2_X1 U9096 ( .A1(n6666), .A2(n10444), .ZN(n6670) );
  NAND2_X1 U9097 ( .A1(n10545), .A2(n10429), .ZN(n6666) );
  NOR2_X1 U9098 ( .A1(n10444), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6669) );
  AND2_X1 U9099 ( .A1(n9677), .A2(n6477), .ZN(n6674) );
  NAND2_X1 U9100 ( .A1(n6676), .A2(n12558), .ZN(n12191) );
  NAND2_X1 U9101 ( .A1(n6676), .A2(n6487), .ZN(n6675) );
  INV_X1 U9102 ( .A(n12190), .ZN(n6676) );
  NAND2_X1 U9103 ( .A1(n9676), .A2(n9677), .ZN(n12190) );
  NAND2_X1 U9104 ( .A1(n11684), .A2(n6680), .ZN(n6679) );
  NAND2_X1 U9105 ( .A1(n6679), .A2(n6677), .ZN(n9659) );
  OAI21_X1 U9106 ( .B1(n12132), .B2(n6689), .A(n6687), .ZN(n9692) );
  NAND2_X1 U9107 ( .A1(n6687), .A2(n6689), .ZN(n6685) );
  NAND2_X1 U9108 ( .A1(n12132), .A2(n6687), .ZN(n6686) );
  AOI21_X1 U9109 ( .B1(n12228), .B2(n6688), .A(n9689), .ZN(n6687) );
  INV_X1 U9110 ( .A(n9687), .ZN(n6688) );
  INV_X1 U9111 ( .A(n12228), .ZN(n6689) );
  NAND2_X1 U9112 ( .A1(n12226), .A2(n12228), .ZN(n12227) );
  NAND2_X1 U9113 ( .A1(n12132), .A2(n9687), .ZN(n12226) );
  NAND3_X1 U9114 ( .A1(n6959), .A2(n6690), .A3(n6958), .ZN(n6692) );
  NAND3_X1 U9115 ( .A1(n6959), .A2(n6958), .A3(n6961), .ZN(n10892) );
  INV_X1 U9116 ( .A(n6692), .ZN(n10891) );
  NAND2_X2 U9117 ( .A1(n7411), .A2(n7410), .ZN(n7932) );
  NAND2_X1 U9118 ( .A1(n6701), .A2(n6702), .ZN(n14634) );
  NAND2_X1 U9119 ( .A1(n14620), .A2(n6543), .ZN(n6701) );
  OAI21_X1 U9120 ( .B1(n10164), .B2(n6717), .A(n6714), .ZN(n13018) );
  MUX2_X1 U9121 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9112), .S(n12985), .Z(n12982) );
  XNOR2_X1 U9122 ( .A(n6729), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  INV_X1 U9123 ( .A(n14205), .ZN(n6731) );
  INV_X1 U9124 ( .A(n14264), .ZN(n6734) );
  NAND2_X1 U9125 ( .A1(n6526), .A2(n14223), .ZN(n6737) );
  AOI21_X1 U9126 ( .B1(n14217), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6741), .ZN(
        n6744) );
  NAND2_X1 U9127 ( .A1(n6742), .A2(n6745), .ZN(n6741) );
  NAND2_X1 U9128 ( .A1(n9013), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6742) );
  NOR2_X1 U9129 ( .A1(n14217), .A2(n9013), .ZN(n9015) );
  NOR2_X1 U9130 ( .A1(n9013), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6747) );
  INV_X1 U9131 ( .A(n14217), .ZN(n6748) );
  NOR2_X1 U9132 ( .A1(n15171), .A2(n15172), .ZN(n15170) );
  NAND2_X1 U9133 ( .A1(n15169), .A2(n15168), .ZN(n15167) );
  XNOR2_X1 U9134 ( .A(n9001), .B(n6750), .ZN(n15169) );
  OR2_X1 U9135 ( .A1(n12344), .A2(n12740), .ZN(n6753) );
  NAND2_X1 U9136 ( .A1(n12325), .A2(n12324), .ZN(n12343) );
  OAI22_X1 U9137 ( .A1(n12323), .A2(n12744), .B1(n6851), .B2(n12322), .ZN(
        n12325) );
  NAND2_X2 U9138 ( .A1(n7322), .A2(n9048), .ZN(n9162) );
  AND3_X2 U9139 ( .A1(n9074), .A2(n9075), .A3(n9057), .ZN(n9062) );
  NAND2_X1 U9140 ( .A1(n11388), .A2(n6772), .ZN(n13236) );
  INV_X1 U9141 ( .A(n6776), .ZN(n13235) );
  MUX2_X1 U9142 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9737), .Z(n8144) );
  OAI21_X2 U9143 ( .B1(n8668), .B2(n10886), .A(n8224), .ZN(n8225) );
  NAND2_X1 U9144 ( .A1(n8668), .A2(n8224), .ZN(n6785) );
  NAND2_X1 U9145 ( .A1(n8450), .A2(n6437), .ZN(n6797) );
  NAND2_X1 U9146 ( .A1(n6797), .A2(n6798), .ZN(n8177) );
  INV_X1 U9147 ( .A(n10561), .ZN(n6818) );
  OR2_X1 U9148 ( .A1(n6827), .A2(n6824), .ZN(n6822) );
  NAND3_X1 U9149 ( .A1(n6827), .A2(n6826), .A3(n6824), .ZN(n6823) );
  INV_X1 U9150 ( .A(n10502), .ZN(n6824) );
  NAND2_X1 U9151 ( .A1(n11538), .A2(n6829), .ZN(n6828) );
  OAI21_X1 U9152 ( .B1(n14780), .B2(n6843), .A(n6842), .ZN(n14804) );
  NAND2_X1 U9153 ( .A1(n6841), .A2(n6839), .ZN(n14802) );
  NAND2_X1 U9154 ( .A1(n14780), .A2(n6842), .ZN(n6841) );
  NAND4_X1 U9155 ( .A1(n6857), .A2(n6855), .A3(n6554), .A4(n6854), .ZN(n8116)
         );
  NAND3_X1 U9156 ( .A1(n6622), .A2(n6858), .A3(n7431), .ZN(n6857) );
  XNOR2_X1 U9157 ( .A(n6859), .B(n12391), .ZN(n12401) );
  XNOR2_X1 U9158 ( .A(n12386), .B(n14230), .ZN(n12369) );
  XNOR2_X2 U9159 ( .A(n6860), .B(n8256), .ZN(n8937) );
  NAND3_X1 U9160 ( .A1(n8250), .A2(n8252), .A3(n7390), .ZN(n6861) );
  AND3_X2 U9161 ( .A1(n7141), .A2(n6513), .A3(n8131), .ZN(n8250) );
  OR2_X2 U9162 ( .A1(n13868), .A2(n13844), .ZN(n13845) );
  NAND3_X1 U9163 ( .A1(n11614), .A2(n6862), .A3(n14245), .ZN(n14054) );
  INV_X1 U9164 ( .A(n6865), .ZN(n11615) );
  NOR2_X1 U9165 ( .A1(n14573), .A2(n6869), .ZN(n11132) );
  NAND2_X1 U9166 ( .A1(n7852), .A2(n8072), .ZN(n12493) );
  INV_X1 U9167 ( .A(n6873), .ZN(n12409) );
  OAI21_X1 U9168 ( .B1(n11399), .B2(n11644), .A(n6881), .ZN(n14835) );
  NAND2_X1 U9169 ( .A1(n6880), .A2(n6879), .ZN(n7550) );
  NAND2_X1 U9170 ( .A1(n11399), .A2(n6881), .ZN(n6879) );
  NAND2_X2 U9171 ( .A1(n10424), .A2(n9771), .ZN(n7758) );
  OAI22_X1 U9172 ( .A1(n7758), .A2(n9746), .B1(n10424), .B2(n10502), .ZN(n7455) );
  NAND3_X1 U9173 ( .A1(n6508), .A2(n7469), .A3(n7468), .ZN(n14885) );
  OAI21_X2 U9174 ( .B1(n11652), .B2(n7588), .A(n8001), .ZN(n14285) );
  OAI21_X2 U9175 ( .B1(n12672), .B2(n7694), .A(n7693), .ZN(n12625) );
  OAI21_X2 U9176 ( .B1(n14278), .B2(n7939), .A(n8017), .ZN(n12672) );
  XNOR2_X2 U9177 ( .A(n6897), .B(n9098), .ZN(n11773) );
  NAND3_X1 U9178 ( .A1(n7363), .A2(n9062), .A3(n7366), .ZN(n6898) );
  NAND2_X1 U9179 ( .A1(n10857), .A2(n10856), .ZN(n10859) );
  AND2_X1 U9180 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6904), .ZN(n9130) );
  OAI21_X1 U9181 ( .B1(n11001), .B2(n6908), .A(n6907), .ZN(n11067) );
  AOI21_X1 U9182 ( .B1(n13218), .B2(n6527), .A(n6912), .ZN(n13169) );
  NAND2_X1 U9183 ( .A1(n13627), .A2(n14532), .ZN(n10313) );
  AND3_X4 U9184 ( .A1(n8538), .A2(n6468), .A3(n6926), .ZN(n14532) );
  NAND2_X1 U9185 ( .A1(n10811), .A2(n6931), .ZN(n6928) );
  NAND2_X1 U9186 ( .A1(n6928), .A2(n6929), .ZN(n11130) );
  NAND2_X1 U9187 ( .A1(n11101), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U9188 ( .A1(n10795), .A2(n6937), .ZN(n6939) );
  NAND2_X1 U9189 ( .A1(n10795), .A2(n10796), .ZN(n10794) );
  NAND2_X1 U9190 ( .A1(n11608), .A2(n6529), .ZN(n11611) );
  NAND2_X2 U9191 ( .A1(n8269), .A2(n8260), .ZN(n8691) );
  XNOR2_X2 U9192 ( .A(n6957), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U9193 ( .A1(n9613), .A2(n14918), .ZN(n9617) );
  NAND2_X1 U9194 ( .A1(n6960), .A2(n10640), .ZN(n6959) );
  INV_X1 U9195 ( .A(n10633), .ZN(n6960) );
  NAND3_X1 U9196 ( .A1(n6965), .A2(n9607), .A3(n9606), .ZN(n9610) );
  NAND2_X1 U9197 ( .A1(n9604), .A2(n9605), .ZN(n9694) );
  INV_X1 U9198 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U9199 ( .A1(n9690), .A2(n6970), .ZN(n6968) );
  NAND2_X1 U9200 ( .A1(n6968), .A2(n6967), .ZN(P3_U3154) );
  NAND2_X1 U9201 ( .A1(n12083), .A2(n12164), .ZN(n6971) );
  NAND2_X1 U9202 ( .A1(n6971), .A2(n6972), .ZN(n12128) );
  NAND4_X1 U9203 ( .A1(n6986), .A2(n6478), .A3(n6987), .A4(n6985), .ZN(n7934)
         );
  NAND3_X1 U9204 ( .A1(n6478), .A2(n7560), .A3(n6988), .ZN(n7719) );
  NAND2_X1 U9205 ( .A1(n11340), .A2(n7398), .ZN(n11547) );
  NAND2_X1 U9206 ( .A1(n9670), .A2(n9669), .ZN(n12107) );
  OAI21_X1 U9207 ( .B1(n9624), .B2(n14890), .A(n12173), .ZN(n12150) );
  AOI21_X2 U9208 ( .B1(n12117), .B2(n9642), .A(n9641), .ZN(n11684) );
  NAND2_X1 U9209 ( .A1(n12107), .A2(n9671), .ZN(n9675) );
  NAND2_X1 U9210 ( .A1(n11342), .A2(n11341), .ZN(n11340) );
  AND2_X2 U9211 ( .A1(n8928), .A2(n8249), .ZN(n7390) );
  NAND2_X1 U9212 ( .A1(n10127), .A2(n10128), .ZN(n10144) );
  NAND2_X1 U9213 ( .A1(n13506), .A2(n6998), .ZN(n6995) );
  NAND2_X1 U9214 ( .A1(n6995), .A2(n6996), .ZN(n13558) );
  OAI21_X1 U9215 ( .B1(n11284), .B2(n7006), .A(n7003), .ZN(n13387) );
  NAND2_X1 U9216 ( .A1(n11284), .A2(n7003), .ZN(n7002) );
  NAND2_X1 U9217 ( .A1(n7007), .A2(n7009), .ZN(n13437) );
  NAND3_X1 U9218 ( .A1(n6445), .A2(n14411), .A3(n7017), .ZN(n7007) );
  NAND2_X1 U9219 ( .A1(n14411), .A2(n13416), .ZN(n14383) );
  INV_X1 U9220 ( .A(n10771), .ZN(n7019) );
  INV_X1 U9221 ( .A(n14372), .ZN(n7032) );
  AOI21_X2 U9222 ( .B1(n7032), .B2(n7035), .A(n7031), .ZN(n13415) );
  NAND2_X1 U9223 ( .A1(n10144), .A2(n10130), .ZN(n7038) );
  NAND2_X1 U9224 ( .A1(n10144), .A2(n10129), .ZN(n7039) );
  NAND3_X1 U9225 ( .A1(n7039), .A2(n7038), .A3(n7037), .ZN(n7041) );
  INV_X1 U9226 ( .A(n7041), .ZN(n10685) );
  INV_X2 U9227 ( .A(n10283), .ZN(n12978) );
  XNOR2_X2 U9228 ( .A(n10283), .B(n11784), .ZN(n11990) );
  AND2_X2 U9229 ( .A1(n7046), .A2(n9116), .ZN(n10283) );
  NAND2_X1 U9230 ( .A1(n13259), .A2(n7053), .ZN(n7047) );
  NAND2_X1 U9231 ( .A1(n13259), .A2(n13287), .ZN(n7058) );
  NAND2_X1 U9232 ( .A1(n7047), .A2(n6498), .ZN(P2_U3528) );
  INV_X4 U9233 ( .A(n9134), .ZN(n9433) );
  NAND2_X1 U9234 ( .A1(n9433), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U9235 ( .A1(n10822), .A2(n7059), .ZN(n7060) );
  NAND2_X1 U9236 ( .A1(n7060), .A2(n7061), .ZN(n10849) );
  NAND2_X1 U9237 ( .A1(n10852), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U9238 ( .A1(n13123), .A2(n7071), .ZN(n7070) );
  OAI21_X1 U9239 ( .B1(n13201), .B2(n7083), .A(n7080), .ZN(n13172) );
  OAI21_X1 U9240 ( .B1(n13201), .B2(n11751), .A(n11752), .ZN(n13186) );
  NAND2_X1 U9241 ( .A1(n11753), .A2(n7084), .ZN(n7083) );
  NAND2_X1 U9242 ( .A1(n13244), .A2(n7085), .ZN(n11750) );
  NOR2_X2 U9243 ( .A1(n14219), .A2(n14218), .ZN(n14217) );
  INV_X1 U9244 ( .A(n7089), .ZN(n9034) );
  NAND2_X1 U9245 ( .A1(n14473), .A2(n14474), .ZN(n14470) );
  AOI21_X1 U9246 ( .B1(n14467), .B2(n14468), .A(n7091), .ZN(n7090) );
  NOR2_X1 U9247 ( .A1(n14467), .A2(n14468), .ZN(n14466) );
  INV_X1 U9248 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U9249 ( .A1(n11522), .A2(n7102), .ZN(n7098) );
  NAND2_X1 U9250 ( .A1(n7098), .A2(n7097), .ZN(n12260) );
  NAND3_X1 U9251 ( .A1(n7101), .A2(n7100), .A3(n11520), .ZN(n7097) );
  INV_X1 U9252 ( .A(n12300), .ZN(n7107) );
  NAND2_X1 U9253 ( .A1(n7128), .A2(n7129), .ZN(n8828) );
  NAND2_X1 U9254 ( .A1(n8807), .A2(n7131), .ZN(n7128) );
  INV_X1 U9255 ( .A(n8361), .ZN(n7141) );
  NAND4_X1 U9256 ( .A1(n8125), .A2(n8123), .A3(n8124), .A4(n8421), .ZN(n8361)
         );
  NAND2_X1 U9257 ( .A1(n7142), .A2(n7143), .ZN(n8788) );
  NAND3_X1 U9258 ( .A1(n8782), .A2(n6539), .A3(n8781), .ZN(n7142) );
  OAI22_X1 U9259 ( .A1(n8795), .A2(n7145), .B1(n8796), .B2(n7144), .ZN(n8800)
         );
  NAND2_X1 U9260 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NAND2_X1 U9261 ( .A1(n7146), .A2(n7147), .ZN(n8917) );
  NAND3_X1 U9262 ( .A1(n8879), .A2(n6549), .A3(n8878), .ZN(n7146) );
  NAND2_X1 U9263 ( .A1(n7149), .A2(n7150), .ZN(n8777) );
  NAND3_X1 U9264 ( .A1(n8772), .A2(n6550), .A3(n8771), .ZN(n7149) );
  NAND2_X1 U9265 ( .A1(n7152), .A2(n7153), .ZN(n8863) );
  NAND3_X1 U9266 ( .A1(n8858), .A2(n6548), .A3(n8857), .ZN(n7152) );
  NAND2_X1 U9267 ( .A1(n7155), .A2(n7156), .ZN(n8845) );
  NAND3_X1 U9268 ( .A1(n8840), .A2(n6536), .A3(n8839), .ZN(n7155) );
  NAND2_X1 U9269 ( .A1(n7158), .A2(n7159), .ZN(n8767) );
  NAND3_X1 U9270 ( .A1(n8760), .A2(n6540), .A3(n8759), .ZN(n7158) );
  NAND2_X1 U9271 ( .A1(n7161), .A2(n7162), .ZN(n8874) );
  NAND3_X1 U9272 ( .A1(n8868), .A2(n6535), .A3(n8867), .ZN(n7161) );
  NAND2_X1 U9273 ( .A1(n7164), .A2(n7433), .ZN(n7464) );
  OAI21_X1 U9274 ( .B1(n7451), .B2(n7452), .A(n7164), .ZN(n7453) );
  NAND2_X1 U9275 ( .A1(n7451), .A2(n7452), .ZN(n7164) );
  INV_X1 U9276 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U9277 ( .A1(n7165), .A2(n8122), .ZN(P3_U3296) );
  NAND2_X1 U9278 ( .A1(n7166), .A2(n8101), .ZN(n7165) );
  INV_X1 U9279 ( .A(n8096), .ZN(n7167) );
  NAND2_X1 U9280 ( .A1(n8097), .A2(n9607), .ZN(n7168) );
  NAND2_X1 U9281 ( .A1(n7173), .A2(n7170), .ZN(n7169) );
  INV_X1 U9282 ( .A(n7769), .ZN(n7170) );
  INV_X1 U9283 ( .A(n7756), .ZN(n7172) );
  NAND2_X1 U9284 ( .A1(n7715), .A2(n7178), .ZN(n7174) );
  NAND2_X1 U9285 ( .A1(n7174), .A2(n7175), .ZN(n7738) );
  NAND2_X1 U9286 ( .A1(n7642), .A2(n7184), .ZN(n7181) );
  NAND2_X1 U9287 ( .A1(n7181), .A2(n7182), .ZN(n7696) );
  OAI21_X1 U9288 ( .B1(n7530), .B2(n7192), .A(n7190), .ZN(n7556) );
  OAI21_X1 U9289 ( .B1(n7530), .B2(n7529), .A(n7531), .ZN(n7547) );
  NAND2_X1 U9290 ( .A1(n7529), .A2(n7531), .ZN(n7194) );
  NAND2_X1 U9291 ( .A1(n7613), .A2(n6555), .ZN(n7197) );
  NAND2_X1 U9292 ( .A1(n7857), .A2(n7204), .ZN(n7200) );
  OAI21_X1 U9293 ( .B1(n7857), .B2(n7203), .A(n7201), .ZN(n7897) );
  NAND2_X1 U9294 ( .A1(n7857), .A2(n7856), .ZN(n7873) );
  INV_X1 U9295 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7206) );
  OAI21_X1 U9296 ( .B1(n13833), .B2(n7222), .A(n7221), .ZN(n13932) );
  NAND2_X2 U9297 ( .A1(n7220), .A2(n7219), .ZN(n13930) );
  NAND2_X1 U9298 ( .A1(n13833), .A2(n7221), .ZN(n7220) );
  NAND2_X1 U9299 ( .A1(n7234), .A2(n7232), .ZN(n10805) );
  NAND3_X1 U9300 ( .A1(n10793), .A2(n7235), .A3(n6439), .ZN(n7234) );
  OAI21_X1 U9301 ( .B1(n10793), .B2(n7236), .A(n7235), .ZN(n14563) );
  AND2_X1 U9302 ( .A1(n7238), .A2(n8250), .ZN(n8258) );
  NAND2_X1 U9303 ( .A1(n8250), .A2(n7239), .ZN(n14182) );
  XNOR2_X2 U9304 ( .A(n8223), .B(n8222), .ZN(n8668) );
  NAND2_X1 U9305 ( .A1(n8532), .A2(n8531), .ZN(n8138) );
  NAND2_X1 U9306 ( .A1(n8479), .A2(n8155), .ZN(n7259) );
  NAND2_X1 U9307 ( .A1(n8479), .A2(n6531), .ZN(n7256) );
  NAND2_X1 U9308 ( .A1(n8418), .A2(n7267), .ZN(n7264) );
  NAND2_X1 U9309 ( .A1(n7264), .A2(n7265), .ZN(n8405) );
  OAI21_X1 U9310 ( .B1(n8656), .B2(n7276), .A(n8226), .ZN(n8313) );
  AOI21_X1 U9311 ( .B1(n8226), .B2(n7273), .A(n7272), .ZN(n7271) );
  NAND3_X1 U9312 ( .A1(n11937), .A2(n11942), .A3(n11946), .ZN(n11943) );
  NAND2_X1 U9313 ( .A1(n7281), .A2(n7280), .ZN(n11953) );
  NAND2_X1 U9314 ( .A1(n10329), .A2(n7282), .ZN(n10330) );
  NAND2_X1 U9315 ( .A1(n12849), .A2(n7294), .ZN(n9465) );
  INV_X1 U9316 ( .A(n7293), .ZN(n12903) );
  NAND2_X1 U9317 ( .A1(n12823), .A2(n7297), .ZN(n7296) );
  NAND3_X1 U9318 ( .A1(n7304), .A2(n11992), .A3(n9932), .ZN(n7301) );
  NAND2_X2 U9319 ( .A1(n10917), .A2(n12028), .ZN(n9137) );
  NAND2_X1 U9320 ( .A1(n7309), .A2(n6533), .ZN(n12931) );
  NAND2_X1 U9321 ( .A1(n12863), .A2(n7316), .ZN(n7313) );
  NAND2_X1 U9322 ( .A1(n7313), .A2(n7314), .ZN(n12843) );
  NOR2_X2 U9323 ( .A1(n7320), .A2(n7345), .ZN(n9250) );
  NAND2_X1 U9324 ( .A1(n12464), .A2(n12463), .ZN(n12683) );
  NAND2_X1 U9325 ( .A1(n14824), .A2(n7327), .ZN(n7325) );
  NAND2_X1 U9326 ( .A1(n7325), .A2(n7326), .ZN(n14286) );
  NAND2_X1 U9327 ( .A1(n7332), .A2(n7330), .ZN(n12437) );
  NAND4_X1 U9328 ( .A1(n7403), .A2(n6649), .A3(n7333), .A4(n6758), .ZN(n7479)
         );
  NAND2_X1 U9329 ( .A1(n11402), .A2(n11311), .ZN(n11645) );
  NAND2_X1 U9330 ( .A1(n12455), .A2(n12454), .ZN(n12471) );
  NAND2_X1 U9331 ( .A1(n12455), .A2(n7336), .ZN(n12472) );
  NAND2_X1 U9332 ( .A1(n12422), .A2(n12664), .ZN(n7341) );
  NOR2_X1 U9333 ( .A1(n7932), .A2(n7413), .ZN(n8105) );
  NAND4_X2 U9334 ( .A1(n9117), .A2(n9118), .A3(n9120), .A4(n9119), .ZN(n12979)
         );
  NAND2_X1 U9335 ( .A1(n12979), .A2(n7346), .ZN(n11782) );
  INV_X2 U9336 ( .A(n11797), .ZN(n7348) );
  NAND2_X1 U9337 ( .A1(n7349), .A2(n7350), .ZN(n11800) );
  OR2_X1 U9338 ( .A1(n11795), .A2(n7351), .ZN(n7350) );
  NAND2_X1 U9339 ( .A1(n7355), .A2(n7356), .ZN(n11861) );
  NAND3_X1 U9340 ( .A1(n11855), .A2(n6542), .A3(n11854), .ZN(n7355) );
  NAND2_X1 U9341 ( .A1(n7357), .A2(n6544), .ZN(n11837) );
  NAND3_X1 U9342 ( .A1(n11830), .A2(n6551), .A3(n11829), .ZN(n7357) );
  NAND2_X1 U9343 ( .A1(n7359), .A2(n6545), .ZN(n11825) );
  NAND3_X1 U9344 ( .A1(n11818), .A2(n6541), .A3(n11817), .ZN(n7359) );
  NAND2_X1 U9345 ( .A1(n7361), .A2(n6546), .ZN(n11850) );
  NAND3_X1 U9346 ( .A1(n11842), .A2(n6552), .A3(n11841), .ZN(n7361) );
  NOR2_X1 U9347 ( .A1(n9162), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7363) );
  NAND3_X1 U9348 ( .A1(n7366), .A2(n9062), .A3(n7364), .ZN(n13360) );
  NAND2_X1 U9349 ( .A1(n7367), .A2(n7368), .ZN(n11917) );
  NAND3_X1 U9350 ( .A1(n11912), .A2(n6547), .A3(n11911), .ZN(n7367) );
  NAND2_X1 U9351 ( .A1(n7370), .A2(n7371), .ZN(n11907) );
  NAND3_X1 U9352 ( .A1(n11901), .A2(n6537), .A3(n11900), .ZN(n7370) );
  NAND2_X1 U9353 ( .A1(n7372), .A2(n7374), .ZN(n11813) );
  NAND3_X1 U9354 ( .A1(n11805), .A2(n11804), .A3(n7373), .ZN(n7372) );
  AOI21_X1 U9355 ( .B1(n13628), .B2(n10123), .A(n10032), .ZN(n10036) );
  INV_X1 U9356 ( .A(n13790), .ZN(n14068) );
  NAND2_X1 U9357 ( .A1(n7825), .A2(n7815), .ZN(n7824) );
  NAND2_X1 U9358 ( .A1(n7637), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9359 ( .A1(n9069), .A2(n9068), .ZN(n9969) );
  NOR2_X1 U9360 ( .A1(n8691), .A2(n9830), .ZN(n8515) );
  NAND2_X1 U9361 ( .A1(n7639), .A2(n7638), .ZN(n7642) );
  NAND2_X1 U9362 ( .A1(n7624), .A2(n10055), .ZN(n7638) );
  NAND2_X1 U9363 ( .A1(n9127), .A2(n9126), .ZN(n10270) );
  NAND2_X1 U9364 ( .A1(n7577), .A2(n7576), .ZN(n7579) );
  NAND2_X1 U9365 ( .A1(n7597), .A2(n7596), .ZN(n7599) );
  INV_X1 U9366 ( .A(n9793), .ZN(n8934) );
  NAND4_X2 U9367 ( .A1(n9142), .A2(n9141), .A3(n9140), .A4(n9139), .ZN(n12977)
         );
  INV_X1 U9368 ( .A(n10185), .ZN(n11991) );
  NAND2_X1 U9369 ( .A1(n7894), .A2(n8086), .ZN(n7929) );
  NAND2_X1 U9370 ( .A1(n9509), .A2(n9508), .ZN(n12863) );
  NAND2_X1 U9371 ( .A1(n7811), .A2(n7810), .ZN(n7813) );
  AND2_X1 U9372 ( .A1(n12038), .A2(n9932), .ZN(n11968) );
  NOR2_X1 U9373 ( .A1(n14761), .A2(n9932), .ZN(n9592) );
  AND2_X1 U9374 ( .A1(n9932), .A2(n12040), .ZN(n9954) );
  NAND2_X1 U9375 ( .A1(n7836), .A2(n7835), .ZN(n7838) );
  NAND2_X1 U9376 ( .A1(n13074), .A2(n11760), .ZN(n11762) );
  NAND2_X1 U9377 ( .A1(n9539), .A2(n9538), .ZN(n9572) );
  AND2_X1 U9378 ( .A1(n9121), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7451) );
  NAND4_X2 U9379 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n12975)
         );
  INV_X1 U9380 ( .A(n9379), .ZN(n9394) );
  OR2_X1 U9381 ( .A1(n13415), .A2(n13414), .ZN(n13416) );
  INV_X1 U9382 ( .A(n11730), .ZN(n11962) );
  INV_X1 U9383 ( .A(n7925), .ZN(n12754) );
  AND2_X1 U9384 ( .A1(n13877), .A2(n13876), .ZN(n13879) );
  INV_X1 U9385 ( .A(n8260), .ZN(n8270) );
  NAND2_X1 U9386 ( .A1(n9077), .A2(n9078), .ZN(n9086) );
  OAI21_X1 U9387 ( .B1(n10805), .B2(n10810), .A(n10804), .ZN(n10809) );
  OR2_X1 U9388 ( .A1(n6477), .A2(n9677), .ZN(n9678) );
  NOR2_X1 U9389 ( .A1(n12259), .A2(n10668), .ZN(n7940) );
  XNOR2_X1 U9390 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7452) );
  INV_X1 U9391 ( .A(n7420), .ZN(n7421) );
  INV_X1 U9392 ( .A(n14914), .ZN(n7968) );
  OAI211_X2 U9393 ( .C1(n9148), .C2(n9977), .A(n9136), .B(n9135), .ZN(n11793)
         );
  CLKBUF_X1 U9394 ( .A(n14866), .Z(n14868) );
  CLKBUF_X1 U9395 ( .A(n11645), .Z(n11312) );
  OR2_X1 U9396 ( .A1(n7428), .A2(n8112), .ZN(n7417) );
  INV_X1 U9397 ( .A(n14893), .ZN(n11301) );
  INV_X1 U9398 ( .A(n8026), .ZN(n7692) );
  NOR2_X1 U9399 ( .A1(n9653), .A2(n12141), .ZN(n7377) );
  AND2_X1 U9400 ( .A1(n7654), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7378) );
  OR2_X1 U9401 ( .A1(n11492), .A2(n13617), .ZN(n7379) );
  OR2_X1 U9402 ( .A1(n11719), .A2(n13206), .ZN(n7381) );
  NOR2_X1 U9403 ( .A1(n12634), .A2(n12640), .ZN(n7382) );
  AND2_X1 U9404 ( .A1(n12692), .A2(n14972), .ZN(n7383) );
  AND2_X1 U9405 ( .A1(n11980), .A2(n11979), .ZN(n7384) );
  OR2_X1 U9406 ( .A1(n9481), .A2(n9480), .ZN(n7387) );
  AND2_X1 U9407 ( .A1(n9650), .A2(n12416), .ZN(n7388) );
  AND2_X1 U9408 ( .A1(n9066), .A2(n9065), .ZN(n7389) );
  NAND2_X1 U9409 ( .A1(n9931), .A2(n12038), .ZN(n14764) );
  INV_X1 U9410 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8707) );
  AND2_X1 U9411 ( .A1(n8539), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7391) );
  INV_X1 U9412 ( .A(n12523), .ZN(n7823) );
  AND2_X1 U9413 ( .A1(n8195), .A2(n8194), .ZN(n7392) );
  AND2_X1 U9414 ( .A1(n8176), .A2(n8175), .ZN(n7393) );
  AND2_X1 U9415 ( .A1(n10121), .A2(n13395), .ZN(n7394) );
  INV_X1 U9416 ( .A(n9125), .ZN(n9126) );
  AND2_X1 U9417 ( .A1(n11672), .A2(n14292), .ZN(n7395) );
  INV_X1 U9418 ( .A(P3_U3897), .ZN(n12258) );
  AND2_X1 U9419 ( .A1(n8183), .A2(n8182), .ZN(n7396) );
  INV_X1 U9420 ( .A(n13851), .ZN(n13880) );
  INV_X1 U9421 ( .A(n8117), .ZN(n10437) );
  INV_X1 U9422 ( .A(n12525), .ZN(n12547) );
  AND2_X1 U9423 ( .A1(n7809), .A2(n7808), .ZN(n12525) );
  INV_X1 U9424 ( .A(n13282), .ZN(n12016) );
  OR2_X1 U9425 ( .A1(n13290), .A2(n12953), .ZN(n7397) );
  INV_X1 U9426 ( .A(n13924), .ZN(n13788) );
  INV_X1 U9427 ( .A(n11401), .ZN(n11310) );
  OR2_X1 U9428 ( .A1(n9631), .A2(n11647), .ZN(n7398) );
  AND4_X1 U9429 ( .A1(n9520), .A2(n9519), .A3(n9518), .A4(n9517), .ZN(n11929)
         );
  INV_X1 U9430 ( .A(n11929), .ZN(n12952) );
  INV_X1 U9431 ( .A(n13159), .ZN(n11763) );
  AND2_X1 U9432 ( .A1(n14112), .A2(n13934), .ZN(n7399) );
  AND2_X1 U9433 ( .A1(n13296), .A2(n12954), .ZN(n7400) );
  OAI21_X1 U9434 ( .B1(n11396), .B2(n11395), .A(n11394), .ZN(n11568) );
  NAND2_X1 U9435 ( .A1(n9938), .A2(n10824), .ZN(n14769) );
  OAI21_X1 U9436 ( .B1(n8733), .B2(n8729), .A(n8728), .ZN(n8742) );
  NAND2_X1 U9437 ( .A1(n8745), .A2(n8744), .ZN(n8751) );
  OAI21_X1 U9438 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8755) );
  MUX2_X1 U9439 ( .A(n12975), .B(n11806), .S(n11967), .Z(n11808) );
  INV_X1 U9440 ( .A(n11808), .ZN(n11809) );
  MUX2_X1 U9441 ( .A(n12974), .B(n11810), .S(n11797), .Z(n11811) );
  MUX2_X1 U9442 ( .A(n12972), .B(n14746), .S(n11967), .Z(n11823) );
  INV_X1 U9443 ( .A(n11832), .ZN(n11833) );
  MUX2_X1 U9444 ( .A(n12969), .B(n11834), .S(n11967), .Z(n11835) );
  MUX2_X1 U9445 ( .A(n12967), .B(n11847), .S(n11967), .Z(n11848) );
  OAI21_X1 U9446 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8802) );
  INV_X1 U9447 ( .A(n11857), .ZN(n11858) );
  MUX2_X1 U9448 ( .A(n12965), .B(n14339), .S(n11967), .Z(n11859) );
  MUX2_X1 U9449 ( .A(n12963), .B(n14332), .S(n11967), .Z(n11874) );
  NAND2_X1 U9450 ( .A1(n11893), .A2(n11892), .ZN(n11896) );
  NAND2_X1 U9451 ( .A1(n8848), .A2(n8847), .ZN(n8849) );
  MUX2_X1 U9452 ( .A(n12957), .B(n13195), .S(n11967), .Z(n11905) );
  MUX2_X1 U9453 ( .A(n12955), .B(n13159), .S(n11967), .Z(n11915) );
  INV_X1 U9454 ( .A(n11948), .ZN(n11935) );
  NAND2_X1 U9455 ( .A1(n11936), .A2(n11935), .ZN(n11937) );
  NAND2_X1 U9456 ( .A1(n11941), .A2(n11940), .ZN(n11942) );
  OR2_X1 U9457 ( .A1(n12427), .A2(n12426), .ZN(n12428) );
  AND2_X1 U9458 ( .A1(n7937), .A2(n7925), .ZN(n7926) );
  INV_X1 U9459 ( .A(n14854), .ZN(n11306) );
  NOR2_X1 U9460 ( .A1(n10038), .A2(n14476), .ZN(n10040) );
  INV_X1 U9461 ( .A(n13412), .ZN(n11614) );
  INV_X1 U9462 ( .A(n10355), .ZN(n8525) );
  INV_X1 U9463 ( .A(n11098), .ZN(n10806) );
  INV_X1 U9464 ( .A(n8344), .ZN(n8215) );
  INV_X1 U9465 ( .A(n9674), .ZN(n9672) );
  OR2_X1 U9466 ( .A1(n8092), .A2(n7926), .ZN(n7927) );
  INV_X1 U9467 ( .A(n14821), .ZN(n11649) );
  AND2_X1 U9468 ( .A1(n9496), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9513) );
  NOR2_X1 U9469 ( .A1(n9385), .A2(n9091), .ZN(n9386) );
  NAND2_X1 U9470 ( .A1(n13282), .A2(n12952), .ZN(n11726) );
  INV_X1 U9471 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15122) );
  INV_X1 U9472 ( .A(n14332), .ZN(n11387) );
  INV_X1 U9473 ( .A(n11388), .ZN(n11389) );
  INV_X1 U9474 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U9475 ( .A1(n10034), .A2(n10033), .ZN(n10124) );
  NOR2_X1 U9476 ( .A1(n10040), .A2(n10039), .ZN(n10041) );
  AND2_X1 U9477 ( .A1(n14399), .A2(n14400), .ZN(n13403) );
  AND2_X1 U9478 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  AND2_X1 U9479 ( .A1(n8208), .A2(n8637), .ZN(n8209) );
  INV_X1 U9480 ( .A(SI_17_), .ZN(n8197) );
  INV_X1 U9481 ( .A(SI_11_), .ZN(n8168) );
  NAND2_X1 U9482 ( .A1(n12257), .A2(n10644), .ZN(n7969) );
  OR2_X1 U9483 ( .A1(n9634), .A2(n14290), .ZN(n9635) );
  OR2_X1 U9484 ( .A1(n7761), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7776) );
  NOR2_X1 U9485 ( .A1(n10564), .A2(n10563), .ZN(n10562) );
  NOR2_X1 U9486 ( .A1(n12485), .A2(n14915), .ZN(n12488) );
  INV_X1 U9487 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7489) );
  INV_X1 U9488 ( .A(n7455), .ZN(n7457) );
  INV_X1 U9489 ( .A(n9524), .ZN(n9525) );
  INV_X1 U9490 ( .A(n11986), .ZN(n11987) );
  NOR2_X1 U9491 ( .A1(n9442), .A2(n9093), .ZN(n9457) );
  AND2_X1 U9492 ( .A1(n9386), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9398) );
  INV_X1 U9493 ( .A(n12006), .ZN(n11068) );
  OR2_X1 U9494 ( .A1(n9218), .A2(n9217), .ZN(n9257) );
  INV_X1 U9495 ( .A(n14764), .ZN(n13261) );
  OR2_X1 U9496 ( .A1(n9305), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n9307) );
  INV_X1 U9497 ( .A(n13552), .ZN(n13456) );
  AND2_X1 U9498 ( .A1(n11497), .A2(n11498), .ZN(n11496) );
  INV_X1 U9499 ( .A(n10689), .ZN(n13537) );
  NAND2_X1 U9500 ( .A1(n8910), .A2(n7385), .ZN(n8911) );
  INV_X1 U9501 ( .A(n8349), .ZN(n8328) );
  INV_X1 U9502 ( .A(n8539), .ZN(n8268) );
  INV_X1 U9503 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9882) );
  NOR2_X1 U9504 ( .A1(n13881), .A2(n13949), .ZN(n13882) );
  INV_X1 U9505 ( .A(n13974), .ZN(n13832) );
  OR2_X1 U9506 ( .A1(n8487), .A2(n8271), .ZN(n8608) );
  NAND2_X1 U9507 ( .A1(n10310), .A2(n10309), .ZN(n10354) );
  AND2_X1 U9508 ( .A1(n8189), .A2(n8378), .ZN(n8190) );
  NAND2_X1 U9509 ( .A1(n8178), .A2(n9752), .ZN(n8133) );
  INV_X1 U9510 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8955) );
  OR2_X1 U9511 ( .A1(n7523), .A2(n7522), .ZN(n7538) );
  INV_X1 U9512 ( .A(n12668), .ZN(n9644) );
  NAND2_X1 U9513 ( .A1(n7746), .A2(n7745), .ZN(n7761) );
  OR2_X1 U9514 ( .A1(n12064), .A2(n14840), .ZN(n9629) );
  INV_X1 U9515 ( .A(n12575), .ZN(n9667) );
  AND2_X1 U9516 ( .A1(n9687), .A2(n9685), .ZN(n12130) );
  OR2_X1 U9517 ( .A1(n7801), .A2(n7788), .ZN(n7789) );
  INV_X1 U9518 ( .A(n11520), .ZN(n11522) );
  NAND2_X1 U9519 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  INV_X1 U9520 ( .A(n12390), .ZN(n12391) );
  NAND2_X1 U9521 ( .A1(n7805), .A2(n7804), .ZN(n7819) );
  INV_X1 U9522 ( .A(n12572), .ZN(n12568) );
  NAND2_X1 U9523 ( .A1(n7590), .A2(n7589), .ZN(n7605) );
  INV_X1 U9524 ( .A(n12392), .ZN(n10617) );
  OR2_X1 U9525 ( .A1(n7801), .A2(n12819), .ZN(n7876) );
  OR2_X1 U9526 ( .A1(n7801), .A2(n11431), .ZN(n7841) );
  INV_X1 U9527 ( .A(n12252), .ZN(n11672) );
  NAND2_X1 U9528 ( .A1(n9523), .A2(n9525), .ZN(n9526) );
  OR2_X1 U9529 ( .A1(n9426), .A2(n9425), .ZN(n9442) );
  INV_X1 U9530 ( .A(n12862), .ZN(n9508) );
  INV_X1 U9531 ( .A(n12898), .ZN(n12940) );
  AND2_X1 U9532 ( .A1(n9457), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9468) );
  OR2_X1 U9533 ( .A1(n9350), .A2(n11661), .ZN(n9385) );
  INV_X1 U9534 ( .A(n12019), .ZN(n11761) );
  OR2_X1 U9535 ( .A1(n9593), .A2(n9592), .ZN(n9943) );
  AND2_X1 U9536 ( .A1(n9548), .A2(n9552), .ZN(n14717) );
  INV_X1 U9537 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U9538 ( .A1(n9307), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9346) );
  INV_X1 U9539 ( .A(n13619), .ZN(n11366) );
  INV_X1 U9540 ( .A(n13521), .ZN(n13442) );
  INV_X1 U9541 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8428) );
  OR2_X1 U9542 ( .A1(n10302), .A2(n10303), .ZN(n10048) );
  NOR2_X1 U9543 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  NOR2_X1 U9544 ( .A1(n8647), .A2(n13584), .ZN(n8348) );
  INV_X1 U9545 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13659) );
  INV_X1 U9546 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U9547 ( .A1(n13985), .A2(n13809), .ZN(n13975) );
  INV_X1 U9548 ( .A(n14005), .ZN(n14017) );
  INV_X1 U9549 ( .A(n14141), .ZN(n14045) );
  INV_X1 U9550 ( .A(n13782), .ZN(n11138) );
  INV_X1 U9551 ( .A(n14576), .ZN(n10321) );
  AND2_X1 U9552 ( .A1(n10304), .A2(n10303), .ZN(n10347) );
  NAND2_X1 U9553 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  INV_X1 U9554 ( .A(n10689), .ZN(n13395) );
  AND2_X1 U9555 ( .A1(n8201), .A2(n8200), .ZN(n8394) );
  AOI22_X1 U9556 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n8955), .B1(n9011), .B2(
        n8954), .ZN(n8957) );
  OAI21_X1 U9557 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n8972), .A(n8971), .ZN(
        n8976) );
  OAI21_X1 U9558 ( .B1(n12762), .B2(n12245), .A(n9730), .ZN(n9731) );
  AOI21_X1 U9559 ( .B1(n12480), .B2(n7886), .A(n7882), .ZN(n12485) );
  AND4_X1 U9560 ( .A1(n7731), .A2(n7730), .A3(n7729), .A4(n7728), .ZN(n12622)
         );
  INV_X1 U9561 ( .A(n12399), .ZN(n14809) );
  AND2_X1 U9562 ( .A1(n10345), .A2(n10617), .ZN(n12684) );
  NAND2_X1 U9563 ( .A1(n10626), .A2(n10533), .ZN(n11176) );
  AND2_X1 U9564 ( .A1(n10526), .A2(n10525), .ZN(n10626) );
  INV_X1 U9565 ( .A(n14955), .ZN(n14966) );
  NOR2_X1 U9566 ( .A1(n10091), .A2(n12803), .ZN(n10093) );
  OR2_X1 U9567 ( .A1(n9694), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9696) );
  INV_X1 U9568 ( .A(n11474), .ZN(n11057) );
  OAI21_X1 U9569 ( .B1(n13092), .B2(n12924), .A(n9598), .ZN(n9599) );
  AND2_X1 U9570 ( .A1(n14764), .A2(n9570), .ZN(n9571) );
  INV_X1 U9571 ( .A(n9530), .ZN(n11966) );
  AND4_X1 U9572 ( .A1(n9586), .A2(n9585), .A3(n9584), .A4(n9583), .ZN(n11933)
         );
  INV_X1 U9573 ( .A(n14700), .ZN(n14683) );
  AND2_X1 U9574 ( .A1(n14616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14694) );
  INV_X1 U9575 ( .A(n12011), .ZN(n11744) );
  INV_X1 U9576 ( .A(n13115), .ZN(n13199) );
  INV_X1 U9577 ( .A(n14721), .ZN(n9945) );
  INV_X1 U9578 ( .A(n13287), .ZN(n14749) );
  NOR2_X1 U9579 ( .A1(n9944), .A2(n9937), .ZN(n10824) );
  AND2_X1 U9580 ( .A1(n9568), .A2(n9567), .ZN(n9944) );
  OR2_X1 U9581 ( .A1(n8592), .A2(n10016), .ZN(n8594) );
  OR2_X1 U9582 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  AND2_X1 U9583 ( .A1(n14369), .A2(n14588), .ZN(n14407) );
  AND2_X1 U9584 ( .A1(n8373), .A2(n8372), .ZN(n13568) );
  NAND2_X1 U9585 ( .A1(n8625), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8528) );
  INV_X1 U9586 ( .A(n14522), .ZN(n14486) );
  INV_X1 U9587 ( .A(n14524), .ZN(n14494) );
  NAND2_X1 U9588 ( .A1(n10306), .A2(n10305), .ZN(n15144) );
  INV_X1 U9589 ( .A(n14260), .ZN(n15149) );
  AND2_X1 U9590 ( .A1(n10347), .A2(n13782), .ZN(n14247) );
  NAND2_X1 U9591 ( .A1(n9914), .A2(n9913), .ZN(n10303) );
  INV_X1 U9592 ( .A(n14554), .ZN(n14571) );
  NAND2_X1 U9593 ( .A1(n13395), .A2(n9917), .ZN(n14578) );
  INV_X1 U9594 ( .A(n14592), .ZN(n14588) );
  AND2_X1 U9595 ( .A1(n10038), .A2(n9797), .ZN(n10306) );
  AND2_X1 U9596 ( .A1(n10456), .A2(n10455), .ZN(n14799) );
  INV_X1 U9597 ( .A(n12229), .ZN(n12237) );
  NAND2_X1 U9598 ( .A1(n9717), .A2(n9716), .ZN(n12245) );
  INV_X1 U9599 ( .A(n12502), .ZN(n12452) );
  INV_X1 U9600 ( .A(n12622), .ZN(n12589) );
  INV_X1 U9601 ( .A(n14799), .ZN(n14797) );
  OR2_X1 U9602 ( .A1(n10438), .A2(n10436), .ZN(n14815) );
  NAND2_X1 U9603 ( .A1(n14902), .A2(n14907), .ZN(n12677) );
  AND2_X1 U9604 ( .A1(n12591), .A2(n12590), .ZN(n12727) );
  AND2_X1 U9605 ( .A1(n12670), .A2(n12669), .ZN(n12748) );
  OR2_X1 U9606 ( .A1(n11176), .A2(n12684), .ZN(n12466) );
  NAND2_X1 U9607 ( .A1(n11176), .A2(n14910), .ZN(n14927) );
  INV_X1 U9608 ( .A(n14993), .ZN(n14990) );
  INV_X1 U9609 ( .A(n12415), .ZN(n12801) );
  INV_X1 U9610 ( .A(n12278), .ZN(n14216) );
  INV_X1 U9611 ( .A(n14227), .ZN(n12821) );
  INV_X1 U9612 ( .A(n12911), .ZN(n12924) );
  INV_X1 U9613 ( .A(n11951), .ZN(n12949) );
  INV_X1 U9614 ( .A(n14694), .ZN(n14658) );
  NAND2_X1 U9615 ( .A1(n14714), .A2(n13053), .ZN(n13197) );
  AND2_X1 U9616 ( .A1(n13171), .A2(n13170), .ZN(n13309) );
  INV_X1 U9617 ( .A(n14714), .ZN(n13253) );
  INV_X1 U9618 ( .A(n13183), .ZN(n13248) );
  NAND2_X1 U9619 ( .A1(n14723), .A2(n14718), .ZN(n14720) );
  AND2_X1 U9620 ( .A1(n9594), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14723) );
  INV_X1 U9621 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13376) );
  INV_X1 U9622 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10500) );
  INV_X1 U9623 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9824) );
  INV_X1 U9624 ( .A(n14120), .ZN(n13599) );
  INV_X1 U9625 ( .A(n14407), .ZN(n14419) );
  NAND2_X1 U9626 ( .A1(n10710), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14425) );
  INV_X1 U9627 ( .A(n13568), .ZN(n14021) );
  OR2_X1 U9628 ( .A1(n8393), .A2(n8392), .ZN(n14386) );
  OR2_X1 U9629 ( .A1(n14479), .A2(n9846), .ZN(n14520) );
  OR2_X1 U9630 ( .A1(n14479), .A2(n13642), .ZN(n14524) );
  AND2_X1 U9631 ( .A1(n13850), .A2(n15144), .ZN(n14042) );
  INV_X1 U9632 ( .A(n14247), .ZN(n13998) );
  INV_X1 U9633 ( .A(n15146), .ZN(n14258) );
  OR2_X1 U9634 ( .A1(n9924), .A2(n10303), .ZN(n14613) );
  OR2_X1 U9635 ( .A1(n9924), .A2(n9915), .ZN(n14599) );
  AND2_X1 U9636 ( .A1(n9793), .A2(n14194), .ZN(n10025) );
  INV_X1 U9637 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10203) );
  AND2_X1 U9638 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9956), .ZN(P2_U3947) );
  NOR2_X1 U9639 ( .A1(n10038), .A2(n9804), .ZN(P1_U4016) );
  NOR2_X2 U9640 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7406) );
  INV_X2 U9641 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7481) );
  NAND4_X1 U9642 ( .A1(n7406), .A2(n7405), .A3(n7481), .A4(n7404), .ZN(n7407)
         );
  NOR2_X1 U9643 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n7412) );
  NAND4_X1 U9644 ( .A1(n7412), .A2(n8102), .A3(n6993), .A4(n8109), .ZN(n7413)
         );
  INV_X1 U9645 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U9646 ( .A1(n7428), .A2(n7415), .ZN(n7418) );
  INV_X1 U9647 ( .A(n12062), .ZN(n7422) );
  AND2_X2 U9648 ( .A1(n7422), .A2(n7421), .ZN(n7488) );
  NAND2_X1 U9649 ( .A1(n7488), .A2(n14900), .ZN(n7426) );
  AND2_X2 U9650 ( .A1(n12062), .A2(n7420), .ZN(n7458) );
  NAND2_X1 U9651 ( .A1(n7458), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9652 ( .A1(n7671), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U9653 ( .A1(n7509), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7423) );
  INV_X1 U9654 ( .A(n7428), .ZN(n7429) );
  NAND2_X4 U9655 ( .A1(n8118), .A2(n8116), .ZN(n10424) );
  OR2_X1 U9656 ( .A1(n7816), .A2(SI_3_), .ZN(n7440) );
  INV_X2 U9657 ( .A(n8324), .ZN(n9771) );
  NAND2_X1 U9658 ( .A1(n9777), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7433) );
  XNOR2_X1 U9659 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7463) );
  NAND2_X1 U9660 ( .A1(n7464), .A2(n7463), .ZN(n7435) );
  NAND2_X1 U9661 ( .A1(n9779), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9662 ( .A1(n7435), .A2(n7434), .ZN(n7476) );
  XNOR2_X1 U9663 ( .A(n7476), .B(n7475), .ZN(n9763) );
  OR2_X1 U9664 ( .A1(n7758), .A2(n9763), .ZN(n7439) );
  NAND2_X1 U9665 ( .A1(n7436), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7437) );
  XNOR2_X1 U9666 ( .A(n7437), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10586) );
  OR2_X1 U9667 ( .A1(n10424), .A2(n10586), .ZN(n7438) );
  INV_X1 U9668 ( .A(n11302), .ZN(n14899) );
  NAND2_X1 U9669 ( .A1(n7458), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U9670 ( .A1(n7488), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U9671 ( .A1(n7671), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9672 ( .A1(n7509), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7441) );
  NAND4_X1 U9673 ( .A1(n7444), .A2(n7443), .A3(n7442), .A4(n7441), .ZN(n12259)
         );
  INV_X1 U9674 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15037) );
  INV_X1 U9675 ( .A(SI_0_), .ZN(n9741) );
  XNOR2_X1 U9676 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .ZN(n9740) );
  OAI211_X1 U9677 ( .C1(n15037), .C2(n10424), .A(n7446), .B(n7445), .ZN(n9612)
         );
  INV_X1 U9678 ( .A(n9612), .ZN(n10668) );
  NAND2_X1 U9679 ( .A1(n7458), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9680 ( .A1(n7509), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7449) );
  NAND2_X1 U9681 ( .A1(n7671), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7447) );
  INV_X1 U9682 ( .A(n7453), .ZN(n9746) );
  INV_X1 U9683 ( .A(n7465), .ZN(n7454) );
  INV_X1 U9684 ( .A(SI_1_), .ZN(n9745) );
  NAND2_X1 U9685 ( .A1(n7457), .A2(n7456), .ZN(n10517) );
  INV_X1 U9686 ( .A(n10517), .ZN(n10644) );
  NAND2_X1 U9687 ( .A1(n7940), .A2(n7969), .ZN(n9616) );
  NAND2_X1 U9688 ( .A1(n9616), .A2(n7966), .ZN(n14906) );
  NAND2_X1 U9689 ( .A1(n7488), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U9690 ( .A1(n7458), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9691 ( .A1(n7671), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U9692 ( .A1(n7509), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7459) );
  AND4_X2 U9693 ( .A1(n7462), .A2(n7461), .A3(n7460), .A4(n7459), .ZN(n11299)
         );
  INV_X1 U9694 ( .A(n11299), .ZN(n14891) );
  XNOR2_X1 U9695 ( .A(n7464), .B(n7463), .ZN(n9765) );
  OR2_X1 U9696 ( .A1(n7758), .A2(n9765), .ZN(n7469) );
  OR2_X1 U9697 ( .A1(n6434), .A2(SI_2_), .ZN(n7468) );
  INV_X1 U9698 ( .A(n7436), .ZN(n7466) );
  OR2_X1 U9699 ( .A1(n10424), .A2(n10557), .ZN(n7467) );
  NAND2_X1 U9700 ( .A1(n14906), .A2(n7968), .ZN(n14886) );
  NAND2_X1 U9701 ( .A1(n14916), .A2(n11302), .ZN(n7976) );
  AND2_X1 U9702 ( .A1(n14885), .A2(n7976), .ZN(n7970) );
  NAND2_X1 U9703 ( .A1(n14886), .A2(n7970), .ZN(n14870) );
  NAND2_X1 U9704 ( .A1(n7458), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U9705 ( .A1(n7509), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U9706 ( .A1(n7671), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7472) );
  AND2_X1 U9707 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7470) );
  NOR2_X1 U9708 ( .A1(n7490), .A2(n7470), .ZN(n14884) );
  INV_X1 U9709 ( .A(n14884), .ZN(n12178) );
  NAND2_X1 U9710 ( .A1(n7488), .A2(n12178), .ZN(n7471) );
  NAND2_X1 U9711 ( .A1(n7476), .A2(n7475), .ZN(n7478) );
  NAND2_X1 U9712 ( .A1(n9773), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7477) );
  XNOR2_X1 U9713 ( .A(n7497), .B(n7496), .ZN(n9769) );
  OR2_X1 U9714 ( .A1(n7758), .A2(n9769), .ZN(n7484) );
  NAND2_X1 U9715 ( .A1(n7480), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7482) );
  XNOR2_X1 U9716 ( .A(n7482), .B(n7481), .ZN(n10439) );
  INV_X1 U9717 ( .A(n10439), .ZN(n10573) );
  OR2_X1 U9718 ( .A1(n10424), .A2(n10573), .ZN(n7483) );
  NAND2_X1 U9719 ( .A1(n10890), .A2(n14864), .ZN(n7977) );
  INV_X1 U9720 ( .A(n14864), .ZN(n7486) );
  NAND2_X1 U9721 ( .A1(n14890), .A2(n7486), .ZN(n7978) );
  NAND2_X1 U9722 ( .A1(n7977), .A2(n7978), .ZN(n14867) );
  INV_X1 U9723 ( .A(n14867), .ZN(n14871) );
  NAND3_X1 U9724 ( .A1(n14869), .A2(n14870), .A3(n14871), .ZN(n7487) );
  NAND2_X1 U9725 ( .A1(n7487), .A2(n7977), .ZN(n14850) );
  NAND2_X1 U9726 ( .A1(n7509), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9727 ( .A1(n7458), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9728 ( .A1(n7490), .A2(n7489), .ZN(n7523) );
  OR2_X1 U9729 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  NAND2_X1 U9730 ( .A1(n7523), .A2(n7491), .ZN(n14860) );
  NAND2_X1 U9731 ( .A1(n7488), .A2(n14860), .ZN(n7493) );
  NAND2_X1 U9732 ( .A1(n7671), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7492) );
  NAND4_X1 U9733 ( .A1(n7495), .A2(n7494), .A3(n7493), .A4(n7492), .ZN(n12255)
         );
  OR2_X1 U9734 ( .A1(n7801), .A2(SI_5_), .ZN(n7507) );
  NAND2_X1 U9735 ( .A1(n7497), .A2(n7496), .ZN(n7499) );
  NAND2_X1 U9736 ( .A1(n9781), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7498) );
  XNOR2_X1 U9737 ( .A(n7516), .B(n7515), .ZN(n9767) );
  OR2_X1 U9738 ( .A1(n7758), .A2(n9767), .ZN(n7506) );
  NOR2_X1 U9739 ( .A1(n7480), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7502) );
  NOR2_X1 U9740 ( .A1(n7502), .A2(n8112), .ZN(n7500) );
  MUX2_X1 U9741 ( .A(n8112), .B(n7500), .S(P3_IR_REG_5__SCAN_IN), .Z(n7504) );
  INV_X1 U9742 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7501) );
  NAND2_X1 U9743 ( .A1(n7502), .A2(n7501), .ZN(n7533) );
  INV_X1 U9744 ( .A(n7533), .ZN(n7503) );
  INV_X1 U9745 ( .A(n10448), .ZN(n10756) );
  OR2_X1 U9746 ( .A1(n10424), .A2(n10756), .ZN(n7505) );
  XNOR2_X1 U9747 ( .A(n12255), .B(n14859), .ZN(n14854) );
  NAND2_X1 U9748 ( .A1(n14850), .A2(n14854), .ZN(n7508) );
  INV_X1 U9749 ( .A(n12255), .ZN(n14873) );
  NAND2_X1 U9750 ( .A1(n14873), .A2(n14859), .ZN(n7961) );
  NAND2_X1 U9751 ( .A1(n7508), .A2(n7961), .ZN(n11400) );
  NAND2_X1 U9752 ( .A1(n7509), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U9753 ( .A1(n7906), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7512) );
  XNOR2_X1 U9754 ( .A(n7523), .B(P3_REG3_REG_6__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U9755 ( .A1(n7488), .A2(n12221), .ZN(n7511) );
  NAND2_X1 U9756 ( .A1(n7911), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9757 ( .A1(n7533), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7514) );
  XNOR2_X1 U9758 ( .A(n7514), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10488) );
  INV_X1 U9759 ( .A(n10488), .ZN(n10451) );
  NAND2_X1 U9760 ( .A1(n7516), .A2(n7515), .ZN(n7518) );
  NAND2_X1 U9761 ( .A1(n9775), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7517) );
  XNOR2_X1 U9762 ( .A(n9786), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7519) );
  XNOR2_X1 U9763 ( .A(n7530), .B(n7519), .ZN(n9754) );
  OR2_X1 U9764 ( .A1(n7758), .A2(n9754), .ZN(n7521) );
  INV_X1 U9765 ( .A(SI_6_), .ZN(n9753) );
  OR2_X1 U9766 ( .A1(n7801), .A2(n9753), .ZN(n7520) );
  OAI211_X1 U9767 ( .C1(n10424), .C2(n10451), .A(n7521), .B(n7520), .ZN(n12218) );
  NAND2_X1 U9768 ( .A1(n11315), .A2(n12218), .ZN(n7987) );
  INV_X1 U9769 ( .A(n12218), .ZN(n9626) );
  NAND2_X1 U9770 ( .A1(n14855), .A2(n9626), .ZN(n7985) );
  NAND2_X1 U9771 ( .A1(n11400), .A2(n11401), .ZN(n11399) );
  NAND2_X1 U9772 ( .A1(n7906), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9773 ( .A1(n7912), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7527) );
  OAI21_X1 U9774 ( .B1(n7523), .B2(P3_REG3_REG_6__SCAN_IN), .A(
        P3_REG3_REG_7__SCAN_IN), .ZN(n7524) );
  INV_X1 U9775 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15130) );
  INV_X1 U9776 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U9777 ( .A1(n15130), .A2(n10491), .ZN(n7522) );
  NAND2_X1 U9778 ( .A1(n7524), .A2(n7538), .ZN(n12068) );
  NAND2_X1 U9779 ( .A1(n7488), .A2(n12068), .ZN(n7526) );
  NAND2_X1 U9780 ( .A1(n7911), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7525) );
  OR2_X1 U9781 ( .A1(n7801), .A2(SI_7_), .ZN(n7537) );
  NAND2_X1 U9782 ( .A1(n9784), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7531) );
  INV_X1 U9783 ( .A(n7546), .ZN(n7532) );
  XNOR2_X1 U9784 ( .A(n7547), .B(n7532), .ZN(n9759) );
  OR2_X1 U9785 ( .A1(n7758), .A2(n9759), .ZN(n7536) );
  NAND2_X1 U9786 ( .A1(n7544), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7534) );
  XNOR2_X1 U9787 ( .A(n7534), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10489) );
  OR2_X1 U9788 ( .A1(n10424), .A2(n10489), .ZN(n7535) );
  NAND2_X1 U9789 ( .A1(n14840), .A2(n12067), .ZN(n7988) );
  INV_X1 U9790 ( .A(n12067), .ZN(n14953) );
  NAND2_X1 U9791 ( .A1(n12254), .A2(n14953), .ZN(n7989) );
  NAND2_X1 U9792 ( .A1(n7509), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7543) );
  NAND2_X1 U9793 ( .A1(n7458), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7542) );
  AND2_X1 U9794 ( .A1(n7538), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7539) );
  OR2_X1 U9795 ( .A1(n7539), .A2(n7570), .ZN(n14846) );
  NAND2_X1 U9796 ( .A1(n7886), .A2(n14846), .ZN(n7541) );
  NAND2_X1 U9797 ( .A1(n7911), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7540) );
  OAI21_X1 U9798 ( .B1(n7544), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7545) );
  XNOR2_X1 U9799 ( .A(n7545), .B(P3_IR_REG_8__SCAN_IN), .ZN(n14789) );
  XNOR2_X1 U9800 ( .A(n7556), .B(n7555), .ZN(n9739) );
  OR2_X1 U9801 ( .A1(n7758), .A2(n9739), .ZN(n7549) );
  INV_X1 U9802 ( .A(SI_8_), .ZN(n9738) );
  OR2_X1 U9803 ( .A1(n7801), .A2(n9738), .ZN(n7548) );
  OAI211_X1 U9804 ( .C1(n10424), .C2(n11056), .A(n7549), .B(n7548), .ZN(n14845) );
  NAND2_X1 U9805 ( .A1(n11647), .A2(n14845), .ZN(n7994) );
  INV_X1 U9806 ( .A(n11647), .ZN(n14826) );
  INV_X1 U9807 ( .A(n14845), .ZN(n11646) );
  NAND2_X1 U9808 ( .A1(n14826), .A2(n11646), .ZN(n7995) );
  NAND2_X1 U9809 ( .A1(n7994), .A2(n7995), .ZN(n14837) );
  INV_X1 U9810 ( .A(n14837), .ZN(n7991) );
  NAND2_X1 U9811 ( .A1(n7912), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9812 ( .A1(n7906), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7553) );
  INV_X1 U9813 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11051) );
  XNOR2_X1 U9814 ( .A(n7570), .B(n11051), .ZN(n14831) );
  NAND2_X1 U9815 ( .A1(n7886), .A2(n14831), .ZN(n7552) );
  NAND2_X1 U9816 ( .A1(n7911), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9817 ( .A1(n9801), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7557) );
  XNOR2_X1 U9818 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7576) );
  INV_X1 U9819 ( .A(n7576), .ZN(n7559) );
  XNOR2_X1 U9820 ( .A(n7577), .B(n7559), .ZN(n9757) );
  OR2_X1 U9821 ( .A1(n7758), .A2(n9757), .ZN(n7566) );
  OR2_X1 U9822 ( .A1(n7801), .A2(SI_9_), .ZN(n7565) );
  NOR2_X1 U9823 ( .A1(n7560), .A2(n8112), .ZN(n7561) );
  MUX2_X1 U9824 ( .A(n8112), .B(n7561), .S(P3_IR_REG_9__SCAN_IN), .Z(n7563) );
  OR2_X1 U9825 ( .A1(n7563), .A2(n7562), .ZN(n11474) );
  OR2_X1 U9826 ( .A1(n10424), .A2(n11057), .ZN(n7564) );
  NAND2_X1 U9827 ( .A1(n14839), .A2(n14830), .ZN(n8002) );
  INV_X1 U9828 ( .A(n8002), .ZN(n7568) );
  INV_X1 U9829 ( .A(n14830), .ZN(n7567) );
  NAND2_X1 U9830 ( .A1(n12253), .A2(n7567), .ZN(n8000) );
  NAND2_X1 U9831 ( .A1(n7912), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9832 ( .A1(n7458), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7574) );
  NOR2_X1 U9833 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_REG3_REG_10__SCAN_IN), 
        .ZN(n7569) );
  INV_X1 U9834 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15065) );
  AOI21_X1 U9835 ( .B1(n7570), .B2(n11051), .A(n15065), .ZN(n7571) );
  OR2_X1 U9836 ( .A1(n7590), .A2(n7571), .ZN(n12097) );
  NAND2_X1 U9837 ( .A1(n7886), .A2(n12097), .ZN(n7573) );
  NAND2_X1 U9838 ( .A1(n7911), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U9839 ( .A1(n9807), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7578) );
  XNOR2_X1 U9840 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7596) );
  INV_X1 U9841 ( .A(n7596), .ZN(n7580) );
  XNOR2_X1 U9842 ( .A(n7597), .B(n7580), .ZN(n9750) );
  OR2_X1 U9843 ( .A1(n7758), .A2(n9750), .ZN(n7587) );
  OR2_X1 U9844 ( .A1(n7801), .A2(SI_10_), .ZN(n7586) );
  NOR2_X1 U9845 ( .A1(n7562), .A2(n8112), .ZN(n7581) );
  MUX2_X1 U9846 ( .A(n8112), .B(n7581), .S(P3_IR_REG_10__SCAN_IN), .Z(n7584)
         );
  INV_X1 U9847 ( .A(n7582), .ZN(n7583) );
  INV_X1 U9848 ( .A(n11475), .ZN(n14800) );
  OR2_X1 U9849 ( .A1(n10424), .A2(n14800), .ZN(n7585) );
  INV_X1 U9850 ( .A(n11671), .ZN(n12090) );
  NAND2_X1 U9851 ( .A1(n14825), .A2(n12090), .ZN(n7999) );
  INV_X1 U9852 ( .A(n7999), .ZN(n7588) );
  NAND2_X1 U9853 ( .A1(n14290), .A2(n11671), .ZN(n8001) );
  NAND2_X1 U9854 ( .A1(n7912), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9855 ( .A1(n7458), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7594) );
  INV_X1 U9856 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7589) );
  OR2_X1 U9857 ( .A1(n7590), .A2(n7589), .ZN(n7591) );
  NAND2_X1 U9858 ( .A1(n7605), .A2(n7591), .ZN(n14293) );
  NAND2_X1 U9859 ( .A1(n7886), .A2(n14293), .ZN(n7593) );
  NAND2_X1 U9860 ( .A1(n7911), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U9861 ( .A1(n15124), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7598) );
  XNOR2_X1 U9862 ( .A(n9824), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7600) );
  XNOR2_X1 U9863 ( .A(n7613), .B(n7600), .ZN(n9761) );
  OR2_X1 U9864 ( .A1(n7758), .A2(n9761), .ZN(n7604) );
  OR2_X1 U9865 ( .A1(n7801), .A2(SI_11_), .ZN(n7603) );
  NAND2_X1 U9866 ( .A1(n7582), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7601) );
  XNOR2_X1 U9867 ( .A(n7601), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11526) );
  OR2_X1 U9868 ( .A1(n10424), .A2(n11526), .ZN(n7602) );
  XNOR2_X1 U9869 ( .A(n12252), .B(n12201), .ZN(n14284) );
  NAND2_X1 U9870 ( .A1(n11672), .A2(n12201), .ZN(n8007) );
  NAND2_X1 U9871 ( .A1(n7912), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7610) );
  NAND2_X1 U9872 ( .A1(n7458), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9873 ( .A1(n7605), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7606) );
  NAND2_X1 U9874 ( .A1(n7631), .A2(n7606), .ZN(n12123) );
  NAND2_X1 U9875 ( .A1(n7886), .A2(n12123), .ZN(n7608) );
  NAND2_X1 U9876 ( .A1(n7911), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7607) );
  OR2_X1 U9877 ( .A1(n7582), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U9878 ( .A1(n7626), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7611) );
  XNOR2_X1 U9879 ( .A(n7611), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U9880 ( .A1(n9824), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U9881 ( .A1(n9951), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9882 ( .A1(n9950), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9883 ( .A1(n7622), .A2(n7615), .ZN(n7616) );
  NAND2_X1 U9884 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  NAND2_X1 U9885 ( .A1(n7623), .A2(n7618), .ZN(n9782) );
  OR2_X1 U9886 ( .A1(n7758), .A2(n9782), .ZN(n7620) );
  OR2_X1 U9887 ( .A1(n7801), .A2(n15112), .ZN(n7619) );
  OAI211_X1 U9888 ( .C1(n10424), .C2(n12263), .A(n7620), .B(n7619), .ZN(n12410) );
  NAND2_X1 U9889 ( .A1(n14289), .A2(n12410), .ZN(n8012) );
  INV_X1 U9890 ( .A(n12410), .ZN(n9636) );
  NAND2_X1 U9891 ( .A1(n14272), .A2(n9636), .ZN(n8010) );
  NAND2_X1 U9892 ( .A1(n8012), .A2(n8010), .ZN(n11674) );
  INV_X1 U9893 ( .A(n11674), .ZN(n7946) );
  NAND2_X1 U9894 ( .A1(n11668), .A2(n7946), .ZN(n7621) );
  XNOR2_X1 U9895 ( .A(n7637), .B(n10057), .ZN(n14214) );
  NAND2_X1 U9896 ( .A1(n14214), .A2(n7923), .ZN(n7630) );
  NAND2_X1 U9897 ( .A1(n7644), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7627) );
  XNOR2_X1 U9898 ( .A(n7627), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12278) );
  OAI22_X1 U9899 ( .A1(n7801), .A2(n8179), .B1(n10424), .B2(n14216), .ZN(n7628) );
  INV_X1 U9900 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U9901 ( .A1(n7630), .A2(n7629), .ZN(n12413) );
  NAND2_X1 U9902 ( .A1(n7631), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7632) );
  AND2_X1 U9903 ( .A1(n7654), .A2(n7632), .ZN(n14275) );
  INV_X1 U9904 ( .A(n14275), .ZN(n11689) );
  NAND2_X1 U9905 ( .A1(n7886), .A2(n11689), .ZN(n7636) );
  NAND2_X1 U9906 ( .A1(n7458), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U9907 ( .A1(n7911), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9908 ( .A1(n7912), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7633) );
  AND2_X1 U9909 ( .A1(n12413), .A2(n9644), .ZN(n7939) );
  OR2_X1 U9910 ( .A1(n12413), .A2(n9644), .ZN(n8017) );
  NAND2_X1 U9911 ( .A1(n10206), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U9912 ( .A1(n10237), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7640) );
  OR2_X1 U9913 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  NAND2_X1 U9914 ( .A1(n7660), .A2(n7643), .ZN(n9818) );
  NAND2_X1 U9915 ( .A1(n9818), .A2(n7923), .ZN(n7653) );
  NOR2_X1 U9916 ( .A1(n7644), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7648) );
  NOR2_X1 U9917 ( .A1(n7648), .A2(n8112), .ZN(n7645) );
  MUX2_X1 U9918 ( .A(n8112), .B(n7645), .S(P3_IR_REG_14__SCAN_IN), .Z(n7646)
         );
  INV_X1 U9919 ( .A(n7646), .ZN(n7649) );
  NAND2_X1 U9920 ( .A1(n7648), .A2(n7647), .ZN(n7681) );
  NAND2_X1 U9921 ( .A1(n7649), .A2(n7681), .ZN(n12309) );
  INV_X1 U9922 ( .A(n12309), .ZN(n7650) );
  OAI22_X1 U9923 ( .A1(n7801), .A2(SI_14_), .B1(n7650), .B2(n10424), .ZN(n7651) );
  INV_X1 U9924 ( .A(n7651), .ZN(n7652) );
  NAND2_X1 U9925 ( .A1(n7458), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9926 ( .A1(n7911), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7657) );
  OR2_X1 U9927 ( .A1(n7378), .A2(n7669), .ZN(n12675) );
  NAND2_X1 U9928 ( .A1(n7886), .A2(n12675), .ZN(n7656) );
  NAND2_X1 U9929 ( .A1(n7912), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U9930 ( .A1(n12415), .A2(n12652), .ZN(n12655) );
  NAND2_X1 U9931 ( .A1(n12801), .A2(n14273), .ZN(n8020) );
  INV_X1 U9932 ( .A(n12664), .ZN(n12671) );
  NAND2_X1 U9933 ( .A1(n10261), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7678) );
  INV_X1 U9934 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U9935 ( .A1(n10260), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7661) );
  INV_X1 U9936 ( .A(n7676), .ZN(n7662) );
  XNOR2_X1 U9937 ( .A(n7677), .B(n7662), .ZN(n9927) );
  NAND2_X1 U9938 ( .A1(n9927), .A2(n7923), .ZN(n7667) );
  NAND2_X1 U9939 ( .A1(n7681), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7664) );
  XNOR2_X1 U9940 ( .A(n7664), .B(n7663), .ZN(n12332) );
  OAI22_X1 U9941 ( .A1(n7801), .A2(n9928), .B1(n10424), .B2(n12332), .ZN(n7665) );
  INV_X1 U9942 ( .A(n7665), .ZN(n7666) );
  NAND2_X1 U9943 ( .A1(n7667), .A2(n7666), .ZN(n12424) );
  NAND2_X1 U9944 ( .A1(n7912), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9945 ( .A1(n7906), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7674) );
  INV_X1 U9946 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7668) );
  OR2_X1 U9947 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  NAND2_X1 U9948 ( .A1(n7686), .A2(n7670), .ZN(n12659) );
  NAND2_X1 U9949 ( .A1(n7886), .A2(n12659), .ZN(n7673) );
  NAND2_X1 U9950 ( .A1(n7911), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7672) );
  NAND4_X1 U9951 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n12667)
         );
  XNOR2_X1 U9952 ( .A(n12424), .B(n12667), .ZN(n12649) );
  INV_X1 U9953 ( .A(n12649), .ZN(n12656) );
  OR2_X1 U9954 ( .A1(n12671), .A2(n12656), .ZN(n12639) );
  NAND2_X1 U9955 ( .A1(n10203), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9956 ( .A1(n10161), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7679) );
  INV_X1 U9957 ( .A(n7695), .ZN(n7680) );
  XNOR2_X1 U9958 ( .A(n7696), .B(n7680), .ZN(n14220) );
  NAND2_X1 U9959 ( .A1(n14220), .A2(n7923), .ZN(n7685) );
  OR2_X1 U9960 ( .A1(n7681), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U9961 ( .A1(n7682), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U9962 ( .A(n7702), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12344) );
  OAI22_X1 U9963 ( .A1(n7801), .A2(n8191), .B1(n10424), .B2(n14222), .ZN(n7683) );
  INV_X1 U9964 ( .A(n7683), .ZN(n7684) );
  NAND2_X1 U9965 ( .A1(n7685), .A2(n7684), .ZN(n12417) );
  NAND2_X1 U9966 ( .A1(n7912), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9967 ( .A1(n7458), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U9968 ( .A1(n7686), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U9969 ( .A1(n7708), .A2(n7687), .ZN(n12643) );
  NAND2_X1 U9970 ( .A1(n7886), .A2(n12643), .ZN(n7689) );
  NAND2_X1 U9971 ( .A1(n7911), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7688) );
  OR2_X1 U9972 ( .A1(n12417), .A2(n12651), .ZN(n7960) );
  NAND2_X1 U9973 ( .A1(n12417), .A2(n12651), .ZN(n8026) );
  NAND2_X1 U9974 ( .A1(n7960), .A2(n8026), .ZN(n12634) );
  INV_X1 U9975 ( .A(n12634), .ZN(n12641) );
  OR2_X1 U9976 ( .A1(n12639), .A2(n12634), .ZN(n7694) );
  INV_X1 U9977 ( .A(n12667), .ZN(n12638) );
  NAND2_X1 U9978 ( .A1(n12424), .A2(n12638), .ZN(n8025) );
  OR2_X1 U9979 ( .A1(n12656), .A2(n12655), .ZN(n12653) );
  AND2_X1 U9980 ( .A1(n8025), .A2(n12653), .ZN(n12640) );
  NAND2_X1 U9981 ( .A1(n10240), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U9982 ( .A1(n10239), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7699) );
  INV_X1 U9983 ( .A(n7714), .ZN(n7700) );
  XNOR2_X1 U9984 ( .A(n7715), .B(n7700), .ZN(n14208) );
  NAND2_X1 U9985 ( .A1(n14208), .A2(n7923), .ZN(n7707) );
  NAND2_X1 U9986 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  NAND2_X1 U9987 ( .A1(n7703), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7704) );
  XNOR2_X1 U9988 ( .A(n7704), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12359) );
  OAI22_X1 U9989 ( .A1(n7801), .A2(n8197), .B1(n10424), .B2(n14210), .ZN(n7705) );
  INV_X1 U9990 ( .A(n7705), .ZN(n7706) );
  NAND2_X1 U9991 ( .A1(n7707), .A2(n7706), .ZN(n12430) );
  NAND2_X1 U9992 ( .A1(n7912), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9993 ( .A1(n7906), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7712) );
  AND2_X1 U9994 ( .A1(n7708), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7709) );
  OR2_X1 U9995 ( .A1(n7709), .A2(n7726), .ZN(n12626) );
  NAND2_X1 U9996 ( .A1(n7886), .A2(n12626), .ZN(n7711) );
  NAND2_X1 U9997 ( .A1(n7911), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7710) );
  OR2_X1 U9998 ( .A1(n12430), .A2(n12637), .ZN(n8031) );
  NAND2_X1 U9999 ( .A1(n12430), .A2(n12637), .ZN(n8035) );
  NAND2_X1 U10000 ( .A1(n8031), .A2(n8035), .ZN(n12619) );
  INV_X1 U10001 ( .A(n12619), .ZN(n12624) );
  NAND2_X1 U10002 ( .A1(n12625), .A2(n12624), .ZN(n12623) );
  NAND2_X1 U10003 ( .A1(n12623), .A2(n8035), .ZN(n12607) );
  INV_X1 U10004 ( .A(n12607), .ZN(n7732) );
  NAND2_X1 U10005 ( .A1(n15099), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U10006 ( .A1(n10500), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7717) );
  INV_X1 U10007 ( .A(n7733), .ZN(n7718) );
  XNOR2_X1 U10008 ( .A(n7734), .B(n7718), .ZN(n14228) );
  NAND2_X1 U10009 ( .A1(n14228), .A2(n7923), .ZN(n7724) );
  INV_X1 U10010 ( .A(SI_18_), .ZN(n8633) );
  NAND2_X1 U10011 ( .A1(n7719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7721) );
  INV_X1 U10012 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7720) );
  XNOR2_X1 U10013 ( .A(n7721), .B(n7720), .ZN(n14230) );
  OAI22_X1 U10014 ( .A1(n7801), .A2(n8633), .B1(n10424), .B2(n14230), .ZN(
        n7722) );
  INV_X1 U10015 ( .A(n7722), .ZN(n7723) );
  NAND2_X1 U10016 ( .A1(n7912), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10017 ( .A1(n7906), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7730) );
  INV_X1 U10018 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7725) );
  NOR2_X1 U10019 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  OR2_X1 U10020 ( .A1(n7746), .A2(n7727), .ZN(n12610) );
  NAND2_X1 U10021 ( .A1(n7886), .A2(n12610), .ZN(n7729) );
  NAND2_X1 U10022 ( .A1(n7911), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U10023 ( .A1(n12609), .A2(n12622), .ZN(n8037) );
  NAND2_X1 U10024 ( .A1(n12605), .A2(n8034), .ZN(n12593) );
  INV_X1 U10025 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U10026 ( .A1(n10597), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7752) );
  INV_X1 U10027 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U10028 ( .A1(n10596), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7736) );
  OR2_X1 U10029 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U10030 ( .A1(n7753), .A2(n7739), .ZN(n10156) );
  NAND2_X1 U10031 ( .A1(n10156), .A2(n7923), .ZN(n7744) );
  NAND2_X1 U10032 ( .A1(n6511), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7741) );
  OAI22_X1 U10033 ( .A1(n7801), .A2(SI_19_), .B1(n10617), .B2(n10424), .ZN(
        n7742) );
  INV_X1 U10034 ( .A(n7742), .ZN(n7743) );
  NAND2_X1 U10035 ( .A1(n7912), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10036 ( .A1(n7906), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7750) );
  INV_X1 U10037 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7745) );
  OR2_X1 U10038 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  NAND2_X1 U10039 ( .A1(n7761), .A2(n7747), .ZN(n12594) );
  NAND2_X1 U10040 ( .A1(n7886), .A2(n12594), .ZN(n7749) );
  NAND2_X1 U10041 ( .A1(n7911), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7748) );
  NAND4_X1 U10042 ( .A1(n7751), .A2(n7750), .A3(n7749), .A4(n7748), .ZN(n12574) );
  NAND2_X1 U10043 ( .A1(n12782), .A2(n12574), .ZN(n8042) );
  NAND2_X1 U10044 ( .A1(n7756), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10045 ( .A1(n7770), .A2(n7757), .ZN(n10343) );
  OR2_X1 U10046 ( .A1(n10343), .A2(n7758), .ZN(n7760) );
  INV_X1 U10047 ( .A(SI_20_), .ZN(n10344) );
  NAND2_X1 U10048 ( .A1(n7906), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10049 ( .A1(n7911), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10050 ( .A1(n7761), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U10051 ( .A1(n7776), .A2(n7762), .ZN(n12577) );
  NAND2_X1 U10052 ( .A1(n7886), .A2(n12577), .ZN(n7764) );
  NAND2_X1 U10053 ( .A1(n7912), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7763) );
  NAND4_X1 U10054 ( .A1(n7766), .A2(n7765), .A3(n7764), .A4(n7763), .ZN(n12588) );
  XNOR2_X1 U10055 ( .A(n12721), .B(n12588), .ZN(n12572) );
  NAND2_X1 U10056 ( .A1(n7767), .A2(n12572), .ZN(n12571) );
  INV_X1 U10057 ( .A(n12588), .ZN(n12559) );
  OR2_X1 U10058 ( .A1(n12721), .A2(n12559), .ZN(n7768) );
  NAND2_X1 U10059 ( .A1(n12571), .A2(n7768), .ZN(n12561) );
  INV_X1 U10060 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U10061 ( .A1(n10737), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7787) );
  INV_X1 U10062 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U10063 ( .A1(n10740), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U10064 ( .A1(n7787), .A2(n7771), .ZN(n7785) );
  XNOR2_X1 U10065 ( .A(n7786), .B(n7785), .ZN(n10589) );
  NAND2_X1 U10066 ( .A1(n10589), .A2(n7923), .ZN(n7773) );
  INV_X1 U10067 ( .A(SI_21_), .ZN(n10590) );
  NAND2_X1 U10068 ( .A1(n7912), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10069 ( .A1(n7906), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7780) );
  INV_X1 U10070 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10071 ( .A1(n7776), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U10072 ( .A1(n7791), .A2(n7777), .ZN(n12563) );
  NAND2_X1 U10073 ( .A1(n7886), .A2(n12563), .ZN(n7779) );
  NAND2_X1 U10074 ( .A1(n7911), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U10075 ( .A1(n12562), .A2(n9667), .ZN(n7782) );
  NAND2_X1 U10076 ( .A1(n12561), .A2(n7782), .ZN(n7784) );
  OR2_X1 U10077 ( .A1(n12562), .A2(n9667), .ZN(n7783) );
  NAND2_X1 U10078 ( .A1(n7784), .A2(n7783), .ZN(n12550) );
  INV_X1 U10079 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11097) );
  XNOR2_X1 U10080 ( .A(n11097), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n7798) );
  XNOR2_X1 U10081 ( .A(n7799), .B(n7798), .ZN(n10651) );
  NAND2_X1 U10082 ( .A1(n10651), .A2(n7923), .ZN(n7790) );
  INV_X1 U10083 ( .A(SI_22_), .ZN(n7788) );
  NAND2_X1 U10084 ( .A1(n7791), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10085 ( .A1(n7806), .A2(n7792), .ZN(n12551) );
  NAND2_X1 U10086 ( .A1(n7886), .A2(n12551), .ZN(n7796) );
  NAND2_X1 U10087 ( .A1(n7906), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10088 ( .A1(n7911), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10089 ( .A1(n7912), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7793) );
  NAND4_X1 U10090 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n12535) );
  NAND2_X1 U10091 ( .A1(n12714), .A2(n12558), .ZN(n8055) );
  NAND2_X1 U10092 ( .A1(n12550), .A2(n8055), .ZN(n7797) );
  NAND2_X1 U10093 ( .A1(n7797), .A2(n8054), .ZN(n12541) );
  NAND2_X1 U10094 ( .A1(n11097), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U10095 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n7810) );
  XNOR2_X1 U10096 ( .A(n7811), .B(n7810), .ZN(n10883) );
  NAND2_X1 U10097 ( .A1(n10883), .A2(n7923), .ZN(n7803) );
  INV_X1 U10098 ( .A(SI_23_), .ZN(n10886) );
  INV_X1 U10099 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10100 ( .A1(n7806), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10101 ( .A1(n7819), .A2(n7807), .ZN(n12539) );
  AOI22_X1 U10102 ( .A1(n12539), .A2(n7886), .B1(n7911), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n7809) );
  AOI22_X1 U10103 ( .A1(n7912), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n7906), .B2(
        P3_REG0_REG_23__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U10104 ( .A(n12709), .B(n12525), .ZN(n12439) );
  OR2_X1 U10105 ( .A1(n12709), .A2(n12525), .ZN(n8059) );
  INV_X1 U10106 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11273) );
  NAND2_X1 U10107 ( .A1(n11273), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7812) );
  INV_X1 U10108 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U10109 ( .A1(n7814), .A2(n11559), .ZN(n7815) );
  INV_X1 U10110 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11555) );
  XNOR2_X1 U10111 ( .A(n7824), .B(n11555), .ZN(n11268) );
  NAND2_X1 U10112 ( .A1(n11268), .A2(n7923), .ZN(n7818) );
  INV_X1 U10113 ( .A(SI_24_), .ZN(n11269) );
  INV_X1 U10114 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U10115 ( .A1(n7819), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10116 ( .A1(n7829), .A2(n7820), .ZN(n12528) );
  NAND2_X1 U10117 ( .A1(n12528), .A2(n7886), .ZN(n7822) );
  AOI22_X1 U10118 ( .A1(n7912), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n7906), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n7821) );
  INV_X1 U10119 ( .A(n12536), .ZN(n12136) );
  OR2_X1 U10120 ( .A1(n12443), .A2(n12136), .ZN(n8060) );
  NAND2_X1 U10121 ( .A1(n12443), .A2(n12136), .ZN(n8062) );
  NAND2_X1 U10122 ( .A1(n8060), .A2(n8062), .ZN(n12523) );
  INV_X1 U10123 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U10124 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13376), .B2(n14196), .ZN(n7826) );
  XNOR2_X1 U10125 ( .A(n7836), .B(n7826), .ZN(n11325) );
  NAND2_X1 U10126 ( .A1(n11325), .A2(n7923), .ZN(n7828) );
  INV_X1 U10127 ( .A(SI_25_), .ZN(n11327) );
  NAND2_X1 U10128 ( .A1(n7829), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10129 ( .A1(n7845), .A2(n7830), .ZN(n12516) );
  NAND2_X1 U10130 ( .A1(n12516), .A2(n7886), .ZN(n7833) );
  AOI22_X1 U10131 ( .A1(n7912), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n7906), .B2(
        P3_REG0_REG_25__SCAN_IN), .ZN(n7832) );
  NAND2_X1 U10132 ( .A1(n7911), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7831) );
  OR2_X1 U10133 ( .A1(n12699), .A2(n12526), .ZN(n8066) );
  NAND2_X1 U10134 ( .A1(n12699), .A2(n12526), .ZN(n8067) );
  NAND2_X1 U10135 ( .A1(n12515), .A2(n12514), .ZN(n7834) );
  NAND2_X1 U10136 ( .A1(n7834), .A2(n8067), .ZN(n12499) );
  NAND2_X1 U10137 ( .A1(n13376), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10138 ( .A1(n14196), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7837) );
  INV_X1 U10139 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14192) );
  INV_X1 U10140 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U10141 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14192), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n15097), .ZN(n7839) );
  INV_X1 U10142 ( .A(n7839), .ZN(n7840) );
  XNOR2_X1 U10143 ( .A(n7853), .B(n7840), .ZN(n11430) );
  NAND2_X1 U10144 ( .A1(n11430), .A2(n7923), .ZN(n7842) );
  INV_X1 U10145 ( .A(SI_26_), .ZN(n11431) );
  INV_X1 U10146 ( .A(n7845), .ZN(n7844) );
  INV_X1 U10147 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U10148 ( .A1(n7844), .A2(n7843), .ZN(n7864) );
  NAND2_X1 U10149 ( .A1(n7845), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10150 ( .A1(n7864), .A2(n7846), .ZN(n12506) );
  NAND2_X1 U10151 ( .A1(n12506), .A2(n7886), .ZN(n7851) );
  INV_X1 U10152 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U10153 ( .A1(n7912), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10154 ( .A1(n7906), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7847) );
  OAI211_X1 U10155 ( .C1(n12697), .C2(n7891), .A(n7848), .B(n7847), .ZN(n7849)
         );
  INV_X1 U10156 ( .A(n7849), .ZN(n7850) );
  NAND2_X1 U10157 ( .A1(n12499), .A2(n8071), .ZN(n7852) );
  NAND2_X1 U10158 ( .A1(n12507), .A2(n12486), .ZN(n8072) );
  INV_X1 U10159 ( .A(n7853), .ZN(n7855) );
  NAND2_X1 U10160 ( .A1(n14192), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U10161 ( .A1(n15097), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7856) );
  INV_X1 U10162 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11776) );
  INV_X1 U10163 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U10164 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n11776), .B2(n14189), .ZN(n7858) );
  INV_X1 U10165 ( .A(n7858), .ZN(n7859) );
  XNOR2_X1 U10166 ( .A(n7873), .B(n7859), .ZN(n11517) );
  NAND2_X1 U10167 ( .A1(n11517), .A2(n7923), .ZN(n7861) );
  INV_X1 U10168 ( .A(SI_27_), .ZN(n11518) );
  NAND2_X2 U10169 ( .A1(n7861), .A2(n7860), .ZN(n12453) );
  INV_X1 U10170 ( .A(n7864), .ZN(n7863) );
  INV_X1 U10171 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10172 ( .A1(n7863), .A2(n7862), .ZN(n7878) );
  NAND2_X1 U10173 ( .A1(n7864), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10174 ( .A1(n7878), .A2(n7865), .ZN(n12494) );
  NAND2_X1 U10175 ( .A1(n12494), .A2(n7886), .ZN(n7870) );
  INV_X1 U10176 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n15058) );
  NAND2_X1 U10177 ( .A1(n7912), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10178 ( .A1(n7906), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7866) );
  OAI211_X1 U10179 ( .C1(n15058), .C2(n7891), .A(n7867), .B(n7866), .ZN(n7868)
         );
  INV_X1 U10180 ( .A(n7868), .ZN(n7869) );
  NAND2_X1 U10181 ( .A1(n12453), .A2(n12502), .ZN(n12476) );
  NOR2_X1 U10182 ( .A1(n14189), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10183 ( .A1(n14189), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7874) );
  INV_X1 U10184 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13370) );
  INV_X1 U10185 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U10186 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13370), .B2(n11701), .ZN(n7875) );
  XNOR2_X1 U10187 ( .A(n7883), .B(n7875), .ZN(n12818) );
  NAND2_X1 U10188 ( .A1(n12818), .A2(n7923), .ZN(n7877) );
  INV_X1 U10189 ( .A(SI_28_), .ZN(n12819) );
  NAND2_X1 U10190 ( .A1(n7878), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10191 ( .A1(n12407), .A2(n7879), .ZN(n12480) );
  INV_X1 U10192 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U10193 ( .A1(n7906), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U10194 ( .A1(n7912), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7880) );
  OAI211_X1 U10195 ( .C1(n12691), .C2(n7891), .A(n7881), .B(n7880), .ZN(n7882)
         );
  NAND2_X1 U10196 ( .A1(n12479), .A2(n12485), .ZN(n7938) );
  XNOR2_X1 U10197 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n7895) );
  XNOR2_X1 U10198 ( .A(n7897), .B(n7895), .ZN(n12814) );
  NAND2_X1 U10199 ( .A1(n12814), .A2(n7923), .ZN(n7885) );
  INV_X1 U10200 ( .A(SI_29_), .ZN(n12816) );
  OR2_X1 U10201 ( .A1(n7801), .A2(n12816), .ZN(n7884) );
  NAND2_X1 U10202 ( .A1(n7885), .A2(n7884), .ZN(n12465) );
  INV_X1 U10203 ( .A(n12407), .ZN(n7887) );
  NAND2_X1 U10204 ( .A1(n7887), .A2(n7886), .ZN(n7917) );
  INV_X1 U10205 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10206 ( .A1(n7906), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10207 ( .A1(n7912), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7888) );
  OAI211_X1 U10208 ( .C1(n7891), .C2(n7890), .A(n7889), .B(n7888), .ZN(n7892)
         );
  INV_X1 U10209 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U10210 ( .A1(n12465), .A2(n12473), .ZN(n8081) );
  NAND2_X1 U10211 ( .A1(n12409), .A2(n12457), .ZN(n7894) );
  INV_X1 U10212 ( .A(n7895), .ZN(n7896) );
  INV_X1 U10213 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U10214 ( .A1(n11771), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7898) );
  INV_X1 U10215 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U10216 ( .A1(n13364), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7901) );
  INV_X1 U10217 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U10218 ( .A1(n14187), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10219 ( .A1(n7901), .A2(n7900), .ZN(n7918) );
  NAND2_X1 U10220 ( .A1(n7921), .A2(n7901), .ZN(n7903) );
  XNOR2_X1 U10221 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n7902) );
  XNOR2_X1 U10222 ( .A(n7903), .B(n7902), .ZN(n12812) );
  NAND2_X1 U10223 ( .A1(n12812), .A2(n7923), .ZN(n7905) );
  INV_X1 U10224 ( .A(SI_31_), .ZN(n12808) );
  OR2_X1 U10225 ( .A1(n7801), .A2(n12808), .ZN(n7904) );
  NAND2_X1 U10226 ( .A1(n7911), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U10227 ( .A1(n7912), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10228 ( .A1(n7906), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n7907) );
  AND3_X1 U10229 ( .A1(n7909), .A2(n7908), .A3(n7907), .ZN(n7910) );
  AND2_X1 U10230 ( .A1(n7917), .A2(n7910), .ZN(n12406) );
  NOR2_X1 U10231 ( .A1(n7925), .A2(n12406), .ZN(n8088) );
  NAND2_X1 U10232 ( .A1(n7911), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10233 ( .A1(n7912), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10234 ( .A1(n7458), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n7913) );
  AND3_X1 U10235 ( .A1(n7915), .A2(n7914), .A3(n7913), .ZN(n7916) );
  NAND2_X1 U10236 ( .A1(n7917), .A2(n7916), .ZN(n12461) );
  INV_X1 U10237 ( .A(n12406), .ZN(n12251) );
  NAND2_X1 U10238 ( .A1(n7919), .A2(n7918), .ZN(n7920) );
  NAND2_X1 U10239 ( .A1(n7921), .A2(n7920), .ZN(n12059) );
  INV_X1 U10240 ( .A(SI_30_), .ZN(n12060) );
  NOR2_X1 U10241 ( .A1(n7801), .A2(n12060), .ZN(n7922) );
  AOI21_X1 U10242 ( .B1(n12059), .B2(n7923), .A(n7922), .ZN(n7953) );
  AOI21_X1 U10243 ( .B1(n12461), .B2(n12251), .A(n7953), .ZN(n7924) );
  NOR2_X1 U10244 ( .A1(n8088), .A2(n7924), .ZN(n7928) );
  AND2_X1 U10245 ( .A1(n7953), .A2(n12461), .ZN(n7937) );
  XNOR2_X1 U10246 ( .A(n7930), .B(n10617), .ZN(n8098) );
  NAND2_X1 U10247 ( .A1(n7932), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7931) );
  MUX2_X1 U10248 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7931), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7933) );
  NAND2_X1 U10249 ( .A1(n7935), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10250 ( .A1(n10540), .A2(n10618), .ZN(n10518) );
  INV_X1 U10251 ( .A(n12457), .ZN(n7956) );
  INV_X1 U10252 ( .A(n7937), .ZN(n8085) );
  AND2_X2 U10253 ( .A1(n8079), .A2(n7938), .ZN(n12477) );
  AND2_X2 U10254 ( .A1(n8071), .A2(n8072), .ZN(n12501) );
  INV_X1 U10255 ( .A(n12584), .ZN(n12592) );
  INV_X1 U10256 ( .A(n7939), .ZN(n8016) );
  NAND2_X1 U10257 ( .A1(n8016), .A2(n8017), .ZN(n14279) );
  NAND2_X1 U10258 ( .A1(n8001), .A2(n7999), .ZN(n11669) );
  NOR2_X1 U10259 ( .A1(n10638), .A2(n7962), .ZN(n10628) );
  NAND4_X1 U10260 ( .A1(n14871), .A2(n7991), .A3(n14893), .A4(n10628), .ZN(
        n7944) );
  NOR2_X1 U10261 ( .A1(n11644), .A2(n14914), .ZN(n7942) );
  NAND2_X1 U10262 ( .A1(n7966), .A2(n7969), .ZN(n11295) );
  INV_X1 U10263 ( .A(n7941), .ZN(n10639) );
  NAND4_X1 U10264 ( .A1(n7942), .A2(n14821), .A3(n11401), .A4(n10639), .ZN(
        n7943) );
  NOR4_X1 U10265 ( .A1(n11669), .A2(n11306), .A3(n7944), .A4(n7943), .ZN(n7945) );
  NAND4_X1 U10266 ( .A1(n12664), .A2(n7946), .A3(n14284), .A4(n7945), .ZN(
        n7947) );
  OR4_X1 U10267 ( .A1(n12656), .A2(n12634), .A3(n14279), .A4(n7947), .ZN(n7948) );
  NOR4_X1 U10268 ( .A1(n12592), .A2(n12608), .A3(n12619), .A4(n7948), .ZN(
        n7949) );
  XNOR2_X1 U10269 ( .A(n12562), .B(n12575), .ZN(n12560) );
  NAND4_X1 U10270 ( .A1(n12549), .A2(n12572), .A3(n7949), .A4(n12560), .ZN(
        n7950) );
  NOR2_X1 U10271 ( .A1(n12439), .A2(n7950), .ZN(n7951) );
  NAND4_X1 U10272 ( .A1(n12501), .A2(n12514), .A3(n7823), .A4(n7951), .ZN(
        n7952) );
  NOR2_X1 U10273 ( .A1(n12451), .A2(n7952), .ZN(n7955) );
  INV_X1 U10274 ( .A(n12461), .ZN(n7954) );
  XNOR2_X1 U10275 ( .A(n7957), .B(n12392), .ZN(n8097) );
  NAND2_X1 U10276 ( .A1(n10592), .A2(n10618), .ZN(n9712) );
  NAND2_X1 U10277 ( .A1(n10345), .A2(n12392), .ZN(n10620) );
  INV_X1 U10278 ( .A(n10620), .ZN(n10536) );
  NAND2_X1 U10279 ( .A1(n6525), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7958) );
  MUX2_X1 U10280 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7958), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7959) );
  OAI21_X1 U10281 ( .B1(n12638), .B2(n12424), .A(n7960), .ZN(n8024) );
  AND2_X1 U10282 ( .A1(n7987), .A2(n7961), .ZN(n7983) );
  OAI21_X1 U10283 ( .B1(n7962), .B2(n10592), .A(n10529), .ZN(n7965) );
  INV_X1 U10284 ( .A(n7962), .ZN(n7963) );
  NAND3_X1 U10285 ( .A1(n7969), .A2(n7963), .A3(n10652), .ZN(n7964) );
  AOI22_X1 U10286 ( .A1(n7965), .A2(n7964), .B1(n10638), .B2(n10592), .ZN(
        n7967) );
  MUX2_X1 U10287 ( .A(n10619), .B(n7967), .S(n7966), .Z(n7972) );
  OAI21_X1 U10288 ( .B1(n10619), .B2(n7969), .A(n7968), .ZN(n7971) );
  OAI22_X1 U10289 ( .A1(n7972), .A2(n7971), .B1(n10619), .B2(n7970), .ZN(n7975) );
  AOI21_X1 U10290 ( .B1(n14869), .B2(n7973), .A(n10529), .ZN(n7974) );
  AOI21_X1 U10291 ( .B1(n7975), .B2(n14869), .A(n7974), .ZN(n7981) );
  OAI21_X1 U10292 ( .B1(n10529), .B2(n7976), .A(n14871), .ZN(n7980) );
  MUX2_X1 U10293 ( .A(n7978), .B(n7977), .S(n10529), .Z(n7979) );
  OAI211_X1 U10294 ( .C1(n7981), .C2(n7980), .A(n14854), .B(n7979), .ZN(n7982)
         );
  OAI21_X1 U10295 ( .B1(n7983), .B2(n10529), .A(n7982), .ZN(n7986) );
  OAI21_X1 U10296 ( .B1(n14873), .B2(n14859), .A(n7985), .ZN(n7984) );
  AOI22_X1 U10297 ( .A1(n7986), .A2(n7985), .B1(n10529), .B2(n7984), .ZN(n7993) );
  OAI21_X1 U10298 ( .B1(n10619), .B2(n7987), .A(n11313), .ZN(n7992) );
  MUX2_X1 U10299 ( .A(n7989), .B(n7988), .S(n10619), .Z(n7990) );
  OAI211_X1 U10300 ( .C1(n7993), .C2(n7992), .A(n7991), .B(n7990), .ZN(n7998)
         );
  INV_X1 U10301 ( .A(n11669), .ZN(n7997) );
  MUX2_X1 U10302 ( .A(n7995), .B(n7994), .S(n10529), .Z(n7996) );
  AND4_X1 U10303 ( .A1(n7998), .A2(n14821), .A3(n7997), .A4(n7996), .ZN(n8006)
         );
  OAI21_X1 U10304 ( .B1(n11669), .B2(n8000), .A(n7999), .ZN(n8004) );
  OAI21_X1 U10305 ( .B1(n11669), .B2(n8002), .A(n8001), .ZN(n8003) );
  MUX2_X1 U10306 ( .A(n8004), .B(n8003), .S(n10619), .Z(n8005) );
  INV_X1 U10307 ( .A(n14284), .ZN(n14287) );
  NOR3_X1 U10308 ( .A1(n8006), .A2(n8005), .A3(n14287), .ZN(n8009) );
  AOI21_X1 U10309 ( .B1(n8012), .B2(n8007), .A(n10619), .ZN(n8008) );
  OAI21_X1 U10310 ( .B1(n8009), .B2(n8008), .A(n8010), .ZN(n8015) );
  OAI21_X1 U10311 ( .B1(n11672), .B2(n12201), .A(n8010), .ZN(n8011) );
  NAND2_X1 U10312 ( .A1(n8011), .A2(n10619), .ZN(n8014) );
  INV_X1 U10313 ( .A(n8012), .ZN(n8013) );
  AOI22_X1 U10314 ( .A1(n8015), .A2(n8014), .B1(n10619), .B2(n8013), .ZN(n8019) );
  MUX2_X1 U10315 ( .A(n8017), .B(n8016), .S(n10619), .Z(n8018) );
  OAI211_X1 U10316 ( .C1(n8019), .C2(n14279), .A(n12664), .B(n8018), .ZN(n8022) );
  MUX2_X1 U10317 ( .A(n8020), .B(n12655), .S(n10529), .Z(n8021) );
  AND3_X1 U10318 ( .A1(n8022), .A2(n12649), .A3(n8021), .ZN(n8023) );
  AOI21_X1 U10319 ( .B1(n10529), .B2(n8024), .A(n8023), .ZN(n8028) );
  AND2_X1 U10320 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  OAI22_X1 U10321 ( .A1(n8028), .A2(n7692), .B1(n8027), .B2(n10529), .ZN(n8030) );
  INV_X1 U10322 ( .A(n12417), .ZN(n12794) );
  NAND3_X1 U10323 ( .A1(n12794), .A2(n10619), .A3(n12416), .ZN(n8029) );
  AOI211_X1 U10324 ( .C1(n8030), .C2(n8029), .A(n12619), .B(n12608), .ZN(n8045) );
  INV_X1 U10325 ( .A(n8031), .ZN(n8032) );
  NAND2_X1 U10326 ( .A1(n8037), .A2(n8032), .ZN(n8033) );
  NAND3_X1 U10327 ( .A1(n8042), .A2(n8034), .A3(n8033), .ZN(n8040) );
  INV_X1 U10328 ( .A(n8035), .ZN(n8036) );
  NAND2_X1 U10329 ( .A1(n12602), .A2(n8036), .ZN(n8038) );
  NAND3_X1 U10330 ( .A1(n8038), .A2(n8041), .A3(n8037), .ZN(n8039) );
  MUX2_X1 U10331 ( .A(n8040), .B(n8039), .S(n10529), .Z(n8044) );
  MUX2_X1 U10332 ( .A(n8042), .B(n8041), .S(n10619), .Z(n8043) );
  OAI211_X1 U10333 ( .C1(n8045), .C2(n8044), .A(n12572), .B(n8043), .ZN(n8049)
         );
  NAND2_X1 U10334 ( .A1(n12588), .A2(n10619), .ZN(n8047) );
  NAND2_X1 U10335 ( .A1(n12559), .A2(n10529), .ZN(n8046) );
  MUX2_X1 U10336 ( .A(n8047), .B(n8046), .S(n12721), .Z(n8048) );
  NAND3_X1 U10337 ( .A1(n8049), .A2(n12560), .A3(n8048), .ZN(n8053) );
  NAND2_X1 U10338 ( .A1(n12575), .A2(n10529), .ZN(n8051) );
  NAND2_X1 U10339 ( .A1(n9667), .A2(n10619), .ZN(n8050) );
  MUX2_X1 U10340 ( .A(n8051), .B(n8050), .S(n12562), .Z(n8052) );
  NAND3_X1 U10341 ( .A1(n8053), .A2(n12549), .A3(n8052), .ZN(n8057) );
  MUX2_X1 U10342 ( .A(n8055), .B(n8054), .S(n10619), .Z(n8056) );
  NAND3_X1 U10343 ( .A1(n8057), .A2(n12540), .A3(n8056), .ZN(n8058) );
  OAI21_X1 U10344 ( .B1(n8058), .B2(n12523), .A(n12514), .ZN(n8070) );
  NAND2_X1 U10345 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  AND2_X1 U10346 ( .A1(n8061), .A2(n8062), .ZN(n8065) );
  NAND2_X1 U10347 ( .A1(n12709), .A2(n12525), .ZN(n8063) );
  OAI21_X1 U10348 ( .B1(n12523), .B2(n8063), .A(n8062), .ZN(n8064) );
  MUX2_X1 U10349 ( .A(n8065), .B(n8064), .S(n10619), .Z(n8069) );
  MUX2_X1 U10350 ( .A(n8067), .B(n8066), .S(n10619), .Z(n8068) );
  OAI211_X1 U10351 ( .C1(n8070), .C2(n8069), .A(n12501), .B(n8068), .ZN(n8074)
         );
  MUX2_X1 U10352 ( .A(n8072), .B(n8071), .S(n10529), .Z(n8073) );
  AOI21_X1 U10353 ( .B1(n8074), .B2(n8073), .A(n12451), .ZN(n8076) );
  NOR3_X1 U10354 ( .A1(n12453), .A2(n12502), .A3(n10619), .ZN(n8075) );
  NOR2_X1 U10355 ( .A1(n8076), .A2(n8075), .ZN(n8084) );
  NAND2_X1 U10356 ( .A1(n12477), .A2(n10619), .ZN(n8083) );
  INV_X1 U10357 ( .A(n12477), .ZN(n8080) );
  NAND2_X1 U10358 ( .A1(n8077), .A2(n10619), .ZN(n8078) );
  OAI211_X1 U10359 ( .C1(n8084), .C2(n8080), .A(n8079), .B(n8078), .ZN(n8082)
         );
  OAI211_X1 U10360 ( .C1(n8084), .C2(n8083), .A(n8082), .B(n8081), .ZN(n8087)
         );
  NAND3_X1 U10361 ( .A1(n8087), .A2(n8086), .A3(n8085), .ZN(n8091) );
  INV_X1 U10362 ( .A(n8088), .ZN(n8090) );
  NAND3_X1 U10363 ( .A1(n8091), .A2(n8090), .A3(n8089), .ZN(n8094) );
  INV_X1 U10364 ( .A(n8092), .ZN(n8093) );
  NAND2_X1 U10365 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  MUX2_X1 U10366 ( .A(n10536), .B(n12684), .S(n8095), .Z(n8096) );
  OR2_X1 U10367 ( .A1(n10422), .A2(P3_U3151), .ZN(n10884) );
  INV_X1 U10368 ( .A(n10884), .ZN(n8101) );
  OAI21_X1 U10369 ( .B1(n8108), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8104) );
  MUX2_X1 U10370 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8104), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8107) );
  INV_X1 U10371 ( .A(n8105), .ZN(n8106) );
  NAND2_X1 U10372 ( .A1(n8107), .A2(n8106), .ZN(n11328) );
  INV_X1 U10373 ( .A(n9602), .ZN(n8114) );
  NOR2_X1 U10374 ( .A1(n8105), .A2(n8112), .ZN(n8111) );
  MUX2_X1 U10375 ( .A(n8112), .B(n8111), .S(P3_IR_REG_26__SCAN_IN), .Z(n8113)
         );
  NAND2_X1 U10376 ( .A1(n8114), .A2(n9605), .ZN(n8115) );
  NOR2_X1 U10377 ( .A1(n10529), .A2(n10620), .ZN(n10627) );
  NAND2_X1 U10378 ( .A1(n10660), .A2(n10627), .ZN(n10662) );
  NOR3_X1 U10379 ( .A1(n10662), .A2(n10437), .A3(n8119), .ZN(n8121) );
  OAI21_X1 U10380 ( .B1(n10884), .B2(n10652), .A(P3_B_REG_SCAN_IN), .ZN(n8120)
         );
  OR2_X1 U10381 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  NOR2_X1 U10382 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8125) );
  NOR2_X2 U10383 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8124) );
  NOR2_X1 U10384 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8129) );
  INV_X1 U10385 ( .A(n8358), .ZN(n8131) );
  NAND2_X1 U10386 ( .A1(n8708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8132) );
  XNOR2_X2 U10387 ( .A(n8132), .B(n8707), .ZN(n13782) );
  INV_X1 U10388 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9752) );
  XNOR2_X1 U10389 ( .A(n8135), .B(SI_1_), .ZN(n8532) );
  AND2_X1 U10390 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10391 ( .A1(n9737), .A2(n8134), .ZN(n9123) );
  INV_X1 U10392 ( .A(n8135), .ZN(n8136) );
  NAND2_X1 U10393 ( .A1(n8136), .A2(SI_1_), .ZN(n8137) );
  NAND2_X1 U10394 ( .A1(n8138), .A2(n8137), .ZN(n8519) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n8178), .Z(n8140) );
  XNOR2_X1 U10396 ( .A(n8140), .B(SI_2_), .ZN(n8518) );
  INV_X1 U10397 ( .A(n8518), .ZN(n8139) );
  NAND2_X1 U10398 ( .A1(n8519), .A2(n8139), .ZN(n8142) );
  NAND2_X1 U10399 ( .A1(n8140), .A2(SI_2_), .ZN(n8141) );
  NAND2_X1 U10400 ( .A1(n8508), .A2(n8143), .ZN(n8146) );
  NAND2_X1 U10401 ( .A1(n8144), .A2(SI_3_), .ZN(n8145) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8178), .Z(n8148) );
  XNOR2_X1 U10403 ( .A(n8148), .B(SI_4_), .ZN(n8492) );
  INV_X1 U10404 ( .A(n8492), .ZN(n8147) );
  NAND2_X1 U10405 ( .A1(n8493), .A2(n8147), .ZN(n8150) );
  NAND2_X1 U10406 ( .A1(n8148), .A2(SI_4_), .ZN(n8149) );
  NAND2_X1 U10407 ( .A1(n8150), .A2(n8149), .ZN(n8568) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8178), .Z(n8152) );
  XNOR2_X1 U10409 ( .A(n8152), .B(SI_5_), .ZN(n8567) );
  INV_X1 U10410 ( .A(n8567), .ZN(n8151) );
  NAND2_X1 U10411 ( .A1(n8152), .A2(SI_5_), .ZN(n8153) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8231), .Z(n8154) );
  XNOR2_X1 U10413 ( .A(n8154), .B(SI_6_), .ZN(n8555) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9771), .Z(n8156) );
  XNOR2_X1 U10415 ( .A(n8156), .B(SI_7_), .ZN(n8478) );
  INV_X1 U10416 ( .A(n8478), .ZN(n8155) );
  NAND2_X1 U10417 ( .A1(n8156), .A2(SI_7_), .ZN(n8157) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n9771), .Z(n8159) );
  XNOR2_X1 U10419 ( .A(n8159), .B(SI_8_), .ZN(n8464) );
  INV_X1 U10420 ( .A(n8464), .ZN(n8158) );
  NAND2_X1 U10421 ( .A1(n8159), .A2(SI_8_), .ZN(n8160) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n8231), .Z(n8162) );
  XNOR2_X1 U10423 ( .A(n8162), .B(SI_9_), .ZN(n8449) );
  INV_X1 U10424 ( .A(n8449), .ZN(n8161) );
  NAND2_X1 U10425 ( .A1(n8162), .A2(SI_9_), .ZN(n8163) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n8178), .Z(n8165) );
  XNOR2_X1 U10427 ( .A(n8165), .B(SI_10_), .ZN(n8600) );
  INV_X1 U10428 ( .A(n8600), .ZN(n8164) );
  NAND2_X1 U10429 ( .A1(n8165), .A2(SI_10_), .ZN(n8166) );
  MUX2_X1 U10430 ( .A(n9824), .B(n9820), .S(n9771), .Z(n8169) );
  NAND2_X1 U10431 ( .A1(n8169), .A2(n8168), .ZN(n8172) );
  INV_X1 U10432 ( .A(n8169), .ZN(n8170) );
  NAND2_X1 U10433 ( .A1(n8170), .A2(SI_11_), .ZN(n8171) );
  NAND2_X1 U10434 ( .A1(n8172), .A2(n8171), .ZN(n8435) );
  MUX2_X1 U10435 ( .A(n9950), .B(n9951), .S(n8178), .Z(n8173) );
  NAND2_X1 U10436 ( .A1(n8173), .A2(n15112), .ZN(n8176) );
  INV_X1 U10437 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U10438 ( .A1(n8174), .A2(SI_12_), .ZN(n8175) );
  MUX2_X1 U10439 ( .A(n10057), .B(n10055), .S(n8178), .Z(n8180) );
  NAND2_X1 U10440 ( .A1(n8180), .A2(n8179), .ZN(n8183) );
  INV_X1 U10441 ( .A(n8180), .ZN(n8181) );
  NAND2_X1 U10442 ( .A1(n8181), .A2(SI_13_), .ZN(n8182) );
  MUX2_X1 U10443 ( .A(n10237), .B(n10206), .S(n8231), .Z(n8616) );
  INV_X1 U10444 ( .A(SI_14_), .ZN(n9817) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n8231), .Z(n8187) );
  NAND2_X1 U10446 ( .A1(n8187), .A2(SI_15_), .ZN(n8379) );
  OAI21_X1 U10447 ( .B1(n8616), .B2(n9817), .A(n8379), .ZN(n8184) );
  INV_X1 U10448 ( .A(n8184), .ZN(n8185) );
  INV_X1 U10449 ( .A(n8616), .ZN(n8374) );
  NOR2_X1 U10450 ( .A1(n8374), .A2(SI_14_), .ZN(n8186) );
  NAND2_X1 U10451 ( .A1(n8186), .A2(n8379), .ZN(n8189) );
  INV_X1 U10452 ( .A(n8187), .ZN(n8188) );
  NAND2_X1 U10453 ( .A1(n8188), .A2(n9928), .ZN(n8378) );
  MUX2_X1 U10454 ( .A(n10161), .B(n10203), .S(n8231), .Z(n8192) );
  INV_X1 U10455 ( .A(n8192), .ZN(n8193) );
  NAND2_X1 U10456 ( .A1(n8193), .A2(SI_16_), .ZN(n8194) );
  MUX2_X1 U10457 ( .A(n10239), .B(n10240), .S(n8231), .Z(n8198) );
  INV_X1 U10458 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10459 ( .A1(n8199), .A2(SI_17_), .ZN(n8200) );
  MUX2_X1 U10460 ( .A(n10500), .B(n15099), .S(n8231), .Z(n8357) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n8231), .Z(n8206) );
  NAND2_X1 U10462 ( .A1(n8206), .A2(SI_19_), .ZN(n8638) );
  OAI21_X1 U10463 ( .B1(n8633), .B2(n8357), .A(n8638), .ZN(n8203) );
  INV_X1 U10464 ( .A(n8203), .ZN(n8204) );
  INV_X1 U10465 ( .A(n8357), .ZN(n8631) );
  NOR2_X1 U10466 ( .A1(n8631), .A2(SI_18_), .ZN(n8205) );
  NAND2_X1 U10467 ( .A1(n8205), .A2(n8638), .ZN(n8208) );
  INV_X1 U10468 ( .A(n8206), .ZN(n8207) );
  INV_X1 U10469 ( .A(SI_19_), .ZN(n10157) );
  NAND2_X1 U10470 ( .A1(n8207), .A2(n10157), .ZN(n8637) );
  INV_X1 U10471 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10594) );
  INV_X1 U10472 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10600) );
  MUX2_X1 U10473 ( .A(n10594), .B(n10600), .S(n8231), .Z(n8334) );
  INV_X1 U10474 ( .A(n8334), .ZN(n8210) );
  NAND2_X1 U10475 ( .A1(n8335), .A2(n8210), .ZN(n8214) );
  INV_X1 U10476 ( .A(n8211), .ZN(n8212) );
  NAND2_X1 U10477 ( .A1(n8214), .A2(n8213), .ZN(n8345) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8231), .Z(n8216) );
  XNOR2_X1 U10479 ( .A(n8216), .B(SI_21_), .ZN(n8344) );
  NAND2_X1 U10480 ( .A1(n8345), .A2(n8215), .ZN(n8218) );
  NAND2_X1 U10481 ( .A1(n8216), .A2(SI_21_), .ZN(n8217) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n8231), .Z(n9453) );
  INV_X1 U10483 ( .A(n9453), .ZN(n8221) );
  NAND2_X1 U10484 ( .A1(n8219), .A2(SI_22_), .ZN(n8220) );
  OAI21_X2 U10485 ( .B1(n9454), .B2(n8221), .A(n8220), .ZN(n8223) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n8231), .Z(n8222) );
  NAND2_X1 U10487 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n8231), .Z(n8655) );
  MUX2_X1 U10489 ( .A(n13376), .B(n14196), .S(n8231), .Z(n8227) );
  NAND2_X1 U10490 ( .A1(n8227), .A2(n11327), .ZN(n8230) );
  INV_X1 U10491 ( .A(n8227), .ZN(n8228) );
  NAND2_X1 U10492 ( .A1(n8228), .A2(SI_25_), .ZN(n8229) );
  NAND2_X1 U10493 ( .A1(n8230), .A2(n8229), .ZN(n8312) );
  MUX2_X1 U10494 ( .A(n15097), .B(n14192), .S(n8231), .Z(n8298) );
  OAI21_X1 U10495 ( .B1(n8300), .B2(n11431), .A(n8298), .ZN(n8233) );
  NAND2_X1 U10496 ( .A1(n8300), .A2(n11431), .ZN(n8232) );
  NAND2_X1 U10497 ( .A1(n8233), .A2(n8232), .ZN(n8288) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n9771), .Z(n8285) );
  NOR2_X1 U10499 ( .A1(n8285), .A2(SI_27_), .ZN(n8235) );
  NAND2_X1 U10500 ( .A1(n8285), .A2(SI_27_), .ZN(n8234) );
  OAI21_X2 U10501 ( .B1(n8288), .B2(n8235), .A(n8234), .ZN(n8265) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n9771), .Z(n8236) );
  XNOR2_X1 U10503 ( .A(n8236), .B(SI_28_), .ZN(n8264) );
  INV_X1 U10504 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U10505 ( .A1(n8237), .A2(n12819), .ZN(n8238) );
  OAI21_X2 U10506 ( .B1(n8265), .B2(n8264), .A(n8238), .ZN(n8693) );
  INV_X1 U10507 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11772) );
  MUX2_X1 U10508 ( .A(n11772), .B(n11771), .S(n9771), .Z(n8239) );
  XNOR2_X1 U10509 ( .A(n8239), .B(SI_29_), .ZN(n8692) );
  NAND2_X1 U10510 ( .A1(n8693), .A2(n8692), .ZN(n8241) );
  NAND2_X1 U10511 ( .A1(n8239), .A2(n12816), .ZN(n8240) );
  MUX2_X1 U10512 ( .A(n13364), .B(n14187), .S(n9771), .Z(n8242) );
  XNOR2_X1 U10513 ( .A(n8242), .B(SI_30_), .ZN(n8683) );
  INV_X1 U10514 ( .A(n8683), .ZN(n8243) );
  MUX2_X1 U10515 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n9771), .Z(n8244) );
  XNOR2_X1 U10516 ( .A(n8244), .B(SI_31_), .ZN(n8245) );
  NOR2_X1 U10517 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8248) );
  NOR3_X1 U10518 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .ZN(n8249) );
  XNOR2_X2 U10519 ( .A(n8253), .B(n8252), .ZN(n14191) );
  AND2_X2 U10520 ( .A1(n8326), .A2(n9771), .ZN(n8534) );
  NAND2_X1 U10521 ( .A1(n14185), .A2(n8534), .ZN(n8255) );
  NAND2_X4 U10522 ( .A1(n8326), .A2(n9737), .ZN(n8694) );
  INV_X1 U10523 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14180) );
  OR2_X1 U10524 ( .A1(n8694), .A2(n14180), .ZN(n8254) );
  XNOR2_X2 U10525 ( .A(n8257), .B(n14179), .ZN(n8260) );
  INV_X1 U10526 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15083) );
  NAND2_X2 U10527 ( .A1(n8270), .A2(n8261), .ZN(n8542) );
  NAND2_X1 U10528 ( .A1(n8687), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10529 ( .A1(n8539), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8262) );
  OAI211_X1 U10530 ( .C1(n8691), .C2(n15083), .A(n8263), .B(n8262), .ZN(n13793) );
  XNOR2_X1 U10531 ( .A(n13790), .B(n13793), .ZN(n8908) );
  NAND2_X1 U10532 ( .A1(n13367), .A2(n8534), .ZN(n8267) );
  OR2_X1 U10533 ( .A1(n8694), .A2(n11701), .ZN(n8266) );
  NAND2_X1 U10534 ( .A1(n8539), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8284) );
  INV_X1 U10535 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13867) );
  OR2_X1 U10536 ( .A1(n8542), .A2(n13867), .ZN(n8283) );
  NAND2_X1 U10537 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8577) );
  INV_X1 U10538 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8576) );
  NOR2_X1 U10539 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U10540 ( .A1(n8578), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10541 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n8271) );
  NAND2_X1 U10542 ( .A1(n8607), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8592) );
  INV_X1 U10543 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8412) );
  INV_X1 U10544 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10545 ( .A1(n8400), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8645) );
  INV_X1 U10546 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8644) );
  INV_X1 U10547 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13584) );
  NAND2_X1 U10548 ( .A1(n8348), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10549 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n8328), .ZN(n8673) );
  INV_X1 U10550 ( .A(n8673), .ZN(n8272) );
  NAND2_X1 U10551 ( .A1(n8272), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8675) );
  INV_X1 U10552 ( .A(n8675), .ZN(n8273) );
  NAND2_X1 U10553 ( .A1(n8273), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8662) );
  INV_X1 U10554 ( .A(n8662), .ZN(n8274) );
  NAND2_X1 U10555 ( .A1(n8274), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8319) );
  INV_X1 U10556 ( .A(n8319), .ZN(n8275) );
  NAND2_X1 U10557 ( .A1(n8275), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8306) );
  INV_X1 U10558 ( .A(n8306), .ZN(n8276) );
  NAND2_X1 U10559 ( .A1(n8276), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8292) );
  INV_X1 U10560 ( .A(n8292), .ZN(n8277) );
  NAND2_X1 U10561 ( .A1(n8277), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13849) );
  INV_X1 U10562 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10563 ( .A1(n8292), .A2(n8278), .ZN(n8279) );
  NAND2_X1 U10564 ( .A1(n13849), .A2(n8279), .ZN(n13864) );
  OR2_X1 U10565 ( .A1(n8676), .A2(n13864), .ZN(n8282) );
  INV_X1 U10566 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8280) );
  OR2_X1 U10567 ( .A1(n8691), .A2(n8280), .ZN(n8281) );
  NAND4_X1 U10568 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n13851) );
  XNOR2_X1 U10569 ( .A(n14085), .B(n13880), .ZN(n13862) );
  INV_X1 U10570 ( .A(n8285), .ZN(n8286) );
  XNOR2_X1 U10571 ( .A(n8286), .B(SI_27_), .ZN(n8287) );
  OR2_X1 U10572 ( .A1(n8694), .A2(n14189), .ZN(n8289) );
  NAND2_X1 U10573 ( .A1(n8539), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8297) );
  INV_X1 U10574 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8290) );
  OR2_X1 U10575 ( .A1(n8691), .A2(n8290), .ZN(n8296) );
  INV_X1 U10576 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n15068) );
  NAND2_X1 U10577 ( .A1(n8306), .A2(n15068), .ZN(n8291) );
  NAND2_X1 U10578 ( .A1(n8292), .A2(n8291), .ZN(n13889) );
  OR2_X1 U10579 ( .A1(n8698), .A2(n13889), .ZN(n8295) );
  INV_X1 U10580 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8293) );
  OR2_X1 U10581 ( .A1(n8542), .A2(n8293), .ZN(n8294) );
  NAND4_X1 U10582 ( .A1(n8297), .A2(n8296), .A3(n8295), .A4(n8294), .ZN(n13817) );
  INV_X1 U10583 ( .A(n13817), .ZN(n13840) );
  XNOR2_X1 U10584 ( .A(n8298), .B(SI_26_), .ZN(n8299) );
  XNOR2_X1 U10585 ( .A(n8300), .B(n8299), .ZN(n13371) );
  NAND2_X1 U10586 ( .A1(n13371), .A2(n8534), .ZN(n8302) );
  OR2_X1 U10587 ( .A1(n8694), .A2(n14192), .ZN(n8301) );
  NAND2_X1 U10588 ( .A1(n8697), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8311) );
  INV_X1 U10589 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8303) );
  OR2_X1 U10590 ( .A1(n8268), .A2(n8303), .ZN(n8310) );
  INV_X1 U10591 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U10592 ( .A1(n8319), .A2(n8304), .ZN(n8305) );
  NAND2_X1 U10593 ( .A1(n8306), .A2(n8305), .ZN(n13898) );
  OR2_X1 U10594 ( .A1(n8698), .A2(n13898), .ZN(n8309) );
  INV_X1 U10595 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8307) );
  OR2_X1 U10596 ( .A1(n8542), .A2(n8307), .ZN(n8308) );
  NAND4_X1 U10597 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n13839) );
  XNOR2_X1 U10598 ( .A(n14098), .B(n13881), .ZN(n13904) );
  XNOR2_X1 U10599 ( .A(n8313), .B(n8312), .ZN(n13374) );
  NAND2_X1 U10600 ( .A1(n13374), .A2(n8534), .ZN(n8315) );
  OR2_X1 U10601 ( .A1(n8694), .A2(n14196), .ZN(n8314) );
  NAND2_X1 U10602 ( .A1(n8697), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8323) );
  INV_X1 U10603 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8316) );
  OR2_X1 U10604 ( .A1(n8268), .A2(n8316), .ZN(n8322) );
  INV_X1 U10605 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10606 ( .A1(n8662), .A2(n8317), .ZN(n8318) );
  NAND2_X1 U10607 ( .A1(n8319), .A2(n8318), .ZN(n13921) );
  OR2_X1 U10608 ( .A1(n8676), .A2(n13921), .ZN(n8321) );
  INV_X1 U10609 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n13922) );
  OR2_X1 U10610 ( .A1(n8542), .A2(n13922), .ZN(n8320) );
  NAND4_X1 U10611 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n13933) );
  XNOR2_X1 U10612 ( .A(n13924), .B(n13933), .ZN(n13812) );
  OR2_X1 U10613 ( .A1(n9454), .A2(n8324), .ZN(n8325) );
  XNOR2_X1 U10614 ( .A(n8325), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U10615 ( .A1(n8539), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8333) );
  INV_X1 U10616 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8327) );
  OR2_X1 U10617 ( .A1(n8542), .A2(n8327), .ZN(n8332) );
  OAI21_X1 U10618 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8328), .A(n8673), .ZN(
        n13593) );
  OR2_X1 U10619 ( .A1(n8676), .A2(n13593), .ZN(n8331) );
  INV_X1 U10620 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8329) );
  OR2_X1 U10621 ( .A1(n8691), .A2(n8329), .ZN(n8330) );
  NAND4_X1 U10622 ( .A1(n8333), .A2(n8332), .A3(n8331), .A4(n8330), .ZN(n13984) );
  XNOR2_X1 U10623 ( .A(n13599), .B(n13984), .ZN(n13974) );
  XNOR2_X1 U10624 ( .A(n8335), .B(n8334), .ZN(n10593) );
  NAND2_X1 U10625 ( .A1(n10593), .A2(n8534), .ZN(n8337) );
  OR2_X1 U10626 ( .A1(n8694), .A2(n10600), .ZN(n8336) );
  AND2_X1 U10627 ( .A1(n8647), .A2(n13584), .ZN(n8338) );
  OR2_X1 U10628 ( .A1(n8348), .A2(n8338), .ZN(n14008) );
  INV_X1 U10629 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10630 ( .A1(n8687), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10631 ( .A1(n8539), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8339) );
  OAI211_X1 U10632 ( .C1(n8691), .C2(n8341), .A(n8340), .B(n8339), .ZN(n8342)
         );
  INV_X1 U10633 ( .A(n8342), .ZN(n8343) );
  OAI21_X1 U10634 ( .B1(n14008), .B2(n8698), .A(n8343), .ZN(n14022) );
  INV_X1 U10635 ( .A(n14022), .ZN(n13828) );
  XNOR2_X1 U10636 ( .A(n14130), .B(n13828), .ZN(n14013) );
  XNOR2_X1 U10637 ( .A(n8345), .B(n8344), .ZN(n10736) );
  NAND2_X1 U10638 ( .A1(n10736), .A2(n8534), .ZN(n8347) );
  OR2_X1 U10639 ( .A1(n8694), .A2(n10737), .ZN(n8346) );
  OR2_X1 U10640 ( .A1(n8348), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10641 ( .A1(n8350), .A2(n8349), .ZN(n13994) );
  OR2_X1 U10642 ( .A1(n13994), .A2(n8698), .ZN(n8356) );
  INV_X1 U10643 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10644 ( .A1(n8687), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10645 ( .A1(n8539), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8351) );
  OAI211_X1 U10646 ( .C1(n8691), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8354)
         );
  INV_X1 U10647 ( .A(n8354), .ZN(n8355) );
  NAND2_X1 U10648 ( .A1(n8356), .A2(n8355), .ZN(n14002) );
  INV_X1 U10649 ( .A(n14002), .ZN(n13830) );
  XNOR2_X1 U10650 ( .A(n14125), .B(n13830), .ZN(n13986) );
  XNOR2_X1 U10651 ( .A(n8634), .B(SI_18_), .ZN(n8632) );
  XNOR2_X1 U10652 ( .A(n8632), .B(n8357), .ZN(n10475) );
  NAND2_X1 U10653 ( .A1(n10475), .A2(n8534), .ZN(n8365) );
  INV_X1 U10654 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8359) );
  INV_X1 U10655 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10656 ( .A1(n8571), .A2(n8360), .ZN(n8480) );
  NOR2_X1 U10657 ( .A1(n8466), .A2(n8361), .ZN(n8382) );
  INV_X1 U10658 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10659 ( .A1(n8382), .A2(n8383), .ZN(n8406) );
  OAI21_X1 U10660 ( .B1(n8408), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10661 ( .A(n8362), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13775) );
  NOR2_X1 U10662 ( .A1(n8694), .A2(n15099), .ZN(n8363) );
  AOI21_X1 U10663 ( .B1(n13775), .B2(n9815), .A(n8363), .ZN(n8364) );
  OR2_X1 U10664 ( .A1(n8400), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8366) );
  AND2_X1 U10665 ( .A1(n8645), .A2(n8366), .ZN(n14041) );
  NAND2_X1 U10666 ( .A1(n14041), .A2(n8625), .ZN(n8373) );
  INV_X1 U10667 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10668 ( .A1(n8539), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8369) );
  INV_X1 U10669 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8367) );
  OR2_X1 U10670 ( .A1(n8542), .A2(n8367), .ZN(n8368) );
  OAI211_X1 U10671 ( .C1(n8370), .C2(n8691), .A(n8369), .B(n8368), .ZN(n8371)
         );
  INV_X1 U10672 ( .A(n8371), .ZN(n8372) );
  NAND2_X1 U10673 ( .A1(n14141), .A2(n13568), .ZN(n8823) );
  XNOR2_X1 U10674 ( .A(n8375), .B(SI_14_), .ZN(n8617) );
  NAND2_X1 U10675 ( .A1(n8617), .A2(n8374), .ZN(n8377) );
  OR2_X1 U10676 ( .A1(n8375), .A2(n9817), .ZN(n8376) );
  NAND2_X1 U10677 ( .A1(n8377), .A2(n8376), .ZN(n8381) );
  NAND2_X1 U10678 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  NAND2_X1 U10679 ( .A1(n10259), .A2(n8534), .ZN(n8387) );
  OR2_X1 U10680 ( .A1(n8382), .A2(n8251), .ZN(n8384) );
  MUX2_X1 U10681 ( .A(n8384), .B(P1_IR_REG_31__SCAN_IN), .S(n8383), .Z(n8385)
         );
  AND2_X1 U10682 ( .A1(n8385), .A2(n8406), .ZN(n11259) );
  AOI22_X1 U10683 ( .A1(n11259), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n8386) );
  OR2_X1 U10684 ( .A1(n8624), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10685 ( .A1(n8413), .A2(n8388), .ZN(n14424) );
  NAND2_X1 U10686 ( .A1(n8539), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8389) );
  OAI21_X1 U10687 ( .B1(n14424), .B2(n8698), .A(n8389), .ZN(n8393) );
  INV_X1 U10688 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10689 ( .A1(n8687), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8390) );
  OAI21_X1 U10690 ( .B1(n8691), .B2(n8391), .A(n8390), .ZN(n8392) );
  INV_X1 U10691 ( .A(n14386), .ZN(n11604) );
  NAND2_X1 U10692 ( .A1(n13412), .A2(n11604), .ZN(n8805) );
  XNOR2_X1 U10693 ( .A(n8395), .B(n8394), .ZN(n10238) );
  NAND2_X1 U10694 ( .A1(n10238), .A2(n8534), .ZN(n8398) );
  NAND2_X1 U10695 ( .A1(n8408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10696 ( .A(n8396), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U10697 ( .A1(n11254), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n8397) );
  AND2_X1 U10698 ( .A1(n8415), .A2(n8399), .ZN(n8401) );
  OR2_X1 U10699 ( .A1(n8401), .A2(n8400), .ZN(n14059) );
  AOI22_X1 U10700 ( .A1(n8697), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n8539), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10701 ( .A1(n8687), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8402) );
  OAI211_X1 U10702 ( .C1(n14059), .C2(n8698), .A(n8403), .B(n8402), .ZN(n14385) );
  INV_X1 U10703 ( .A(n14385), .ZN(n8404) );
  OR2_X1 U10704 ( .A1(n14146), .A2(n8404), .ZN(n13824) );
  NAND2_X1 U10705 ( .A1(n14146), .A2(n8404), .ZN(n8810) );
  NAND2_X1 U10706 ( .A1(n13824), .A2(n8810), .ZN(n13823) );
  XNOR2_X1 U10707 ( .A(n8405), .B(n7392), .ZN(n10160) );
  NAND2_X1 U10708 ( .A1(n10160), .A2(n8534), .ZN(n8411) );
  NAND2_X1 U10709 ( .A1(n8406), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8407) );
  MUX2_X1 U10710 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8407), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8409) );
  AND2_X1 U10711 ( .A1(n8409), .A2(n8408), .ZN(n13756) );
  AOI22_X1 U10712 ( .A1(n13756), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10713 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U10714 ( .A1(n8415), .A2(n8414), .ZN(n14393) );
  AOI22_X1 U10715 ( .A1(n8697), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8687), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10716 ( .A1(n8539), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8416) );
  OAI211_X1 U10717 ( .C1(n14393), .C2(n8698), .A(n8417), .B(n8416), .ZN(n14414) );
  INV_X1 U10718 ( .A(n14414), .ZN(n13820) );
  XNOR2_X1 U10719 ( .A(n14149), .B(n13820), .ZN(n11612) );
  OR2_X1 U10720 ( .A1(n8418), .A2(n7396), .ZN(n8419) );
  NAND2_X1 U10721 ( .A1(n8420), .A2(n8419), .ZN(n10054) );
  NAND2_X1 U10722 ( .A1(n10054), .A2(n8534), .ZN(n8427) );
  NAND2_X1 U10723 ( .A1(n8602), .A2(n8421), .ZN(n8439) );
  OAI21_X1 U10724 ( .B1(n8588), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8423) );
  INV_X1 U10725 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10726 ( .A1(n8423), .A2(n8422), .ZN(n8618) );
  OR2_X1 U10727 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  NAND2_X1 U10728 ( .A1(n8618), .A2(n8424), .ZN(n13743) );
  OAI22_X1 U10729 ( .A1(n13743), .A2(n8326), .B1(n8694), .B2(n10055), .ZN(
        n8425) );
  INV_X1 U10730 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U10731 ( .A1(n8539), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8434) );
  INV_X1 U10732 ( .A(n8622), .ZN(n8430) );
  NAND2_X1 U10733 ( .A1(n8594), .A2(n8428), .ZN(n8429) );
  NAND2_X1 U10734 ( .A1(n8430), .A2(n8429), .ZN(n14410) );
  OR2_X1 U10735 ( .A1(n8676), .A2(n14410), .ZN(n8433) );
  INV_X1 U10736 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10227) );
  OR2_X1 U10737 ( .A1(n8542), .A2(n10227), .ZN(n8432) );
  INV_X1 U10738 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10221) );
  OR2_X1 U10739 ( .A1(n8691), .A2(n10221), .ZN(n8431) );
  NAND4_X1 U10740 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n14361) );
  XNOR2_X1 U10741 ( .A(n14406), .B(n14361), .ZN(n11418) );
  NAND2_X1 U10742 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  NAND2_X1 U10743 ( .A1(n8438), .A2(n8437), .ZN(n9819) );
  NAND2_X1 U10744 ( .A1(n9819), .A2(n8534), .ZN(n8442) );
  NAND2_X1 U10745 ( .A1(n8439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8440) );
  XNOR2_X1 U10746 ( .A(n8440), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U10747 ( .A1(n13731), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10748 ( .A1(n8539), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8448) );
  INV_X1 U10749 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8443) );
  OR2_X1 U10750 ( .A1(n8691), .A2(n8443), .ZN(n8447) );
  OR2_X1 U10751 ( .A1(n8607), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10752 ( .A1(n8592), .A2(n8444), .ZN(n11502) );
  OR2_X1 U10753 ( .A1(n8698), .A2(n11502), .ZN(n8446) );
  INV_X1 U10754 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10004) );
  OR2_X1 U10755 ( .A1(n8542), .A2(n10004), .ZN(n8445) );
  NAND4_X1 U10756 ( .A1(n8448), .A2(n8447), .A3(n8446), .A4(n8445), .ZN(n13617) );
  INV_X1 U10757 ( .A(n13617), .ZN(n11490) );
  XNOR2_X1 U10758 ( .A(n11492), .B(n11490), .ZN(n11110) );
  XNOR2_X1 U10759 ( .A(n8450), .B(n8449), .ZN(n9806) );
  NAND2_X1 U10760 ( .A1(n9806), .A2(n8534), .ZN(n8456) );
  NAND2_X1 U10761 ( .A1(n8468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8451) );
  MUX2_X1 U10762 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8451), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n8453) );
  INV_X1 U10763 ( .A(n8602), .ZN(n8452) );
  NAND2_X1 U10764 ( .A1(n8453), .A2(n8452), .ZN(n13715) );
  OAI22_X1 U10765 ( .A1(n13715), .A2(n8326), .B1(n8694), .B2(n9807), .ZN(n8454) );
  INV_X1 U10766 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U10767 ( .A1(n8539), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8463) );
  INV_X1 U10768 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8457) );
  OR2_X1 U10769 ( .A1(n8691), .A2(n8457), .ZN(n8462) );
  INV_X1 U10770 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8473) );
  INV_X1 U10771 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8458) );
  OAI21_X1 U10772 ( .B1(n8487), .B2(n8473), .A(n8458), .ZN(n8459) );
  NAND2_X1 U10773 ( .A1(n8459), .A2(n8608), .ZN(n11287) );
  OR2_X1 U10774 ( .A1(n8676), .A2(n11287), .ZN(n8461) );
  INV_X1 U10775 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9873) );
  OR2_X1 U10776 ( .A1(n8542), .A2(n9873), .ZN(n8460) );
  NAND4_X1 U10777 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(n13619) );
  XNOR2_X1 U10778 ( .A(n14587), .B(n11366), .ZN(n11098) );
  XNOR2_X1 U10779 ( .A(n8465), .B(n8464), .ZN(n9799) );
  NAND2_X1 U10780 ( .A1(n9799), .A2(n8534), .ZN(n8472) );
  NAND2_X1 U10781 ( .A1(n8466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8467) );
  MUX2_X1 U10782 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8467), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n8469) );
  NAND2_X1 U10783 ( .A1(n8469), .A2(n8468), .ZN(n9869) );
  OAI22_X1 U10784 ( .A1(n8694), .A2(n9801), .B1(n9869), .B2(n8326), .ZN(n8470)
         );
  INV_X1 U10785 ( .A(n8470), .ZN(n8471) );
  NAND2_X1 U10786 ( .A1(n8539), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8477) );
  INV_X1 U10787 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9825) );
  OR2_X1 U10788 ( .A1(n8691), .A2(n9825), .ZN(n8476) );
  XNOR2_X1 U10789 ( .A(n8487), .B(n8473), .ZN(n11197) );
  OR2_X1 U10790 ( .A1(n8698), .A2(n11197), .ZN(n8475) );
  INV_X1 U10791 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10732) );
  OR2_X1 U10792 ( .A1(n8542), .A2(n10732), .ZN(n8474) );
  NAND4_X1 U10793 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n13620) );
  INV_X1 U10794 ( .A(n13620), .ZN(n11186) );
  XNOR2_X1 U10795 ( .A(n11193), .B(n11186), .ZN(n10810) );
  XNOR2_X1 U10796 ( .A(n8479), .B(n8478), .ZN(n9787) );
  NAND2_X1 U10797 ( .A1(n9787), .A2(n8534), .ZN(n8483) );
  NAND2_X1 U10798 ( .A1(n8480), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8481) );
  XNOR2_X1 U10799 ( .A(n8481), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U10800 ( .A1(n8641), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9815), .B2(
        n13696), .ZN(n8482) );
  NAND2_X1 U10801 ( .A1(n8483), .A2(n8482), .ZN(n15148) );
  NAND2_X1 U10802 ( .A1(n8697), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8491) );
  INV_X1 U10803 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n8484) );
  OR2_X1 U10804 ( .A1(n8268), .A2(n8484), .ZN(n8490) );
  NAND2_X1 U10805 ( .A1(n8562), .A2(n8485), .ZN(n8486) );
  NAND2_X1 U10806 ( .A1(n8487), .A2(n8486), .ZN(n15145) );
  OR2_X1 U10807 ( .A1(n8676), .A2(n15145), .ZN(n8489) );
  INV_X1 U10808 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9858) );
  OR2_X1 U10809 ( .A1(n8542), .A2(n9858), .ZN(n8488) );
  NAND4_X1 U10810 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n13621) );
  XNOR2_X1 U10811 ( .A(n15148), .B(n13621), .ZN(n14564) );
  XNOR2_X1 U10812 ( .A(n8493), .B(n8492), .ZN(n9747) );
  NAND2_X1 U10813 ( .A1(n9747), .A2(n8534), .ZN(n8498) );
  NAND2_X1 U10814 ( .A1(n8358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8494) );
  MUX2_X1 U10815 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8494), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8496) );
  INV_X1 U10816 ( .A(n8569), .ZN(n8495) );
  AND2_X1 U10817 ( .A1(n8496), .A2(n8495), .ZN(n14493) );
  AOI22_X1 U10818 ( .A1(n8641), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9815), .B2(
        n14493), .ZN(n8497) );
  NAND2_X1 U10819 ( .A1(n8539), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8502) );
  INV_X1 U10820 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10612) );
  OR2_X1 U10821 ( .A1(n8542), .A2(n10612), .ZN(n8501) );
  OAI21_X1 U10822 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n8577), .ZN(n10969) );
  OR2_X1 U10823 ( .A1(n8676), .A2(n10969), .ZN(n8500) );
  INV_X1 U10824 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9826) );
  OR2_X1 U10825 ( .A1(n8691), .A2(n9826), .ZN(n8499) );
  OR2_X1 U10826 ( .A1(n10693), .A2(n13624), .ZN(n10385) );
  NAND2_X1 U10827 ( .A1(n10693), .A2(n13624), .ZN(n10387) );
  AND2_X1 U10828 ( .A1(n10385), .A2(n10387), .ZN(n10604) );
  NAND2_X1 U10829 ( .A1(n8539), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8506) );
  INV_X1 U10830 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10363) );
  INV_X1 U10831 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9833) );
  OR2_X1 U10832 ( .A1(n8691), .A2(n9833), .ZN(n8504) );
  OR2_X1 U10833 ( .A1(n8676), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U10834 ( .A(n8508), .B(n8507), .ZN(n9742) );
  NAND2_X1 U10835 ( .A1(n9742), .A2(n8534), .ZN(n8512) );
  NAND2_X1 U10836 ( .A1(n8509), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8510) );
  XNOR2_X1 U10837 ( .A(n8510), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U10838 ( .A1(n8641), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n9815), .B2(
        n13663), .ZN(n8511) );
  NAND2_X1 U10839 ( .A1(n10375), .A2(n8732), .ZN(n10381) );
  INV_X1 U10840 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8514) );
  INV_X1 U10841 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9830) );
  XNOR2_X1 U10842 ( .A(n8519), .B(n8518), .ZN(n9735) );
  NAND2_X1 U10843 ( .A1(n9735), .A2(n8534), .ZN(n8524) );
  OR2_X1 U10844 ( .A1(n7208), .A2(n8251), .ZN(n8521) );
  XNOR2_X1 U10845 ( .A(n8521), .B(n8520), .ZN(n13650) );
  OR2_X1 U10846 ( .A1(n8326), .A2(n13650), .ZN(n8523) );
  INV_X1 U10847 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9736) );
  OR2_X1 U10848 ( .A1(n8694), .A2(n9736), .ZN(n8522) );
  AND3_X2 U10849 ( .A1(n8524), .A2(n8523), .A3(n8522), .ZN(n10355) );
  NAND2_X1 U10850 ( .A1(n13626), .A2(n10355), .ZN(n8527) );
  NAND2_X1 U10851 ( .A1(n8539), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8530) );
  INV_X1 U10852 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9847) );
  OR2_X1 U10853 ( .A1(n8542), .A2(n9847), .ZN(n8529) );
  XNOR2_X1 U10854 ( .A(n8532), .B(n8531), .ZN(n9776) );
  INV_X1 U10855 ( .A(n9776), .ZN(n8533) );
  NAND2_X1 U10856 ( .A1(n8534), .A2(n8533), .ZN(n8538) );
  NAND2_X1 U10857 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8535) );
  MUX2_X1 U10858 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8535), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8537) );
  INV_X1 U10859 ( .A(n7208), .ZN(n8536) );
  NAND2_X1 U10860 ( .A1(n8537), .A2(n8536), .ZN(n13631) );
  INV_X1 U10861 ( .A(n10308), .ZN(n8719) );
  NAND2_X1 U10862 ( .A1(n8539), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8547) );
  INV_X1 U10863 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8540) );
  OR2_X1 U10864 ( .A1(n8676), .A2(n8540), .ZN(n8546) );
  INV_X1 U10865 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8541) );
  OR2_X1 U10866 ( .A1(n8542), .A2(n8541), .ZN(n8545) );
  INV_X1 U10867 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8543) );
  OR2_X1 U10868 ( .A1(n8691), .A2(n8543), .ZN(n8544) );
  INV_X1 U10869 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U10870 ( .A1(n9771), .A2(SI_0_), .ZN(n8549) );
  INV_X1 U10871 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10872 ( .A1(n8549), .A2(n8548), .ZN(n8551) );
  NAND2_X1 U10873 ( .A1(n8551), .A2(n8550), .ZN(n14201) );
  MUX2_X1 U10874 ( .A(n14476), .B(n14201), .S(n8326), .Z(n10669) );
  NAND2_X1 U10875 ( .A1(n13628), .A2(n10669), .ZN(n8552) );
  NAND2_X1 U10876 ( .A1(n10312), .A2(n8552), .ZN(n10405) );
  INV_X1 U10877 ( .A(n10405), .ZN(n8553) );
  NAND2_X1 U10878 ( .A1(n8719), .A2(n8553), .ZN(n8554) );
  NOR4_X1 U10879 ( .A1(n10604), .A2(n10381), .A3(n10353), .A4(n8554), .ZN(
        n8585) );
  XNOR2_X1 U10880 ( .A(n8556), .B(n8555), .ZN(n9783) );
  NAND2_X1 U10881 ( .A1(n9783), .A2(n8534), .ZN(n8559) );
  OR2_X1 U10882 ( .A1(n8571), .A2(n8251), .ZN(n8557) );
  XNOR2_X1 U10883 ( .A(n8557), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U10884 ( .A1(n8641), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9815), .B2(
        n9888), .ZN(n8558) );
  NAND2_X1 U10885 ( .A1(n8559), .A2(n8558), .ZN(n10786) );
  NAND2_X1 U10886 ( .A1(n8697), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8566) );
  INV_X1 U10887 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8560) );
  OR2_X1 U10888 ( .A1(n8268), .A2(n8560), .ZN(n8565) );
  OR2_X1 U10889 ( .A1(n8578), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10890 ( .A1(n8562), .A2(n8561), .ZN(n10784) );
  OR2_X1 U10891 ( .A1(n8676), .A2(n10784), .ZN(n8564) );
  INV_X1 U10892 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10397) );
  OR2_X1 U10893 ( .A1(n8542), .A2(n10397), .ZN(n8563) );
  NAND4_X1 U10894 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n13622) );
  XNOR2_X1 U10895 ( .A(n10786), .B(n13622), .ZN(n10396) );
  XNOR2_X1 U10896 ( .A(n8568), .B(n8567), .ZN(n9755) );
  NAND2_X1 U10897 ( .A1(n9755), .A2(n8534), .ZN(n8574) );
  NOR2_X1 U10898 ( .A1(n8569), .A2(n8251), .ZN(n8570) );
  MUX2_X1 U10899 ( .A(n8251), .B(n8570), .S(P1_IR_REG_5__SCAN_IN), .Z(n8572)
         );
  OR2_X1 U10900 ( .A1(n8572), .A2(n8571), .ZN(n13679) );
  INV_X1 U10901 ( .A(n13679), .ZN(n13674) );
  AOI22_X1 U10902 ( .A1(n8641), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9815), .B2(
        n13674), .ZN(n8573) );
  NAND2_X1 U10903 ( .A1(n8539), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8583) );
  INV_X1 U10904 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8575) );
  OR2_X1 U10905 ( .A1(n8691), .A2(n8575), .ZN(n8582) );
  AND2_X1 U10906 ( .A1(n8577), .A2(n8576), .ZN(n8579) );
  OR2_X1 U10907 ( .A1(n8579), .A2(n8578), .ZN(n10791) );
  OR2_X1 U10908 ( .A1(n8676), .A2(n10791), .ZN(n8581) );
  INV_X1 U10909 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9853) );
  OR2_X1 U10910 ( .A1(n8542), .A2(n9853), .ZN(n8580) );
  NAND4_X1 U10911 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n13623) );
  NAND2_X1 U10912 ( .A1(n14557), .A2(n13623), .ZN(n8584) );
  NAND2_X1 U10913 ( .A1(n10390), .A2(n8584), .ZN(n10389) );
  NAND4_X1 U10914 ( .A1(n14564), .A2(n8585), .A3(n10396), .A4(n10389), .ZN(
        n8586) );
  NOR4_X1 U10915 ( .A1(n11110), .A2(n11098), .A3(n10810), .A4(n8586), .ZN(
        n8615) );
  XNOR2_X1 U10916 ( .A(n8587), .B(n7393), .ZN(n9949) );
  NAND2_X1 U10917 ( .A1(n9949), .A2(n8534), .ZN(n8591) );
  NAND2_X1 U10918 ( .A1(n8588), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10919 ( .A(n8589), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U10920 ( .A1(n10228), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U10921 ( .A1(n8539), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10922 ( .A1(n8592), .A2(n10016), .ZN(n8593) );
  NAND2_X1 U10923 ( .A1(n8594), .A2(n8593), .ZN(n14382) );
  OR2_X1 U10924 ( .A1(n8676), .A2(n14382), .ZN(n8597) );
  INV_X1 U10925 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11223) );
  OR2_X1 U10926 ( .A1(n8542), .A2(n11223), .ZN(n8596) );
  INV_X1 U10927 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10012) );
  OR2_X1 U10928 ( .A1(n8691), .A2(n10012), .ZN(n8595) );
  NAND4_X1 U10929 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n14253) );
  OR2_X1 U10930 ( .A1(n14238), .A2(n14253), .ZN(n11416) );
  NAND2_X1 U10931 ( .A1(n14238), .A2(n14253), .ZN(n8599) );
  NAND2_X1 U10932 ( .A1(n11416), .A2(n8599), .ZN(n11410) );
  XNOR2_X1 U10933 ( .A(n8601), .B(n8600), .ZN(n9810) );
  NAND2_X1 U10934 ( .A1(n9810), .A2(n8534), .ZN(n8605) );
  OR2_X1 U10935 ( .A1(n8602), .A2(n8251), .ZN(n8603) );
  XNOR2_X1 U10936 ( .A(n8603), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U10937 ( .A1(n10011), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10938 ( .A1(n8539), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8614) );
  INV_X1 U10939 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8606) );
  OR2_X1 U10940 ( .A1(n8691), .A2(n8606), .ZN(n8613) );
  INV_X1 U10941 ( .A(n8607), .ZN(n8610) );
  NAND2_X1 U10942 ( .A1(n8608), .A2(n9882), .ZN(n8609) );
  NAND2_X1 U10943 ( .A1(n8610), .A2(n8609), .ZN(n11139) );
  OR2_X1 U10944 ( .A1(n8676), .A2(n11139), .ZN(n8612) );
  INV_X1 U10945 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9876) );
  OR2_X1 U10946 ( .A1(n8542), .A2(n9876), .ZN(n8611) );
  NAND4_X1 U10947 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n13618) );
  XNOR2_X1 U10948 ( .A(n11358), .B(n13618), .ZN(n11137) );
  NAND4_X1 U10949 ( .A1(n11418), .A2(n8615), .A3(n11410), .A4(n11137), .ZN(
        n8630) );
  XNOR2_X1 U10950 ( .A(n8617), .B(n8616), .ZN(n10205) );
  NAND2_X1 U10951 ( .A1(n10205), .A2(n8534), .ZN(n8621) );
  NAND2_X1 U10952 ( .A1(n8618), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8619) );
  XNOR2_X1 U10953 ( .A(n8619), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U10954 ( .A1(n11249), .A2(n9815), .B1(n8641), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8620) );
  NOR2_X1 U10955 ( .A1(n8622), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8623) );
  OR2_X1 U10956 ( .A1(n8624), .A2(n8623), .ZN(n14368) );
  INV_X1 U10957 ( .A(n14368), .ZN(n11423) );
  NAND2_X1 U10958 ( .A1(n11423), .A2(n8625), .ZN(n8629) );
  NAND2_X1 U10959 ( .A1(n8697), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10960 ( .A1(n8539), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8627) );
  INV_X1 U10961 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10226) );
  OR2_X1 U10962 ( .A1(n8542), .A2(n10226), .ZN(n8626) );
  NAND4_X1 U10963 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(n14416) );
  INV_X1 U10964 ( .A(n14416), .ZN(n14396) );
  OR2_X1 U10965 ( .A1(n14428), .A2(n14396), .ZN(n11595) );
  NAND2_X1 U10966 ( .A1(n14428), .A2(n14396), .ZN(n11596) );
  NOR4_X1 U10967 ( .A1(n13823), .A2(n11612), .A3(n8630), .A4(n11419), .ZN(
        n8653) );
  NAND2_X1 U10968 ( .A1(n8632), .A2(n8631), .ZN(n8636) );
  OR2_X1 U10969 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10970 ( .A1(n8636), .A2(n8635), .ZN(n8640) );
  NAND2_X1 U10971 ( .A1(n8638), .A2(n8637), .ZN(n8639) );
  NAND2_X1 U10972 ( .A1(n10595), .A2(n8534), .ZN(n8643) );
  AOI22_X1 U10973 ( .A1(n8641), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11138), 
        .B2(n9815), .ZN(n8642) );
  NAND2_X1 U10974 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U10975 ( .A1(n8647), .A2(n8646), .ZN(n14026) );
  OR2_X1 U10976 ( .A1(n14026), .A2(n8698), .ZN(n8652) );
  INV_X1 U10977 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13770) );
  NAND2_X1 U10978 ( .A1(n8687), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U10979 ( .A1(n8539), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8648) );
  OAI211_X1 U10980 ( .C1(n8691), .C2(n13770), .A(n8649), .B(n8648), .ZN(n8650)
         );
  INV_X1 U10981 ( .A(n8650), .ZN(n8651) );
  NAND2_X1 U10982 ( .A1(n8652), .A2(n8651), .ZN(n14001) );
  XNOR2_X1 U10983 ( .A(n14134), .B(n14001), .ZN(n14019) );
  NAND4_X1 U10984 ( .A1(n6521), .A2(n11625), .A3(n8653), .A4(n14019), .ZN(
        n8654) );
  NOR4_X1 U10985 ( .A1(n13974), .A2(n14013), .A3(n13986), .A4(n8654), .ZN(
        n8681) );
  XNOR2_X1 U10986 ( .A(n8656), .B(n8655), .ZN(n11554) );
  NAND2_X1 U10987 ( .A1(n11554), .A2(n8534), .ZN(n8658) );
  OR2_X1 U10988 ( .A1(n8694), .A2(n11555), .ZN(n8657) );
  NAND2_X1 U10989 ( .A1(n8697), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8667) );
  INV_X1 U10990 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8659) );
  OR2_X1 U10991 ( .A1(n8268), .A2(n8659), .ZN(n8666) );
  INV_X1 U10992 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10993 ( .A1(n8675), .A2(n8660), .ZN(n8661) );
  NAND2_X1 U10994 ( .A1(n8662), .A2(n8661), .ZN(n13940) );
  OR2_X1 U10995 ( .A1(n8698), .A2(n13940), .ZN(n8665) );
  INV_X1 U10996 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8663) );
  OR2_X1 U10997 ( .A1(n8542), .A2(n8663), .ZN(n8664) );
  NAND4_X1 U10998 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n13837) );
  XNOR2_X1 U10999 ( .A(n14106), .B(n13837), .ZN(n13931) );
  XNOR2_X1 U11000 ( .A(n8668), .B(SI_23_), .ZN(n11274) );
  NAND2_X1 U11001 ( .A1(n11274), .A2(n8534), .ZN(n8670) );
  INV_X1 U11002 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11277) );
  OR2_X1 U11003 ( .A1(n8694), .A2(n11277), .ZN(n8669) );
  NAND2_X1 U11004 ( .A1(n8697), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8680) );
  INV_X1 U11005 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11006 ( .A1(n8268), .A2(n8671), .ZN(n8679) );
  INV_X1 U11007 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11008 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U11009 ( .A1(n8675), .A2(n8674), .ZN(n13953) );
  OR2_X1 U11010 ( .A1(n8676), .A2(n13953), .ZN(n8678) );
  INV_X1 U11011 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13957) );
  OR2_X1 U11012 ( .A1(n8542), .A2(n13957), .ZN(n8677) );
  NAND4_X1 U11013 ( .A1(n8680), .A2(n8679), .A3(n8678), .A4(n8677), .ZN(n13934) );
  XNOR2_X1 U11014 ( .A(n14112), .B(n13934), .ZN(n13961) );
  NAND4_X1 U11015 ( .A1(n13812), .A2(n8681), .A3(n13931), .A4(n13961), .ZN(
        n8682) );
  NOR4_X1 U11016 ( .A1(n13862), .A2(n13876), .A3(n13904), .A4(n8682), .ZN(
        n8705) );
  NAND2_X1 U11017 ( .A1(n13363), .A2(n8534), .ZN(n8686) );
  OR2_X1 U11018 ( .A1(n8694), .A2(n14187), .ZN(n8685) );
  INV_X1 U11019 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11020 ( .A1(n8687), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11021 ( .A1(n8539), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8688) );
  OAI211_X1 U11022 ( .C1(n8691), .C2(n8690), .A(n8689), .B(n8688), .ZN(n13847)
         );
  XNOR2_X1 U11023 ( .A(n13789), .B(n13847), .ZN(n8704) );
  NAND2_X1 U11024 ( .A1(n11770), .A2(n8534), .ZN(n8696) );
  OR2_X1 U11025 ( .A1(n8694), .A2(n11771), .ZN(n8695) );
  NAND2_X1 U11026 ( .A1(n8539), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11027 ( .A1(n8697), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11028 ( .A1(n8698), .A2(n13849), .ZN(n8701) );
  INV_X1 U11029 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8699) );
  OR2_X1 U11030 ( .A1(n8542), .A2(n8699), .ZN(n8700) );
  NAND4_X1 U11031 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n13616) );
  XNOR2_X1 U11032 ( .A(n13844), .B(n13616), .ZN(n13842) );
  NAND4_X1 U11033 ( .A1(n8908), .A2(n8705), .A3(n8704), .A4(n13842), .ZN(n8706) );
  XOR2_X1 U11034 ( .A(n11138), .B(n8706), .Z(n8715) );
  NAND2_X1 U11035 ( .A1(n8711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8710) );
  INV_X1 U11036 ( .A(n8921), .ZN(n8712) );
  NAND2_X1 U11037 ( .A1(n6512), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11038 ( .A1(n10738), .A2(n9908), .ZN(n8887) );
  NAND2_X1 U11039 ( .A1(n14200), .A2(n10738), .ZN(n8716) );
  MUX2_X2 U11040 ( .A(n10323), .B(n8716), .S(n13782), .Z(n8893) );
  XNOR2_X1 U11041 ( .A(n14200), .B(n11138), .ZN(n8717) );
  NAND2_X1 U11042 ( .A1(n8717), .A2(n9908), .ZN(n8718) );
  NAND2_X1 U11043 ( .A1(n8893), .A2(n8718), .ZN(n8726) );
  XNOR2_X1 U11044 ( .A(n10312), .B(n8815), .ZN(n8720) );
  OAI211_X1 U11045 ( .C1(n10405), .C2(n10033), .A(n8720), .B(n8719), .ZN(n8725) );
  INV_X1 U11046 ( .A(n10313), .ZN(n8722) );
  INV_X1 U11047 ( .A(n10311), .ZN(n8721) );
  MUX2_X1 U11048 ( .A(n8722), .B(n8721), .S(n8726), .Z(n8723) );
  INV_X1 U11049 ( .A(n8723), .ZN(n8724) );
  NAND2_X1 U11050 ( .A1(n8725), .A2(n8724), .ZN(n8733) );
  INV_X1 U11051 ( .A(n8726), .ZN(n8815) );
  INV_X4 U11052 ( .A(n8815), .ZN(n8892) );
  AND2_X1 U11053 ( .A1(n8892), .A2(n8525), .ZN(n8729) );
  OAI211_X1 U11054 ( .C1(n10355), .C2(n8892), .A(n8732), .B(n8526), .ZN(n8727)
         );
  INV_X1 U11055 ( .A(n8727), .ZN(n8728) );
  INV_X1 U11056 ( .A(n8764), .ZN(n8891) );
  NAND2_X1 U11057 ( .A1(n13626), .A2(n8891), .ZN(n8734) );
  INV_X1 U11058 ( .A(n8729), .ZN(n8730) );
  NAND2_X1 U11059 ( .A1(n8734), .A2(n8730), .ZN(n8731) );
  NAND3_X1 U11060 ( .A1(n8733), .A2(n8732), .A3(n8731), .ZN(n8741) );
  INV_X1 U11061 ( .A(n8734), .ZN(n8739) );
  NAND2_X1 U11062 ( .A1(n13625), .A2(n8891), .ZN(n8736) );
  NAND2_X1 U11063 ( .A1(n8736), .A2(n8735), .ZN(n8738) );
  INV_X1 U11064 ( .A(n8735), .ZN(n13516) );
  NAND2_X1 U11065 ( .A1(n13625), .A2(n13516), .ZN(n8737) );
  AOI22_X1 U11066 ( .A1(n10355), .A2(n8739), .B1(n8738), .B2(n8737), .ZN(n8740) );
  MUX2_X1 U11067 ( .A(n10712), .B(n10967), .S(n8892), .Z(n8747) );
  MUX2_X1 U11069 ( .A(n13624), .B(n10693), .S(n8891), .Z(n8746) );
  NAND2_X1 U11070 ( .A1(n8747), .A2(n8746), .ZN(n8745) );
  INV_X1 U11071 ( .A(n10375), .ZN(n8743) );
  NAND2_X1 U11072 ( .A1(n8743), .A2(n8891), .ZN(n8744) );
  INV_X1 U11073 ( .A(n8746), .ZN(n8749) );
  INV_X1 U11074 ( .A(n8747), .ZN(n8748) );
  NAND2_X1 U11075 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  MUX2_X1 U11076 ( .A(n13623), .B(n14557), .S(n8892), .Z(n8756) );
  NAND2_X1 U11077 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  MUX2_X1 U11078 ( .A(n13623), .B(n14557), .S(n8891), .Z(n8753) );
  NAND2_X1 U11079 ( .A1(n8754), .A2(n8753), .ZN(n8760) );
  INV_X1 U11080 ( .A(n8755), .ZN(n8758) );
  INV_X1 U11081 ( .A(n8756), .ZN(n8757) );
  NAND2_X1 U11082 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  MUX2_X1 U11083 ( .A(n13622), .B(n10786), .S(n8880), .Z(n8762) );
  MUX2_X1 U11084 ( .A(n13622), .B(n10786), .S(n8892), .Z(n8761) );
  INV_X1 U11085 ( .A(n8762), .ZN(n8763) );
  MUX2_X1 U11086 ( .A(n13621), .B(n15148), .S(n8892), .Z(n8768) );
  NAND2_X1 U11087 ( .A1(n8767), .A2(n8768), .ZN(n8766) );
  INV_X1 U11088 ( .A(n8764), .ZN(n8880) );
  MUX2_X1 U11089 ( .A(n13621), .B(n15148), .S(n8880), .Z(n8765) );
  NAND2_X1 U11090 ( .A1(n8766), .A2(n8765), .ZN(n8772) );
  INV_X1 U11091 ( .A(n8767), .ZN(n8770) );
  INV_X1 U11092 ( .A(n8768), .ZN(n8769) );
  NAND2_X1 U11093 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  MUX2_X1 U11094 ( .A(n13620), .B(n11193), .S(n8880), .Z(n8774) );
  MUX2_X1 U11095 ( .A(n13620), .B(n11193), .S(n8892), .Z(n8773) );
  MUX2_X1 U11096 ( .A(n13619), .B(n14587), .S(n8892), .Z(n8778) );
  NAND2_X1 U11097 ( .A1(n8777), .A2(n8778), .ZN(n8776) );
  MUX2_X1 U11098 ( .A(n13619), .B(n14587), .S(n8880), .Z(n8775) );
  NAND2_X1 U11099 ( .A1(n8776), .A2(n8775), .ZN(n8782) );
  INV_X1 U11100 ( .A(n8777), .ZN(n8780) );
  INV_X1 U11101 ( .A(n8778), .ZN(n8779) );
  NAND2_X1 U11102 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  MUX2_X1 U11103 ( .A(n13618), .B(n11358), .S(n8880), .Z(n8784) );
  MUX2_X1 U11104 ( .A(n13618), .B(n11358), .S(n8892), .Z(n8783) );
  INV_X1 U11105 ( .A(n8784), .ZN(n8785) );
  MUX2_X1 U11106 ( .A(n13617), .B(n11492), .S(n8892), .Z(n8789) );
  NAND2_X1 U11107 ( .A1(n8788), .A2(n8789), .ZN(n8787) );
  MUX2_X1 U11108 ( .A(n13617), .B(n11492), .S(n8880), .Z(n8786) );
  NAND2_X1 U11109 ( .A1(n8787), .A2(n8786), .ZN(n8793) );
  INV_X1 U11110 ( .A(n8788), .ZN(n8791) );
  INV_X1 U11111 ( .A(n8789), .ZN(n8790) );
  NAND2_X1 U11112 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  NAND2_X1 U11113 ( .A1(n8793), .A2(n8792), .ZN(n8795) );
  MUX2_X1 U11114 ( .A(n14253), .B(n14238), .S(n8880), .Z(n8796) );
  MUX2_X1 U11115 ( .A(n14253), .B(n14238), .S(n8892), .Z(n8794) );
  INV_X1 U11116 ( .A(n8796), .ZN(n8797) );
  MUX2_X1 U11117 ( .A(n14361), .B(n14406), .S(n8892), .Z(n8799) );
  INV_X1 U11118 ( .A(n14361), .ZN(n13397) );
  INV_X1 U11119 ( .A(n14406), .ZN(n14434) );
  MUX2_X1 U11120 ( .A(n13397), .B(n14434), .S(n8880), .Z(n8798) );
  AOI21_X1 U11121 ( .B1(n8802), .B2(n8801), .A(n11419), .ZN(n8804) );
  AOI21_X1 U11122 ( .B1(n11598), .B2(n11595), .A(n8892), .ZN(n8803) );
  OAI21_X1 U11123 ( .B1(n8804), .B2(n8803), .A(n8805), .ZN(n8807) );
  NAND2_X1 U11124 ( .A1(n8805), .A2(n11596), .ZN(n8806) );
  AND2_X1 U11125 ( .A1(n14414), .A2(n8892), .ZN(n8808) );
  AOI21_X1 U11126 ( .B1(n14149), .B2(n8891), .A(n8808), .ZN(n8809) );
  NAND3_X1 U11127 ( .A1(n13824), .A2(n8810), .A3(n8809), .ZN(n8820) );
  XNOR2_X1 U11128 ( .A(n14146), .B(n14385), .ZN(n8811) );
  MUX2_X1 U11129 ( .A(n14414), .B(n14149), .S(n8892), .Z(n8814) );
  NAND2_X1 U11130 ( .A1(n8811), .A2(n8814), .ZN(n8813) );
  INV_X1 U11131 ( .A(n11598), .ZN(n8812) );
  AOI22_X1 U11132 ( .A1(n8820), .A2(n8813), .B1(n8812), .B2(n8892), .ZN(n8822)
         );
  INV_X1 U11133 ( .A(n8814), .ZN(n8819) );
  AND2_X1 U11134 ( .A1(n14385), .A2(n8891), .ZN(n8817) );
  OAI21_X1 U11135 ( .B1(n8815), .B2(n14385), .A(n14146), .ZN(n8816) );
  OAI21_X1 U11136 ( .B1(n8817), .B2(n14146), .A(n8816), .ZN(n8818) );
  OAI21_X1 U11137 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  MUX2_X1 U11138 ( .A(n8823), .B(n13825), .S(n8880), .Z(n8824) );
  NAND2_X1 U11139 ( .A1(n14001), .A2(n8891), .ZN(n8826) );
  INV_X1 U11140 ( .A(n14001), .ZN(n13826) );
  NAND2_X1 U11141 ( .A1(n13826), .A2(n8892), .ZN(n8825) );
  MUX2_X1 U11142 ( .A(n8826), .B(n8825), .S(n14134), .Z(n8827) );
  NAND2_X1 U11143 ( .A1(n8828), .A2(n8827), .ZN(n8830) );
  MUX2_X1 U11144 ( .A(n14022), .B(n14130), .S(n8892), .Z(n8831) );
  MUX2_X1 U11145 ( .A(n14022), .B(n14130), .S(n8880), .Z(n8829) );
  INV_X1 U11146 ( .A(n8831), .ZN(n8832) );
  MUX2_X1 U11147 ( .A(n14002), .B(n14125), .S(n8880), .Z(n8836) );
  MUX2_X1 U11148 ( .A(n14002), .B(n14125), .S(n8892), .Z(n8833) );
  NAND2_X1 U11149 ( .A1(n8834), .A2(n8833), .ZN(n8840) );
  INV_X1 U11150 ( .A(n8835), .ZN(n8838) );
  INV_X1 U11151 ( .A(n8836), .ZN(n8837) );
  NAND2_X1 U11152 ( .A1(n8838), .A2(n8837), .ZN(n8839) );
  MUX2_X1 U11153 ( .A(n13984), .B(n14120), .S(n8892), .Z(n8842) );
  MUX2_X1 U11154 ( .A(n13984), .B(n14120), .S(n8880), .Z(n8841) );
  MUX2_X1 U11155 ( .A(n13934), .B(n14112), .S(n8891), .Z(n8846) );
  NAND2_X1 U11156 ( .A1(n8845), .A2(n8846), .ZN(n8844) );
  MUX2_X1 U11157 ( .A(n13934), .B(n14112), .S(n8892), .Z(n8843) );
  NAND2_X1 U11158 ( .A1(n8844), .A2(n8843), .ZN(n8850) );
  INV_X1 U11159 ( .A(n8845), .ZN(n8848) );
  INV_X1 U11160 ( .A(n8846), .ZN(n8847) );
  NAND2_X1 U11161 ( .A1(n8850), .A2(n8849), .ZN(n8853) );
  MUX2_X1 U11162 ( .A(n13837), .B(n14106), .S(n8892), .Z(n8854) );
  NAND2_X1 U11163 ( .A1(n8853), .A2(n8854), .ZN(n8852) );
  MUX2_X1 U11164 ( .A(n13837), .B(n14106), .S(n8880), .Z(n8851) );
  NAND2_X1 U11165 ( .A1(n8852), .A2(n8851), .ZN(n8858) );
  INV_X1 U11166 ( .A(n8853), .ZN(n8856) );
  INV_X1 U11167 ( .A(n8854), .ZN(n8855) );
  NAND2_X1 U11168 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  MUX2_X1 U11169 ( .A(n13933), .B(n13924), .S(n8880), .Z(n8860) );
  MUX2_X1 U11170 ( .A(n13933), .B(n13924), .S(n8892), .Z(n8859) );
  MUX2_X1 U11171 ( .A(n13839), .B(n14098), .S(n8892), .Z(n8864) );
  NAND2_X1 U11172 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  MUX2_X1 U11173 ( .A(n13839), .B(n14098), .S(n8891), .Z(n8861) );
  NAND2_X1 U11174 ( .A1(n8862), .A2(n8861), .ZN(n8868) );
  INV_X1 U11175 ( .A(n8863), .ZN(n8866) );
  INV_X1 U11176 ( .A(n8864), .ZN(n8865) );
  NAND2_X1 U11177 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  MUX2_X1 U11178 ( .A(n13817), .B(n14093), .S(n8891), .Z(n8870) );
  MUX2_X1 U11179 ( .A(n13817), .B(n14093), .S(n8892), .Z(n8869) );
  MUX2_X1 U11180 ( .A(n13851), .B(n14085), .S(n8892), .Z(n8875) );
  NAND2_X1 U11181 ( .A1(n8874), .A2(n8875), .ZN(n8873) );
  MUX2_X1 U11182 ( .A(n13851), .B(n14085), .S(n8880), .Z(n8872) );
  NAND2_X1 U11183 ( .A1(n8873), .A2(n8872), .ZN(n8879) );
  INV_X1 U11184 ( .A(n8874), .ZN(n8877) );
  INV_X1 U11185 ( .A(n8875), .ZN(n8876) );
  NAND2_X1 U11186 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  MUX2_X1 U11187 ( .A(n13616), .B(n13844), .S(n8880), .Z(n8882) );
  MUX2_X1 U11188 ( .A(n13616), .B(n13844), .S(n8892), .Z(n8881) );
  INV_X1 U11189 ( .A(n13793), .ZN(n8884) );
  MUX2_X1 U11190 ( .A(n13790), .B(n13793), .S(n8892), .Z(n8883) );
  NAND2_X1 U11191 ( .A1(n14200), .A2(n8889), .ZN(n10043) );
  OAI21_X1 U11192 ( .B1(n9908), .B2(n14200), .A(n10043), .ZN(n8886) );
  NAND2_X1 U11193 ( .A1(n10031), .A2(n11138), .ZN(n8885) );
  AND2_X1 U11194 ( .A1(n8886), .A2(n8885), .ZN(n8907) );
  INV_X1 U11195 ( .A(n8907), .ZN(n8888) );
  NAND2_X1 U11196 ( .A1(n8888), .A2(n8887), .ZN(n8900) );
  NOR2_X1 U11197 ( .A1(n8901), .A2(n8900), .ZN(n8906) );
  NAND2_X1 U11198 ( .A1(n8889), .A2(n9908), .ZN(n9918) );
  OAI21_X1 U11199 ( .B1(n13793), .B2(n9918), .A(n13847), .ZN(n8890) );
  MUX2_X1 U11200 ( .A(n8890), .B(n14071), .S(n8892), .Z(n8905) );
  INV_X1 U11201 ( .A(n8905), .ZN(n8899) );
  NAND2_X1 U11202 ( .A1(n13789), .A2(n8891), .ZN(n8897) );
  NAND2_X1 U11203 ( .A1(n13793), .A2(n8892), .ZN(n8894) );
  NAND2_X1 U11204 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  NAND2_X1 U11205 ( .A1(n8895), .A2(n13847), .ZN(n8896) );
  NAND2_X1 U11206 ( .A1(n8897), .A2(n8896), .ZN(n8904) );
  INV_X1 U11207 ( .A(n8904), .ZN(n8898) );
  OR2_X1 U11208 ( .A1(n8899), .A2(n8898), .ZN(n8909) );
  NAND3_X1 U11209 ( .A1(n8917), .A2(n8906), .A3(n8909), .ZN(n8914) );
  NOR2_X1 U11210 ( .A1(n8908), .A2(n8900), .ZN(n8903) );
  INV_X1 U11211 ( .A(n8901), .ZN(n8902) );
  MUX2_X1 U11212 ( .A(n8907), .B(n8903), .S(n8902), .Z(n8912) );
  NOR2_X1 U11213 ( .A1(n8905), .A2(n8904), .ZN(n8916) );
  NAND2_X1 U11214 ( .A1(n8906), .A2(n8916), .ZN(n8910) );
  NAND2_X1 U11215 ( .A1(n8908), .A2(n8907), .ZN(n8915) );
  NAND3_X1 U11216 ( .A1(n7386), .A2(n8914), .A3(n8913), .ZN(n8919) );
  NOR3_X1 U11217 ( .A1(n8917), .A2(n8916), .A3(n8915), .ZN(n8918) );
  NOR2_X1 U11218 ( .A1(n8919), .A2(n8918), .ZN(n8941) );
  NAND2_X1 U11219 ( .A1(n8921), .A2(n8920), .ZN(n8925) );
  NAND2_X1 U11220 ( .A1(n8925), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8923) );
  XNOR2_X1 U11221 ( .A(n8923), .B(n8922), .ZN(n10706) );
  INV_X1 U11222 ( .A(n10706), .ZN(n8924) );
  NAND2_X1 U11223 ( .A1(n8924), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11275) );
  INV_X1 U11224 ( .A(n8925), .ZN(n8926) );
  NAND2_X1 U11225 ( .A1(n8926), .A2(n8922), .ZN(n8931) );
  INV_X1 U11226 ( .A(n8928), .ZN(n8929) );
  OAI21_X1 U11227 ( .B1(n8711), .B2(n8929), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8930) );
  XNOR2_X1 U11228 ( .A(n8930), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9803) );
  INV_X1 U11229 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8932) );
  INV_X1 U11230 ( .A(n10043), .ZN(n9916) );
  NAND2_X1 U11231 ( .A1(n10602), .A2(n13782), .ZN(n10029) );
  NAND2_X1 U11232 ( .A1(n9916), .A2(n10029), .ZN(n8936) );
  NAND2_X1 U11233 ( .A1(n10707), .A2(n9797), .ZN(n10301) );
  INV_X1 U11234 ( .A(n8937), .ZN(n13642) );
  NAND2_X1 U11235 ( .A1(n9916), .A2(n13642), .ZN(n13949) );
  NOR3_X1 U11236 ( .A1(n10301), .A2(n14191), .A3(n13949), .ZN(n8939) );
  OAI21_X1 U11237 ( .B1(n11275), .B2(n14200), .A(P1_B_REG_SCAN_IN), .ZN(n8938)
         );
  OR2_X1 U11238 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  OAI21_X1 U11239 ( .B1(n8941), .B2(n11275), .A(n8940), .ZN(P1_U3242) );
  INV_X1 U11240 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U11241 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12328), .ZN(n8975) );
  INV_X1 U11242 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8942) );
  AOI22_X1 U11243 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n8942), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n12328), .ZN(n9033) );
  INV_X1 U11244 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14514) );
  INV_X1 U11245 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12306) );
  XOR2_X1 U11246 ( .A(n14514), .B(n12306), .Z(n8977) );
  INV_X1 U11247 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n8972) );
  INV_X1 U11248 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8969) );
  INV_X1 U11249 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U11250 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n8967), .ZN(n8981) );
  INV_X1 U11251 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13729) );
  XNOR2_X1 U11252 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n13712), .ZN(n8987) );
  INV_X1 U11253 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8961) );
  XOR2_X1 U11254 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n8961), .Z(n9017) );
  XNOR2_X1 U11255 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n8996) );
  NAND2_X1 U11256 ( .A1(n8996), .A2(n8997), .ZN(n8943) );
  NAND2_X1 U11257 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8945), .ZN(n8946) );
  NAND2_X1 U11258 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8947), .ZN(n8950) );
  INV_X1 U11259 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U11260 ( .A1(n8988), .A2(n8948), .ZN(n8949) );
  NAND2_X1 U11261 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8951), .ZN(n8953) );
  INV_X1 U11262 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U11263 ( .A1(n9005), .A2(n13672), .ZN(n8952) );
  INV_X1 U11264 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U11265 ( .A1(n8957), .A2(n8956), .ZN(n8959) );
  XNOR2_X1 U11266 ( .A(n8957), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11267 ( .A1(n9014), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11268 ( .A1(n8959), .A2(n8958), .ZN(n9018) );
  NAND2_X1 U11269 ( .A1(n9017), .A2(n9018), .ZN(n8960) );
  NAND2_X1 U11270 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8984), .ZN(n8964) );
  NOR2_X1 U11271 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8984), .ZN(n8963) );
  XNOR2_X1 U11272 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8982) );
  NAND2_X1 U11273 ( .A1(n8983), .A2(n8982), .ZN(n8965) );
  XNOR2_X1 U11274 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(n8969), .ZN(n9027) );
  NOR2_X1 U11275 ( .A1(n9028), .A2(n9027), .ZN(n8968) );
  AOI21_X1 U11276 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n8969), .A(n8968), .ZN(
        n8979) );
  INV_X1 U11277 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U11278 ( .A(n8970), .B(n8972), .ZN(n8978) );
  NAND2_X1 U11279 ( .A1(n8979), .A2(n8978), .ZN(n8971) );
  NOR2_X1 U11280 ( .A1(n8977), .A2(n8976), .ZN(n8973) );
  AOI21_X1 U11281 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n14514), .A(n8973), .ZN(
        n9032) );
  NAND2_X1 U11282 ( .A1(n9033), .A2(n9032), .ZN(n8974) );
  NAND2_X1 U11283 ( .A1(n8975), .A2(n8974), .ZN(n9037) );
  XNOR2_X1 U11284 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9037), .ZN(n9038) );
  XNOR2_X1 U11285 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9038), .ZN(n14266) );
  XOR2_X1 U11286 ( .A(n8977), .B(n8976), .Z(n14468) );
  XNOR2_X1 U11287 ( .A(n8979), .B(n8978), .ZN(n14464) );
  XNOR2_X1 U11288 ( .A(n8981), .B(n8980), .ZN(n9025) );
  XNOR2_X1 U11289 ( .A(n8983), .B(n8982), .ZN(n14452) );
  XNOR2_X1 U11290 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n8984), .ZN(n8985) );
  XNOR2_X1 U11291 ( .A(n8985), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14236) );
  XOR2_X1 U11292 ( .A(n8987), .B(n8986), .Z(n9022) );
  XNOR2_X1 U11293 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n8988), .ZN(n8990) );
  INV_X1 U11294 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11295 ( .A1(n8990), .A2(n8989), .ZN(n9004) );
  XNOR2_X1 U11296 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8990), .ZN(n15159) );
  XNOR2_X1 U11297 ( .A(n8991), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n9002) );
  AND2_X1 U11298 ( .A1(n8994), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n8995) );
  OAI21_X1 U11299 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n8993), .A(n8992), .ZN(
        n15163) );
  NAND2_X1 U11300 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15163), .ZN(n15172) );
  XOR2_X1 U11301 ( .A(n8997), .B(n8996), .Z(n8998) );
  NOR2_X1 U11302 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  XNOR2_X1 U11303 ( .A(n8999), .B(n8998), .ZN(n14213) );
  INV_X1 U11304 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14212) );
  NOR2_X1 U11305 ( .A1(n14213), .A2(n14212), .ZN(n14211) );
  NAND2_X1 U11306 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  INV_X1 U11307 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15168) );
  NAND2_X1 U11308 ( .A1(n15159), .A2(n15158), .ZN(n15157) );
  INV_X1 U11309 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15161) );
  NAND2_X1 U11310 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  INV_X1 U11311 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9009) );
  NOR2_X1 U11312 ( .A1(n9010), .A2(n9009), .ZN(n9013) );
  XNOR2_X1 U11313 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n9012) );
  XOR2_X1 U11314 ( .A(n9012), .B(n9011), .Z(n14218) );
  INV_X1 U11315 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9016) );
  XNOR2_X1 U11316 ( .A(n9014), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15166) );
  XNOR2_X1 U11317 ( .A(n9018), .B(n9017), .ZN(n9020) );
  NAND2_X1 U11318 ( .A1(n9019), .A2(n9020), .ZN(n9021) );
  INV_X1 U11319 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14224) );
  NOR2_X1 U11320 ( .A1(n9022), .A2(n9023), .ZN(n9024) );
  INV_X1 U11321 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14654) );
  INV_X1 U11322 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U11323 ( .A1(n9026), .A2(n9025), .ZN(n14457) );
  XOR2_X1 U11324 ( .A(n9028), .B(n9027), .Z(n9030) );
  INV_X1 U11325 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14460) );
  NAND2_X1 U11326 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  XNOR2_X1 U11327 ( .A(n9033), .B(n9032), .ZN(n9035) );
  NAND2_X1 U11328 ( .A1(n9034), .A2(n9035), .ZN(n14472) );
  INV_X1 U11329 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U11330 ( .A1(n14472), .A2(n14470), .ZN(n14265) );
  NAND2_X1 U11331 ( .A1(n14266), .A2(n14265), .ZN(n9036) );
  NOR2_X1 U11332 ( .A1(n14266), .A2(n14265), .ZN(n14264) );
  XNOR2_X1 U11333 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n9042) );
  NOR2_X1 U11334 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9037), .ZN(n9040) );
  INV_X1 U11335 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n12349) );
  NOR2_X1 U11336 ( .A1(n12349), .A2(n9038), .ZN(n9039) );
  NOR2_X1 U11337 ( .A1(n9040), .A2(n9039), .ZN(n9041) );
  XNOR2_X1 U11338 ( .A(n9042), .B(n9041), .ZN(n14205) );
  INV_X1 U11339 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U11340 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  OAI21_X1 U11341 ( .B1(n14529), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n9043), .ZN(
        n9045) );
  XNOR2_X1 U11342 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9044) );
  XNOR2_X1 U11343 ( .A(n9045), .B(n9044), .ZN(n9046) );
  NOR2_X1 U11344 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n9053) );
  NOR2_X1 U11345 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9056) );
  NOR2_X1 U11346 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n9055) );
  NOR2_X1 U11347 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9057) );
  NAND2_X1 U11348 ( .A1(n9250), .A2(n9062), .ZN(n9553) );
  NAND3_X1 U11349 ( .A1(n9541), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n9069) );
  NOR2_X1 U11350 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n9059) );
  NAND4_X1 U11351 ( .A1(n9060), .A2(n9059), .A3(n9554), .A4(n9058), .ZN(n9061)
         );
  INV_X1 U11352 ( .A(n9096), .ZN(n9067) );
  INV_X1 U11353 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9064) );
  INV_X1 U11354 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9544) );
  INV_X1 U11355 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9063) );
  NAND4_X1 U11356 ( .A1(n9064), .A2(n9544), .A3(n9063), .A4(
        P2_IR_REG_27__SCAN_IN), .ZN(n9066) );
  XNOR2_X1 U11357 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_27__SCAN_IN), .ZN(
        n9065) );
  NOR2_X1 U11358 ( .A1(n9067), .A2(n7389), .ZN(n9068) );
  XNOR2_X2 U11359 ( .A(n9071), .B(n9070), .ZN(n9967) );
  NAND2_X1 U11360 ( .A1(n9148), .A2(n9737), .ZN(n9111) );
  INV_X1 U11361 ( .A(n9111), .ZN(n9191) );
  NAND2_X1 U11362 ( .A1(n10736), .A2(n11959), .ZN(n9073) );
  INV_X1 U11363 ( .A(n9075), .ZN(n9076) );
  INV_X1 U11364 ( .A(n9077), .ZN(n9083) );
  INV_X1 U11365 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9078) );
  INV_X1 U11366 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9081) );
  INV_X1 U11367 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9247) );
  XNOR2_X1 U11368 ( .A(n9247), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U11369 ( .A1(n9083), .A2(n9082), .ZN(n9084) );
  AND2_X2 U11370 ( .A1(n9085), .A2(n9084), .ZN(n11992) );
  AOI21_X1 U11371 ( .B1(n7401), .B2(n9080), .A(n9247), .ZN(n9088) );
  INV_X2 U11372 ( .A(n9573), .ZN(n13053) );
  XNOR2_X1 U11373 ( .A(n13195), .B(n12840), .ZN(n9451) );
  NAND2_X1 U11374 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9180) );
  INV_X1 U11375 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9179) );
  NOR2_X1 U11376 ( .A1(n9180), .A2(n9179), .ZN(n9178) );
  NAND2_X1 U11377 ( .A1(n9178), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9218) );
  INV_X1 U11378 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11379 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n9090) );
  INV_X1 U11380 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U11381 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n9091) );
  NAND2_X1 U11382 ( .A1(n9398), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9426) );
  INV_X1 U11383 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9425) );
  INV_X1 U11384 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9092) );
  INV_X1 U11385 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U11386 ( .B1(n9442), .B2(n9092), .A(n12854), .ZN(n9095) );
  NAND2_X1 U11387 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n9093) );
  INV_X1 U11388 ( .A(n9457), .ZN(n9094) );
  NAND2_X1 U11389 ( .A1(n9095), .A2(n9094), .ZN(n13192) );
  XNOR2_X2 U11390 ( .A(n9097), .B(n13357), .ZN(n13365) );
  NAND2_X4 U11391 ( .A1(n9100), .A2(n9099), .ZN(n11731) );
  OR2_X1 U11392 ( .A1(n13192), .A2(n11731), .ZN(n9106) );
  NAND2_X1 U11393 ( .A1(n13365), .A2(n9099), .ZN(n9236) );
  INV_X1 U11394 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11395 ( .A1(n9530), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9102) );
  NAND2_X4 U11396 ( .A1(n9100), .A2(n11773), .ZN(n11730) );
  NAND2_X1 U11397 ( .A1(n11962), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9101) );
  OAI211_X1 U11398 ( .C1(n11741), .C2(n9103), .A(n9102), .B(n9101), .ZN(n9104)
         );
  INV_X1 U11399 ( .A(n9104), .ZN(n9105) );
  NAND2_X1 U11400 ( .A1(n9106), .A2(n9105), .ZN(n12957) );
  AND2_X1 U11401 ( .A1(n11992), .A2(n12023), .ZN(n9108) );
  NAND2_X1 U11402 ( .A1(n12957), .A2(n13221), .ZN(n9452) );
  INV_X1 U11403 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9976) );
  OR2_X1 U11404 ( .A1(n9148), .A2(n12985), .ZN(n9110) );
  XNOR2_X2 U11405 ( .A(n10931), .B(n9137), .ZN(n10282) );
  INV_X1 U11406 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10930) );
  OR2_X1 U11407 ( .A1(n11731), .A2(n10930), .ZN(n9116) );
  NAND2_X1 U11408 ( .A1(n9138), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9115) );
  INV_X1 U11409 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n12986) );
  OR2_X1 U11410 ( .A1(n9236), .A2(n12986), .ZN(n9114) );
  INV_X1 U11411 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9112) );
  OR2_X1 U11412 ( .A1(n11730), .A2(n9112), .ZN(n9113) );
  NAND2_X1 U11413 ( .A1(n12978), .A2(n9477), .ZN(n9128) );
  INV_X1 U11414 ( .A(n10277), .ZN(n9127) );
  NAND2_X1 U11415 ( .A1(n9138), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9120) );
  INV_X1 U11416 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10136) );
  OR2_X1 U11417 ( .A1(n9236), .A2(n10136), .ZN(n9119) );
  INV_X1 U11418 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9975) );
  OR2_X1 U11419 ( .A1(n11730), .A2(n9975), .ZN(n9118) );
  INV_X1 U11420 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10292) );
  INV_X1 U11421 ( .A(n12979), .ZN(n9124) );
  OAI21_X1 U11422 ( .B1(n9771), .B2(n9741), .A(n9121), .ZN(n9122) );
  NAND2_X1 U11423 ( .A1(n9123), .A2(n9122), .ZN(n13378) );
  MUX2_X1 U11424 ( .A(n9976), .B(n13378), .S(n9148), .Z(n11780) );
  OR2_X1 U11425 ( .A1(n9124), .A2(n11780), .ZN(n10276) );
  INV_X1 U11426 ( .A(n11780), .ZN(n10297) );
  OR2_X1 U11427 ( .A1(n9137), .A2(n10297), .ZN(n10269) );
  OAI21_X1 U11428 ( .B1(n13206), .B2(n10276), .A(n10269), .ZN(n9125) );
  NAND2_X1 U11429 ( .A1(n10282), .A2(n9128), .ZN(n9129) );
  NAND2_X1 U11430 ( .A1(n10270), .A2(n9129), .ZN(n9143) );
  MUX2_X1 U11431 ( .A(n9247), .B(n9130), .S(P2_IR_REG_2__SCAN_IN), .Z(n9131)
         );
  INV_X1 U11432 ( .A(n9131), .ZN(n9133) );
  NAND2_X1 U11433 ( .A1(n9133), .A2(n9132), .ZN(n9977) );
  NAND2_X1 U11434 ( .A1(n9191), .A2(n9735), .ZN(n9136) );
  OR2_X1 U11435 ( .A1(n9134), .A2(n9779), .ZN(n9135) );
  NAND2_X1 U11436 ( .A1(n9530), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9142) );
  INV_X1 U11437 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10874) );
  OR2_X1 U11438 ( .A1(n11731), .A2(n10874), .ZN(n9141) );
  OR2_X1 U11439 ( .A1(n11730), .A2(n10875), .ZN(n9140) );
  INV_X1 U11440 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9959) );
  OR2_X1 U11441 ( .A1(n9236), .A2(n9959), .ZN(n9139) );
  NAND2_X1 U11442 ( .A1(n12977), .A2(n9477), .ZN(n9145) );
  XNOR2_X1 U11443 ( .A(n9144), .B(n9145), .ZN(n10284) );
  INV_X1 U11444 ( .A(n9144), .ZN(n9146) );
  NAND2_X1 U11445 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND2_X1 U11446 ( .A1(n9132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U11447 ( .A(n9149), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U11448 ( .A1(n9433), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6435), .B2(
        n13010), .ZN(n9151) );
  NAND2_X1 U11449 ( .A1(n9742), .A2(n11959), .ZN(n9150) );
  XNOR2_X1 U11450 ( .A(n9137), .B(n14730), .ZN(n9157) );
  NAND2_X1 U11451 ( .A1(n9530), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9156) );
  OR2_X1 U11452 ( .A1(n11731), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9155) );
  INV_X1 U11453 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9152) );
  OR2_X1 U11454 ( .A1(n11730), .A2(n9152), .ZN(n9154) );
  INV_X1 U11455 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9960) );
  OR2_X1 U11456 ( .A1(n9236), .A2(n9960), .ZN(n9153) );
  NAND4_X1 U11457 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n12976) );
  AND2_X1 U11458 ( .A1(n12976), .A2(n9477), .ZN(n9158) );
  NAND2_X1 U11459 ( .A1(n9157), .A2(n9158), .ZN(n9171) );
  INV_X1 U11460 ( .A(n9157), .ZN(n10337) );
  INV_X1 U11461 ( .A(n9158), .ZN(n9159) );
  NAND2_X1 U11462 ( .A1(n10337), .A2(n9159), .ZN(n9160) );
  NAND2_X1 U11463 ( .A1(n9747), .A2(n9191), .ZN(n9166) );
  NAND2_X1 U11464 ( .A1(n9162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9161) );
  MUX2_X1 U11465 ( .A(n9161), .B(P2_IR_REG_31__SCAN_IN), .S(n9163), .Z(n9164)
         );
  NAND2_X1 U11466 ( .A1(n6766), .A2(n9163), .ZN(n9192) );
  NAND2_X1 U11467 ( .A1(n9164), .A2(n9192), .ZN(n14617) );
  INV_X1 U11468 ( .A(n14617), .ZN(n9963) );
  AOI22_X1 U11469 ( .A1(n9433), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6435), .B2(
        n9963), .ZN(n9165) );
  NAND2_X1 U11470 ( .A1(n9530), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9170) );
  INV_X1 U11471 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9962) );
  OAI21_X1 U11472 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9180), .ZN(n10907) );
  OR2_X1 U11473 ( .A1(n11731), .A2(n10907), .ZN(n9168) );
  INV_X1 U11474 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9978) );
  OR2_X1 U11475 ( .A1(n11730), .A2(n9978), .ZN(n9167) );
  NAND2_X1 U11476 ( .A1(n12975), .A2(n9477), .ZN(n9172) );
  INV_X1 U11477 ( .A(n9172), .ZN(n9173) );
  OR2_X1 U11478 ( .A1(n10467), .A2(n9173), .ZN(n9174) );
  NAND2_X1 U11479 ( .A1(n9755), .A2(n11959), .ZN(n9177) );
  NAND2_X1 U11480 ( .A1(n9192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9175) );
  XNOR2_X1 U11481 ( .A(n9175), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11482 ( .A1(n9433), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6435), .B2(
        n9979), .ZN(n9176) );
  NAND2_X1 U11483 ( .A1(n9177), .A2(n9176), .ZN(n11810) );
  XNOR2_X1 U11484 ( .A(n11810), .B(n12840), .ZN(n9187) );
  NAND2_X1 U11485 ( .A1(n9530), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9185) );
  INV_X1 U11486 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9964) );
  OR2_X1 U11487 ( .A1(n11741), .A2(n9964), .ZN(n9184) );
  INV_X1 U11488 ( .A(n9178), .ZN(n9200) );
  NAND2_X1 U11489 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U11490 ( .A1(n9200), .A2(n9181), .ZN(n10949) );
  OR2_X1 U11491 ( .A1(n11731), .A2(n10949), .ZN(n9183) );
  INV_X1 U11492 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10947) );
  OR2_X1 U11493 ( .A1(n11730), .A2(n10947), .ZN(n9182) );
  NAND4_X1 U11494 ( .A1(n9185), .A2(n9184), .A3(n9183), .A4(n9182), .ZN(n12974) );
  NAND2_X1 U11495 ( .A1(n12974), .A2(n13221), .ZN(n9188) );
  XNOR2_X1 U11496 ( .A(n9187), .B(n9188), .ZN(n10468) );
  INV_X1 U11497 ( .A(n9187), .ZN(n9189) );
  NAND2_X1 U11498 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  NAND2_X1 U11499 ( .A1(n9783), .A2(n11974), .ZN(n9197) );
  INV_X1 U11500 ( .A(n9192), .ZN(n9194) );
  INV_X1 U11501 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11502 ( .A1(n9194), .A2(n9193), .ZN(n9213) );
  NAND2_X1 U11503 ( .A1(n9213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9195) );
  XNOR2_X1 U11504 ( .A(n9195), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11505 ( .A1(n9433), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6435), .B2(
        n9991), .ZN(n9196) );
  NAND2_X1 U11506 ( .A1(n9197), .A2(n9196), .ZN(n11819) );
  XNOR2_X1 U11507 ( .A(n11819), .B(n12840), .ZN(n9207) );
  NAND2_X1 U11508 ( .A1(n9198), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9206) );
  INV_X1 U11509 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10940) );
  OR2_X1 U11510 ( .A1(n11730), .A2(n10940), .ZN(n9205) );
  INV_X1 U11511 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U11512 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  NAND2_X1 U11513 ( .A1(n9218), .A2(n9201), .ZN(n10979) );
  OR2_X1 U11514 ( .A1(n11731), .A2(n10979), .ZN(n9204) );
  INV_X1 U11515 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9202) );
  OR2_X1 U11516 ( .A1(n11966), .A2(n9202), .ZN(n9203) );
  NAND4_X1 U11517 ( .A1(n9206), .A2(n9205), .A3(n9204), .A4(n9203), .ZN(n12973) );
  INV_X2 U11518 ( .A(n9477), .ZN(n13206) );
  AND2_X1 U11519 ( .A1(n12973), .A2(n13221), .ZN(n9208) );
  NAND2_X1 U11520 ( .A1(n9207), .A2(n9208), .ZN(n9212) );
  INV_X1 U11521 ( .A(n9207), .ZN(n10760) );
  INV_X1 U11522 ( .A(n9208), .ZN(n9209) );
  NAND2_X1 U11523 ( .A1(n10760), .A2(n9209), .ZN(n9210) );
  NAND2_X1 U11524 ( .A1(n9212), .A2(n9210), .ZN(n10987) );
  INV_X1 U11525 ( .A(n10987), .ZN(n9211) );
  NAND2_X1 U11526 ( .A1(n10984), .A2(n9212), .ZN(n9229) );
  NAND2_X1 U11527 ( .A1(n9787), .A2(n11974), .ZN(n9216) );
  NAND2_X1 U11528 ( .A1(n9230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11529 ( .A(n9214), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14633) );
  AOI22_X1 U11530 ( .A1(n9433), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6435), .B2(
        n14633), .ZN(n9215) );
  NAND2_X1 U11531 ( .A1(n9216), .A2(n9215), .ZN(n14746) );
  XNOR2_X1 U11532 ( .A(n14746), .B(n12840), .ZN(n9225) );
  NAND2_X1 U11533 ( .A1(n11962), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9224) );
  INV_X1 U11534 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9966) );
  OR2_X1 U11535 ( .A1(n11741), .A2(n9966), .ZN(n9223) );
  NAND2_X1 U11536 ( .A1(n9218), .A2(n9217), .ZN(n9219) );
  NAND2_X1 U11537 ( .A1(n9257), .A2(n9219), .ZN(n11031) );
  OR2_X1 U11538 ( .A1(n11731), .A2(n11031), .ZN(n9222) );
  INV_X1 U11539 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9220) );
  OR2_X1 U11540 ( .A1(n11966), .A2(n9220), .ZN(n9221) );
  NAND4_X1 U11541 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(n12972) );
  AND2_X1 U11542 ( .A1(n12972), .A2(n9477), .ZN(n9226) );
  NAND2_X1 U11543 ( .A1(n9225), .A2(n9226), .ZN(n9242) );
  INV_X1 U11544 ( .A(n9225), .ZN(n11121) );
  INV_X1 U11545 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U11546 ( .A1(n11121), .A2(n9227), .ZN(n9228) );
  AND2_X1 U11547 ( .A1(n9242), .A2(n9228), .ZN(n10758) );
  NAND2_X1 U11548 ( .A1(n9229), .A2(n10758), .ZN(n11119) );
  NAND2_X1 U11549 ( .A1(n9799), .A2(n11974), .ZN(n9235) );
  OAI21_X1 U11550 ( .B1(n9230), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11551 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9231), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9233) );
  INV_X1 U11552 ( .A(n9248), .ZN(n9232) );
  AOI22_X1 U11553 ( .A1(n9433), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6435), .B2(
        n10166), .ZN(n9234) );
  XNOR2_X1 U11554 ( .A(n14755), .B(n12840), .ZN(n9244) );
  NAND2_X1 U11555 ( .A1(n9198), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9241) );
  INV_X1 U11556 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9237) );
  OR2_X1 U11557 ( .A1(n11966), .A2(n9237), .ZN(n9240) );
  INV_X1 U11558 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9256) );
  XNOR2_X1 U11559 ( .A(n9257), .B(n9256), .ZN(n11113) );
  OR2_X1 U11560 ( .A1(n11731), .A2(n11113), .ZN(n9239) );
  INV_X1 U11561 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10842) );
  OR2_X1 U11562 ( .A1(n11730), .A2(n10842), .ZN(n9238) );
  NAND4_X1 U11563 ( .A1(n9241), .A2(n9240), .A3(n9239), .A4(n9238), .ZN(n12971) );
  NAND2_X1 U11564 ( .A1(n12971), .A2(n13221), .ZN(n9245) );
  XNOR2_X1 U11565 ( .A(n9244), .B(n9245), .ZN(n11124) );
  AND2_X1 U11566 ( .A1(n11124), .A2(n9242), .ZN(n9243) );
  INV_X1 U11567 ( .A(n9244), .ZN(n11017) );
  NAND2_X1 U11568 ( .A1(n11017), .A2(n9245), .ZN(n9246) );
  NAND2_X1 U11569 ( .A1(n11129), .A2(n9246), .ZN(n9264) );
  NAND2_X1 U11570 ( .A1(n9806), .A2(n11974), .ZN(n9253) );
  NOR2_X1 U11571 ( .A1(n9248), .A2(n9247), .ZN(n9249) );
  MUX2_X1 U11572 ( .A(n9247), .B(n9249), .S(P2_IR_REG_9__SCAN_IN), .Z(n9251)
         );
  OR2_X1 U11573 ( .A1(n9251), .A2(n9287), .ZN(n10167) );
  INV_X1 U11574 ( .A(n10167), .ZN(n14650) );
  AOI22_X1 U11575 ( .A1(n9433), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6435), .B2(
        n14650), .ZN(n9252) );
  NAND2_X1 U11576 ( .A1(n9253), .A2(n9252), .ZN(n11834) );
  XNOR2_X1 U11577 ( .A(n11834), .B(n12840), .ZN(n9265) );
  NAND2_X1 U11578 ( .A1(n9530), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9263) );
  INV_X1 U11579 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9254) );
  OR2_X1 U11580 ( .A1(n11741), .A2(n9254), .ZN(n9262) );
  INV_X1 U11581 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9255) );
  OAI21_X1 U11582 ( .B1(n9257), .B2(n9256), .A(n9255), .ZN(n9258) );
  NAND2_X1 U11583 ( .A1(n9258), .A2(n9274), .ZN(n11011) );
  OR2_X1 U11584 ( .A1(n11731), .A2(n11011), .ZN(n9261) );
  INV_X1 U11585 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9259) );
  OR2_X1 U11586 ( .A1(n11730), .A2(n9259), .ZN(n9260) );
  NAND4_X1 U11587 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n12969) );
  NAND2_X1 U11588 ( .A1(n12969), .A2(n13221), .ZN(n9266) );
  XNOR2_X1 U11589 ( .A(n9265), .B(n9266), .ZN(n11015) );
  INV_X1 U11590 ( .A(n9265), .ZN(n9267) );
  NAND2_X1 U11591 ( .A1(n9267), .A2(n9266), .ZN(n9268) );
  NAND2_X1 U11592 ( .A1(n9810), .A2(n11974), .ZN(n9271) );
  OR2_X1 U11593 ( .A1(n9287), .A2(n9247), .ZN(n9269) );
  XNOR2_X1 U11594 ( .A(n9269), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U11595 ( .A1(n9433), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6435), 
        .B2(n10210), .ZN(n9270) );
  NAND2_X1 U11596 ( .A1(n9271), .A2(n9270), .ZN(n11843) );
  XNOR2_X1 U11597 ( .A(n11843), .B(n9529), .ZN(n9281) );
  NAND2_X1 U11598 ( .A1(n9138), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9279) );
  INV_X1 U11599 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9272) );
  OR2_X1 U11600 ( .A1(n11741), .A2(n9272), .ZN(n9278) );
  INV_X1 U11601 ( .A(n9273), .ZN(n9294) );
  NAND2_X1 U11602 ( .A1(n9274), .A2(n15122), .ZN(n9275) );
  NAND2_X1 U11603 ( .A1(n9294), .A2(n9275), .ZN(n11206) );
  OR2_X1 U11604 ( .A1(n11731), .A2(n11206), .ZN(n9277) );
  INV_X1 U11605 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10867) );
  OR2_X1 U11606 ( .A1(n11730), .A2(n10867), .ZN(n9276) );
  NAND4_X1 U11607 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n12968) );
  NAND2_X1 U11608 ( .A1(n12968), .A2(n13221), .ZN(n9282) );
  XNOR2_X1 U11609 ( .A(n9281), .B(n9282), .ZN(n11201) );
  INV_X1 U11610 ( .A(n11201), .ZN(n9280) );
  INV_X1 U11611 ( .A(n9281), .ZN(n9284) );
  INV_X1 U11612 ( .A(n9282), .ZN(n9283) );
  NAND2_X1 U11613 ( .A1(n9284), .A2(n9283), .ZN(n9285) );
  NAND2_X1 U11614 ( .A1(n9819), .A2(n11974), .ZN(n9290) );
  INV_X1 U11615 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11616 ( .A1(n9287), .A2(n9286), .ZN(n9305) );
  NAND2_X1 U11617 ( .A1(n9305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9288) );
  XNOR2_X1 U11618 ( .A(n9288), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U11619 ( .A1(n9433), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6435), 
        .B2(n11446), .ZN(n9289) );
  XNOR2_X1 U11620 ( .A(n11847), .B(n9529), .ZN(n9300) );
  NAND2_X1 U11621 ( .A1(n9198), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9299) );
  INV_X1 U11622 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9291) );
  OR2_X1 U11623 ( .A1(n11966), .A2(n9291), .ZN(n9298) );
  INV_X1 U11624 ( .A(n9292), .ZN(n9313) );
  INV_X1 U11625 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11626 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  NAND2_X1 U11627 ( .A1(n9313), .A2(n9295), .ZN(n11333) );
  OR2_X1 U11628 ( .A1(n11731), .A2(n11333), .ZN(n9297) );
  OR2_X1 U11629 ( .A1(n11730), .A2(n10208), .ZN(n9296) );
  NAND4_X1 U11630 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n12967) );
  NAND2_X1 U11631 ( .A1(n12967), .A2(n13221), .ZN(n9301) );
  NAND2_X1 U11632 ( .A1(n9300), .A2(n9301), .ZN(n11330) );
  NAND2_X1 U11633 ( .A1(n11331), .A2(n11330), .ZN(n9304) );
  INV_X1 U11634 ( .A(n9300), .ZN(n9303) );
  INV_X1 U11635 ( .A(n9301), .ZN(n9302) );
  NAND2_X1 U11636 ( .A1(n9303), .A2(n9302), .ZN(n11329) );
  NAND2_X1 U11637 ( .A1(n9304), .A2(n11329), .ZN(n11509) );
  INV_X1 U11638 ( .A(n11509), .ZN(n9326) );
  NAND2_X1 U11639 ( .A1(n9949), .A2(n11974), .ZN(n9310) );
  NAND2_X1 U11640 ( .A1(n9307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9306) );
  MUX2_X1 U11641 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9306), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9308) );
  INV_X1 U11642 ( .A(n9346), .ZN(n9328) );
  NAND2_X1 U11643 ( .A1(n9308), .A2(n9328), .ZN(n11447) );
  INV_X1 U11644 ( .A(n11447), .ZN(n13026) );
  AOI22_X1 U11645 ( .A1(n9433), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6435), 
        .B2(n13026), .ZN(n9309) );
  XNOR2_X1 U11646 ( .A(n14345), .B(n9529), .ZN(n9320) );
  NAND2_X1 U11647 ( .A1(n9198), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9319) );
  INV_X1 U11648 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11081) );
  OR2_X1 U11649 ( .A1(n11730), .A2(n11081), .ZN(n9318) );
  INV_X1 U11650 ( .A(n9311), .ZN(n9333) );
  INV_X1 U11651 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11652 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  NAND2_X1 U11653 ( .A1(n9333), .A2(n9314), .ZN(n11513) );
  OR2_X1 U11654 ( .A1(n11731), .A2(n11513), .ZN(n9317) );
  INV_X1 U11655 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9315) );
  OR2_X1 U11656 ( .A1(n11966), .A2(n9315), .ZN(n9316) );
  NAND4_X1 U11657 ( .A1(n9319), .A2(n9318), .A3(n9317), .A4(n9316), .ZN(n12966) );
  NAND2_X1 U11658 ( .A1(n12966), .A2(n13221), .ZN(n9321) );
  NAND2_X1 U11659 ( .A1(n9320), .A2(n9321), .ZN(n9327) );
  INV_X1 U11660 ( .A(n9320), .ZN(n9323) );
  INV_X1 U11661 ( .A(n9321), .ZN(n9322) );
  NAND2_X1 U11662 ( .A1(n9323), .A2(n9322), .ZN(n9324) );
  NAND2_X1 U11663 ( .A1(n9327), .A2(n9324), .ZN(n11510) );
  INV_X1 U11664 ( .A(n11510), .ZN(n9325) );
  NAND2_X1 U11665 ( .A1(n9326), .A2(n9325), .ZN(n11507) );
  NAND2_X1 U11666 ( .A1(n10054), .A2(n11974), .ZN(n9331) );
  NAND2_X1 U11667 ( .A1(n9328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9329) );
  XNOR2_X1 U11668 ( .A(n9329), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U11669 ( .A1(n9433), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11448), 
        .B2(n6435), .ZN(n9330) );
  XNOR2_X1 U11670 ( .A(n14339), .B(n9529), .ZN(n9340) );
  NAND2_X1 U11671 ( .A1(n11962), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9339) );
  INV_X1 U11672 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U11673 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  NAND2_X1 U11674 ( .A1(n9350), .A2(n9334), .ZN(n11562) );
  OR2_X1 U11675 ( .A1(n11731), .A2(n11562), .ZN(n9338) );
  INV_X1 U11676 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11449) );
  OR2_X1 U11677 ( .A1(n11741), .A2(n11449), .ZN(n9337) );
  INV_X1 U11678 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9335) );
  OR2_X1 U11679 ( .A1(n11966), .A2(n9335), .ZN(n9336) );
  NAND4_X1 U11680 ( .A1(n9339), .A2(n9338), .A3(n9337), .A4(n9336), .ZN(n12965) );
  NAND2_X1 U11681 ( .A1(n12965), .A2(n13221), .ZN(n9341) );
  XNOR2_X1 U11682 ( .A(n9340), .B(n9341), .ZN(n11560) );
  INV_X1 U11683 ( .A(n9340), .ZN(n9343) );
  INV_X1 U11684 ( .A(n9341), .ZN(n9342) );
  NAND2_X1 U11685 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  NAND2_X1 U11686 ( .A1(n10205), .A2(n11974), .ZN(n9349) );
  INV_X1 U11687 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U11688 ( .A1(n9346), .A2(n9345), .ZN(n9363) );
  NAND2_X1 U11689 ( .A1(n9363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9347) );
  XNOR2_X1 U11690 ( .A(n9347), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14672) );
  AOI22_X1 U11691 ( .A1(n14672), .A2(n6435), .B1(n9433), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9348) );
  XNOR2_X1 U11692 ( .A(n11867), .B(n9529), .ZN(n9357) );
  NAND2_X1 U11693 ( .A1(n9350), .A2(n11661), .ZN(n9351) );
  NAND2_X1 U11694 ( .A1(n9385), .A2(n9351), .ZN(n11662) );
  INV_X1 U11695 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11450) );
  OR2_X1 U11696 ( .A1(n11741), .A2(n11450), .ZN(n9354) );
  INV_X1 U11697 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9352) );
  OR2_X1 U11698 ( .A1(n11730), .A2(n9352), .ZN(n9353) );
  AND2_X1 U11699 ( .A1(n9354), .A2(n9353), .ZN(n9356) );
  NAND2_X1 U11700 ( .A1(n9530), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U11701 ( .C1(n11731), .C2(n11662), .A(n9356), .B(n9355), .ZN(
        n12964) );
  NAND2_X1 U11702 ( .A1(n12964), .A2(n13221), .ZN(n9358) );
  NAND2_X1 U11703 ( .A1(n9357), .A2(n9358), .ZN(n12930) );
  INV_X1 U11704 ( .A(n9357), .ZN(n9360) );
  INV_X1 U11705 ( .A(n9358), .ZN(n9359) );
  NAND2_X1 U11706 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  NAND2_X1 U11707 ( .A1(n12930), .A2(n9361), .ZN(n11660) );
  INV_X1 U11708 ( .A(n11660), .ZN(n9362) );
  NAND2_X1 U11709 ( .A1(n10259), .A2(n11974), .ZN(n9366) );
  OAI21_X1 U11710 ( .B1(n9363), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U11711 ( .A(n9364), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U11712 ( .A1(n14681), .A2(n6435), .B1(n9433), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9365) );
  XNOR2_X1 U11713 ( .A(n14332), .B(n12840), .ZN(n9374) );
  INV_X1 U11714 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11715 ( .A1(n9138), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11716 ( .A1(n11962), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9367) );
  OAI211_X1 U11717 ( .C1(n11741), .C2(n9369), .A(n9368), .B(n9367), .ZN(n9370)
         );
  INV_X1 U11718 ( .A(n9370), .ZN(n9372) );
  XNOR2_X1 U11719 ( .A(n9385), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n12938) );
  INV_X1 U11720 ( .A(n11731), .ZN(n9470) );
  NAND2_X1 U11721 ( .A1(n12938), .A2(n9470), .ZN(n9371) );
  NAND2_X1 U11722 ( .A1(n9372), .A2(n9371), .ZN(n12963) );
  AND2_X1 U11723 ( .A1(n12963), .A2(n13221), .ZN(n9375) );
  NAND2_X1 U11724 ( .A1(n9373), .A2(n12930), .ZN(n9376) );
  INV_X1 U11725 ( .A(n9374), .ZN(n12932) );
  INV_X1 U11726 ( .A(n9375), .ZN(n12936) );
  NAND2_X1 U11727 ( .A1(n10160), .A2(n11974), .ZN(n9382) );
  NAND2_X1 U11728 ( .A1(n9377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9378) );
  MUX2_X1 U11729 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9378), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9380) );
  AND2_X1 U11730 ( .A1(n9380), .A2(n9394), .ZN(n11444) );
  AOI22_X1 U11731 ( .A1(n9433), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6435), 
        .B2(n11444), .ZN(n9381) );
  XNOR2_X1 U11732 ( .A(n14321), .B(n9529), .ZN(n9391) );
  INV_X1 U11733 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11439) );
  INV_X1 U11734 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9384) );
  INV_X1 U11735 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9383) );
  OAI21_X1 U11736 ( .B1(n9385), .B2(n9384), .A(n9383), .ZN(n9387) );
  INV_X1 U11737 ( .A(n9386), .ZN(n9400) );
  NAND2_X1 U11738 ( .A1(n9387), .A2(n9400), .ZN(n11696) );
  OR2_X1 U11739 ( .A1(n11696), .A2(n11731), .ZN(n9389) );
  AOI22_X1 U11740 ( .A1(n9198), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9530), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n9388) );
  OAI211_X1 U11741 ( .C1(n11730), .C2(n11439), .A(n9389), .B(n9388), .ZN(
        n12962) );
  NAND2_X1 U11742 ( .A1(n12962), .A2(n13221), .ZN(n9390) );
  NAND2_X1 U11743 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  OAI21_X1 U11744 ( .B1(n9391), .B2(n9390), .A(n9392), .ZN(n11694) );
  INV_X1 U11745 ( .A(n9392), .ZN(n9393) );
  NAND2_X1 U11746 ( .A1(n10238), .A2(n11959), .ZN(n9397) );
  NAND2_X1 U11747 ( .A1(n9394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9395) );
  XNOR2_X1 U11748 ( .A(n9395), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U11749 ( .A1(n9433), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6435), 
        .B2(n11589), .ZN(n9396) );
  XNOR2_X1 U11750 ( .A(n12876), .B(n9529), .ZN(n9406) );
  INV_X1 U11751 ( .A(n9398), .ZN(n9414) );
  INV_X1 U11752 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U11753 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U11754 ( .A1(n9414), .A2(n9401), .ZN(n12873) );
  AOI22_X1 U11755 ( .A1(n9198), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9138), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n9404) );
  INV_X1 U11756 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9402) );
  OR2_X1 U11757 ( .A1(n11730), .A2(n9402), .ZN(n9403) );
  OAI211_X1 U11758 ( .C1(n12873), .C2(n11731), .A(n9404), .B(n9403), .ZN(
        n12961) );
  NAND2_X1 U11759 ( .A1(n12961), .A2(n13221), .ZN(n9405) );
  NAND2_X1 U11760 ( .A1(n9406), .A2(n9405), .ZN(n9407) );
  OAI21_X1 U11761 ( .B1(n9406), .B2(n9405), .A(n9407), .ZN(n12871) );
  INV_X1 U11762 ( .A(n9407), .ZN(n9408) );
  NOR2_X2 U11763 ( .A1(n12870), .A2(n9408), .ZN(n12905) );
  NAND2_X1 U11764 ( .A1(n10475), .A2(n11959), .ZN(n9412) );
  INV_X1 U11765 ( .A(n7401), .ZN(n9409) );
  NAND2_X1 U11766 ( .A1(n9409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9410) );
  XNOR2_X1 U11767 ( .A(n9410), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U11768 ( .A1(n9433), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n14693), 
        .B2(n6435), .ZN(n9411) );
  XNOR2_X1 U11769 ( .A(n13330), .B(n12840), .ZN(n9423) );
  INV_X1 U11770 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11771 ( .A1(n9414), .A2(n9413), .ZN(n9415) );
  NAND2_X1 U11772 ( .A1(n9426), .A2(n9415), .ZN(n13238) );
  OR2_X1 U11773 ( .A1(n13238), .A2(n11731), .ZN(n9421) );
  INV_X1 U11774 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U11775 ( .A1(n11962), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U11776 ( .A1(n9530), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9416) );
  OAI211_X1 U11777 ( .C1(n11741), .C2(n9418), .A(n9417), .B(n9416), .ZN(n9419)
         );
  INV_X1 U11778 ( .A(n9419), .ZN(n9420) );
  NAND2_X1 U11779 ( .A1(n9421), .A2(n9420), .ZN(n12960) );
  NAND2_X1 U11780 ( .A1(n12960), .A2(n13221), .ZN(n9422) );
  XNOR2_X1 U11781 ( .A(n9423), .B(n9422), .ZN(n12904) );
  INV_X1 U11782 ( .A(n9422), .ZN(n9424) );
  NAND2_X1 U11783 ( .A1(n9426), .A2(n9425), .ZN(n9427) );
  AND2_X1 U11784 ( .A1(n9442), .A2(n9427), .ZN(n13224) );
  NAND2_X1 U11785 ( .A1(n13224), .A2(n9470), .ZN(n9432) );
  INV_X1 U11786 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U11787 ( .A1(n11962), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9429) );
  INV_X1 U11788 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15042) );
  OR2_X1 U11789 ( .A1(n11966), .A2(n15042), .ZN(n9428) );
  OAI211_X1 U11790 ( .C1(n11741), .C2(n15050), .A(n9429), .B(n9428), .ZN(n9430) );
  INV_X1 U11791 ( .A(n9430), .ZN(n9431) );
  NAND2_X1 U11792 ( .A1(n9432), .A2(n9431), .ZN(n12959) );
  AND2_X1 U11793 ( .A1(n12959), .A2(n13221), .ZN(n9437) );
  NAND2_X1 U11794 ( .A1(n10595), .A2(n11959), .ZN(n9435) );
  AOI22_X1 U11795 ( .A1(n12027), .A2(n6435), .B1(n9433), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n9434) );
  XNOR2_X1 U11796 ( .A(n13326), .B(n12840), .ZN(n9436) );
  NOR2_X1 U11797 ( .A1(n9436), .A2(n9437), .ZN(n9438) );
  AOI21_X1 U11798 ( .B1(n9437), .B2(n9436), .A(n9438), .ZN(n12830) );
  INV_X1 U11799 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U11800 ( .A1(n12829), .A2(n9439), .ZN(n12891) );
  NAND2_X1 U11801 ( .A1(n10593), .A2(n11959), .ZN(n9441) );
  XNOR2_X1 U11802 ( .A(n13321), .B(n12840), .ZN(n9450) );
  XNOR2_X1 U11803 ( .A(n9442), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U11804 ( .A1(n13210), .A2(n9470), .ZN(n9448) );
  INV_X1 U11805 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11806 ( .A1(n11962), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11807 ( .A1(n9530), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9443) );
  OAI211_X1 U11808 ( .C1(n11741), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9446)
         );
  INV_X1 U11809 ( .A(n9446), .ZN(n9447) );
  NAND2_X1 U11810 ( .A1(n9448), .A2(n9447), .ZN(n12958) );
  AND2_X1 U11811 ( .A1(n12958), .A2(n9477), .ZN(n9449) );
  NOR2_X1 U11812 ( .A1(n9450), .A2(n9449), .ZN(n12887) );
  NAND2_X1 U11813 ( .A1(n9450), .A2(n9449), .ZN(n12888) );
  XNOR2_X1 U11814 ( .A(n9451), .B(n9452), .ZN(n12850) );
  XNOR2_X1 U11815 ( .A(n9454), .B(n9453), .ZN(n11095) );
  NAND2_X1 U11816 ( .A1(n11095), .A2(n11959), .ZN(n9456) );
  XNOR2_X1 U11817 ( .A(n13307), .B(n12840), .ZN(n9464) );
  NOR2_X1 U11818 ( .A1(n9457), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9458) );
  OR2_X1 U11819 ( .A1(n9468), .A2(n9458), .ZN(n12897) );
  INV_X1 U11820 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U11821 ( .A1(n9530), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11822 ( .A1(n11962), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9459) );
  OAI211_X1 U11823 ( .C1(n11741), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9462)
         );
  INV_X1 U11824 ( .A(n9462), .ZN(n9463) );
  OAI21_X1 U11825 ( .B1(n12897), .B2(n11731), .A(n9463), .ZN(n12956) );
  INV_X1 U11826 ( .A(n12956), .ZN(n11719) );
  NAND2_X1 U11827 ( .A1(n11274), .A2(n11959), .ZN(n9467) );
  XNOR2_X1 U11828 ( .A(n13159), .B(n12840), .ZN(n9479) );
  OR2_X1 U11829 ( .A1(n9468), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U11830 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n9468), .ZN(n9485) );
  AND2_X1 U11831 ( .A1(n9469), .A2(n9485), .ZN(n13160) );
  NAND2_X1 U11832 ( .A1(n13160), .A2(n9470), .ZN(n9476) );
  INV_X1 U11833 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U11834 ( .A1(n9138), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11835 ( .A1(n11962), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9471) );
  OAI211_X1 U11836 ( .C1(n11741), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9474)
         );
  INV_X1 U11837 ( .A(n9474), .ZN(n9475) );
  NAND2_X1 U11838 ( .A1(n9476), .A2(n9475), .ZN(n12955) );
  AND2_X1 U11839 ( .A1(n12955), .A2(n9477), .ZN(n9478) );
  INV_X1 U11840 ( .A(n9479), .ZN(n9480) );
  NAND2_X1 U11841 ( .A1(n11554), .A2(n11959), .ZN(n9483) );
  NAND2_X2 U11842 ( .A1(n9483), .A2(n9482), .ZN(n13296) );
  XNOR2_X1 U11843 ( .A(n13296), .B(n9529), .ZN(n12860) );
  NAND2_X1 U11844 ( .A1(n9530), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9490) );
  INV_X1 U11845 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9484) );
  OR2_X1 U11846 ( .A1(n11741), .A2(n9484), .ZN(n9489) );
  INV_X1 U11847 ( .A(n9485), .ZN(n9486) );
  NAND2_X1 U11848 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n9486), .ZN(n9498) );
  OAI21_X1 U11849 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n9486), .A(n9498), .ZN(
        n13147) );
  OR2_X1 U11850 ( .A1(n11731), .A2(n13147), .ZN(n9488) );
  INV_X1 U11851 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13148) );
  OR2_X1 U11852 ( .A1(n11730), .A2(n13148), .ZN(n9487) );
  NAND4_X1 U11853 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n12954) );
  NAND2_X1 U11854 ( .A1(n12954), .A2(n13221), .ZN(n9491) );
  NOR2_X1 U11855 ( .A1(n12860), .A2(n9491), .ZN(n9492) );
  AOI21_X1 U11856 ( .B1(n12860), .B2(n9491), .A(n9492), .ZN(n12879) );
  NAND2_X1 U11857 ( .A1(n13374), .A2(n11959), .ZN(n9494) );
  AND2_X2 U11858 ( .A1(n9494), .A2(n9493), .ZN(n13290) );
  XNOR2_X1 U11859 ( .A(n13290), .B(n9529), .ZN(n12914) );
  NAND2_X1 U11860 ( .A1(n9138), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9503) );
  INV_X1 U11861 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9495) );
  OR2_X1 U11862 ( .A1(n11741), .A2(n9495), .ZN(n9502) );
  INV_X1 U11863 ( .A(n9498), .ZN(n9496) );
  INV_X1 U11864 ( .A(n9513), .ZN(n9514) );
  INV_X1 U11865 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11866 ( .A1(n9498), .A2(n9497), .ZN(n9499) );
  NAND2_X1 U11867 ( .A1(n9514), .A2(n9499), .ZN(n13128) );
  OR2_X1 U11868 ( .A1(n11731), .A2(n13128), .ZN(n9501) );
  INV_X1 U11869 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13129) );
  OR2_X1 U11870 ( .A1(n11730), .A2(n13129), .ZN(n9500) );
  NOR2_X1 U11871 ( .A1(n12918), .A2(n13206), .ZN(n9504) );
  NAND2_X1 U11872 ( .A1(n12914), .A2(n9504), .ZN(n9521) );
  INV_X1 U11873 ( .A(n12914), .ZN(n9506) );
  INV_X1 U11874 ( .A(n9504), .ZN(n9505) );
  NAND2_X1 U11875 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  NAND2_X1 U11876 ( .A1(n9521), .A2(n9507), .ZN(n12862) );
  NAND2_X1 U11877 ( .A1(n13371), .A2(n11959), .ZN(n9511) );
  XNOR2_X1 U11878 ( .A(n13282), .B(n12840), .ZN(n9523) );
  NAND2_X1 U11879 ( .A1(n9530), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9520) );
  INV_X1 U11880 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9512) );
  OR2_X1 U11881 ( .A1(n11741), .A2(n9512), .ZN(n9519) );
  NAND2_X1 U11882 ( .A1(n9513), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9578) );
  INV_X1 U11883 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15039) );
  NAND2_X1 U11884 ( .A1(n9514), .A2(n15039), .ZN(n9515) );
  NAND2_X1 U11885 ( .A1(n9578), .A2(n9515), .ZN(n13105) );
  OR2_X1 U11886 ( .A1(n11731), .A2(n13105), .ZN(n9518) );
  INV_X1 U11887 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9516) );
  OR2_X1 U11888 ( .A1(n11730), .A2(n9516), .ZN(n9517) );
  NOR2_X1 U11889 ( .A1(n11929), .A2(n13206), .ZN(n9524) );
  XNOR2_X1 U11890 ( .A(n9523), .B(n9524), .ZN(n12916) );
  NAND2_X1 U11891 ( .A1(n11775), .A2(n11974), .ZN(n9528) );
  XNOR2_X1 U11892 ( .A(n13092), .B(n9529), .ZN(n9537) );
  NAND2_X1 U11893 ( .A1(n9530), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9535) );
  INV_X1 U11894 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9531) );
  OR2_X1 U11895 ( .A1(n11741), .A2(n9531), .ZN(n9534) );
  INV_X1 U11896 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9596) );
  XNOR2_X1 U11897 ( .A(n9578), .B(n9596), .ZN(n13088) );
  OR2_X1 U11898 ( .A1(n11731), .A2(n13088), .ZN(n9533) );
  INV_X1 U11899 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13091) );
  OR2_X1 U11900 ( .A1(n11730), .A2(n13091), .ZN(n9532) );
  NOR2_X1 U11901 ( .A1(n11934), .A2(n13206), .ZN(n9536) );
  NAND2_X1 U11902 ( .A1(n9537), .A2(n9536), .ZN(n12837) );
  OAI21_X1 U11903 ( .B1(n9537), .B2(n9536), .A(n12837), .ZN(n9538) );
  XNOR2_X1 U11904 ( .A(n9545), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9550) );
  INV_X1 U11905 ( .A(n9550), .ZN(n13375) );
  NAND2_X1 U11906 ( .A1(n9541), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9542) );
  XNOR2_X1 U11907 ( .A(n9542), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9566) );
  XOR2_X1 U11908 ( .A(n9566), .B(P2_B_REG_SCAN_IN), .Z(n9543) );
  NAND2_X1 U11909 ( .A1(n13375), .A2(n9543), .ZN(n9548) );
  NAND2_X1 U11910 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  NAND2_X1 U11911 ( .A1(n9546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9547) );
  INV_X1 U11912 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9549) );
  INV_X1 U11913 ( .A(n9552), .ZN(n13372) );
  AOI22_X1 U11914 ( .A1(n14717), .A2(n9549), .B1(n13372), .B2(n13375), .ZN(
        n9593) );
  AND2_X1 U11915 ( .A1(n9550), .A2(n9566), .ZN(n9551) );
  NAND2_X1 U11916 ( .A1(n9552), .A2(n9551), .ZN(n9733) );
  NAND2_X1 U11917 ( .A1(n9553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9555) );
  XNOR2_X1 U11918 ( .A(n9555), .B(n9554), .ZN(n11271) );
  AND2_X1 U11919 ( .A1(n9733), .A2(n11271), .ZN(n9594) );
  AND2_X1 U11920 ( .A1(n9593), .A2(n14723), .ZN(n14724) );
  NOR4_X1 U11921 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9559) );
  NOR4_X1 U11922 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9558) );
  NOR4_X1 U11923 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9557) );
  NOR4_X1 U11924 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9556) );
  NAND4_X1 U11925 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9565)
         );
  NOR2_X1 U11926 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .ZN(
        n9563) );
  NOR4_X1 U11927 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9562) );
  NOR4_X1 U11928 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9561) );
  NOR4_X1 U11929 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n9560) );
  NAND4_X1 U11930 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9564)
         );
  OAI21_X1 U11931 ( .B1(n9565), .B2(n9564), .A(n14717), .ZN(n9941) );
  NAND2_X1 U11932 ( .A1(n14724), .A2(n9941), .ZN(n10826) );
  INV_X1 U11933 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U11934 ( .A1(n14717), .A2(n14722), .ZN(n9568) );
  INV_X1 U11935 ( .A(n9566), .ZN(n11557) );
  NAND2_X1 U11936 ( .A1(n13372), .A2(n11557), .ZN(n9567) );
  INV_X1 U11937 ( .A(n9944), .ZN(n9569) );
  NOR2_X1 U11938 ( .A1(n12040), .A2(n9932), .ZN(n9931) );
  NAND2_X1 U11939 ( .A1(n13053), .A2(n11992), .ZN(n12038) );
  INV_X1 U11940 ( .A(n9954), .ZN(n9570) );
  INV_X1 U11941 ( .A(n9576), .ZN(n9574) );
  INV_X1 U11942 ( .A(n11992), .ZN(n11969) );
  AND2_X1 U11943 ( .A1(n12023), .A2(n11969), .ZN(n12026) );
  NAND2_X1 U11944 ( .A1(n12031), .A2(n12026), .ZN(n10840) );
  AND2_X2 U11945 ( .A1(n9573), .A2(n11992), .ZN(n11779) );
  NAND2_X2 U11946 ( .A1(n9592), .A2(n14723), .ZN(n14716) );
  INV_X1 U11947 ( .A(n12038), .ZN(n9575) );
  INV_X1 U11948 ( .A(n12908), .ZN(n12942) );
  NAND2_X1 U11949 ( .A1(n9198), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9586) );
  INV_X1 U11950 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13081) );
  OR2_X1 U11951 ( .A1(n11730), .A2(n13081), .ZN(n9585) );
  INV_X1 U11952 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9577) );
  OAI21_X1 U11953 ( .B1(n9578), .B2(n9596), .A(n9577), .ZN(n9581) );
  INV_X1 U11954 ( .A(n9578), .ZN(n9580) );
  AND2_X1 U11955 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9579) );
  NAND2_X1 U11956 ( .A1(n9580), .A2(n9579), .ZN(n11764) );
  NAND2_X1 U11957 ( .A1(n9581), .A2(n11764), .ZN(n13080) );
  OR2_X1 U11958 ( .A1(n11731), .A2(n13080), .ZN(n9584) );
  INV_X1 U11959 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9582) );
  OR2_X1 U11960 ( .A1(n11966), .A2(n9582), .ZN(n9583) );
  NAND2_X1 U11961 ( .A1(n12950), .A2(n6433), .ZN(n9589) );
  INV_X1 U11962 ( .A(n9967), .ZN(n9587) );
  NAND2_X1 U11963 ( .A1(n9954), .A2(n9587), .ZN(n12919) );
  OR2_X1 U11964 ( .A1(n12919), .A2(n11929), .ZN(n9588) );
  NAND2_X1 U11965 ( .A1(n9589), .A2(n9588), .ZN(n13271) );
  INV_X1 U11966 ( .A(n9592), .ZN(n9591) );
  NAND2_X1 U11967 ( .A1(n9944), .A2(n9941), .ZN(n9590) );
  NAND2_X1 U11968 ( .A1(n9591), .A2(n9590), .ZN(n9595) );
  NAND2_X1 U11969 ( .A1(n11968), .A2(n12040), .ZN(n9940) );
  NAND4_X1 U11970 ( .A1(n9595), .A2(n9594), .A3(n9940), .A4(n9943), .ZN(n10273) );
  OAI22_X1 U11971 ( .A1(n12940), .A2(n13088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9596), .ZN(n9597) );
  AOI21_X1 U11972 ( .B1(n12942), .B2(n13271), .A(n9597), .ZN(n9598) );
  INV_X1 U11973 ( .A(n9599), .ZN(n9600) );
  XNOR2_X1 U11974 ( .A(n9602), .B(P3_B_REG_SCAN_IN), .ZN(n9603) );
  NAND2_X1 U11975 ( .A1(n9603), .A2(n11328), .ZN(n9604) );
  INV_X1 U11976 ( .A(n9605), .ZN(n11433) );
  NAND2_X1 U11977 ( .A1(n9602), .A2(n11433), .ZN(n9606) );
  INV_X1 U11978 ( .A(n9712), .ZN(n9607) );
  OAI21_X1 U11979 ( .B1(n10592), .B2(n10618), .A(n10620), .ZN(n9608) );
  INV_X1 U11980 ( .A(n9608), .ZN(n9609) );
  XNOR2_X1 U11981 ( .A(n9682), .B(n14864), .ZN(n9623) );
  INV_X1 U11982 ( .A(n9623), .ZN(n9624) );
  XNOR2_X1 U11983 ( .A(n9682), .B(n11302), .ZN(n9621) );
  INV_X1 U11984 ( .A(n9621), .ZN(n9622) );
  NAND2_X1 U11985 ( .A1(n11294), .A2(n12045), .ZN(n9615) );
  XNOR2_X1 U11986 ( .A(n10517), .B(n9619), .ZN(n9613) );
  NAND3_X1 U11987 ( .A1(n10517), .A2(n12257), .A3(n12045), .ZN(n9614) );
  INV_X1 U11988 ( .A(n9617), .ZN(n9618) );
  XNOR2_X1 U11989 ( .A(n9620), .B(n11299), .ZN(n10633) );
  XNOR2_X1 U11990 ( .A(n9621), .B(n14916), .ZN(n10893) );
  XNOR2_X1 U11991 ( .A(n9623), .B(n14890), .ZN(n12175) );
  XNOR2_X1 U11992 ( .A(n9682), .B(n14859), .ZN(n9625) );
  XNOR2_X1 U11993 ( .A(n9625), .B(n12255), .ZN(n12149) );
  XNOR2_X1 U11994 ( .A(n9682), .B(n9626), .ZN(n9627) );
  XNOR2_X1 U11995 ( .A(n9627), .B(n11315), .ZN(n12215) );
  NAND2_X1 U11996 ( .A1(n9627), .A2(n14855), .ZN(n9628) );
  XNOR2_X1 U11997 ( .A(n11644), .B(n12045), .ZN(n12064) );
  XNOR2_X1 U11998 ( .A(n9682), .B(n11646), .ZN(n9630) );
  XNOR2_X1 U11999 ( .A(n9630), .B(n11647), .ZN(n11341) );
  INV_X1 U12000 ( .A(n9630), .ZN(n9631) );
  XNOR2_X1 U12001 ( .A(n9682), .B(n14830), .ZN(n9632) );
  XNOR2_X1 U12002 ( .A(n9632), .B(n14839), .ZN(n11548) );
  NAND2_X1 U12003 ( .A1(n9632), .A2(n14839), .ZN(n9633) );
  XNOR2_X1 U12004 ( .A(n9682), .B(n11671), .ZN(n9634) );
  XNOR2_X1 U12005 ( .A(n9634), .B(n14290), .ZN(n12094) );
  XNOR2_X1 U12006 ( .A(n9682), .B(n12201), .ZN(n9638) );
  XNOR2_X1 U12007 ( .A(n9682), .B(n9636), .ZN(n9639) );
  NOR2_X1 U12008 ( .A1(n9639), .A2(n14272), .ZN(n9637) );
  AOI21_X1 U12009 ( .B1(n9638), .B2(n11672), .A(n9637), .ZN(n9642) );
  INV_X1 U12010 ( .A(n9637), .ZN(n12116) );
  INV_X1 U12011 ( .A(n9638), .ZN(n12118) );
  NAND3_X1 U12012 ( .A1(n12116), .A2(n12118), .A3(n12252), .ZN(n9640) );
  NAND2_X1 U12013 ( .A1(n9639), .A2(n14272), .ZN(n12115) );
  NAND2_X1 U12014 ( .A1(n9640), .A2(n12115), .ZN(n9641) );
  XNOR2_X1 U12015 ( .A(n12413), .B(n12045), .ZN(n11682) );
  NOR2_X1 U12016 ( .A1(n11682), .A2(n12668), .ZN(n9645) );
  INV_X1 U12017 ( .A(n11682), .ZN(n9643) );
  XNOR2_X1 U12018 ( .A(n12415), .B(n9682), .ZN(n9646) );
  XNOR2_X1 U12019 ( .A(n9646), .B(n12652), .ZN(n12075) );
  XNOR2_X1 U12020 ( .A(n12424), .B(n9682), .ZN(n9651) );
  XNOR2_X1 U12021 ( .A(n9651), .B(n12638), .ZN(n12238) );
  INV_X1 U12022 ( .A(n12238), .ZN(n9647) );
  NAND2_X1 U12023 ( .A1(n9646), .A2(n12652), .ZN(n12235) );
  AND2_X1 U12024 ( .A1(n9647), .A2(n12235), .ZN(n12140) );
  XNOR2_X1 U12025 ( .A(n12417), .B(n9682), .ZN(n9649) );
  XNOR2_X1 U12026 ( .A(n9649), .B(n12416), .ZN(n12142) );
  AND2_X1 U12027 ( .A1(n12140), .A2(n12142), .ZN(n9648) );
  INV_X1 U12028 ( .A(n9649), .ZN(n9650) );
  INV_X1 U12029 ( .A(n12142), .ZN(n9653) );
  INV_X1 U12030 ( .A(n9651), .ZN(n9652) );
  NAND2_X1 U12031 ( .A1(n9652), .A2(n12667), .ZN(n12141) );
  XNOR2_X1 U12032 ( .A(n12430), .B(n9682), .ZN(n9654) );
  XNOR2_X1 U12033 ( .A(n9654), .B(n12429), .ZN(n12158) );
  INV_X1 U12034 ( .A(n9654), .ZN(n9655) );
  XNOR2_X1 U12035 ( .A(n12609), .B(n9682), .ZN(n9656) );
  XNOR2_X1 U12036 ( .A(n9656), .B(n12589), .ZN(n12207) );
  INV_X1 U12037 ( .A(n9656), .ZN(n9657) );
  NAND2_X1 U12038 ( .A1(n9657), .A2(n12589), .ZN(n9658) );
  NAND2_X1 U12039 ( .A1(n9659), .A2(n9658), .ZN(n12099) );
  XNOR2_X1 U12040 ( .A(n12782), .B(n9682), .ZN(n9660) );
  INV_X1 U12041 ( .A(n12574), .ZN(n12604) );
  XNOR2_X1 U12042 ( .A(n9660), .B(n12604), .ZN(n12100) );
  NAND2_X1 U12043 ( .A1(n12099), .A2(n12100), .ZN(n9662) );
  NAND2_X1 U12044 ( .A1(n9660), .A2(n12574), .ZN(n9661) );
  NAND2_X1 U12045 ( .A1(n9662), .A2(n9661), .ZN(n12183) );
  XNOR2_X1 U12046 ( .A(n12721), .B(n9682), .ZN(n9663) );
  XNOR2_X1 U12047 ( .A(n9663), .B(n12588), .ZN(n12184) );
  NAND2_X1 U12048 ( .A1(n12183), .A2(n12184), .ZN(n9666) );
  INV_X1 U12049 ( .A(n9663), .ZN(n9664) );
  NAND2_X1 U12050 ( .A1(n9664), .A2(n12588), .ZN(n9665) );
  NAND2_X1 U12051 ( .A1(n9666), .A2(n9665), .ZN(n12106) );
  INV_X1 U12052 ( .A(n12106), .ZN(n9670) );
  XNOR2_X1 U12053 ( .A(n12562), .B(n9682), .ZN(n9668) );
  NAND2_X1 U12054 ( .A1(n9668), .A2(n9667), .ZN(n9671) );
  OAI21_X1 U12055 ( .B1(n9668), .B2(n9667), .A(n9671), .ZN(n12109) );
  INV_X1 U12056 ( .A(n12109), .ZN(n9669) );
  INV_X1 U12057 ( .A(n9675), .ZN(n9673) );
  XNOR2_X1 U12058 ( .A(n12714), .B(n9682), .ZN(n9674) );
  NAND2_X1 U12059 ( .A1(n9673), .A2(n9672), .ZN(n9676) );
  NAND2_X1 U12060 ( .A1(n9675), .A2(n9674), .ZN(n9677) );
  XNOR2_X1 U12061 ( .A(n12443), .B(n9682), .ZN(n9679) );
  NAND2_X1 U12062 ( .A1(n9679), .A2(n12136), .ZN(n12129) );
  INV_X1 U12063 ( .A(n9679), .ZN(n9680) );
  NAND2_X1 U12064 ( .A1(n9680), .A2(n12536), .ZN(n9681) );
  NAND2_X1 U12065 ( .A1(n12128), .A2(n12129), .ZN(n9686) );
  XNOR2_X1 U12066 ( .A(n12699), .B(n9682), .ZN(n9683) );
  NAND2_X1 U12067 ( .A1(n9683), .A2(n12526), .ZN(n9687) );
  INV_X1 U12068 ( .A(n9683), .ZN(n9684) );
  INV_X1 U12069 ( .A(n12526), .ZN(n12447) );
  NAND2_X1 U12070 ( .A1(n9684), .A2(n12447), .ZN(n9685) );
  NAND2_X1 U12071 ( .A1(n9686), .A2(n12130), .ZN(n12132) );
  XNOR2_X1 U12072 ( .A(n12507), .B(n12045), .ZN(n9688) );
  NOR2_X1 U12073 ( .A1(n9688), .A2(n12512), .ZN(n9689) );
  AOI21_X1 U12074 ( .B1(n9688), .B2(n12512), .A(n9689), .ZN(n12228) );
  INV_X1 U12075 ( .A(n9692), .ZN(n9690) );
  XNOR2_X1 U12076 ( .A(n12453), .B(n12045), .ZN(n12051) );
  NOR2_X1 U12077 ( .A1(n12051), .A2(n12452), .ZN(n12047) );
  AOI21_X1 U12078 ( .B1(n12051), .B2(n12452), .A(n12047), .ZN(n9691) );
  INV_X1 U12079 ( .A(n9693), .ZN(n12806) );
  NAND2_X1 U12080 ( .A1(n11328), .A2(n11433), .ZN(n9695) );
  NOR2_X1 U12081 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .ZN(
        n9700) );
  NOR4_X1 U12082 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_6__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9699) );
  NOR4_X1 U12083 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9698) );
  NOR4_X1 U12084 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n9697) );
  NAND4_X1 U12085 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n9706)
         );
  NOR4_X1 U12086 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9704) );
  NOR4_X1 U12087 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9703) );
  NOR4_X1 U12088 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9702) );
  NOR4_X1 U12089 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9701) );
  NAND4_X1 U12090 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n9705)
         );
  NOR2_X1 U12091 ( .A1(n9706), .A2(n9705), .ZN(n9707) );
  NAND3_X1 U12092 ( .A1(n12806), .A2(n12804), .A3(n10524), .ZN(n10664) );
  AND2_X1 U12093 ( .A1(n10592), .A2(n10345), .ZN(n9708) );
  XNOR2_X1 U12094 ( .A(n12685), .B(n9708), .ZN(n9710) );
  NAND2_X1 U12095 ( .A1(n10592), .A2(n12392), .ZN(n9709) );
  NAND2_X1 U12096 ( .A1(n9710), .A2(n9709), .ZN(n10656) );
  NAND2_X1 U12097 ( .A1(n12685), .A2(n10592), .ZN(n14954) );
  NAND2_X1 U12098 ( .A1(n10656), .A2(n14954), .ZN(n9714) );
  NAND2_X1 U12099 ( .A1(n9693), .A2(n10524), .ZN(n9711) );
  NAND2_X1 U12100 ( .A1(n10652), .A2(n10617), .ZN(n10519) );
  NOR2_X1 U12101 ( .A1(n10519), .A2(n9712), .ZN(n10659) );
  INV_X1 U12102 ( .A(n10659), .ZN(n9713) );
  OAI22_X1 U12103 ( .A1(n10664), .A2(n9714), .B1(n10655), .B2(n9713), .ZN(
        n9715) );
  INV_X1 U12104 ( .A(n12684), .ZN(n14908) );
  NAND2_X1 U12105 ( .A1(n10664), .A2(n14908), .ZN(n9717) );
  AND2_X1 U12106 ( .A1(n10660), .A2(n14907), .ZN(n9716) );
  NAND2_X1 U12107 ( .A1(n10664), .A2(n10656), .ZN(n9721) );
  OAI211_X1 U12108 ( .C1(n10536), .C2(n10529), .A(n9734), .B(n10422), .ZN(
        n9718) );
  INV_X1 U12109 ( .A(n9718), .ZN(n9720) );
  NAND2_X1 U12110 ( .A1(n10655), .A2(n10659), .ZN(n9719) );
  NAND3_X1 U12111 ( .A1(n9721), .A2(n9720), .A3(n9719), .ZN(n9722) );
  NAND2_X1 U12112 ( .A1(n9722), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9725) );
  INV_X1 U12113 ( .A(n10662), .ZN(n9723) );
  NAND2_X1 U12114 ( .A1(n10655), .A2(n9723), .ZN(n9724) );
  NAND2_X2 U12115 ( .A1(n9725), .A2(n9724), .ZN(n12248) );
  NOR2_X1 U12116 ( .A1(n10655), .A2(n10662), .ZN(n9727) );
  OR2_X1 U12117 ( .A1(n8119), .A2(n8117), .ZN(n10436) );
  NAND2_X1 U12118 ( .A1(n10436), .A2(n10424), .ZN(n10521) );
  NAND2_X1 U12119 ( .A1(n9727), .A2(n10521), .ZN(n12244) );
  INV_X1 U12120 ( .A(n10521), .ZN(n9726) );
  AOI22_X1 U12121 ( .A1(n12512), .A2(n12242), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9728) );
  OAI21_X1 U12122 ( .B1(n12485), .B2(n12244), .A(n9728), .ZN(n9729) );
  AOI21_X1 U12123 ( .B1(n12494), .B2(n12248), .A(n9729), .ZN(n9730) );
  INV_X1 U12124 ( .A(n11271), .ZN(n9732) );
  NOR2_X1 U12125 ( .A1(n9733), .A2(n9732), .ZN(n9956) );
  INV_X1 U12126 ( .A(n9797), .ZN(n9804) );
  NOR2_X4 U12127 ( .A1(n9734), .A2(n12803), .ZN(P3_U3897) );
  AND2_X1 U12128 ( .A1(n8178), .A2(P1_U3086), .ZN(n14184) );
  INV_X1 U12129 ( .A(n9735), .ZN(n9778) );
  AND2_X1 U12130 ( .A1(n9737), .A2(P1_U3086), .ZN(n9811) );
  OAI222_X1 U12131 ( .A1(n13650), .A2(P1_U3086), .B1(n14198), .B2(n9778), .C1(
        n9736), .C2(n14195), .ZN(P1_U3353) );
  AND2_X1 U12132 ( .A1(n8231), .A2(P3_U3151), .ZN(n14227) );
  NAND2_X1 U12133 ( .A1(n9737), .A2(P3_U3151), .ZN(n12817) );
  OAI222_X1 U12134 ( .A1(n12821), .A2(n9739), .B1(n12817), .B2(n9738), .C1(
        n11056), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12135 ( .A1(P3_U3151), .A2(n15037), .B1(n12817), .B2(n9741), .C1(
        n12821), .C2(n9740), .ZN(P3_U3295) );
  INV_X1 U12136 ( .A(n13663), .ZN(n9744) );
  INV_X1 U12137 ( .A(n9742), .ZN(n9772) );
  INV_X1 U12138 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9743) );
  OAI222_X1 U12139 ( .A1(n9744), .A2(P1_U3086), .B1(n14198), .B2(n9772), .C1(
        n9743), .C2(n14195), .ZN(P1_U3352) );
  OAI222_X1 U12140 ( .A1(n10502), .A2(P3_U3151), .B1(n12821), .B2(n9746), .C1(
        n9745), .C2(n12817), .ZN(P3_U3294) );
  INV_X1 U12141 ( .A(n14493), .ZN(n9749) );
  INV_X1 U12142 ( .A(n9747), .ZN(n9780) );
  INV_X1 U12143 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9748) );
  OAI222_X1 U12144 ( .A1(n9749), .A2(P1_U3086), .B1(n14198), .B2(n9780), .C1(
        n9748), .C2(n14195), .ZN(P1_U3351) );
  INV_X1 U12145 ( .A(n9750), .ZN(n9751) );
  INV_X1 U12146 ( .A(SI_10_), .ZN(n15116) );
  OAI222_X1 U12147 ( .A1(n12821), .A2(n9751), .B1(n12817), .B2(n15116), .C1(
        n11475), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X2 U12148 ( .A(n9811), .ZN(n14195) );
  OAI222_X1 U12149 ( .A1(n13631), .A2(P1_U3086), .B1(n14198), .B2(n9776), .C1(
        n9752), .C2(n14195), .ZN(P1_U3354) );
  OAI222_X1 U12150 ( .A1(n10451), .A2(P3_U3151), .B1(n12821), .B2(n9754), .C1(
        n9753), .C2(n12817), .ZN(P3_U3289) );
  INV_X1 U12151 ( .A(n9755), .ZN(n9774) );
  INV_X1 U12152 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9756) );
  OAI222_X1 U12153 ( .A1(n13679), .A2(P1_U3086), .B1(n14198), .B2(n9774), .C1(
        n9756), .C2(n14195), .ZN(P1_U3350) );
  INV_X1 U12154 ( .A(n12817), .ZN(n14226) );
  AOI222_X1 U12155 ( .A1(n9757), .A2(n14227), .B1(SI_9_), .B2(n14226), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11057), .ZN(n9758) );
  INV_X1 U12156 ( .A(n9758), .ZN(P3_U3286) );
  AOI222_X1 U12157 ( .A1(n9759), .A2(n14227), .B1(SI_7_), .B2(n14226), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10489), .ZN(n9760) );
  INV_X1 U12158 ( .A(n9760), .ZN(P3_U3288) );
  AOI222_X1 U12159 ( .A1(n9761), .A2(n14227), .B1(SI_11_), .B2(n14226), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11526), .ZN(n9762) );
  INV_X1 U12160 ( .A(n9762), .ZN(P3_U3284) );
  AOI222_X1 U12161 ( .A1(n9763), .A2(n14227), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10586), .C1(SI_3_), .C2(n14226), .ZN(n9764) );
  INV_X1 U12162 ( .A(n9764), .ZN(P3_U3292) );
  AOI222_X1 U12163 ( .A1(n9765), .A2(n14227), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10557), .C1(SI_2_), .C2(n14226), .ZN(n9766) );
  INV_X1 U12164 ( .A(n9766), .ZN(P3_U3293) );
  AOI222_X1 U12165 ( .A1(n9767), .A2(n14227), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10756), .C1(SI_5_), .C2(n14226), .ZN(n9768) );
  INV_X1 U12166 ( .A(n9768), .ZN(P3_U3290) );
  AOI222_X1 U12167 ( .A1(n9769), .A2(n14227), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10573), .C1(SI_4_), .C2(n14226), .ZN(n9770) );
  INV_X1 U12168 ( .A(n9770), .ZN(P3_U3291) );
  NOR2_X1 U12169 ( .A1(n9771), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13366) );
  INV_X1 U12170 ( .A(n13010), .ZN(n9961) );
  OAI222_X1 U12171 ( .A1(n13377), .A2(n9773), .B1(n13373), .B2(n9772), .C1(
        P2_U3088), .C2(n9961), .ZN(P2_U3324) );
  INV_X1 U12172 ( .A(n9979), .ZN(n10090) );
  OAI222_X1 U12173 ( .A1(n13377), .A2(n9775), .B1(n13373), .B2(n9774), .C1(
        P2_U3088), .C2(n10090), .ZN(P2_U3322) );
  OAI222_X1 U12174 ( .A1(n13377), .A2(n9777), .B1(n13373), .B2(n9776), .C1(
        P2_U3088), .C2(n12985), .ZN(P2_U3326) );
  OAI222_X1 U12175 ( .A1(n13377), .A2(n9779), .B1(n13373), .B2(n9778), .C1(
        P2_U3088), .C2(n9977), .ZN(P2_U3325) );
  OAI222_X1 U12176 ( .A1(n13377), .A2(n9781), .B1(n13373), .B2(n9780), .C1(
        P2_U3088), .C2(n14617), .ZN(P2_U3323) );
  OAI222_X1 U12177 ( .A1(n12821), .A2(n9782), .B1(n12817), .B2(n15112), .C1(
        n12263), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12178 ( .A(n9888), .ZN(n9895) );
  INV_X1 U12179 ( .A(n9783), .ZN(n9785) );
  OAI222_X1 U12180 ( .A1(n9895), .A2(P1_U3086), .B1(n14198), .B2(n9785), .C1(
        n9784), .C2(n14195), .ZN(P1_U3349) );
  INV_X1 U12181 ( .A(n9991), .ZN(n10003) );
  OAI222_X1 U12182 ( .A1(n13377), .A2(n9786), .B1(n13373), .B2(n9785), .C1(
        P2_U3088), .C2(n10003), .ZN(P2_U3321) );
  INV_X1 U12183 ( .A(n13696), .ZN(n9840) );
  INV_X1 U12184 ( .A(n9787), .ZN(n9790) );
  OAI222_X1 U12185 ( .A1(n9840), .A2(P1_U3086), .B1(n14198), .B2(n9790), .C1(
        n9788), .C2(n14195), .ZN(P1_U3348) );
  INV_X1 U12186 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9791) );
  INV_X1 U12187 ( .A(n14633), .ZN(n9789) );
  OAI222_X1 U12188 ( .A1(n13377), .A2(n9791), .B1(n13373), .B2(n9790), .C1(
        P2_U3088), .C2(n9789), .ZN(P2_U3320) );
  INV_X1 U12189 ( .A(n9792), .ZN(n11556) );
  NAND3_X1 U12190 ( .A1(n11556), .A2(n9793), .A3(P1_B_REG_SCAN_IN), .ZN(n9796)
         );
  INV_X1 U12191 ( .A(P1_B_REG_SCAN_IN), .ZN(n9794) );
  INV_X1 U12192 ( .A(n9803), .ZN(n14194) );
  AOI21_X1 U12193 ( .B1(n9792), .B2(n9794), .A(n14194), .ZN(n9795) );
  NAND2_X1 U12194 ( .A1(n9912), .A2(n10306), .ZN(n14531) );
  INV_X1 U12195 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9798) );
  AOI22_X1 U12196 ( .A1(n14531), .A2(n9798), .B1(n9797), .B2(n10025), .ZN(
        P1_U3446) );
  INV_X1 U12197 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9800) );
  INV_X1 U12198 ( .A(n9799), .ZN(n9802) );
  INV_X1 U12199 ( .A(n10166), .ZN(n9989) );
  OAI222_X1 U12200 ( .A1(n13377), .A2(n9800), .B1(n13373), .B2(n9802), .C1(
        P2_U3088), .C2(n9989), .ZN(P2_U3319) );
  OAI222_X1 U12201 ( .A1(n9869), .A2(P1_U3086), .B1(n14198), .B2(n9802), .C1(
        n9801), .C2(n14195), .ZN(P1_U3347) );
  INV_X1 U12202 ( .A(n14531), .ZN(n14530) );
  OR2_X1 U12203 ( .A1(n9792), .A2(n9803), .ZN(n9913) );
  OAI22_X1 U12204 ( .A1(n14530), .A2(P1_D_REG_0__SCAN_IN), .B1(n9804), .B2(
        n9913), .ZN(n9805) );
  INV_X1 U12205 ( .A(n9805), .ZN(P1_U3445) );
  INV_X1 U12206 ( .A(n9806), .ZN(n9808) );
  OAI222_X1 U12207 ( .A1(n13715), .A2(P1_U3086), .B1(n14198), .B2(n9808), .C1(
        n9807), .C2(n14195), .ZN(P1_U3346) );
  INV_X1 U12208 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9809) );
  OAI222_X1 U12209 ( .A1(n13377), .A2(n9809), .B1(n13373), .B2(n9808), .C1(
        P2_U3088), .C2(n10167), .ZN(P2_U3318) );
  INV_X1 U12210 ( .A(n9810), .ZN(n9813) );
  AOI22_X1 U12211 ( .A1(n10011), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9811), .ZN(n9812) );
  OAI21_X1 U12212 ( .B1(n9813), .B2(n14198), .A(n9812), .ZN(P1_U3345) );
  INV_X1 U12213 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9814) );
  INV_X1 U12214 ( .A(n10210), .ZN(n10172) );
  OAI222_X1 U12215 ( .A1(n13377), .A2(n9814), .B1(n13373), .B2(n9813), .C1(
        P2_U3088), .C2(n10172), .ZN(P2_U3317) );
  INV_X1 U12216 ( .A(n10306), .ZN(n10045) );
  NAND2_X1 U12217 ( .A1(n10045), .A2(n11275), .ZN(n9844) );
  AOI21_X1 U12218 ( .B1(n9916), .B2(n10706), .A(n9815), .ZN(n9843) );
  INV_X1 U12219 ( .A(n9843), .ZN(n9816) );
  AND2_X1 U12220 ( .A1(n9844), .A2(n9816), .ZN(n14497) );
  CLKBUF_X2 U12221 ( .A(P1_U4016), .Z(n13644) );
  NOR2_X1 U12222 ( .A1(n14497), .A2(n13644), .ZN(P1_U3085) );
  OAI222_X1 U12223 ( .A1(n12821), .A2(n9818), .B1(n12817), .B2(n9817), .C1(
        n12309), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12224 ( .A(n13731), .ZN(n9821) );
  INV_X1 U12225 ( .A(n9819), .ZN(n9823) );
  OAI222_X1 U12226 ( .A1(n9821), .A2(P1_U3086), .B1(n14198), .B2(n9823), .C1(
        n9820), .C2(n14195), .ZN(P1_U3344) );
  INV_X1 U12227 ( .A(n11446), .ZN(n9822) );
  OAI222_X1 U12228 ( .A1(n13377), .A2(n9824), .B1(n13373), .B2(n9823), .C1(
        P2_U3088), .C2(n9822), .ZN(P2_U3316) );
  MUX2_X1 U12229 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9825), .S(n9869), .Z(n9842)
         );
  INV_X1 U12230 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14609) );
  MUX2_X1 U12231 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9826), .S(n14493), .Z(n9837) );
  INV_X1 U12232 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9827) );
  MUX2_X1 U12233 ( .A(n9827), .B(P1_REG1_REG_1__SCAN_IN), .S(n13631), .Z(n9829) );
  AND2_X1 U12234 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9828) );
  NAND2_X1 U12235 ( .A1(n9829), .A2(n9828), .ZN(n13653) );
  INV_X1 U12236 ( .A(n13631), .ZN(n13634) );
  NAND2_X1 U12237 ( .A1(n13634), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U12238 ( .A1(n13653), .A2(n13652), .ZN(n9832) );
  MUX2_X1 U12239 ( .A(n9830), .B(P1_REG1_REG_2__SCAN_IN), .S(n13650), .Z(n9831) );
  NAND2_X1 U12240 ( .A1(n9832), .A2(n9831), .ZN(n13666) );
  INV_X1 U12241 ( .A(n13650), .ZN(n9848) );
  NAND2_X1 U12242 ( .A1(n9848), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13665) );
  NAND2_X1 U12243 ( .A1(n13666), .A2(n13665), .ZN(n9835) );
  MUX2_X1 U12244 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9833), .S(n13663), .Z(n9834) );
  NAND2_X1 U12245 ( .A1(n9835), .A2(n9834), .ZN(n14482) );
  NAND2_X1 U12246 ( .A1(n13663), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U12247 ( .A1(n14482), .A2(n14481), .ZN(n9836) );
  NAND2_X1 U12248 ( .A1(n9837), .A2(n9836), .ZN(n14485) );
  INV_X1 U12249 ( .A(n14485), .ZN(n9838) );
  AOI21_X1 U12250 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n14493), .A(n9838), .ZN(
        n13676) );
  MUX2_X1 U12251 ( .A(n8575), .B(P1_REG1_REG_5__SCAN_IN), .S(n13679), .Z(
        n13677) );
  NAND2_X1 U12252 ( .A1(n13676), .A2(n13677), .ZN(n13675) );
  OAI21_X1 U12253 ( .B1(n13674), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13675), .ZN(
        n9893) );
  INV_X1 U12254 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14607) );
  MUX2_X1 U12255 ( .A(n14607), .B(P1_REG1_REG_6__SCAN_IN), .S(n9888), .Z(n9892) );
  NOR2_X1 U12256 ( .A1(n9893), .A2(n9892), .ZN(n13701) );
  NOR2_X1 U12257 ( .A1(n9895), .A2(n14607), .ZN(n13695) );
  MUX2_X1 U12258 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14609), .S(n13696), .Z(
        n9839) );
  OAI21_X1 U12259 ( .B1(n13701), .B2(n13695), .A(n9839), .ZN(n13699) );
  OAI21_X1 U12260 ( .B1(n14609), .B2(n9840), .A(n13699), .ZN(n9841) );
  NOR2_X1 U12261 ( .A1(n9841), .A2(n9842), .ZN(n13708) );
  AOI21_X1 U12262 ( .B1(n9842), .B2(n9841), .A(n13708), .ZN(n9868) );
  NAND2_X1 U12263 ( .A1(n9844), .A2(n9843), .ZN(n14479) );
  INV_X1 U12264 ( .A(n14191), .ZN(n14475) );
  OR2_X1 U12265 ( .A1(n14479), .A2(n14475), .ZN(n14522) );
  AND2_X1 U12266 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11194) );
  NOR2_X1 U12267 ( .A1(n14524), .A2(n9869), .ZN(n9845) );
  AOI211_X1 U12268 ( .C1(n14497), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11194), .B(
        n9845), .ZN(n9867) );
  OR2_X1 U12269 ( .A1(n8937), .A2(n14191), .ZN(n9846) );
  INV_X1 U12270 ( .A(n14520), .ZN(n14492) );
  MUX2_X1 U12271 ( .A(n9847), .B(P1_REG2_REG_1__SCAN_IN), .S(n13631), .Z(
        n13630) );
  AND2_X1 U12272 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13641) );
  NAND2_X1 U12273 ( .A1(n13630), .A2(n13641), .ZN(n13629) );
  OAI21_X1 U12274 ( .B1(n9847), .B2(n13631), .A(n13629), .ZN(n13647) );
  XNOR2_X1 U12275 ( .A(n13650), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n13646) );
  NAND2_X1 U12276 ( .A1(n13647), .A2(n13646), .ZN(n9850) );
  NAND2_X1 U12277 ( .A1(n9848), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12278 ( .A1(n9850), .A2(n9849), .ZN(n13661) );
  MUX2_X1 U12279 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10363), .S(n13663), .Z(
        n13662) );
  NAND2_X1 U12280 ( .A1(n13661), .A2(n13662), .ZN(n14488) );
  NAND2_X1 U12281 ( .A1(n13663), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U12282 ( .A1(n14488), .A2(n14487), .ZN(n9852) );
  MUX2_X1 U12283 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10612), .S(n14493), .Z(
        n9851) );
  NAND2_X1 U12284 ( .A1(n9852), .A2(n9851), .ZN(n14491) );
  NAND2_X1 U12285 ( .A1(n14493), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U12286 ( .A1(n14491), .A2(n13680), .ZN(n9855) );
  MUX2_X1 U12287 ( .A(n9853), .B(P1_REG2_REG_5__SCAN_IN), .S(n13679), .Z(n9854) );
  NAND2_X1 U12288 ( .A1(n9855), .A2(n9854), .ZN(n13683) );
  NAND2_X1 U12289 ( .A1(n13674), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12290 ( .A1(n13683), .A2(n9890), .ZN(n9857) );
  MUX2_X1 U12291 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10397), .S(n9888), .Z(n9856) );
  NAND2_X1 U12292 ( .A1(n9857), .A2(n9856), .ZN(n13692) );
  NAND2_X1 U12293 ( .A1(n9888), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13691) );
  NAND2_X1 U12294 ( .A1(n13692), .A2(n13691), .ZN(n9860) );
  MUX2_X1 U12295 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9858), .S(n13696), .Z(n9859) );
  NAND2_X1 U12296 ( .A1(n9860), .A2(n9859), .ZN(n13694) );
  NAND2_X1 U12297 ( .A1(n13696), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12298 ( .A1(n13694), .A2(n9864), .ZN(n9862) );
  MUX2_X1 U12299 ( .A(n10732), .B(P1_REG2_REG_8__SCAN_IN), .S(n9869), .Z(n9861) );
  NAND2_X1 U12300 ( .A1(n9862), .A2(n9861), .ZN(n13718) );
  MUX2_X1 U12301 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10732), .S(n9869), .Z(n9863) );
  NAND3_X1 U12302 ( .A1(n13694), .A2(n9864), .A3(n9863), .ZN(n9865) );
  NAND3_X1 U12303 ( .A1(n14492), .A2(n13718), .A3(n9865), .ZN(n9866) );
  OAI211_X1 U12304 ( .C1(n9868), .C2(n14522), .A(n9867), .B(n9866), .ZN(
        P1_U3251) );
  INV_X1 U12305 ( .A(n13715), .ZN(n13714) );
  INV_X1 U12306 ( .A(n9869), .ZN(n9872) );
  NOR2_X1 U12307 ( .A1(n9872), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13706) );
  MUX2_X1 U12308 ( .A(n8457), .B(P1_REG1_REG_9__SCAN_IN), .S(n13715), .Z(
        n13707) );
  OAI21_X1 U12309 ( .B1(n13708), .B2(n13706), .A(n13707), .ZN(n13705) );
  OAI21_X1 U12310 ( .B1(n13714), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13705), .ZN(
        n9871) );
  MUX2_X1 U12311 ( .A(n8606), .B(P1_REG1_REG_10__SCAN_IN), .S(n10011), .Z(
        n9870) );
  NOR2_X1 U12312 ( .A1(n9871), .A2(n9870), .ZN(n10010) );
  AOI211_X1 U12313 ( .C1(n9871), .C2(n9870), .A(n14522), .B(n10010), .ZN(n9887) );
  INV_X1 U12314 ( .A(n10011), .ZN(n9885) );
  NAND2_X1 U12315 ( .A1(n9872), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U12316 ( .A1(n13718), .A2(n13717), .ZN(n9875) );
  MUX2_X1 U12317 ( .A(n9873), .B(P1_REG2_REG_9__SCAN_IN), .S(n13715), .Z(n9874) );
  NAND2_X1 U12318 ( .A1(n9875), .A2(n9874), .ZN(n13720) );
  NAND2_X1 U12319 ( .A1(n13714), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U12320 ( .A1(n13720), .A2(n9880), .ZN(n9878) );
  MUX2_X1 U12321 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9876), .S(n10011), .Z(
        n9877) );
  NAND2_X1 U12322 ( .A1(n9878), .A2(n9877), .ZN(n13734) );
  MUX2_X1 U12323 ( .A(n9876), .B(P1_REG2_REG_10__SCAN_IN), .S(n10011), .Z(
        n9879) );
  NAND3_X1 U12324 ( .A1(n13720), .A2(n9880), .A3(n9879), .ZN(n9881) );
  NAND3_X1 U12325 ( .A1(n14492), .A2(n13734), .A3(n9881), .ZN(n9884) );
  NOR2_X1 U12326 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9882), .ZN(n11364) );
  AOI21_X1 U12327 ( .B1(n14497), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11364), 
        .ZN(n9883) );
  OAI211_X1 U12328 ( .C1(n14524), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9886)
         );
  OR2_X1 U12329 ( .A1(n9887), .A2(n9886), .ZN(P1_U3253) );
  MUX2_X1 U12330 ( .A(n10397), .B(P1_REG2_REG_6__SCAN_IN), .S(n9888), .Z(n9889) );
  NAND3_X1 U12331 ( .A1(n13683), .A2(n9890), .A3(n9889), .ZN(n9891) );
  AND3_X1 U12332 ( .A1(n14492), .A2(n13692), .A3(n9891), .ZN(n9898) );
  AOI211_X1 U12333 ( .C1(n9893), .C2(n9892), .A(n13701), .B(n14522), .ZN(n9897) );
  NAND2_X1 U12334 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U12335 ( .A1(n14497), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9894) );
  OAI211_X1 U12336 ( .C1(n14524), .C2(n9895), .A(n10781), .B(n9894), .ZN(n9896) );
  OR3_X1 U12337 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(P1_U3249) );
  NOR2_X1 U12338 ( .A1(n9912), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9911) );
  INV_X1 U12339 ( .A(n10301), .ZN(n10049) );
  NOR4_X1 U12340 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9907) );
  NOR4_X1 U12341 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9906) );
  INV_X1 U12342 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15085) );
  INV_X1 U12343 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15123) );
  INV_X1 U12344 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15131) );
  INV_X1 U12345 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15108) );
  NAND4_X1 U12346 ( .A1(n15085), .A2(n15123), .A3(n15131), .A4(n15108), .ZN(
        n9904) );
  NOR4_X1 U12347 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9902) );
  NOR4_X1 U12348 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9901) );
  NOR4_X1 U12349 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9900) );
  NOR4_X1 U12350 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9899) );
  NAND4_X1 U12351 ( .A1(n9902), .A2(n9901), .A3(n9900), .A4(n9899), .ZN(n9903)
         );
  NOR4_X1 U12352 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n9904), .A4(n9903), .ZN(n9905) );
  AND3_X1 U12353 ( .A1(n9907), .A2(n9906), .A3(n9905), .ZN(n10022) );
  INV_X1 U12354 ( .A(n10022), .ZN(n9909) );
  AOI21_X1 U12355 ( .B1(n10024), .B2(n9909), .A(n10305), .ZN(n9910) );
  OAI211_X1 U12356 ( .C1(n9911), .C2(n10025), .A(n10049), .B(n9910), .ZN(n9924) );
  OR2_X1 U12357 ( .A1(n9912), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9914) );
  INV_X1 U12358 ( .A(n10303), .ZN(n9915) );
  INV_X1 U12359 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12360 ( .A1(n9916), .A2(n8937), .ZN(n13951) );
  NOR2_X1 U12361 ( .A1(n10125), .A2(n13951), .ZN(n10404) );
  INV_X1 U12362 ( .A(n10404), .ZN(n9921) );
  OAI21_X1 U12363 ( .B1(n9919), .B2(n11138), .A(n10033), .ZN(n10774) );
  INV_X1 U12364 ( .A(n10774), .ZN(n10689) );
  NAND2_X1 U12365 ( .A1(n10031), .A2(n14200), .ZN(n9917) );
  OAI21_X2 U12366 ( .B1(n9919), .B2(n13782), .A(n9918), .ZN(n14554) );
  OAI21_X1 U12367 ( .B1(n14597), .B2(n14554), .A(n10405), .ZN(n9920) );
  OAI211_X1 U12368 ( .C1(n10323), .C2(n10669), .A(n9921), .B(n9920), .ZN(n9925) );
  NAND2_X1 U12369 ( .A1(n14601), .A2(n9925), .ZN(n9922) );
  OAI21_X1 U12370 ( .B1(n14601), .B2(n9923), .A(n9922), .ZN(P1_U3459) );
  NAND2_X1 U12371 ( .A1(n14615), .A2(n9925), .ZN(n9926) );
  OAI21_X1 U12372 ( .B1(n14615), .B2(n8543), .A(n9926), .ZN(P1_U3528) );
  INV_X1 U12373 ( .A(n9927), .ZN(n9929) );
  OAI222_X1 U12374 ( .A1(n12332), .A2(P3_U3151), .B1(n12821), .B2(n9929), .C1(
        n9928), .C2(n12817), .ZN(P3_U3280) );
  INV_X1 U12375 ( .A(n14761), .ZN(n14736) );
  OR2_X1 U12376 ( .A1(n11780), .A2(n12979), .ZN(n10296) );
  AND2_X1 U12377 ( .A1(n11780), .A2(n12979), .ZN(n11783) );
  INV_X1 U12378 ( .A(n11783), .ZN(n9930) );
  NAND2_X1 U12379 ( .A1(n10296), .A2(n9930), .ZN(n14708) );
  AND2_X1 U12380 ( .A1(n10297), .A2(n9931), .ZN(n14710) );
  INV_X1 U12381 ( .A(n10917), .ZN(n13144) );
  NAND2_X1 U12382 ( .A1(n12027), .A2(n12040), .ZN(n9933) );
  NAND2_X1 U12383 ( .A1(n9932), .A2(n11969), .ZN(n12030) );
  OAI21_X1 U12384 ( .B1(n13144), .B2(n14753), .A(n14708), .ZN(n9934) );
  NAND2_X1 U12385 ( .A1(n6433), .A2(n12978), .ZN(n10294) );
  AND2_X1 U12386 ( .A1(n9934), .A2(n10294), .ZN(n14712) );
  INV_X1 U12387 ( .A(n14712), .ZN(n9935) );
  AOI211_X1 U12388 ( .C1(n14736), .C2(n14708), .A(n14710), .B(n9935), .ZN(
        n9948) );
  NAND2_X1 U12389 ( .A1(n14723), .A2(n9941), .ZN(n9936) );
  NOR2_X1 U12390 ( .A1(n9943), .A2(n9936), .ZN(n9938) );
  INV_X1 U12391 ( .A(n9940), .ZN(n9937) );
  NAND2_X1 U12392 ( .A1(n14769), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9939) );
  OAI21_X1 U12393 ( .B1(n9948), .B2(n14769), .A(n9939), .ZN(P2_U3430) );
  NAND2_X1 U12394 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NOR2_X1 U12395 ( .A1(n9943), .A2(n9942), .ZN(n9946) );
  NAND2_X1 U12396 ( .A1(n9944), .A2(n14723), .ZN(n14721) );
  NAND2_X1 U12397 ( .A1(n14776), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9947) );
  OAI21_X1 U12398 ( .B1(n9948), .B2(n14776), .A(n9947), .ZN(P2_U3499) );
  INV_X1 U12399 ( .A(n9949), .ZN(n9952) );
  OAI222_X1 U12400 ( .A1(n13373), .A2(n9952), .B1(n11447), .B2(P2_U3088), .C1(
        n9950), .C2(n13377), .ZN(P2_U3315) );
  INV_X1 U12401 ( .A(n10228), .ZN(n10220) );
  OAI222_X1 U12402 ( .A1(P1_U3086), .A2(n10220), .B1(n14198), .B2(n9952), .C1(
        n9951), .C2(n14195), .ZN(P1_U3343) );
  AOI21_X1 U12403 ( .B1(n9954), .B2(n11271), .A(n6435), .ZN(n9955) );
  OR2_X1 U12404 ( .A1(n9956), .A2(n9955), .ZN(n9974) );
  AND2_X1 U12405 ( .A1(n9974), .A2(n9967), .ZN(n14616) );
  INV_X1 U12406 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12407 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9957) );
  NOR2_X1 U12408 ( .A1(n12985), .A2(n12986), .ZN(n9958) );
  AOI211_X1 U12409 ( .C1(n12986), .C2(n12985), .A(n9957), .B(n9958), .ZN(
        n12987) );
  NOR2_X1 U12410 ( .A1(n12987), .A2(n9958), .ZN(n12994) );
  XOR2_X1 U12411 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9977), .Z(n12995) );
  OAI22_X1 U12412 ( .A1(n12994), .A2(n12995), .B1(n9977), .B2(n9959), .ZN(
        n13013) );
  MUX2_X1 U12413 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9960), .S(n13010), .Z(
        n13014) );
  NAND2_X1 U12414 ( .A1(n13013), .A2(n13014), .ZN(n13012) );
  OAI21_X1 U12415 ( .B1(n9960), .B2(n9961), .A(n13012), .ZN(n14626) );
  MUX2_X1 U12416 ( .A(n9962), .B(P2_REG1_REG_4__SCAN_IN), .S(n14617), .Z(
        n14625) );
  NAND2_X1 U12417 ( .A1(n14626), .A2(n14625), .ZN(n14624) );
  NAND2_X1 U12418 ( .A1(n9963), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U12419 ( .A(n9964), .B(P2_REG1_REG_5__SCAN_IN), .S(n9979), .Z(n10079) );
  AOI21_X1 U12420 ( .B1(n14624), .B2(n10080), .A(n10079), .ZN(n10082) );
  NOR2_X1 U12421 ( .A1(n10090), .A2(n9964), .ZN(n9990) );
  MUX2_X1 U12422 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10265), .S(n9991), .Z(n9965) );
  OAI21_X1 U12423 ( .B1(n10082), .B2(n9990), .A(n9965), .ZN(n9996) );
  OAI21_X1 U12424 ( .B1(n10265), .B2(n10003), .A(n9996), .ZN(n14639) );
  MUX2_X1 U12425 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9966), .S(n14633), .Z(
        n14638) );
  NAND2_X1 U12426 ( .A1(n14639), .A2(n14638), .ZN(n14637) );
  NAND2_X1 U12427 ( .A1(n14633), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9971) );
  INV_X1 U12428 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14774) );
  MUX2_X1 U12429 ( .A(n14774), .B(P2_REG1_REG_8__SCAN_IN), .S(n10166), .Z(
        n9970) );
  AOI21_X1 U12430 ( .B1(n14637), .B2(n9971), .A(n9970), .ZN(n10165) );
  INV_X1 U12431 ( .A(n10165), .ZN(n9973) );
  OR2_X1 U12432 ( .A1(n9967), .A2(P2_U3088), .ZN(n13368) );
  INV_X1 U12433 ( .A(n13368), .ZN(n9968) );
  AND2_X1 U12434 ( .A1(n9974), .A2(n9968), .ZN(n9981) );
  NAND3_X1 U12435 ( .A1(n14637), .A2(n9971), .A3(n9970), .ZN(n9972) );
  NAND3_X1 U12436 ( .A1(n9973), .A2(n14696), .A3(n9972), .ZN(n9988) );
  NOR2_X2 U12437 ( .A1(n9974), .A2(P2_U3088), .ZN(n14680) );
  NAND2_X1 U12438 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11114) );
  INV_X1 U12439 ( .A(n12985), .ZN(n12984) );
  NOR3_X1 U12440 ( .A1(n12982), .A2(n9976), .A3(n9975), .ZN(n12980) );
  AOI21_X1 U12441 ( .B1(n12984), .B2(P2_REG2_REG_1__SCAN_IN), .A(n12980), .ZN(
        n12999) );
  INV_X1 U12442 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10875) );
  MUX2_X1 U12443 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10875), .S(n9977), .Z(
        n12998) );
  OR2_X1 U12444 ( .A1(n12999), .A2(n12998), .ZN(n13006) );
  INV_X1 U12445 ( .A(n9977), .ZN(n12997) );
  NAND2_X1 U12446 ( .A1(n12997), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13005) );
  MUX2_X1 U12447 ( .A(n9152), .B(P2_REG2_REG_3__SCAN_IN), .S(n13010), .Z(
        n13004) );
  AOI21_X1 U12448 ( .B1(n13006), .B2(n13005), .A(n13004), .ZN(n13008) );
  AOI21_X1 U12449 ( .B1(n13010), .B2(P2_REG2_REG_3__SCAN_IN), .A(n13008), .ZN(
        n14622) );
  MUX2_X1 U12450 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9978), .S(n14617), .Z(
        n14621) );
  NOR2_X1 U12451 ( .A1(n14622), .A2(n14621), .ZN(n14620) );
  NOR2_X1 U12452 ( .A1(n14617), .A2(n9978), .ZN(n10085) );
  MUX2_X1 U12453 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10947), .S(n9979), .Z(
        n10084) );
  NAND2_X1 U12454 ( .A1(n9979), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9999) );
  MUX2_X1 U12455 ( .A(n10940), .B(P2_REG2_REG_6__SCAN_IN), .S(n9991), .Z(n9998) );
  INV_X1 U12456 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9980) );
  MUX2_X1 U12457 ( .A(n9980), .B(P2_REG2_REG_7__SCAN_IN), .S(n14633), .Z(
        n14635) );
  AOI21_X1 U12458 ( .B1(n14633), .B2(P2_REG2_REG_7__SCAN_IN), .A(n14634), .ZN(
        n9983) );
  MUX2_X1 U12459 ( .A(n10842), .B(P2_REG2_REG_8__SCAN_IN), .S(n10166), .Z(
        n9982) );
  NOR2_X1 U12460 ( .A1(n9983), .A2(n9982), .ZN(n10162) );
  INV_X1 U12461 ( .A(n12039), .ZN(n11737) );
  NAND2_X1 U12462 ( .A1(n9981), .A2(n11737), .ZN(n14700) );
  AOI211_X1 U12463 ( .C1(n9983), .C2(n9982), .A(n10162), .B(n14700), .ZN(n9984) );
  INV_X1 U12464 ( .A(n9984), .ZN(n9985) );
  NAND2_X1 U12465 ( .A1(n11114), .A2(n9985), .ZN(n9986) );
  AOI21_X1 U12466 ( .B1(n14680), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9986), .ZN(
        n9987) );
  OAI211_X1 U12467 ( .C1(n14658), .C2(n9989), .A(n9988), .B(n9987), .ZN(
        P2_U3222) );
  AND2_X1 U12468 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10980) );
  INV_X1 U12469 ( .A(n10082), .ZN(n9994) );
  INV_X1 U12470 ( .A(n9990), .ZN(n9993) );
  MUX2_X1 U12471 ( .A(n10265), .B(P2_REG1_REG_6__SCAN_IN), .S(n9991), .Z(n9992) );
  NAND3_X1 U12472 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(n9995) );
  AND3_X1 U12473 ( .A1(n14696), .A2(n9996), .A3(n9995), .ZN(n9997) );
  AOI211_X1 U12474 ( .C1(n14680), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10980), .B(
        n9997), .ZN(n10002) );
  NAND3_X1 U12475 ( .A1(n10087), .A2(n9999), .A3(n9998), .ZN(n10000) );
  NAND3_X1 U12476 ( .A1(n6585), .A2(n14683), .A3(n10000), .ZN(n10001) );
  OAI211_X1 U12477 ( .C1(n14658), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        P2_U3220) );
  MUX2_X1 U12478 ( .A(n11223), .B(P1_REG2_REG_12__SCAN_IN), .S(n10228), .Z(
        n10009) );
  NAND2_X1 U12479 ( .A1(n10011), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U12480 ( .A1(n13734), .A2(n13733), .ZN(n10006) );
  MUX2_X1 U12481 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10004), .S(n13731), .Z(
        n10005) );
  NAND2_X1 U12482 ( .A1(n10006), .A2(n10005), .ZN(n13736) );
  NAND2_X1 U12483 ( .A1(n13731), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12484 ( .A1(n13736), .A2(n10007), .ZN(n10008) );
  NOR2_X1 U12485 ( .A1(n10008), .A2(n10009), .ZN(n10230) );
  AOI21_X1 U12486 ( .B1(n10009), .B2(n10008), .A(n10230), .ZN(n10021) );
  AOI21_X1 U12487 ( .B1(n10011), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10010), 
        .ZN(n13725) );
  MUX2_X1 U12488 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n8443), .S(n13731), .Z(
        n13726) );
  NAND2_X1 U12489 ( .A1(n13725), .A2(n13726), .ZN(n13724) );
  OR2_X1 U12490 ( .A1(n13731), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10013) );
  MUX2_X1 U12491 ( .A(n10012), .B(P1_REG1_REG_12__SCAN_IN), .S(n10228), .Z(
        n10014) );
  AOI21_X1 U12492 ( .B1(n13724), .B2(n10013), .A(n10014), .ZN(n10219) );
  AND3_X1 U12493 ( .A1(n13724), .A2(n10014), .A3(n10013), .ZN(n10015) );
  OAI21_X1 U12494 ( .B1(n10219), .B2(n10015), .A(n14486), .ZN(n10020) );
  NOR2_X1 U12495 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10016), .ZN(n10018) );
  NOR2_X1 U12496 ( .A1(n14524), .A2(n10220), .ZN(n10017) );
  AOI211_X1 U12497 ( .C1(n14497), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10018), 
        .B(n10017), .ZN(n10019) );
  OAI211_X1 U12498 ( .C1(n10021), .C2(n14520), .A(n10020), .B(n10019), .ZN(
        P1_U3255) );
  NAND2_X1 U12499 ( .A1(n10022), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12500 ( .A1(n10024), .A2(n10023), .ZN(n10027) );
  INV_X1 U12501 ( .A(n10025), .ZN(n10026) );
  NAND2_X1 U12502 ( .A1(n10027), .A2(n10026), .ZN(n10302) );
  INV_X1 U12503 ( .A(n10305), .ZN(n10028) );
  NAND2_X1 U12504 ( .A1(n10048), .A2(n10028), .ZN(n10709) );
  AND2_X1 U12505 ( .A1(n10709), .A2(n10306), .ZN(n14369) );
  INV_X1 U12506 ( .A(n10029), .ZN(n10030) );
  AND2_X2 U12507 ( .A1(n10034), .A2(n10031), .ZN(n10123) );
  INV_X1 U12508 ( .A(n10669), .ZN(n10307) );
  INV_X1 U12509 ( .A(n13628), .ZN(n10672) );
  OAI21_X1 U12510 ( .B1(n10672), .B2(n13535), .A(n10041), .ZN(n10042) );
  NOR2_X1 U12511 ( .A1(n10042), .A2(n10121), .ZN(n10122) );
  AOI21_X1 U12512 ( .B1(n10121), .B2(n10042), .A(n10122), .ZN(n13640) );
  INV_X1 U12513 ( .A(n13640), .ZN(n10052) );
  INV_X1 U12514 ( .A(n10048), .ZN(n10047) );
  NAND2_X1 U12515 ( .A1(n14592), .A2(n10043), .ZN(n10044) );
  NOR2_X1 U12516 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  INV_X1 U12517 ( .A(n14415), .ZN(n14397) );
  NAND2_X1 U12518 ( .A1(n10709), .A2(n10049), .ZN(n10152) );
  NAND2_X1 U12519 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10152), .ZN(n10050) );
  OAI21_X1 U12520 ( .B1(n14397), .B2(n10125), .A(n10050), .ZN(n10051) );
  AOI21_X1 U12521 ( .B1(n10052), .B2(n14421), .A(n10051), .ZN(n10053) );
  OAI21_X1 U12522 ( .B1(n10669), .B2(n14419), .A(n10053), .ZN(P1_U3232) );
  INV_X1 U12523 ( .A(n10054), .ZN(n10056) );
  OAI222_X1 U12524 ( .A1(n13743), .A2(P1_U3086), .B1(n14198), .B2(n10056), 
        .C1(n10055), .C2(n14195), .ZN(P1_U3342) );
  INV_X1 U12525 ( .A(n11448), .ZN(n14657) );
  OAI222_X1 U12526 ( .A1(n13377), .A2(n10057), .B1(n13373), .B2(n10056), .C1(
        P2_U3088), .C2(n14657), .ZN(P2_U3314) );
  INV_X2 U12527 ( .A(n14769), .ZN(n14754) );
  INV_X1 U12528 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12529 ( .A1(n10917), .A2(n14761), .ZN(n13287) );
  OR2_X1 U12530 ( .A1(n11784), .A2(n12978), .ZN(n10058) );
  NAND2_X1 U12531 ( .A1(n10059), .A2(n10058), .ZN(n10176) );
  INV_X1 U12532 ( .A(n12977), .ZN(n10187) );
  XNOR2_X1 U12533 ( .A(n10176), .B(n10185), .ZN(n10882) );
  NAND2_X1 U12534 ( .A1(n10283), .A2(n11784), .ZN(n10061) );
  XNOR2_X1 U12535 ( .A(n10186), .B(n11991), .ZN(n10064) );
  INV_X2 U12536 ( .A(n12919), .ZN(n12906) );
  NAND2_X1 U12537 ( .A1(n12906), .A2(n12978), .ZN(n10063) );
  NAND2_X1 U12538 ( .A1(n6433), .A2(n12976), .ZN(n10062) );
  AND2_X1 U12539 ( .A1(n10063), .A2(n10062), .ZN(n10287) );
  OAI21_X1 U12540 ( .B1(n10064), .B2(n7052), .A(n10287), .ZN(n10879) );
  INV_X1 U12541 ( .A(n10879), .ZN(n10067) );
  AND2_X1 U12542 ( .A1(n10931), .A2(n11780), .ZN(n10074) );
  NAND2_X1 U12543 ( .A1(n10074), .A2(n10060), .ZN(n10959) );
  OAI211_X1 U12544 ( .C1(n10060), .C2(n10074), .A(n10959), .B(n13206), .ZN(
        n10876) );
  INV_X1 U12545 ( .A(n10876), .ZN(n10065) );
  AOI21_X1 U12546 ( .B1(n13261), .B2(n11793), .A(n10065), .ZN(n10066) );
  OAI211_X1 U12547 ( .C1(n14749), .C2(n10882), .A(n10067), .B(n10066), .ZN(
        n13341) );
  NAND2_X1 U12548 ( .A1(n13341), .A2(n14754), .ZN(n10068) );
  OAI21_X1 U12549 ( .B1(n14754), .B2(n10069), .A(n10068), .ZN(P2_U3436) );
  INV_X1 U12550 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10078) );
  XOR2_X1 U12551 ( .A(n11990), .B(n10296), .Z(n10938) );
  NAND2_X1 U12552 ( .A1(n12906), .A2(n12979), .ZN(n10071) );
  NAND2_X1 U12554 ( .A1(n6433), .A2(n12977), .ZN(n10070) );
  NAND2_X1 U12555 ( .A1(n10071), .A2(n10070), .ZN(n10929) );
  NAND2_X1 U12556 ( .A1(n10297), .A2(n11784), .ZN(n10072) );
  NAND2_X1 U12557 ( .A1(n10072), .A2(n13206), .ZN(n10073) );
  NOR2_X1 U12558 ( .A1(n10074), .A2(n10073), .ZN(n10934) );
  AOI211_X1 U12559 ( .C1(n13261), .C2(n11784), .A(n10929), .B(n10934), .ZN(
        n10076) );
  XNOR2_X1 U12560 ( .A(n11990), .B(n10276), .ZN(n10935) );
  NAND2_X1 U12561 ( .A1(n10935), .A2(n13287), .ZN(n10075) );
  OAI211_X1 U12562 ( .C1(n7052), .C2(n10938), .A(n10076), .B(n10075), .ZN(
        n10158) );
  NAND2_X1 U12563 ( .A1(n10158), .A2(n14754), .ZN(n10077) );
  OAI21_X1 U12564 ( .B1(n14754), .B2(n10078), .A(n10077), .ZN(P2_U3433) );
  AND2_X1 U12565 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10463) );
  INV_X1 U12566 ( .A(n14696), .ZN(n13050) );
  AND3_X1 U12567 ( .A1(n14624), .A2(n10080), .A3(n10079), .ZN(n10081) );
  NOR3_X1 U12568 ( .A1(n13050), .A2(n10082), .A3(n10081), .ZN(n10083) );
  AOI211_X1 U12569 ( .C1(n14680), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10463), .B(
        n10083), .ZN(n10089) );
  OR3_X1 U12570 ( .A1(n14620), .A2(n10085), .A3(n10084), .ZN(n10086) );
  NAND3_X1 U12571 ( .A1(n14683), .A2(n10087), .A3(n10086), .ZN(n10088) );
  OAI211_X1 U12572 ( .C1(n14658), .C2(n10090), .A(n10089), .B(n10088), .ZN(
        P2_U3219) );
  INV_X1 U12573 ( .A(n9694), .ZN(n10091) );
  INV_X1 U12574 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U12575 ( .A1(n10118), .A2(n10092), .ZN(P3_U3244) );
  CLKBUF_X1 U12576 ( .A(n10093), .Z(n10118) );
  INV_X1 U12577 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10094) );
  NOR2_X1 U12578 ( .A1(n10118), .A2(n10094), .ZN(P3_U3263) );
  INV_X1 U12579 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U12580 ( .A1(n10093), .A2(n10095), .ZN(P3_U3262) );
  INV_X1 U12581 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U12582 ( .A1(n10118), .A2(n10096), .ZN(P3_U3261) );
  INV_X1 U12583 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10097) );
  NOR2_X1 U12584 ( .A1(n10093), .A2(n10097), .ZN(P3_U3260) );
  INV_X1 U12585 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U12586 ( .A1(n10093), .A2(n15132), .ZN(P3_U3242) );
  INV_X1 U12587 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15056) );
  NOR2_X1 U12588 ( .A1(n10093), .A2(n15056), .ZN(P3_U3241) );
  INV_X1 U12589 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U12590 ( .A1(n10093), .A2(n10098), .ZN(P3_U3240) );
  INV_X1 U12591 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n15113) );
  NOR2_X1 U12592 ( .A1(n10118), .A2(n15113), .ZN(P3_U3259) );
  INV_X1 U12593 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U12594 ( .A1(n10093), .A2(n10099), .ZN(P3_U3258) );
  INV_X1 U12595 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10100) );
  NOR2_X1 U12596 ( .A1(n10118), .A2(n10100), .ZN(P3_U3257) );
  INV_X1 U12597 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10101) );
  NOR2_X1 U12598 ( .A1(n10118), .A2(n10101), .ZN(P3_U3256) );
  INV_X1 U12599 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U12600 ( .A1(n10118), .A2(n10102), .ZN(P3_U3255) );
  INV_X1 U12601 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U12602 ( .A1(n10118), .A2(n10103), .ZN(P3_U3254) );
  INV_X1 U12603 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10104) );
  NOR2_X1 U12604 ( .A1(n10118), .A2(n10104), .ZN(P3_U3253) );
  INV_X1 U12605 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U12606 ( .A1(n10118), .A2(n10105), .ZN(P3_U3252) );
  INV_X1 U12607 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U12608 ( .A1(n10118), .A2(n10106), .ZN(P3_U3251) );
  INV_X1 U12609 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10107) );
  NOR2_X1 U12610 ( .A1(n10093), .A2(n10107), .ZN(P3_U3245) );
  INV_X1 U12611 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10108) );
  NOR2_X1 U12612 ( .A1(n10093), .A2(n10108), .ZN(P3_U3234) );
  INV_X1 U12613 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U12614 ( .A1(n10118), .A2(n10109), .ZN(P3_U3248) );
  INV_X1 U12615 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U12616 ( .A1(n10118), .A2(n10110), .ZN(P3_U3249) );
  INV_X1 U12617 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10111) );
  NOR2_X1 U12618 ( .A1(n10118), .A2(n10111), .ZN(P3_U3250) );
  INV_X1 U12619 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U12620 ( .A1(n10093), .A2(n10112), .ZN(P3_U3238) );
  INV_X1 U12621 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U12622 ( .A1(n10093), .A2(n10113), .ZN(P3_U3235) );
  INV_X1 U12623 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U12624 ( .A1(n10093), .A2(n10114), .ZN(P3_U3243) );
  INV_X1 U12625 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U12626 ( .A1(n10118), .A2(n10115), .ZN(P3_U3247) );
  INV_X1 U12627 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U12628 ( .A1(n10118), .A2(n10116), .ZN(P3_U3237) );
  INV_X1 U12629 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U12630 ( .A1(n10118), .A2(n10117), .ZN(P3_U3246) );
  INV_X1 U12631 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U12632 ( .A1(n10118), .A2(n10119), .ZN(P3_U3236) );
  INV_X1 U12633 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U12634 ( .A1(n10118), .A2(n10120), .ZN(P3_U3239) );
  NOR2_X1 U12635 ( .A1(n10122), .A2(n7394), .ZN(n10130) );
  OAI22_X1 U12636 ( .A1(n13535), .A2(n10125), .B1(n14532), .B2(n11278), .ZN(
        n10126) );
  INV_X1 U12637 ( .A(n10126), .ZN(n10127) );
  OAI21_X1 U12638 ( .B1(n10128), .B2(n10127), .A(n10144), .ZN(n10129) );
  AOI21_X1 U12639 ( .B1(n10130), .B2(n10129), .A(n10146), .ZN(n10135) );
  INV_X1 U12640 ( .A(n14532), .ZN(n10676) );
  INV_X1 U12641 ( .A(n10152), .ZN(n10132) );
  INV_X1 U12642 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U12643 ( .A1(n14379), .A2(n14252), .ZN(n14394) );
  INV_X1 U12644 ( .A(n14394), .ZN(n14417) );
  AOI22_X1 U12645 ( .A1(n14417), .A2(n13628), .B1(n14415), .B2(n13626), .ZN(
        n10131) );
  OAI21_X1 U12646 ( .B1(n10132), .B2(n10677), .A(n10131), .ZN(n10133) );
  AOI21_X1 U12647 ( .B1(n14407), .B2(n10676), .A(n10133), .ZN(n10134) );
  OAI21_X1 U12648 ( .B1(n10135), .B2(n14401), .A(n10134), .ZN(P1_U3222) );
  AOI22_X1 U12649 ( .A1(n14683), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14696), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U12650 ( .A1(n14696), .A2(n10136), .ZN(n10137) );
  OAI211_X1 U12651 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14700), .A(n14658), .B(
        n10137), .ZN(n10138) );
  INV_X1 U12652 ( .A(n10138), .ZN(n10139) );
  MUX2_X1 U12653 ( .A(n10140), .B(n10139), .S(P2_IR_REG_0__SCAN_IN), .Z(n10143) );
  NOR2_X1 U12654 ( .A1(n10292), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10141) );
  AOI21_X1 U12655 ( .B1(n14680), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n10141), .ZN(
        n10142) );
  NAND2_X1 U12656 ( .A1(n10143), .A2(n10142), .ZN(P2_U3214) );
  INV_X1 U12657 ( .A(n10144), .ZN(n10145) );
  OAI22_X1 U12658 ( .A1(n8526), .A2(n11278), .B1(n10124), .B2(n10355), .ZN(
        n10147) );
  XNOR2_X1 U12659 ( .A(n10147), .B(n13395), .ZN(n10684) );
  OAI22_X1 U12660 ( .A1(n13535), .A2(n8526), .B1(n10355), .B2(n13536), .ZN(
        n10683) );
  XNOR2_X1 U12661 ( .A(n10684), .B(n10683), .ZN(n10148) );
  AOI21_X1 U12662 ( .B1(n10149), .B2(n10148), .A(n10685), .ZN(n10155) );
  NAND2_X1 U12663 ( .A1(n13627), .A2(n14252), .ZN(n10151) );
  NAND2_X1 U12664 ( .A1(n13625), .A2(n14254), .ZN(n10150) );
  NAND2_X1 U12665 ( .A1(n10151), .A2(n10150), .ZN(n10317) );
  AOI22_X1 U12666 ( .A1(n14379), .A2(n10317), .B1(n10152), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10154) );
  NAND2_X1 U12667 ( .A1(n14407), .A2(n8525), .ZN(n10153) );
  OAI211_X1 U12668 ( .C1(n10155), .C2(n14401), .A(n10154), .B(n10153), .ZN(
        P1_U3237) );
  OAI222_X1 U12669 ( .A1(P3_U3151), .A2(n12392), .B1(n12817), .B2(n10157), 
        .C1(n12821), .C2(n10156), .ZN(P3_U3276) );
  NAND2_X1 U12670 ( .A1(n10158), .A2(n6436), .ZN(n10159) );
  OAI21_X1 U12671 ( .B1(n6436), .B2(n12986), .A(n10159), .ZN(P2_U3500) );
  INV_X1 U12672 ( .A(n10160), .ZN(n10204) );
  INV_X1 U12673 ( .A(n11444), .ZN(n11588) );
  OAI222_X1 U12674 ( .A1(n13373), .A2(n10204), .B1(n11588), .B2(P2_U3088), 
        .C1(n10161), .C2(n13377), .ZN(P2_U3311) );
  AOI21_X1 U12675 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10166), .A(n10162), .ZN(
        n14648) );
  MUX2_X1 U12676 ( .A(n9259), .B(P2_REG2_REG_9__SCAN_IN), .S(n10167), .Z(
        n14647) );
  NAND2_X1 U12677 ( .A1(n14648), .A2(n14647), .ZN(n14646) );
  OAI21_X1 U12678 ( .B1(n14650), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14646), .ZN(
        n10164) );
  MUX2_X1 U12679 ( .A(n10867), .B(P2_REG2_REG_10__SCAN_IN), .S(n10210), .Z(
        n10163) );
  AOI211_X1 U12680 ( .C1(n10164), .C2(n10163), .A(n14700), .B(n10207), .ZN(
        n10175) );
  AOI21_X1 U12681 ( .B1(n10166), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10165), .ZN(
        n14645) );
  MUX2_X1 U12682 ( .A(n9254), .B(P2_REG1_REG_9__SCAN_IN), .S(n10167), .Z(
        n14644) );
  NAND2_X1 U12683 ( .A1(n14645), .A2(n14644), .ZN(n14643) );
  OAI21_X1 U12684 ( .B1(n14650), .B2(P2_REG1_REG_9__SCAN_IN), .A(n14643), .ZN(
        n10170) );
  MUX2_X1 U12685 ( .A(n9272), .B(P2_REG1_REG_10__SCAN_IN), .S(n10210), .Z(
        n10169) );
  INV_X1 U12686 ( .A(n10213), .ZN(n10168) );
  AOI211_X1 U12687 ( .C1(n10170), .C2(n10169), .A(n13050), .B(n10168), .ZN(
        n10174) );
  NAND2_X1 U12688 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11205)
         );
  NAND2_X1 U12689 ( .A1(n14680), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10171) );
  OAI211_X1 U12690 ( .C1(n14658), .C2(n10172), .A(n11205), .B(n10171), .ZN(
        n10173) );
  OR3_X1 U12691 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(P2_U3224) );
  INV_X1 U12692 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15024) );
  NAND2_X1 U12693 ( .A1(n10176), .A2(n11991), .ZN(n10178) );
  OR2_X1 U12694 ( .A1(n11793), .A2(n12977), .ZN(n10177) );
  NAND2_X1 U12695 ( .A1(n10178), .A2(n10177), .ZN(n10956) );
  XNOR2_X1 U12696 ( .A(n14730), .B(n12976), .ZN(n11993) );
  INV_X1 U12697 ( .A(n11993), .ZN(n10179) );
  NAND2_X1 U12698 ( .A1(n10956), .A2(n10179), .ZN(n10181) );
  OR2_X1 U12699 ( .A1(n14730), .A2(n12976), .ZN(n10180) );
  NAND2_X1 U12700 ( .A1(n10181), .A2(n10180), .ZN(n10897) );
  XNOR2_X1 U12701 ( .A(n11806), .B(n12975), .ZN(n11994) );
  INV_X1 U12702 ( .A(n11994), .ZN(n10898) );
  NAND2_X1 U12703 ( .A1(n10897), .A2(n10898), .ZN(n10183) );
  OR2_X1 U12704 ( .A1(n11806), .A2(n12975), .ZN(n10182) );
  NAND2_X1 U12705 ( .A1(n10183), .A2(n10182), .ZN(n10243) );
  XNOR2_X1 U12706 ( .A(n11810), .B(n12974), .ZN(n11996) );
  XNOR2_X1 U12707 ( .A(n10243), .B(n11996), .ZN(n10955) );
  INV_X1 U12708 ( .A(n10906), .ZN(n10184) );
  INV_X1 U12709 ( .A(n11810), .ZN(n10950) );
  AOI211_X1 U12710 ( .C1(n11810), .C2(n10184), .A(n13221), .B(n10246), .ZN(
        n10952) );
  AOI21_X1 U12711 ( .B1(n13261), .B2(n11810), .A(n10952), .ZN(n10199) );
  NAND2_X1 U12712 ( .A1(n10186), .A2(n10185), .ZN(n10189) );
  NAND2_X1 U12713 ( .A1(n10187), .A2(n11793), .ZN(n10188) );
  NAND2_X1 U12714 ( .A1(n10960), .A2(n11993), .ZN(n10191) );
  INV_X1 U12715 ( .A(n12976), .ZN(n10338) );
  NAND2_X1 U12716 ( .A1(n14730), .A2(n10338), .ZN(n10190) );
  NAND2_X1 U12717 ( .A1(n10191), .A2(n10190), .ZN(n10899) );
  NAND2_X1 U12718 ( .A1(n10899), .A2(n11994), .ZN(n10194) );
  INV_X1 U12719 ( .A(n12975), .ZN(n10192) );
  NAND2_X1 U12720 ( .A1(n11806), .A2(n10192), .ZN(n10193) );
  XNOR2_X1 U12721 ( .A(n10249), .B(n11996), .ZN(n10198) );
  NAND2_X1 U12722 ( .A1(n12906), .A2(n12975), .ZN(n10196) );
  NAND2_X1 U12723 ( .A1(n6433), .A2(n12973), .ZN(n10195) );
  AND2_X1 U12724 ( .A1(n10196), .A2(n10195), .ZN(n10466) );
  INV_X1 U12725 ( .A(n10466), .ZN(n10197) );
  AOI21_X1 U12726 ( .B1(n10198), .B2(n14753), .A(n10197), .ZN(n10948) );
  OAI211_X1 U12727 ( .C1(n14749), .C2(n10955), .A(n10199), .B(n10948), .ZN(
        n10201) );
  NAND2_X1 U12728 ( .A1(n10201), .A2(n14754), .ZN(n10200) );
  OAI21_X1 U12729 ( .B1(n14754), .B2(n15024), .A(n10200), .ZN(P2_U3445) );
  NAND2_X1 U12730 ( .A1(n10201), .A2(n6436), .ZN(n10202) );
  OAI21_X1 U12731 ( .B1(n6436), .B2(n9964), .A(n10202), .ZN(P2_U3504) );
  INV_X1 U12732 ( .A(n13756), .ZN(n11252) );
  OAI222_X1 U12733 ( .A1(P1_U3086), .A2(n11252), .B1(n14198), .B2(n10204), 
        .C1(n10203), .C2(n14195), .ZN(P1_U3339) );
  INV_X1 U12734 ( .A(n11249), .ZN(n11258) );
  INV_X1 U12735 ( .A(n10205), .ZN(n10236) );
  OAI222_X1 U12736 ( .A1(P1_U3086), .A2(n11258), .B1(n14198), .B2(n10236), 
        .C1(n10206), .C2(n14195), .ZN(P1_U3341) );
  INV_X1 U12737 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10208) );
  MUX2_X1 U12738 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10208), .S(n11446), .Z(
        n10209) );
  AOI21_X1 U12739 ( .B1(n6453), .B2(n6723), .A(n13021), .ZN(n10218) );
  INV_X1 U12740 ( .A(n14680), .ZN(n14705) );
  OAI22_X1 U12741 ( .A1(n14705), .A2(n6752), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9293), .ZN(n10216) );
  NAND2_X1 U12742 ( .A1(n10210), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10212) );
  INV_X1 U12743 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11025) );
  MUX2_X1 U12744 ( .A(n11025), .B(P2_REG1_REG_11__SCAN_IN), .S(n11446), .Z(
        n10211) );
  AOI21_X1 U12745 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n11445) );
  AND3_X1 U12746 ( .A1(n10213), .A2(n10212), .A3(n10211), .ZN(n10214) );
  NOR3_X1 U12747 ( .A1(n11445), .A2(n10214), .A3(n13050), .ZN(n10215) );
  AOI211_X1 U12748 ( .C1(n14694), .C2(n11446), .A(n10216), .B(n10215), .ZN(
        n10217) );
  OAI21_X1 U12749 ( .B1(n10218), .B2(n14700), .A(n10217), .ZN(P2_U3225) );
  INV_X1 U12750 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U12751 ( .A1(n11249), .A2(n15088), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11258), .ZN(n10223) );
  AOI21_X1 U12752 ( .B1(n10012), .B2(n10220), .A(n10219), .ZN(n13742) );
  MUX2_X1 U12753 ( .A(n10221), .B(P1_REG1_REG_13__SCAN_IN), .S(n13743), .Z(
        n13741) );
  NAND2_X1 U12754 ( .A1(n13742), .A2(n13741), .ZN(n13740) );
  OAI21_X1 U12755 ( .B1(n13743), .B2(n10221), .A(n13740), .ZN(n10222) );
  NOR2_X1 U12756 ( .A1(n10223), .A2(n10222), .ZN(n11257) );
  AOI21_X1 U12757 ( .B1(n10223), .B2(n10222), .A(n11257), .ZN(n10235) );
  NAND2_X1 U12758 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14366)
         );
  NAND2_X1 U12759 ( .A1(n14497), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10224) );
  OAI211_X1 U12760 ( .C1(n14524), .C2(n11258), .A(n14366), .B(n10224), .ZN(
        n10225) );
  INV_X1 U12761 ( .A(n10225), .ZN(n10234) );
  MUX2_X1 U12762 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10226), .S(n11249), .Z(
        n10232) );
  MUX2_X1 U12763 ( .A(n10227), .B(P1_REG2_REG_13__SCAN_IN), .S(n13743), .Z(
        n13746) );
  NOR2_X1 U12764 ( .A1(n10228), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U12765 ( .A1(n10230), .A2(n10229), .ZN(n13747) );
  NAND2_X1 U12766 ( .A1(n13746), .A2(n13747), .ZN(n13745) );
  OAI21_X1 U12767 ( .B1(n13743), .B2(n10227), .A(n13745), .ZN(n10231) );
  NAND2_X1 U12768 ( .A1(n10232), .A2(n10231), .ZN(n11247) );
  OAI211_X1 U12769 ( .C1(n10232), .C2(n10231), .A(n11247), .B(n14492), .ZN(
        n10233) );
  OAI211_X1 U12770 ( .C1(n10235), .C2(n14522), .A(n10234), .B(n10233), .ZN(
        P1_U3257) );
  INV_X1 U12771 ( .A(n14672), .ZN(n11451) );
  OAI222_X1 U12772 ( .A1(n13377), .A2(n10237), .B1(n11451), .B2(P2_U3088), 
        .C1(n13373), .C2(n10236), .ZN(P2_U3313) );
  INV_X1 U12773 ( .A(n10238), .ZN(n10241) );
  INV_X1 U12774 ( .A(n11589), .ZN(n13044) );
  OAI222_X1 U12775 ( .A1(n13373), .A2(n10241), .B1(n13044), .B2(P2_U3088), 
        .C1(n10239), .C2(n13377), .ZN(P2_U3310) );
  INV_X1 U12776 ( .A(n11254), .ZN(n13764) );
  OAI222_X1 U12777 ( .A1(P1_U3086), .A2(n13764), .B1(n14198), .B2(n10241), 
        .C1(n10240), .C2(n14195), .ZN(P1_U3338) );
  INV_X1 U12778 ( .A(n11996), .ZN(n10242) );
  NAND2_X1 U12779 ( .A1(n10243), .A2(n10242), .ZN(n10245) );
  OR2_X1 U12780 ( .A1(n11810), .A2(n12974), .ZN(n10244) );
  NAND2_X1 U12781 ( .A1(n10245), .A2(n10244), .ZN(n10822) );
  INV_X1 U12782 ( .A(n12973), .ZN(n10831) );
  XNOR2_X1 U12783 ( .A(n11819), .B(n10831), .ZN(n11998) );
  INV_X1 U12784 ( .A(n11998), .ZN(n10829) );
  XNOR2_X1 U12785 ( .A(n10822), .B(n10829), .ZN(n10946) );
  INV_X1 U12786 ( .A(n10246), .ZN(n10248) );
  INV_X1 U12787 ( .A(n11819), .ZN(n10941) );
  INV_X1 U12788 ( .A(n11028), .ZN(n10247) );
  AOI211_X1 U12789 ( .C1(n11819), .C2(n10248), .A(n13221), .B(n10247), .ZN(
        n10943) );
  AOI21_X1 U12790 ( .B1(n13261), .B2(n11819), .A(n10943), .ZN(n10257) );
  NAND2_X1 U12791 ( .A1(n10249), .A2(n11996), .ZN(n10252) );
  INV_X1 U12792 ( .A(n12974), .ZN(n10250) );
  NAND2_X1 U12793 ( .A1(n11810), .A2(n10250), .ZN(n10251) );
  NAND2_X1 U12794 ( .A1(n10252), .A2(n10251), .ZN(n10830) );
  XNOR2_X1 U12795 ( .A(n10830), .B(n10829), .ZN(n10256) );
  NAND2_X1 U12796 ( .A1(n12906), .A2(n12974), .ZN(n10254) );
  NAND2_X1 U12797 ( .A1(n6433), .A2(n12972), .ZN(n10253) );
  AND2_X1 U12798 ( .A1(n10254), .A2(n10253), .ZN(n10983) );
  INV_X1 U12799 ( .A(n10983), .ZN(n10255) );
  AOI21_X1 U12800 ( .B1(n10256), .B2(n14753), .A(n10255), .ZN(n10939) );
  OAI211_X1 U12801 ( .C1(n14749), .C2(n10946), .A(n10257), .B(n10939), .ZN(
        n10263) );
  NAND2_X1 U12802 ( .A1(n10263), .A2(n14754), .ZN(n10258) );
  OAI21_X1 U12803 ( .B1(n14754), .B2(n9202), .A(n10258), .ZN(P2_U3448) );
  INV_X1 U12804 ( .A(n10259), .ZN(n10262) );
  INV_X1 U12805 ( .A(n14681), .ZN(n11452) );
  OAI222_X1 U12806 ( .A1(n13377), .A2(n10260), .B1(n13373), .B2(n10262), .C1(
        P2_U3088), .C2(n11452), .ZN(P2_U3312) );
  INV_X1 U12807 ( .A(n11259), .ZN(n14510) );
  OAI222_X1 U12808 ( .A1(n14510), .A2(P1_U3086), .B1(n14198), .B2(n10262), 
        .C1(n10261), .C2(n14195), .ZN(P1_U3340) );
  NAND2_X1 U12809 ( .A1(n10263), .A2(n6436), .ZN(n10264) );
  OAI21_X1 U12810 ( .B1(n6436), .B2(n10265), .A(n10264), .ZN(P2_U3505) );
  NOR2_X1 U12811 ( .A1(n12248), .A2(P3_U3151), .ZN(n10646) );
  INV_X1 U12812 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10719) );
  INV_X1 U12813 ( .A(n10628), .ZN(n10267) );
  OAI22_X1 U12814 ( .A1(n12244), .A2(n14918), .B1(n12245), .B2(n10668), .ZN(
        n10266) );
  AOI21_X1 U12815 ( .B1(n12229), .B2(n10267), .A(n10266), .ZN(n10268) );
  OAI21_X1 U12816 ( .B1(n10646), .B2(n10719), .A(n10268), .ZN(P3_U3172) );
  INV_X1 U12817 ( .A(n10269), .ZN(n10272) );
  INV_X1 U12818 ( .A(n10270), .ZN(n10271) );
  AOI21_X1 U12819 ( .B1(n10272), .B2(n10277), .A(n10271), .ZN(n10281) );
  INV_X1 U12820 ( .A(n10929), .ZN(n10274) );
  NOR2_X1 U12821 ( .A1(n10273), .A2(P2_U3088), .ZN(n10293) );
  OAI22_X1 U12822 ( .A1(n12908), .A2(n10274), .B1(n10293), .B2(n10930), .ZN(
        n10275) );
  AOI21_X1 U12823 ( .B1(n11784), .B2(n12943), .A(n10275), .ZN(n10280) );
  NOR2_X1 U12824 ( .A1(n12928), .A2(n13206), .ZN(n12934) );
  INV_X1 U12825 ( .A(n10276), .ZN(n10278) );
  NAND3_X1 U12826 ( .A1(n12934), .A2(n10278), .A3(n10277), .ZN(n10279) );
  OAI211_X1 U12827 ( .C1(n10281), .C2(n12928), .A(n10280), .B(n10279), .ZN(
        P2_U3194) );
  INV_X1 U12828 ( .A(n12934), .ZN(n12858) );
  OAI22_X1 U12829 ( .A1(n12858), .A2(n10283), .B1(n10282), .B2(n12928), .ZN(
        n10286) );
  INV_X1 U12830 ( .A(n10284), .ZN(n10285) );
  NAND3_X1 U12831 ( .A1(n10286), .A2(n10285), .A3(n10270), .ZN(n10290) );
  OAI22_X1 U12832 ( .A1(n12908), .A2(n10287), .B1(n10293), .B2(n10874), .ZN(
        n10288) );
  AOI21_X1 U12833 ( .B1(n11793), .B2(n12943), .A(n10288), .ZN(n10289) );
  OAI211_X1 U12834 ( .C1(n12928), .C2(n10291), .A(n10290), .B(n10289), .ZN(
        P2_U3209) );
  OAI22_X1 U12835 ( .A1(n12908), .A2(n10294), .B1(n10293), .B2(n10292), .ZN(
        n10295) );
  AOI21_X1 U12836 ( .B1(n12934), .B2(n11783), .A(n10295), .ZN(n10300) );
  OAI21_X1 U12837 ( .B1(n11780), .B2(n13221), .A(n10296), .ZN(n10298) );
  AOI22_X1 U12838 ( .A1(n6591), .A2(n10298), .B1(n12943), .B2(n10297), .ZN(
        n10299) );
  NAND2_X1 U12839 ( .A1(n10300), .A2(n10299), .ZN(P2_U3204) );
  NOR2_X1 U12840 ( .A1(n10302), .A2(n10301), .ZN(n10304) );
  INV_X1 U12841 ( .A(n10347), .ZN(n13850) );
  INV_X2 U12842 ( .A(n14042), .ZN(n15146) );
  INV_X1 U12843 ( .A(n10353), .ZN(n10316) );
  NAND2_X1 U12844 ( .A1(n13628), .A2(n10307), .ZN(n10675) );
  NAND2_X1 U12845 ( .A1(n10308), .A2(n10675), .ZN(n10310) );
  NAND2_X1 U12846 ( .A1(n10125), .A2(n14532), .ZN(n10309) );
  XNOR2_X1 U12847 ( .A(n10316), .B(n10354), .ZN(n10320) );
  NAND2_X1 U12848 ( .A1(n10312), .A2(n10311), .ZN(n10314) );
  NAND2_X1 U12849 ( .A1(n10315), .A2(n10316), .ZN(n10351) );
  OAI21_X1 U12850 ( .B1(n10316), .B2(n10315), .A(n10351), .ZN(n10318) );
  AOI21_X1 U12851 ( .B1(n10318), .B2(n14554), .A(n10317), .ZN(n10319) );
  OAI21_X1 U12852 ( .B1(n10320), .B2(n14578), .A(n10319), .ZN(n14539) );
  INV_X1 U12853 ( .A(n14539), .ZN(n10328) );
  AND2_X1 U12854 ( .A1(n14532), .A2(n10669), .ZN(n10671) );
  OAI21_X1 U12855 ( .B1(n10671), .B2(n10355), .A(n14548), .ZN(n10322) );
  NOR2_X1 U12856 ( .A1(n10323), .A2(n10602), .ZN(n10324) );
  INV_X1 U12857 ( .A(n15144), .ZN(n14040) );
  AOI22_X1 U12858 ( .A1(n14042), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14040), .ZN(n10325) );
  OAI21_X1 U12859 ( .B1(n10355), .B2(n14260), .A(n10325), .ZN(n10326) );
  AOI21_X1 U12860 ( .B1(n14247), .B2(n6579), .A(n10326), .ZN(n10327) );
  OAI21_X1 U12861 ( .B1(n14258), .B2(n10328), .A(n10327), .ZN(P1_U3291) );
  INV_X1 U12862 ( .A(n10329), .ZN(n10369) );
  INV_X1 U12863 ( .A(n10336), .ZN(n10331) );
  INV_X1 U12864 ( .A(n10330), .ZN(n10470) );
  AOI21_X1 U12865 ( .B1(n10369), .B2(n10331), .A(n10470), .ZN(n10342) );
  NAND2_X1 U12866 ( .A1(n12906), .A2(n12976), .ZN(n10333) );
  NAND2_X1 U12867 ( .A1(n6433), .A2(n12974), .ZN(n10332) );
  AND2_X1 U12868 ( .A1(n10333), .A2(n10332), .ZN(n10900) );
  INV_X1 U12869 ( .A(n10907), .ZN(n10334) );
  AOI22_X1 U12870 ( .A1(n12898), .A2(n10334), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10335) );
  OAI21_X1 U12871 ( .B1(n12908), .B2(n10900), .A(n10335), .ZN(n10340) );
  NOR4_X1 U12872 ( .A1(n12858), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10339) );
  AOI211_X1 U12873 ( .C1(n11806), .C2(n12943), .A(n10340), .B(n10339), .ZN(
        n10341) );
  OAI21_X1 U12874 ( .B1(n10342), .B2(n12928), .A(n10341), .ZN(P2_U3202) );
  OAI222_X1 U12875 ( .A1(P3_U3151), .A2(n10345), .B1(n12817), .B2(n10344), 
        .C1(n12821), .C2(n10343), .ZN(P3_U3275) );
  INV_X1 U12876 ( .A(n10346), .ZN(n14025) );
  AND2_X1 U12877 ( .A1(n10347), .A2(n14025), .ZN(n13792) );
  INV_X1 U12878 ( .A(n13792), .ZN(n15152) );
  NAND2_X1 U12879 ( .A1(n10348), .A2(n8735), .ZN(n10608) );
  OR2_X1 U12880 ( .A1(n10348), .A2(n8735), .ZN(n10349) );
  NAND2_X1 U12881 ( .A1(n10608), .A2(n10349), .ZN(n14542) );
  INV_X1 U12882 ( .A(n10381), .ZN(n10358) );
  NAND2_X1 U12883 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  NAND2_X1 U12884 ( .A1(n10352), .A2(n10358), .ZN(n10376) );
  OAI21_X1 U12885 ( .B1(n10358), .B2(n10352), .A(n10376), .ZN(n10362) );
  OAI22_X1 U12886 ( .A1(n10712), .A2(n13951), .B1(n8526), .B2(n13949), .ZN(
        n10361) );
  NAND2_X1 U12887 ( .A1(n10354), .A2(n10353), .ZN(n10357) );
  NAND2_X1 U12888 ( .A1(n8526), .A2(n10355), .ZN(n10356) );
  NAND2_X1 U12889 ( .A1(n10357), .A2(n10356), .ZN(n10382) );
  XNOR2_X1 U12890 ( .A(n10382), .B(n10358), .ZN(n10359) );
  NOR2_X1 U12891 ( .A1(n10359), .A2(n14578), .ZN(n10360) );
  MUX2_X1 U12892 ( .A(n10363), .B(n14541), .S(n15146), .Z(n10365) );
  INV_X1 U12893 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U12894 ( .A1(n15149), .A2(n13516), .B1(n14040), .B2(n13658), .ZN(
        n10364) );
  OAI211_X1 U12895 ( .C1(n15152), .C2(n14542), .A(n10365), .B(n10364), .ZN(
        P1_U3290) );
  NAND2_X1 U12896 ( .A1(n12906), .A2(n12977), .ZN(n10367) );
  NAND2_X1 U12897 ( .A1(n6433), .A2(n12975), .ZN(n10366) );
  AND2_X1 U12898 ( .A1(n10367), .A2(n10366), .ZN(n14727) );
  INV_X1 U12899 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U12900 ( .A1(n12898), .A2(n13011), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10368) );
  OAI21_X1 U12901 ( .B1(n12908), .B2(n14727), .A(n10368), .ZN(n10373) );
  AOI211_X1 U12902 ( .C1(n10371), .C2(n10370), .A(n12928), .B(n10369), .ZN(
        n10372) );
  AOI211_X1 U12903 ( .C1(n14730), .C2(n12943), .A(n10373), .B(n10372), .ZN(
        n10374) );
  INV_X1 U12904 ( .A(n10374), .ZN(P2_U3190) );
  OR2_X1 U12905 ( .A1(n10608), .A2(n10693), .ZN(n10790) );
  NOR2_X1 U12906 ( .A1(n10790), .A2(n14557), .ZN(n10789) );
  NAND2_X1 U12907 ( .A1(n10789), .A2(n14561), .ZN(n14572) );
  OAI211_X1 U12908 ( .C1(n10789), .C2(n14561), .A(n14572), .B(n14548), .ZN(
        n14559) );
  NAND2_X1 U12909 ( .A1(n13624), .A2(n10967), .ZN(n10377) );
  NAND2_X1 U12910 ( .A1(n10603), .A2(n10377), .ZN(n10379) );
  OR2_X1 U12911 ( .A1(n13624), .A2(n10967), .ZN(n10378) );
  NAND2_X1 U12912 ( .A1(n10379), .A2(n10378), .ZN(n10793) );
  INV_X1 U12913 ( .A(n13623), .ZN(n10391) );
  NAND2_X1 U12914 ( .A1(n14557), .A2(n10391), .ZN(n10380) );
  NAND2_X1 U12915 ( .A1(n10382), .A2(n10381), .ZN(n10384) );
  INV_X1 U12916 ( .A(n13625), .ZN(n10688) );
  NAND2_X1 U12917 ( .A1(n10688), .A2(n8735), .ZN(n10383) );
  INV_X1 U12918 ( .A(n10385), .ZN(n10386) );
  OAI21_X1 U12919 ( .B1(n10605), .B2(n10386), .A(n10387), .ZN(n10388) );
  INV_X1 U12920 ( .A(n10388), .ZN(n10795) );
  INV_X1 U12921 ( .A(n10389), .ZN(n10796) );
  OAI22_X1 U12922 ( .A1(n14571), .A2(n6570), .B1(n10725), .B2(n14578), .ZN(
        n10395) );
  INV_X1 U12923 ( .A(n13621), .ZN(n11165) );
  OAI22_X1 U12924 ( .A1(n11165), .A2(n13951), .B1(n10391), .B2(n13949), .ZN(
        n10394) );
  AOI22_X1 U12925 ( .A1(n6570), .A2(n14554), .B1(n10725), .B2(n14597), .ZN(
        n10392) );
  NOR2_X1 U12926 ( .A1(n10392), .A2(n10396), .ZN(n10393) );
  AOI211_X1 U12927 ( .C1(n10396), .C2(n10395), .A(n10394), .B(n10393), .ZN(
        n14560) );
  MUX2_X1 U12928 ( .A(n10397), .B(n14560), .S(n15146), .Z(n10400) );
  INV_X1 U12929 ( .A(n10784), .ZN(n10398) );
  AOI22_X1 U12930 ( .A1(n15149), .A2(n10786), .B1(n10398), .B2(n14040), .ZN(
        n10399) );
  OAI211_X1 U12931 ( .C1(n13998), .C2(n14559), .A(n10400), .B(n10399), .ZN(
        P1_U3287) );
  NAND2_X1 U12932 ( .A1(n14042), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10401) );
  OAI21_X1 U12933 ( .B1(n8540), .B2(n15144), .A(n10401), .ZN(n10403) );
  AOI21_X1 U12934 ( .B1(n15152), .B2(n14260), .A(n10669), .ZN(n10402) );
  AOI211_X1 U12935 ( .C1(n10404), .C2(n15146), .A(n10403), .B(n10402), .ZN(
        n10407) );
  OAI21_X1 U12936 ( .B1(n14248), .B2(n13863), .A(n10405), .ZN(n10406) );
  NAND2_X1 U12937 ( .A1(n10407), .A2(n10406), .ZN(P1_U3293) );
  INV_X1 U12938 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11174) );
  INV_X1 U12939 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15087) );
  MUX2_X1 U12940 ( .A(n11174), .B(n15087), .S(n8117), .Z(n10718) );
  NAND2_X1 U12941 ( .A1(n10718), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10717) );
  MUX2_X1 U12942 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n8117), .Z(n10408) );
  XNOR2_X1 U12943 ( .A(n10408), .B(n10557), .ZN(n10543) );
  INV_X1 U12944 ( .A(n10408), .ZN(n10409) );
  AOI22_X1 U12945 ( .A1(n10544), .A2(n10543), .B1(n10557), .B2(n10409), .ZN(
        n10577) );
  MUX2_X1 U12946 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n8117), .Z(n10410) );
  XOR2_X1 U12947 ( .A(n10586), .B(n10410), .Z(n10576) );
  INV_X1 U12948 ( .A(n10586), .ZN(n10444) );
  MUX2_X1 U12949 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n8117), .Z(n10411) );
  XNOR2_X1 U12950 ( .A(n10411), .B(n10573), .ZN(n10561) );
  INV_X1 U12951 ( .A(n10411), .ZN(n10412) );
  INV_X1 U12952 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14862) );
  INV_X1 U12953 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n14982) );
  MUX2_X1 U12954 ( .A(n14862), .B(n14982), .S(n8117), .Z(n10413) );
  NOR2_X1 U12955 ( .A1(n10413), .A2(n10756), .ZN(n10751) );
  AND2_X1 U12956 ( .A1(n10413), .A2(n10756), .ZN(n10750) );
  INV_X1 U12957 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11406) );
  INV_X1 U12958 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10414) );
  MUX2_X1 U12959 ( .A(n11406), .B(n10414), .S(n8117), .Z(n10415) );
  NAND2_X1 U12960 ( .A1(n10415), .A2(n10488), .ZN(n10484) );
  INV_X1 U12961 ( .A(n10415), .ZN(n10416) );
  NAND2_X1 U12962 ( .A1(n10416), .A2(n10451), .ZN(n10417) );
  AND2_X1 U12963 ( .A1(n10484), .A2(n10417), .ZN(n10418) );
  INV_X1 U12964 ( .A(n10485), .ZN(n10420) );
  NOR3_X1 U12965 ( .A1(n6569), .A2(n10750), .A3(n10418), .ZN(n10419) );
  AND2_X1 U12966 ( .A1(P3_U3897), .A2(n8119), .ZN(n14810) );
  OAI21_X1 U12967 ( .B1(n10420), .B2(n10419), .A(n14810), .ZN(n10462) );
  INV_X1 U12968 ( .A(n10660), .ZN(n10421) );
  NAND2_X1 U12969 ( .A1(n10421), .A2(n10884), .ZN(n10456) );
  NAND2_X1 U12970 ( .A1(n10619), .A2(n10422), .ZN(n10423) );
  NAND2_X1 U12971 ( .A1(n10424), .A2(n10423), .ZN(n10455) );
  INV_X1 U12972 ( .A(n10455), .ZN(n10425) );
  NAND2_X1 U12973 ( .A1(n10456), .A2(n10425), .ZN(n10438) );
  INV_X1 U12974 ( .A(n8119), .ZN(n10426) );
  MUX2_X1 U12975 ( .A(n10438), .B(n12258), .S(n10426), .Z(n12393) );
  INV_X1 U12976 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15096) );
  NOR2_X1 U12977 ( .A1(n11174), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U12978 ( .A1(n7465), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10428) );
  OAI21_X1 U12979 ( .B1(n10502), .B2(n10427), .A(n10428), .ZN(n10504) );
  INV_X1 U12980 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10503) );
  OR2_X1 U12981 ( .A1(n10504), .A2(n10503), .ZN(n10506) );
  NAND2_X1 U12982 ( .A1(n10506), .A2(n10428), .ZN(n10546) );
  NAND2_X1 U12983 ( .A1(n10547), .A2(n10546), .ZN(n10545) );
  OR2_X1 U12984 ( .A1(n10557), .A2(n15096), .ZN(n10429) );
  INV_X1 U12985 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U12986 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n10439), .ZN(n10430) );
  OAI21_X1 U12987 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10439), .A(n10430), .ZN(
        n10563) );
  AND2_X1 U12988 ( .A1(n10439), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U12989 ( .A1(n10433), .A2(n10448), .ZN(n10432) );
  INV_X1 U12990 ( .A(n10432), .ZN(n10434) );
  AOI22_X1 U12991 ( .A1(n10488), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11406), 
        .B2(n10451), .ZN(n10435) );
  AOI21_X1 U12992 ( .B1(n6584), .B2(n10435), .A(n10477), .ZN(n10459) );
  OR2_X1 U12993 ( .A1(n10438), .A2(n10437), .ZN(n12399) );
  NAND2_X1 U12994 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n10439), .ZN(n10447) );
  INV_X1 U12995 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n14980) );
  AOI22_X1 U12996 ( .A1(n10573), .A2(n14980), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n10439), .ZN(n10567) );
  INV_X1 U12997 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10440) );
  AND2_X1 U12998 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15037), .ZN(n10441) );
  OR3_X1 U12999 ( .A1(n15087), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        P3_IR_REG_1__SCAN_IN), .ZN(n10442) );
  INV_X1 U13000 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10510) );
  OR2_X1 U13001 ( .A1(n10509), .A2(n10510), .ZN(n10507) );
  NAND2_X1 U13002 ( .A1(n10507), .A2(n10442), .ZN(n10550) );
  OR2_X1 U13003 ( .A1(n10557), .A2(n10440), .ZN(n10443) );
  NAND2_X1 U13004 ( .A1(n10549), .A2(n10443), .ZN(n10445) );
  NAND2_X1 U13005 ( .A1(n10445), .A2(n10444), .ZN(n10446) );
  XNOR2_X1 U13006 ( .A(n10445), .B(n10586), .ZN(n10580) );
  NAND2_X1 U13007 ( .A1(n10567), .A2(n10566), .ZN(n10565) );
  NAND2_X1 U13008 ( .A1(n10447), .A2(n10565), .ZN(n10449) );
  NAND2_X1 U13009 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  XNOR2_X1 U13010 ( .A(n10449), .B(n10756), .ZN(n10744) );
  NAND2_X1 U13011 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n10744), .ZN(n10743) );
  AOI22_X1 U13012 ( .A1(n10488), .A2(n10414), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10451), .ZN(n10452) );
  OAI21_X1 U13013 ( .B1(n10453), .B2(n10452), .A(n10487), .ZN(n10454) );
  NAND2_X1 U13014 ( .A1(n14809), .A2(n10454), .ZN(n10458) );
  NOR2_X1 U13015 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15130), .ZN(n12217) );
  AOI21_X1 U13016 ( .B1(n14799), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12217), .ZN(
        n10457) );
  OAI211_X1 U13017 ( .C1(n10459), .C2(n14815), .A(n10458), .B(n10457), .ZN(
        n10460) );
  AOI21_X1 U13018 ( .B1(n10488), .B2(n14801), .A(n10460), .ZN(n10461) );
  NAND2_X1 U13019 ( .A1(n10462), .A2(n10461), .ZN(P3_U3188) );
  INV_X1 U13020 ( .A(n10949), .ZN(n10464) );
  AOI21_X1 U13021 ( .B1(n12898), .B2(n10464), .A(n10463), .ZN(n10465) );
  OAI21_X1 U13022 ( .B1(n12908), .B2(n10466), .A(n10465), .ZN(n10472) );
  AOI22_X1 U13023 ( .A1(n12934), .A2(n12975), .B1(n6591), .B2(n10467), .ZN(
        n10469) );
  NOR3_X1 U13024 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n10471) );
  AOI211_X1 U13025 ( .C1(n11810), .C2(n12943), .A(n10472), .B(n10471), .ZN(
        n10473) );
  OAI21_X1 U13026 ( .B1(n10474), .B2(n12928), .A(n10473), .ZN(P2_U3199) );
  INV_X1 U13027 ( .A(n13775), .ZN(n14523) );
  INV_X1 U13028 ( .A(n10475), .ZN(n10498) );
  OAI222_X1 U13029 ( .A1(P1_U3086), .A2(n14523), .B1(n14198), .B2(n10498), 
        .C1(n15099), .C2(n14195), .ZN(P1_U3337) );
  NOR2_X1 U13030 ( .A1(n10488), .A2(n11406), .ZN(n10476) );
  INV_X1 U13031 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11324) );
  NOR2_X1 U13032 ( .A1(n11324), .A2(n10478), .ZN(n11054) );
  AOI21_X1 U13033 ( .B1(n10478), .B2(n11324), .A(n11054), .ZN(n10497) );
  INV_X1 U13034 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10479) );
  MUX2_X1 U13035 ( .A(n11324), .B(n10479), .S(n8117), .Z(n10480) );
  NAND2_X1 U13036 ( .A1(n10480), .A2(n10489), .ZN(n11037) );
  INV_X1 U13037 ( .A(n10480), .ZN(n10481) );
  NAND2_X1 U13038 ( .A1(n10481), .A2(n11046), .ZN(n10482) );
  NAND2_X1 U13039 ( .A1(n11037), .A2(n10482), .ZN(n10483) );
  AOI21_X1 U13040 ( .B1(n10485), .B2(n10484), .A(n10483), .ZN(n11039) );
  AND3_X1 U13041 ( .A1(n10485), .A2(n10484), .A3(n10483), .ZN(n10486) );
  OAI21_X1 U13042 ( .B1(n11039), .B2(n10486), .A(n14810), .ZN(n10496) );
  NAND2_X1 U13043 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10490), .ZN(n11048) );
  OAI21_X1 U13044 ( .B1(n10490), .B2(P3_REG1_REG_7__SCAN_IN), .A(n11048), .ZN(
        n10494) );
  NOR2_X1 U13045 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10491), .ZN(n12066) );
  AOI21_X1 U13046 ( .B1(n14799), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12066), .ZN(
        n10492) );
  OAI21_X1 U13047 ( .B1(n12393), .B2(n11046), .A(n10492), .ZN(n10493) );
  AOI21_X1 U13048 ( .B1(n14809), .B2(n10494), .A(n10493), .ZN(n10495) );
  OAI211_X1 U13049 ( .C1(n10497), .C2(n14815), .A(n10496), .B(n10495), .ZN(
        P3_U3189) );
  INV_X1 U13050 ( .A(n14693), .ZN(n10499) );
  OAI222_X1 U13051 ( .A1(n13377), .A2(n10500), .B1(n10499), .B2(P2_U3088), 
        .C1(n13373), .C2(n10498), .ZN(P2_U3309) );
  XOR2_X1 U13052 ( .A(n10501), .B(n10717), .Z(n10516) );
  NAND2_X1 U13053 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  AOI21_X1 U13054 ( .B1(n10506), .B2(n10505), .A(n14815), .ZN(n10514) );
  INV_X1 U13055 ( .A(n10507), .ZN(n10508) );
  AOI21_X1 U13056 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10512) );
  AOI22_X1 U13057 ( .A1(n14799), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10511) );
  OAI21_X1 U13058 ( .B1(n10512), .B2(n12399), .A(n10511), .ZN(n10513) );
  AOI211_X1 U13059 ( .C1(n14801), .C2(n6824), .A(n10514), .B(n10513), .ZN(
        n10515) );
  OAI21_X1 U13060 ( .B1(n14781), .B2(n10516), .A(n10515), .ZN(P3_U3183) );
  AND2_X1 U13061 ( .A1(n10517), .A2(n14907), .ZN(n14930) );
  XNOR2_X1 U13062 ( .A(n7941), .B(n11294), .ZN(n10520) );
  NAND2_X1 U13063 ( .A1(n10520), .A2(n14920), .ZN(n10523) );
  NOR2_X2 U13064 ( .A1(n10521), .A2(n10529), .ZN(n14892) );
  AOI22_X1 U13065 ( .A1(n14891), .A2(n14889), .B1(n14892), .B2(n12259), .ZN(
        n10522) );
  NAND2_X1 U13066 ( .A1(n10523), .A2(n10522), .ZN(n14929) );
  AOI21_X1 U13067 ( .B1(n14930), .B2(n14908), .A(n14929), .ZN(n10535) );
  XNOR2_X1 U13068 ( .A(n9693), .B(n12804), .ZN(n10526) );
  AND2_X1 U13069 ( .A1(n10524), .A2(n10660), .ZN(n10525) );
  AND2_X1 U13070 ( .A1(n10618), .A2(n12392), .ZN(n10527) );
  NAND2_X1 U13071 ( .A1(n10652), .A2(n10527), .ZN(n10538) );
  MUX2_X1 U13072 ( .A(n10620), .B(n10538), .S(n10529), .Z(n10528) );
  INV_X1 U13073 ( .A(n10528), .ZN(n10624) );
  NAND2_X1 U13074 ( .A1(n10529), .A2(n10538), .ZN(n10530) );
  NAND2_X1 U13075 ( .A1(n12804), .A2(n10530), .ZN(n10531) );
  OAI21_X1 U13076 ( .B1(n12804), .B2(n10624), .A(n10531), .ZN(n10532) );
  INV_X1 U13077 ( .A(n10532), .ZN(n10533) );
  NOR2_X1 U13078 ( .A1(n14954), .A2(n14908), .ZN(n10534) );
  MUX2_X1 U13079 ( .A(n10503), .B(n10535), .S(n14927), .Z(n10542) );
  XNOR2_X1 U13080 ( .A(n10639), .B(n10638), .ZN(n14931) );
  AND2_X1 U13081 ( .A1(n14954), .A2(n10536), .ZN(n10537) );
  NAND2_X1 U13082 ( .A1(n10656), .A2(n10537), .ZN(n10539) );
  NAND2_X1 U13083 ( .A1(n10540), .A2(n12684), .ZN(n14879) );
  NAND2_X1 U13084 ( .A1(n14924), .A2(n14879), .ZN(n14291) );
  NAND2_X1 U13085 ( .A1(n14927), .A2(n14291), .ZN(n12583) );
  AOI22_X1 U13086 ( .A1(n14931), .A2(n14281), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14901), .ZN(n10541) );
  NAND2_X1 U13087 ( .A1(n10542), .A2(n10541), .ZN(P3_U3232) );
  XOR2_X1 U13088 ( .A(n10544), .B(n10543), .Z(n10559) );
  OAI21_X1 U13089 ( .B1(n10547), .B2(n10546), .A(n10545), .ZN(n10548) );
  INV_X1 U13090 ( .A(n10548), .ZN(n10555) );
  OAI21_X1 U13091 ( .B1(n10551), .B2(n10550), .A(n10549), .ZN(n10552) );
  NAND2_X1 U13092 ( .A1(n14809), .A2(n10552), .ZN(n10554) );
  AOI22_X1 U13093 ( .A1(n14799), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10553) );
  OAI211_X1 U13094 ( .C1(n10555), .C2(n14815), .A(n10554), .B(n10553), .ZN(
        n10556) );
  AOI21_X1 U13095 ( .B1(n10557), .B2(n14801), .A(n10556), .ZN(n10558) );
  OAI21_X1 U13096 ( .B1(n10559), .B2(n14781), .A(n10558), .ZN(P3_U3184) );
  XOR2_X1 U13097 ( .A(n10561), .B(n10560), .Z(n10575) );
  AOI21_X1 U13098 ( .B1(n10564), .B2(n10563), .A(n10562), .ZN(n10571) );
  OAI21_X1 U13099 ( .B1(n10567), .B2(n10566), .A(n10565), .ZN(n10568) );
  NAND2_X1 U13100 ( .A1(n14809), .A2(n10568), .ZN(n10570) );
  AND2_X1 U13101 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12177) );
  AOI21_X1 U13102 ( .B1(n14799), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n12177), .ZN(
        n10569) );
  OAI211_X1 U13103 ( .C1(n10571), .C2(n14815), .A(n10570), .B(n10569), .ZN(
        n10572) );
  AOI21_X1 U13104 ( .B1(n10573), .B2(n14801), .A(n10572), .ZN(n10574) );
  OAI21_X1 U13105 ( .B1(n10575), .B2(n14781), .A(n10574), .ZN(P3_U3186) );
  XOR2_X1 U13106 ( .A(n10577), .B(n10576), .Z(n10588) );
  XNOR2_X1 U13107 ( .A(n10578), .B(P3_REG2_REG_3__SCAN_IN), .ZN(n10584) );
  OAI21_X1 U13108 ( .B1(n10580), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10579), .ZN(
        n10581) );
  NAND2_X1 U13109 ( .A1(n14809), .A2(n10581), .ZN(n10583) );
  INV_X1 U13110 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U13111 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14900), .ZN(n10887) );
  AOI21_X1 U13112 ( .B1(n14799), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10887), .ZN(
        n10582) );
  OAI211_X1 U13113 ( .C1(n14815), .C2(n10584), .A(n10583), .B(n10582), .ZN(
        n10585) );
  AOI21_X1 U13114 ( .B1(n10586), .B2(n14801), .A(n10585), .ZN(n10587) );
  OAI21_X1 U13115 ( .B1(n10588), .B2(n14781), .A(n10587), .ZN(P3_U3185) );
  INV_X1 U13116 ( .A(n10589), .ZN(n10591) );
  OAI222_X1 U13117 ( .A1(n10592), .A2(P3_U3151), .B1(n12821), .B2(n10591), 
        .C1(n10590), .C2(n12817), .ZN(P3_U3274) );
  INV_X1 U13118 ( .A(n10593), .ZN(n10601) );
  OAI222_X1 U13119 ( .A1(n13373), .A2(n10601), .B1(P2_U3088), .B2(n11992), 
        .C1(n10594), .C2(n13377), .ZN(P2_U3307) );
  INV_X1 U13120 ( .A(n10595), .ZN(n10598) );
  OAI222_X1 U13121 ( .A1(n13377), .A2(n10596), .B1(n13373), .B2(n10598), .C1(
        P2_U3088), .C2(n13053), .ZN(P2_U3308) );
  OAI222_X1 U13122 ( .A1(n13782), .A2(P1_U3086), .B1(n14198), .B2(n10598), 
        .C1(n10597), .C2(n14195), .ZN(P1_U3336) );
  NAND2_X1 U13123 ( .A1(n12258), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10599) );
  OAI21_X1 U13124 ( .B1(n12473), .B2(n12258), .A(n10599), .ZN(P3_U3520) );
  OAI222_X1 U13125 ( .A1(P1_U3086), .A2(n10602), .B1(n14198), .B2(n10601), 
        .C1(n10600), .C2(n14195), .ZN(P1_U3335) );
  XOR2_X1 U13126 ( .A(n10603), .B(n10604), .Z(n14553) );
  INV_X1 U13127 ( .A(n14553), .ZN(n10616) );
  INV_X1 U13128 ( .A(n13863), .ZN(n13978) );
  XOR2_X1 U13129 ( .A(n10605), .B(n10604), .Z(n14551) );
  INV_X1 U13130 ( .A(n14551), .ZN(n10607) );
  OAI22_X1 U13131 ( .A1(n14260), .A2(n10967), .B1(n15144), .B2(n10969), .ZN(
        n10606) );
  AOI21_X1 U13132 ( .B1(n10607), .B2(n14248), .A(n10606), .ZN(n10615) );
  NAND2_X1 U13133 ( .A1(n10608), .A2(n10693), .ZN(n10609) );
  AND2_X1 U13134 ( .A1(n10790), .A2(n10609), .ZN(n14549) );
  NAND2_X1 U13135 ( .A1(n13625), .A2(n14252), .ZN(n10611) );
  NAND2_X1 U13136 ( .A1(n13623), .A2(n14254), .ZN(n10610) );
  NAND2_X1 U13137 ( .A1(n10611), .A2(n10610), .ZN(n14547) );
  AOI21_X1 U13138 ( .B1(n14549), .B2(n14025), .A(n14547), .ZN(n10613) );
  MUX2_X1 U13139 ( .A(n10613), .B(n10612), .S(n14258), .Z(n10614) );
  OAI211_X1 U13140 ( .C1(n10616), .C2(n13978), .A(n10615), .B(n10614), .ZN(
        P1_U3289) );
  OAI22_X1 U13141 ( .A1(n14954), .A2(n10618), .B1(n10617), .B2(n12685), .ZN(
        n10621) );
  AOI21_X1 U13142 ( .B1(n10621), .B2(n10620), .A(n10619), .ZN(n10623) );
  INV_X1 U13143 ( .A(n12804), .ZN(n10622) );
  MUX2_X1 U13144 ( .A(n10624), .B(n10623), .S(n10622), .Z(n10625) );
  NAND2_X1 U13145 ( .A1(n14993), .A2(n14907), .ZN(n12751) );
  OR3_X1 U13146 ( .A1(n10628), .A2(n14907), .A3(n10627), .ZN(n10630) );
  OR2_X1 U13147 ( .A1(n14918), .A2(n14915), .ZN(n10629) );
  AND2_X1 U13148 ( .A1(n10630), .A2(n10629), .ZN(n11175) );
  MUX2_X1 U13149 ( .A(n11175), .B(n15087), .S(n14990), .Z(n10631) );
  OAI21_X1 U13150 ( .B1(n10668), .B2(n12751), .A(n10631), .ZN(P3_U3459) );
  XOR2_X1 U13151 ( .A(n10633), .B(n10632), .Z(n10637) );
  OAI22_X1 U13152 ( .A1(n12244), .A2(n14916), .B1(n12245), .B2(n11298), .ZN(
        n10635) );
  INV_X1 U13153 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n14911) );
  NOR2_X1 U13154 ( .A1(n10646), .A2(n14911), .ZN(n10634) );
  AOI211_X1 U13155 ( .C1(n12242), .C2(n12257), .A(n10635), .B(n10634), .ZN(
        n10636) );
  OAI21_X1 U13156 ( .B1(n10637), .B2(n12237), .A(n10636), .ZN(P3_U3177) );
  INV_X1 U13157 ( .A(n11294), .ZN(n10643) );
  NOR3_X1 U13158 ( .A1(n10639), .A2(n12045), .A3(n10638), .ZN(n10641) );
  AOI211_X1 U13159 ( .C1(n10643), .C2(n10642), .A(n10641), .B(n10640), .ZN(
        n10650) );
  OAI22_X1 U13160 ( .A1(n12244), .A2(n11299), .B1(n12245), .B2(n10644), .ZN(
        n10648) );
  INV_X1 U13161 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10645) );
  NOR2_X1 U13162 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  AOI211_X1 U13163 ( .C1(n12242), .C2(n12259), .A(n10648), .B(n10647), .ZN(
        n10649) );
  OAI21_X1 U13164 ( .B1(n10650), .B2(n12237), .A(n10649), .ZN(P3_U3162) );
  INV_X1 U13165 ( .A(n10651), .ZN(n10654) );
  OAI22_X1 U13166 ( .A1(n10652), .A2(P3_U3151), .B1(SI_22_), .B2(n12817), .ZN(
        n10653) );
  AOI21_X1 U13167 ( .B1(n10654), .B2(n14227), .A(n10653), .ZN(P3_U3273) );
  INV_X1 U13168 ( .A(n10655), .ZN(n10658) );
  AND2_X1 U13169 ( .A1(n10660), .A2(n10656), .ZN(n10657) );
  NAND2_X1 U13170 ( .A1(n10658), .A2(n10657), .ZN(n10666) );
  NAND2_X1 U13171 ( .A1(n10660), .A2(n10659), .ZN(n10661) );
  AND2_X1 U13172 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  OR2_X1 U13173 ( .A1(n10664), .A2(n10663), .ZN(n10665) );
  NAND2_X1 U13174 ( .A1(n14975), .A2(n14907), .ZN(n12802) );
  INV_X1 U13175 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n15055) );
  MUX2_X1 U13176 ( .A(n11175), .B(n15055), .S(n14973), .Z(n10667) );
  OAI21_X1 U13177 ( .B1(n10668), .B2(n12802), .A(n10667), .ZN(P3_U3390) );
  NOR2_X1 U13178 ( .A1(n14532), .A2(n10669), .ZN(n10670) );
  OR2_X1 U13179 ( .A1(n10671), .A2(n10670), .ZN(n14533) );
  XNOR2_X1 U13180 ( .A(n14533), .B(n13627), .ZN(n10673) );
  MUX2_X1 U13181 ( .A(n10308), .B(n10673), .S(n10672), .Z(n10674) );
  AOI222_X1 U13182 ( .A1(n14554), .A2(n10674), .B1(n13626), .B2(n14254), .C1(
        n13628), .C2(n14252), .ZN(n14534) );
  XNOR2_X1 U13183 ( .A(n10308), .B(n10675), .ZN(n14537) );
  NAND2_X1 U13184 ( .A1(n15149), .A2(n10676), .ZN(n10680) );
  NOR2_X1 U13185 ( .A1(n15144), .A2(n10677), .ZN(n10678) );
  AOI21_X1 U13186 ( .B1(n14258), .B2(P1_REG2_REG_1__SCAN_IN), .A(n10678), .ZN(
        n10679) );
  OAI211_X1 U13187 ( .C1(n15152), .C2(n14533), .A(n10680), .B(n10679), .ZN(
        n10681) );
  AOI21_X1 U13188 ( .B1(n14248), .B2(n14537), .A(n10681), .ZN(n10682) );
  OAI21_X1 U13189 ( .B1(n14258), .B2(n14534), .A(n10682), .ZN(P1_U3292) );
  INV_X1 U13190 ( .A(n10683), .ZN(n10687) );
  INV_X1 U13191 ( .A(n10684), .ZN(n10686) );
  OAI22_X1 U13192 ( .A1(n13535), .A2(n10688), .B1(n8735), .B2(n11278), .ZN(
        n10691) );
  OAI22_X1 U13193 ( .A1(n10688), .A2(n13536), .B1(n10124), .B2(n8735), .ZN(
        n10690) );
  XNOR2_X1 U13194 ( .A(n10690), .B(n13537), .ZN(n10692) );
  XOR2_X1 U13195 ( .A(n10691), .B(n10692), .Z(n13514) );
  NAND2_X1 U13196 ( .A1(n13515), .A2(n13514), .ZN(n13513) );
  NAND2_X1 U13197 ( .A1(n10692), .A2(n10691), .ZN(n10695) );
  AOI22_X1 U13198 ( .A1(n13481), .A2(n10693), .B1(n13485), .B2(n13624), .ZN(
        n10696) );
  OAI22_X1 U13199 ( .A1(n10967), .A2(n10124), .B1(n10712), .B2(n11278), .ZN(
        n10694) );
  XNOR2_X1 U13200 ( .A(n10694), .B(n13395), .ZN(n10973) );
  NAND3_X1 U13201 ( .A1(n13513), .A2(n10696), .A3(n10695), .ZN(n10970) );
  INV_X2 U13202 ( .A(n10124), .ZN(n13491) );
  NAND2_X1 U13203 ( .A1(n14557), .A2(n13491), .ZN(n10698) );
  NAND2_X1 U13204 ( .A1(n10123), .A2(n13623), .ZN(n10697) );
  NAND2_X1 U13205 ( .A1(n10698), .A2(n10697), .ZN(n10699) );
  XNOR2_X1 U13206 ( .A(n10699), .B(n13537), .ZN(n10703) );
  NAND2_X1 U13207 ( .A1(n14557), .A2(n13481), .ZN(n10701) );
  NAND2_X1 U13208 ( .A1(n13485), .A2(n13623), .ZN(n10700) );
  NAND2_X1 U13209 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  NOR2_X1 U13210 ( .A1(n10703), .A2(n10702), .ZN(n10770) );
  INV_X1 U13211 ( .A(n10770), .ZN(n10704) );
  NAND2_X1 U13212 ( .A1(n10703), .A2(n10702), .ZN(n10769) );
  NAND2_X1 U13213 ( .A1(n10704), .A2(n10769), .ZN(n10705) );
  XNOR2_X1 U13214 ( .A(n10771), .B(n10705), .ZN(n10716) );
  AND2_X1 U13215 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  NAND2_X1 U13216 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  NOR2_X1 U13217 ( .A1(n14425), .A2(n10791), .ZN(n10714) );
  NAND2_X1 U13218 ( .A1(n14415), .A2(n13622), .ZN(n10711) );
  NAND2_X1 U13219 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n13671) );
  OAI211_X1 U13220 ( .C1(n10712), .C2(n14394), .A(n10711), .B(n13671), .ZN(
        n10713) );
  AOI211_X1 U13221 ( .C1(n14407), .C2(n14557), .A(n10714), .B(n10713), .ZN(
        n10715) );
  OAI21_X1 U13222 ( .B1(n10716), .B2(n14401), .A(n10715), .ZN(P1_U3227) );
  NAND3_X1 U13223 ( .A1(n14815), .A2(n12399), .A3(n14781), .ZN(n10723) );
  OAI21_X1 U13224 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n10718), .A(n10717), .ZN(
        n10722) );
  INV_X1 U13225 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10720) );
  OAI22_X1 U13226 ( .A1(n14797), .A2(n10720), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10719), .ZN(n10721) );
  AOI21_X1 U13227 ( .B1(n10723), .B2(n10722), .A(n10721), .ZN(n10724) );
  OAI21_X1 U13228 ( .B1(n15037), .B2(n12393), .A(n10724), .ZN(P3_U3182) );
  INV_X1 U13229 ( .A(n13622), .ZN(n10776) );
  INV_X1 U13230 ( .A(n14564), .ZN(n14565) );
  NAND2_X1 U13231 ( .A1(n14566), .A2(n14565), .ZN(n10727) );
  OR2_X1 U13232 ( .A1(n15148), .A2(n13621), .ZN(n10726) );
  NAND2_X1 U13233 ( .A1(n10727), .A2(n10726), .ZN(n10811) );
  XOR2_X1 U13234 ( .A(n10811), .B(n10810), .Z(n14579) );
  OR2_X1 U13235 ( .A1(n14572), .A2(n15148), .ZN(n14573) );
  AOI211_X1 U13236 ( .C1(n11193), .C2(n14573), .A(n14576), .B(n10816), .ZN(
        n14582) );
  AND2_X1 U13237 ( .A1(n10786), .A2(n10776), .ZN(n10728) );
  INV_X1 U13238 ( .A(n15148), .ZN(n14575) );
  XNOR2_X1 U13239 ( .A(n10805), .B(n10810), .ZN(n10730) );
  OAI22_X1 U13240 ( .A1(n11366), .A2(n13951), .B1(n11165), .B2(n13949), .ZN(
        n11195) );
  INV_X1 U13241 ( .A(n11195), .ZN(n10729) );
  OAI21_X1 U13242 ( .B1(n10730), .B2(n14571), .A(n10729), .ZN(n14581) );
  AOI21_X1 U13243 ( .B1(n14582), .B2(n13782), .A(n14581), .ZN(n10731) );
  MUX2_X1 U13244 ( .A(n10732), .B(n10731), .S(n15146), .Z(n10735) );
  INV_X1 U13245 ( .A(n11197), .ZN(n10733) );
  AOI22_X1 U13246 ( .A1(n15149), .A2(n11193), .B1(n10733), .B2(n14040), .ZN(
        n10734) );
  OAI211_X1 U13247 ( .C1(n14065), .C2(n14579), .A(n10735), .B(n10734), .ZN(
        P1_U3285) );
  INV_X1 U13248 ( .A(n10736), .ZN(n10739) );
  OAI222_X1 U13249 ( .A1(n10738), .A2(P1_U3086), .B1(n14198), .B2(n10739), 
        .C1(n10737), .C2(n14195), .ZN(P1_U3334) );
  OAI222_X1 U13250 ( .A1(n13377), .A2(n10740), .B1(n13373), .B2(n10739), .C1(
        P2_U3088), .C2(n12023), .ZN(P2_U3306) );
  AOI21_X1 U13251 ( .B1(n10742), .B2(n14862), .A(n10741), .ZN(n10748) );
  OAI21_X1 U13252 ( .B1(n10744), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10743), .ZN(
        n10745) );
  NAND2_X1 U13253 ( .A1(n14809), .A2(n10745), .ZN(n10747) );
  AND2_X1 U13254 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n12152) );
  AOI21_X1 U13255 ( .B1(n14799), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n12152), .ZN(
        n10746) );
  OAI211_X1 U13256 ( .C1(n10748), .C2(n14815), .A(n10747), .B(n10746), .ZN(
        n10755) );
  NAND2_X1 U13257 ( .A1(n6569), .A2(n6820), .ZN(n10753) );
  OAI21_X1 U13258 ( .B1(n10751), .B2(n10750), .A(n10749), .ZN(n10752) );
  AOI21_X1 U13259 ( .B1(n10753), .B2(n10752), .A(n14781), .ZN(n10754) );
  AOI211_X1 U13260 ( .C1(n14801), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10757) );
  INV_X1 U13261 ( .A(n10757), .ZN(P3_U3187) );
  INV_X1 U13262 ( .A(n14746), .ZN(n10768) );
  INV_X1 U13263 ( .A(n10758), .ZN(n10759) );
  AOI21_X1 U13264 ( .B1(n10984), .B2(n10759), .A(n12928), .ZN(n10762) );
  NOR3_X1 U13265 ( .A1(n12858), .A2(n10831), .A3(n10760), .ZN(n10761) );
  OAI21_X1 U13266 ( .B1(n10762), .B2(n10761), .A(n11119), .ZN(n10767) );
  NAND2_X1 U13267 ( .A1(n12906), .A2(n12973), .ZN(n10764) );
  NAND2_X1 U13268 ( .A1(n6433), .A2(n12971), .ZN(n10763) );
  NAND2_X1 U13269 ( .A1(n10764), .A2(n10763), .ZN(n14745) );
  NAND2_X1 U13270 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U13271 ( .B1(n12940), .B2(n11031), .A(n14631), .ZN(n10765) );
  AOI21_X1 U13272 ( .B1(n12942), .B2(n14745), .A(n10765), .ZN(n10766) );
  OAI211_X1 U13273 ( .C1(n10768), .C2(n12924), .A(n10767), .B(n10766), .ZN(
        P2_U3185) );
  NAND2_X1 U13274 ( .A1(n10786), .A2(n13491), .ZN(n10773) );
  NAND2_X1 U13275 ( .A1(n13481), .A2(n13622), .ZN(n10772) );
  NAND2_X1 U13276 ( .A1(n10773), .A2(n10772), .ZN(n10775) );
  XNOR2_X1 U13277 ( .A(n10775), .B(n10689), .ZN(n10779) );
  NOR2_X1 U13278 ( .A1(n13535), .A2(n10776), .ZN(n10777) );
  AOI21_X1 U13279 ( .B1(n10786), .B2(n13481), .A(n10777), .ZN(n10778) );
  NOR2_X1 U13280 ( .A1(n10779), .A2(n10778), .ZN(n11163) );
  NOR2_X1 U13281 ( .A1(n11163), .A2(n6581), .ZN(n10780) );
  XNOR2_X1 U13282 ( .A(n11164), .B(n10780), .ZN(n10788) );
  OAI21_X1 U13283 ( .B1(n14397), .B2(n11165), .A(n10781), .ZN(n10782) );
  AOI21_X1 U13284 ( .B1(n14417), .B2(n13623), .A(n10782), .ZN(n10783) );
  OAI21_X1 U13285 ( .B1(n10784), .B2(n14425), .A(n10783), .ZN(n10785) );
  AOI21_X1 U13286 ( .B1(n14407), .B2(n10786), .A(n10785), .ZN(n10787) );
  OAI21_X1 U13287 ( .B1(n10788), .B2(n14401), .A(n10787), .ZN(P1_U3239) );
  AOI211_X1 U13288 ( .C1(n14557), .C2(n10790), .A(n14576), .B(n10789), .ZN(
        n14556) );
  INV_X1 U13289 ( .A(n14557), .ZN(n10792) );
  OAI22_X1 U13290 ( .A1(n14260), .A2(n10792), .B1(n15144), .B2(n10791), .ZN(
        n10802) );
  XNOR2_X1 U13291 ( .A(n10793), .B(n10796), .ZN(n10800) );
  OAI21_X1 U13292 ( .B1(n10796), .B2(n10795), .A(n10794), .ZN(n10797) );
  NAND2_X1 U13293 ( .A1(n10797), .A2(n14597), .ZN(n10799) );
  AOI22_X1 U13294 ( .A1(n13624), .A2(n14252), .B1(n14254), .B2(n13622), .ZN(
        n10798) );
  OAI211_X1 U13295 ( .C1(n14571), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n14555) );
  MUX2_X1 U13296 ( .A(n14555), .B(P1_REG2_REG_5__SCAN_IN), .S(n14258), .Z(
        n10801) );
  AOI211_X1 U13297 ( .C1(n14247), .C2(n14556), .A(n10802), .B(n10801), .ZN(
        n10803) );
  INV_X1 U13298 ( .A(n10803), .ZN(P1_U3288) );
  OR2_X1 U13299 ( .A1(n11193), .A2(n11186), .ZN(n10804) );
  INV_X1 U13300 ( .A(n10809), .ZN(n10807) );
  INV_X1 U13301 ( .A(n11108), .ZN(n10808) );
  AOI21_X1 U13302 ( .B1(n11098), .B2(n10809), .A(n10808), .ZN(n10815) );
  AOI22_X1 U13303 ( .A1(n14252), .A2(n13620), .B1(n13618), .B2(n14254), .ZN(
        n11288) );
  OR2_X1 U13304 ( .A1(n11193), .A2(n13620), .ZN(n10812) );
  XNOR2_X1 U13305 ( .A(n11099), .B(n11098), .ZN(n10813) );
  NAND2_X1 U13306 ( .A1(n10813), .A2(n14597), .ZN(n10814) );
  OAI211_X1 U13307 ( .C1(n10815), .C2(n14571), .A(n11288), .B(n10814), .ZN(
        n14585) );
  INV_X1 U13308 ( .A(n14585), .ZN(n10821) );
  INV_X1 U13309 ( .A(n10816), .ZN(n10817) );
  INV_X1 U13310 ( .A(n14587), .ZN(n11293) );
  AOI211_X1 U13311 ( .C1(n14587), .C2(n10817), .A(n14576), .B(n11132), .ZN(
        n14586) );
  NOR2_X1 U13312 ( .A1(n11293), .A2(n14260), .ZN(n10819) );
  OAI22_X1 U13313 ( .A1(n15146), .A2(n9873), .B1(n11287), .B2(n15144), .ZN(
        n10818) );
  AOI211_X1 U13314 ( .C1(n14586), .C2(n14247), .A(n10819), .B(n10818), .ZN(
        n10820) );
  OAI21_X1 U13315 ( .B1(n10821), .B2(n14042), .A(n10820), .ZN(P1_U3284) );
  OR2_X1 U13316 ( .A1(n11819), .A2(n12973), .ZN(n10823) );
  INV_X1 U13317 ( .A(n12972), .ZN(n11120) );
  XNOR2_X1 U13318 ( .A(n14746), .B(n11120), .ZN(n11999) );
  INV_X1 U13319 ( .A(n12971), .ZN(n11016) );
  XNOR2_X1 U13320 ( .A(n14755), .B(n11016), .ZN(n12000) );
  XNOR2_X1 U13321 ( .A(n10849), .B(n12000), .ZN(n10835) );
  INV_X1 U13322 ( .A(n10835), .ZN(n14758) );
  INV_X1 U13323 ( .A(n10824), .ZN(n10825) );
  OR2_X1 U13324 ( .A1(n10826), .A2(n10825), .ZN(n10827) );
  INV_X1 U13325 ( .A(n12028), .ZN(n10828) );
  NAND2_X1 U13326 ( .A1(n10828), .A2(n12027), .ZN(n10872) );
  INV_X1 U13327 ( .A(n10872), .ZN(n14707) );
  NAND2_X1 U13328 ( .A1(n14714), .A2(n14707), .ZN(n11077) );
  NAND2_X1 U13329 ( .A1(n11819), .A2(n10831), .ZN(n10832) );
  AND2_X1 U13330 ( .A1(n14746), .A2(n11120), .ZN(n10833) );
  XNOR2_X1 U13331 ( .A(n10857), .B(n12000), .ZN(n10834) );
  NAND2_X1 U13332 ( .A1(n10834), .A2(n14753), .ZN(n10839) );
  NAND2_X1 U13333 ( .A1(n10835), .A2(n13144), .ZN(n10838) );
  NAND2_X1 U13334 ( .A1(n12906), .A2(n12972), .ZN(n10837) );
  NAND2_X1 U13335 ( .A1(n6433), .A2(n12969), .ZN(n10836) );
  AND2_X1 U13336 ( .A1(n10837), .A2(n10836), .ZN(n11118) );
  NAND3_X1 U13337 ( .A1(n10839), .A2(n10838), .A3(n11118), .ZN(n14760) );
  NAND2_X1 U13338 ( .A1(n14760), .A2(n14714), .ZN(n10848) );
  INV_X1 U13339 ( .A(n10840), .ZN(n10841) );
  OAI22_X1 U13340 ( .A1(n14714), .A2(n10842), .B1(n11113), .B2(n14716), .ZN(
        n10846) );
  NAND2_X1 U13341 ( .A1(n11029), .A2(n14755), .ZN(n10843) );
  NAND2_X1 U13342 ( .A1(n10843), .A2(n13206), .ZN(n10844) );
  OR2_X1 U13343 ( .A1(n10920), .A2(n10844), .ZN(n14757) );
  NOR2_X1 U13344 ( .A1(n14757), .A2(n13197), .ZN(n10845) );
  AOI211_X1 U13345 ( .C1(n13194), .C2(n14755), .A(n10846), .B(n10845), .ZN(
        n10847) );
  OAI211_X1 U13346 ( .C1(n14758), .C2(n11077), .A(n10848), .B(n10847), .ZN(
        P2_U3257) );
  INV_X1 U13347 ( .A(n12000), .ZN(n10856) );
  NAND2_X1 U13348 ( .A1(n14755), .A2(n12971), .ZN(n10850) );
  NAND2_X1 U13349 ( .A1(n6509), .A2(n10850), .ZN(n10914) );
  XNOR2_X1 U13350 ( .A(n11834), .B(n12969), .ZN(n12001) );
  INV_X1 U13351 ( .A(n12001), .ZN(n10913) );
  NAND2_X1 U13352 ( .A1(n10914), .A2(n10913), .ZN(n10916) );
  NAND2_X1 U13353 ( .A1(n11834), .A2(n12969), .ZN(n10851) );
  XNOR2_X1 U13354 ( .A(n11843), .B(n12968), .ZN(n12002) );
  INV_X1 U13355 ( .A(n12002), .ZN(n10863) );
  OR2_X1 U13356 ( .A1(n10852), .A2(n10863), .ZN(n10853) );
  NAND2_X1 U13357 ( .A1(n11000), .A2(n10853), .ZN(n14762) );
  NAND2_X1 U13358 ( .A1(n12906), .A2(n12969), .ZN(n10855) );
  NAND2_X1 U13359 ( .A1(n6433), .A2(n12967), .ZN(n10854) );
  NAND2_X1 U13360 ( .A1(n10855), .A2(n10854), .ZN(n11208) );
  INV_X1 U13361 ( .A(n11208), .ZN(n10866) );
  OR2_X1 U13362 ( .A1(n14755), .A2(n11016), .ZN(n10858) );
  NAND2_X1 U13363 ( .A1(n10859), .A2(n10858), .ZN(n10912) );
  NAND2_X1 U13364 ( .A1(n10912), .A2(n12001), .ZN(n10862) );
  INV_X1 U13365 ( .A(n12969), .ZN(n10860) );
  OR2_X1 U13366 ( .A1(n11834), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U13367 ( .A1(n10862), .A2(n10861), .ZN(n11001) );
  XNOR2_X1 U13368 ( .A(n11001), .B(n10863), .ZN(n10864) );
  NAND2_X1 U13369 ( .A1(n10864), .A2(n14753), .ZN(n10865) );
  OAI211_X1 U13370 ( .C1(n14762), .C2(n10917), .A(n10866), .B(n10865), .ZN(
        n14768) );
  NAND2_X1 U13371 ( .A1(n14768), .A2(n14714), .ZN(n10871) );
  OAI22_X1 U13372 ( .A1(n14714), .A2(n10867), .B1(n11206), .B2(n14716), .ZN(
        n10869) );
  INV_X1 U13373 ( .A(n11834), .ZN(n10925) );
  INV_X1 U13374 ( .A(n11843), .ZN(n14765) );
  OAI211_X1 U13375 ( .C1(n10921), .C2(n14765), .A(n13206), .B(n11007), .ZN(
        n14763) );
  NOR2_X1 U13376 ( .A1(n14763), .A2(n13197), .ZN(n10868) );
  AOI211_X1 U13377 ( .C1(n13194), .C2(n11843), .A(n10869), .B(n10868), .ZN(
        n10870) );
  OAI211_X1 U13378 ( .C1(n14762), .C2(n11077), .A(n10871), .B(n10870), .ZN(
        P2_U3255) );
  NAND2_X1 U13379 ( .A1(n10917), .A2(n10872), .ZN(n10873) );
  OAI22_X1 U13380 ( .A1(n14714), .A2(n10875), .B1(n10874), .B2(n14716), .ZN(
        n10878) );
  NOR2_X1 U13381 ( .A1(n13197), .A2(n10876), .ZN(n10877) );
  AOI211_X1 U13382 ( .C1(n13194), .C2(n11793), .A(n10878), .B(n10877), .ZN(
        n10881) );
  NAND2_X1 U13383 ( .A1(n14714), .A2(n10879), .ZN(n10880) );
  OAI211_X1 U13384 ( .C1(n13248), .C2(n10882), .A(n10881), .B(n10880), .ZN(
        P2_U3263) );
  NAND2_X1 U13385 ( .A1(n10883), .A2(n14227), .ZN(n10885) );
  OAI211_X1 U13386 ( .C1(n10886), .C2(n12817), .A(n10885), .B(n10884), .ZN(
        P3_U3272) );
  AOI21_X1 U13387 ( .B1(n12219), .B2(n11302), .A(n10887), .ZN(n10889) );
  NAND2_X1 U13388 ( .A1(n12242), .A2(n14891), .ZN(n10888) );
  OAI211_X1 U13389 ( .C1(n10890), .C2(n12244), .A(n10889), .B(n10888), .ZN(
        n10895) );
  AOI211_X1 U13390 ( .C1(n10893), .C2(n10892), .A(n12237), .B(n10891), .ZN(
        n10894) );
  AOI211_X1 U13391 ( .C1(n14900), .C2(n12248), .A(n10895), .B(n10894), .ZN(
        n10896) );
  INV_X1 U13392 ( .A(n10896), .ZN(P3_U3158) );
  XNOR2_X1 U13393 ( .A(n10897), .B(n10898), .ZN(n14737) );
  INV_X1 U13394 ( .A(n14737), .ZN(n10911) );
  XNOR2_X1 U13395 ( .A(n10899), .B(n10898), .ZN(n10902) );
  NAND2_X1 U13396 ( .A1(n14737), .A2(n13144), .ZN(n10901) );
  OAI211_X1 U13397 ( .C1(n10902), .C2(n7052), .A(n10901), .B(n10900), .ZN(
        n14743) );
  INV_X1 U13398 ( .A(n14714), .ZN(n10962) );
  MUX2_X1 U13399 ( .A(n14743), .B(P2_REG2_REG_4__SCAN_IN), .S(n10962), .Z(
        n10903) );
  INV_X1 U13400 ( .A(n10903), .ZN(n10910) );
  NAND2_X1 U13401 ( .A1(n10957), .A2(n11806), .ZN(n10904) );
  NAND2_X1 U13402 ( .A1(n10904), .A2(n13206), .ZN(n10905) );
  NOR2_X1 U13403 ( .A1(n10906), .A2(n10905), .ZN(n14738) );
  INV_X1 U13404 ( .A(n11806), .ZN(n14741) );
  OAI22_X1 U13405 ( .A1(n13242), .A2(n14741), .B1(n14716), .B2(n10907), .ZN(
        n10908) );
  AOI21_X1 U13406 ( .B1(n13251), .B2(n14738), .A(n10908), .ZN(n10909) );
  OAI211_X1 U13407 ( .C1(n10911), .C2(n11077), .A(n10910), .B(n10909), .ZN(
        P2_U3261) );
  XNOR2_X1 U13408 ( .A(n10912), .B(n10913), .ZN(n10919) );
  OR2_X1 U13409 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  NAND2_X1 U13410 ( .A1(n10916), .A2(n10915), .ZN(n10994) );
  AOI22_X1 U13411 ( .A1(n12906), .A2(n12971), .B1(n6433), .B2(n12968), .ZN(
        n11012) );
  OAI21_X1 U13412 ( .B1(n10994), .B2(n10917), .A(n11012), .ZN(n10918) );
  AOI21_X1 U13413 ( .B1(n10919), .B2(n14753), .A(n10918), .ZN(n10993) );
  INV_X1 U13414 ( .A(n10920), .ZN(n10922) );
  AOI211_X1 U13415 ( .C1(n11834), .C2(n10922), .A(n13221), .B(n10921), .ZN(
        n10991) );
  INV_X1 U13416 ( .A(n11011), .ZN(n10923) );
  INV_X1 U13417 ( .A(n14716), .ZN(n13239) );
  AOI22_X1 U13418 ( .A1(n10962), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10923), 
        .B2(n13239), .ZN(n10924) );
  OAI21_X1 U13419 ( .B1(n10925), .B2(n13242), .A(n10924), .ZN(n10927) );
  NOR2_X1 U13420 ( .A1(n10994), .A2(n11077), .ZN(n10926) );
  AOI211_X1 U13421 ( .C1(n10991), .C2(n13251), .A(n10927), .B(n10926), .ZN(
        n10928) );
  OAI21_X1 U13422 ( .B1(n13253), .B2(n10993), .A(n10928), .ZN(P2_U3256) );
  NAND2_X1 U13423 ( .A1(n14714), .A2(n14753), .ZN(n13115) );
  MUX2_X1 U13424 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10929), .S(n14714), .Z(
        n10933) );
  OAI22_X1 U13425 ( .A1(n13242), .A2(n10931), .B1(n10930), .B2(n14716), .ZN(
        n10932) );
  AOI211_X1 U13426 ( .C1(n10934), .C2(n13251), .A(n10933), .B(n10932), .ZN(
        n10937) );
  NAND2_X1 U13427 ( .A1(n13183), .A2(n10935), .ZN(n10936) );
  OAI211_X1 U13428 ( .C1(n10938), .C2(n13115), .A(n10937), .B(n10936), .ZN(
        P2_U3264) );
  MUX2_X1 U13429 ( .A(n10940), .B(n10939), .S(n14714), .Z(n10945) );
  OAI22_X1 U13430 ( .A1(n13242), .A2(n10941), .B1(n14716), .B2(n10979), .ZN(
        n10942) );
  AOI21_X1 U13431 ( .B1(n10943), .B2(n13251), .A(n10942), .ZN(n10944) );
  OAI211_X1 U13432 ( .C1(n13248), .C2(n10946), .A(n10945), .B(n10944), .ZN(
        P2_U3259) );
  MUX2_X1 U13433 ( .A(n10948), .B(n10947), .S(n10962), .Z(n10954) );
  OAI22_X1 U13434 ( .A1(n13242), .A2(n10950), .B1(n10949), .B2(n14716), .ZN(
        n10951) );
  AOI21_X1 U13435 ( .B1(n10952), .B2(n13251), .A(n10951), .ZN(n10953) );
  OAI211_X1 U13436 ( .C1(n13248), .C2(n10955), .A(n10954), .B(n10953), .ZN(
        P2_U3260) );
  XNOR2_X1 U13437 ( .A(n10956), .B(n11993), .ZN(n14733) );
  INV_X1 U13438 ( .A(n10957), .ZN(n10958) );
  AOI211_X1 U13439 ( .C1(n14730), .C2(n10959), .A(n13221), .B(n10958), .ZN(
        n14728) );
  AOI22_X1 U13440 ( .A1(n14728), .A2(n13251), .B1(n13194), .B2(n14730), .ZN(
        n10966) );
  XNOR2_X1 U13441 ( .A(n10960), .B(n11993), .ZN(n10961) );
  NAND2_X1 U13442 ( .A1(n10961), .A2(n14753), .ZN(n14731) );
  OAI211_X1 U13443 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n14716), .A(n14731), .B(
        n14727), .ZN(n10963) );
  MUX2_X1 U13444 ( .A(n10963), .B(P2_REG2_REG_3__SCAN_IN), .S(n10962), .Z(
        n10964) );
  INV_X1 U13445 ( .A(n10964), .ZN(n10965) );
  OAI211_X1 U13446 ( .C1(n13248), .C2(n14733), .A(n10966), .B(n10965), .ZN(
        P2_U3262) );
  NOR2_X1 U13447 ( .A1(n10967), .A2(n14592), .ZN(n14546) );
  NAND2_X1 U13448 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U13449 ( .A1(n14379), .A2(n14547), .ZN(n10968) );
  OAI211_X1 U13450 ( .C1(n14425), .C2(n10969), .A(n14495), .B(n10968), .ZN(
        n10977) );
  INV_X1 U13451 ( .A(n10970), .ZN(n10972) );
  NOR2_X1 U13452 ( .A1(n10972), .A2(n10971), .ZN(n10974) );
  XNOR2_X1 U13453 ( .A(n10974), .B(n10973), .ZN(n10975) );
  NOR2_X1 U13454 ( .A1(n10975), .A2(n14401), .ZN(n10976) );
  AOI211_X1 U13455 ( .C1(n14369), .C2(n14546), .A(n10977), .B(n10976), .ZN(
        n10978) );
  INV_X1 U13456 ( .A(n10978), .ZN(P1_U3230) );
  INV_X1 U13457 ( .A(n10979), .ZN(n10981) );
  AOI21_X1 U13458 ( .B1(n12898), .B2(n10981), .A(n10980), .ZN(n10982) );
  OAI21_X1 U13459 ( .B1(n12908), .B2(n10983), .A(n10982), .ZN(n10989) );
  INV_X1 U13460 ( .A(n10984), .ZN(n10985) );
  AOI211_X1 U13461 ( .C1(n10987), .C2(n10986), .A(n12928), .B(n10985), .ZN(
        n10988) );
  AOI211_X1 U13462 ( .C1(n11819), .C2(n12911), .A(n10989), .B(n10988), .ZN(
        n10990) );
  INV_X1 U13463 ( .A(n10990), .ZN(P2_U3211) );
  INV_X1 U13464 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10996) );
  AOI21_X1 U13465 ( .B1(n13261), .B2(n11834), .A(n10991), .ZN(n10992) );
  OAI211_X1 U13466 ( .C1(n14761), .C2(n10994), .A(n10993), .B(n10992), .ZN(
        n10997) );
  NAND2_X1 U13467 ( .A1(n10997), .A2(n14754), .ZN(n10995) );
  OAI21_X1 U13468 ( .B1(n14754), .B2(n10996), .A(n10995), .ZN(P2_U3457) );
  NAND2_X1 U13469 ( .A1(n10997), .A2(n6436), .ZN(n10998) );
  OAI21_X1 U13470 ( .B1(n6436), .B2(n9254), .A(n10998), .ZN(P2_U3508) );
  NAND2_X1 U13471 ( .A1(n11843), .A2(n12968), .ZN(n10999) );
  XNOR2_X1 U13472 ( .A(n11847), .B(n12967), .ZN(n12004) );
  INV_X1 U13473 ( .A(n12004), .ZN(n11003) );
  XNOR2_X1 U13474 ( .A(n11074), .B(n11003), .ZN(n11094) );
  INV_X1 U13475 ( .A(n12968), .ZN(n11002) );
  OAI21_X1 U13476 ( .B1(n7376), .B2(n12004), .A(n11066), .ZN(n11092) );
  INV_X1 U13477 ( .A(n11847), .ZN(n11090) );
  NAND2_X1 U13478 ( .A1(n12906), .A2(n12968), .ZN(n11005) );
  NAND2_X1 U13479 ( .A1(n6433), .A2(n12966), .ZN(n11004) );
  AND2_X1 U13480 ( .A1(n11005), .A2(n11004), .ZN(n11336) );
  OAI21_X1 U13481 ( .B1(n11090), .B2(n14764), .A(n11336), .ZN(n11008) );
  INV_X1 U13482 ( .A(n11078), .ZN(n11006) );
  AOI211_X1 U13483 ( .C1(n11847), .C2(n11007), .A(n13221), .B(n11006), .ZN(
        n11086) );
  AOI211_X1 U13484 ( .C1(n11092), .C2(n14753), .A(n11008), .B(n11086), .ZN(
        n11009) );
  OAI21_X1 U13485 ( .B1(n14749), .B2(n11094), .A(n11009), .ZN(n11023) );
  NAND2_X1 U13486 ( .A1(n11023), .A2(n14754), .ZN(n11010) );
  OAI21_X1 U13487 ( .B1(n14754), .B2(n9291), .A(n11010), .ZN(P2_U3463) );
  NAND2_X1 U13488 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14652) );
  OAI21_X1 U13489 ( .B1(n12940), .B2(n11011), .A(n14652), .ZN(n11014) );
  NOR2_X1 U13490 ( .A1(n12908), .A2(n11012), .ZN(n11013) );
  AOI211_X1 U13491 ( .C1(n11834), .C2(n12943), .A(n11014), .B(n11013), .ZN(
        n11021) );
  INV_X1 U13492 ( .A(n11015), .ZN(n11019) );
  OAI22_X1 U13493 ( .A1(n11017), .A2(n12928), .B1(n11016), .B2(n12858), .ZN(
        n11018) );
  NAND3_X1 U13494 ( .A1(n11129), .A2(n11019), .A3(n11018), .ZN(n11020) );
  OAI211_X1 U13495 ( .C1(n11022), .C2(n12928), .A(n11021), .B(n11020), .ZN(
        P2_U3203) );
  NAND2_X1 U13496 ( .A1(n11023), .A2(n6436), .ZN(n11024) );
  OAI21_X1 U13497 ( .B1(n6436), .B2(n11025), .A(n11024), .ZN(P2_U3510) );
  XOR2_X1 U13498 ( .A(n11026), .B(n11999), .Z(n14750) );
  XOR2_X1 U13499 ( .A(n11999), .B(n11027), .Z(n14752) );
  AOI21_X1 U13500 ( .B1(n11028), .B2(n14746), .A(n13221), .ZN(n11030) );
  NAND2_X1 U13501 ( .A1(n11030), .A2(n11029), .ZN(n14747) );
  NOR2_X1 U13502 ( .A1(n14716), .A2(n11031), .ZN(n11033) );
  MUX2_X1 U13503 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n14745), .S(n14714), .Z(
        n11032) );
  AOI211_X1 U13504 ( .C1(n13194), .C2(n14746), .A(n11033), .B(n11032), .ZN(
        n11034) );
  OAI21_X1 U13505 ( .B1(n13197), .B2(n14747), .A(n11034), .ZN(n11035) );
  AOI21_X1 U13506 ( .B1(n14752), .B2(n13199), .A(n11035), .ZN(n11036) );
  OAI21_X1 U13507 ( .B1(n13248), .B2(n14750), .A(n11036), .ZN(P2_U3258) );
  MUX2_X1 U13508 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n8117), .Z(n11040) );
  INV_X1 U13509 ( .A(n11040), .ZN(n11041) );
  INV_X1 U13510 ( .A(n11037), .ZN(n11038) );
  NOR2_X1 U13511 ( .A1(n11039), .A2(n11038), .ZN(n14780) );
  XNOR2_X1 U13512 ( .A(n11040), .B(n11056), .ZN(n14779) );
  MUX2_X1 U13513 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n8117), .Z(n11043) );
  INV_X1 U13514 ( .A(n11043), .ZN(n11042) );
  NAND2_X1 U13515 ( .A1(n11042), .A2(n11057), .ZN(n11462) );
  INV_X1 U13516 ( .A(n11462), .ZN(n11044) );
  AND2_X1 U13517 ( .A1(n11043), .A2(n11474), .ZN(n11461) );
  NOR2_X1 U13518 ( .A1(n11044), .A2(n11461), .ZN(n11045) );
  XNOR2_X1 U13519 ( .A(n11463), .B(n11045), .ZN(n11064) );
  INV_X1 U13520 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U13521 ( .A1(n14789), .A2(n14986), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n11056), .ZN(n14788) );
  NAND2_X1 U13522 ( .A1(n11047), .A2(n11046), .ZN(n11049) );
  NAND2_X1 U13523 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n11050), .ZN(n11468) );
  OAI21_X1 U13524 ( .B1(n11050), .B2(P3_REG1_REG_9__SCAN_IN), .A(n11468), .ZN(
        n11062) );
  NOR2_X1 U13525 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11051), .ZN(n11550) );
  AOI21_X1 U13526 ( .B1(n14799), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11550), .ZN(
        n11052) );
  OAI21_X1 U13527 ( .B1(n12393), .B2(n11474), .A(n11052), .ZN(n11061) );
  INV_X1 U13528 ( .A(n11053), .ZN(n11055) );
  NOR2_X1 U13529 ( .A1(n11055), .A2(n11054), .ZN(n14785) );
  INV_X1 U13530 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U13531 ( .A1(n14789), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n14848), 
        .B2(n11056), .ZN(n14784) );
  NOR2_X1 U13532 ( .A1(n14785), .A2(n14784), .ZN(n14783) );
  INV_X1 U13533 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14833) );
  AOI21_X1 U13534 ( .B1(n11058), .B2(n14833), .A(n11473), .ZN(n11059) );
  NOR2_X1 U13535 ( .A1(n11059), .A2(n14815), .ZN(n11060) );
  AOI211_X1 U13536 ( .C1(n14809), .C2(n11062), .A(n11061), .B(n11060), .ZN(
        n11063) );
  OAI21_X1 U13537 ( .B1(n11064), .B2(n14781), .A(n11063), .ZN(P3_U3191) );
  INV_X1 U13538 ( .A(n12967), .ZN(n11065) );
  INV_X1 U13539 ( .A(n12966), .ZN(n11147) );
  XNOR2_X1 U13540 ( .A(n14345), .B(n11147), .ZN(n12006) );
  AOI21_X1 U13541 ( .B1(n11067), .B2(n12006), .A(n7052), .ZN(n11072) );
  NAND2_X1 U13542 ( .A1(n12906), .A2(n12967), .ZN(n11071) );
  NAND2_X1 U13543 ( .A1(n6433), .A2(n12965), .ZN(n11070) );
  NAND2_X1 U13544 ( .A1(n11071), .A2(n11070), .ZN(n11511) );
  AOI21_X1 U13545 ( .B1(n11072), .B2(n11149), .A(n11511), .ZN(n11076) );
  OR2_X1 U13546 ( .A1(n11847), .A2(n12967), .ZN(n11073) );
  XNOR2_X1 U13547 ( .A(n11146), .B(n11068), .ZN(n14349) );
  NAND2_X1 U13548 ( .A1(n14349), .A2(n13144), .ZN(n11075) );
  AND2_X1 U13549 ( .A1(n11076), .A2(n11075), .ZN(n14351) );
  INV_X1 U13550 ( .A(n11077), .ZN(n13151) );
  NAND2_X1 U13551 ( .A1(n14345), .A2(n11078), .ZN(n11079) );
  NAND2_X1 U13552 ( .A1(n11079), .A2(n13206), .ZN(n11080) );
  OR2_X1 U13553 ( .A1(n11150), .A2(n11080), .ZN(n14346) );
  OAI22_X1 U13554 ( .A1(n14714), .A2(n11081), .B1(n11513), .B2(n14716), .ZN(
        n11082) );
  AOI21_X1 U13555 ( .B1(n14345), .B2(n13194), .A(n11082), .ZN(n11083) );
  OAI21_X1 U13556 ( .B1(n14346), .B2(n13197), .A(n11083), .ZN(n11084) );
  AOI21_X1 U13557 ( .B1(n14349), .B2(n13151), .A(n11084), .ZN(n11085) );
  OAI21_X1 U13558 ( .B1(n14351), .B2(n13253), .A(n11085), .ZN(P2_U3253) );
  NAND2_X1 U13559 ( .A1(n11086), .A2(n13251), .ZN(n11089) );
  OAI22_X1 U13560 ( .A1(n13253), .A2(n11336), .B1(n11333), .B2(n14716), .ZN(
        n11087) );
  AOI21_X1 U13561 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n13253), .A(n11087), 
        .ZN(n11088) );
  OAI211_X1 U13562 ( .C1(n11090), .C2(n13242), .A(n11089), .B(n11088), .ZN(
        n11091) );
  AOI21_X1 U13563 ( .B1(n13199), .B2(n11092), .A(n11091), .ZN(n11093) );
  OAI21_X1 U13564 ( .B1(n11094), .B2(n13248), .A(n11093), .ZN(P2_U3254) );
  INV_X1 U13565 ( .A(n11095), .ZN(n11096) );
  OAI222_X1 U13566 ( .A1(n13377), .A2(n11097), .B1(n13373), .B2(n11096), .C1(
        P2_U3088), .C2(n12031), .ZN(P2_U3305) );
  INV_X1 U13567 ( .A(n11137), .ZN(n11131) );
  NAND2_X1 U13568 ( .A1(n11130), .A2(n11131), .ZN(n11101) );
  OR2_X1 U13569 ( .A1(n11358), .A2(n13618), .ZN(n11100) );
  XOR2_X1 U13570 ( .A(n11216), .B(n11110), .Z(n14440) );
  INV_X1 U13571 ( .A(n11358), .ZN(n14593) );
  AOI21_X1 U13572 ( .B1(n11134), .B2(n11492), .A(n14576), .ZN(n11102) );
  NAND2_X1 U13573 ( .A1(n11102), .A2(n11211), .ZN(n14439) );
  INV_X1 U13574 ( .A(n14439), .ZN(n11106) );
  AOI22_X1 U13575 ( .A1(n14252), .A2(n13618), .B1(n14253), .B2(n14254), .ZN(
        n14438) );
  OAI22_X1 U13576 ( .A1(n14258), .A2(n14438), .B1(n11502), .B2(n15144), .ZN(
        n11103) );
  AOI21_X1 U13577 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n14042), .A(n11103), 
        .ZN(n11104) );
  OAI21_X1 U13578 ( .B1(n6870), .B2(n14260), .A(n11104), .ZN(n11105) );
  AOI21_X1 U13579 ( .B1(n11106), .B2(n14247), .A(n11105), .ZN(n11112) );
  NAND2_X1 U13580 ( .A1(n14587), .A2(n11366), .ZN(n11107) );
  INV_X1 U13581 ( .A(n13618), .ZN(n11356) );
  OR2_X1 U13582 ( .A1(n11358), .A2(n11356), .ZN(n11109) );
  XNOR2_X1 U13583 ( .A(n11213), .B(n11110), .ZN(n14443) );
  NAND2_X1 U13584 ( .A1(n14443), .A2(n13863), .ZN(n11111) );
  OAI211_X1 U13585 ( .C1(n14440), .C2(n14065), .A(n11112), .B(n11111), .ZN(
        P1_U3282) );
  INV_X1 U13586 ( .A(n11113), .ZN(n11116) );
  INV_X1 U13587 ( .A(n11114), .ZN(n11115) );
  AOI21_X1 U13588 ( .B1(n12898), .B2(n11116), .A(n11115), .ZN(n11117) );
  OAI21_X1 U13589 ( .B1(n12908), .B2(n11118), .A(n11117), .ZN(n11127) );
  INV_X1 U13590 ( .A(n11119), .ZN(n11123) );
  NOR3_X1 U13591 ( .A1(n12858), .A2(n11121), .A3(n11120), .ZN(n11122) );
  AOI21_X1 U13592 ( .B1(n11123), .B2(n6591), .A(n11122), .ZN(n11125) );
  NOR2_X1 U13593 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  AOI211_X1 U13594 ( .C1(n14755), .C2(n12911), .A(n11127), .B(n11126), .ZN(
        n11128) );
  OAI21_X1 U13595 ( .B1(n11129), .B2(n12928), .A(n11128), .ZN(P2_U3193) );
  XNOR2_X1 U13596 ( .A(n11130), .B(n11131), .ZN(n14598) );
  INV_X1 U13597 ( .A(n14598), .ZN(n11144) );
  INV_X1 U13598 ( .A(n11132), .ZN(n11133) );
  AOI21_X1 U13599 ( .B1(n11133), .B2(n11358), .A(n14576), .ZN(n11135) );
  AOI22_X1 U13600 ( .A1(n11135), .A2(n11134), .B1(n14254), .B2(n13617), .ZN(
        n14591) );
  OAI211_X1 U13601 ( .C1(n6577), .C2(n11137), .A(n14554), .B(n11136), .ZN(
        n14594) );
  NAND2_X1 U13602 ( .A1(n13619), .A2(n14252), .ZN(n14590) );
  OAI211_X1 U13603 ( .C1(n11138), .C2(n14591), .A(n14594), .B(n14590), .ZN(
        n11142) );
  INV_X1 U13604 ( .A(n11139), .ZN(n11368) );
  AOI22_X1 U13605 ( .A1(n14042), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11368), 
        .B2(n14040), .ZN(n11140) );
  OAI21_X1 U13606 ( .B1(n14593), .B2(n14260), .A(n11140), .ZN(n11141) );
  AOI21_X1 U13607 ( .B1(n11142), .B2(n15146), .A(n11141), .ZN(n11143) );
  OAI21_X1 U13608 ( .B1(n14065), .B2(n11144), .A(n11143), .ZN(P1_U3283) );
  XOR2_X1 U13609 ( .A(n14339), .B(n12965), .Z(n12007) );
  AND2_X1 U13610 ( .A1(n14345), .A2(n12966), .ZN(n11145) );
  OAI22_X1 U13611 ( .A1(n11146), .A2(n11145), .B1(n14345), .B2(n12966), .ZN(
        n11229) );
  XOR2_X1 U13612 ( .A(n12007), .B(n11229), .Z(n14342) );
  OR2_X1 U13613 ( .A1(n14345), .A2(n11147), .ZN(n11148) );
  XNOR2_X1 U13614 ( .A(n11233), .B(n12007), .ZN(n14344) );
  INV_X1 U13615 ( .A(n14339), .ZN(n11154) );
  NAND2_X1 U13616 ( .A1(n11154), .A2(n11150), .ZN(n11236) );
  OAI211_X1 U13617 ( .C1(n11154), .C2(n11150), .A(n13206), .B(n11236), .ZN(
        n14340) );
  NAND2_X1 U13618 ( .A1(n12906), .A2(n12966), .ZN(n11152) );
  NAND2_X1 U13619 ( .A1(n6433), .A2(n12964), .ZN(n11151) );
  NAND2_X1 U13620 ( .A1(n11152), .A2(n11151), .ZN(n14338) );
  INV_X1 U13621 ( .A(n14338), .ZN(n11153) );
  OAI22_X1 U13622 ( .A1(n13253), .A2(n11153), .B1(n11562), .B2(n14716), .ZN(
        n11156) );
  NOR2_X1 U13623 ( .A1(n11154), .A2(n13242), .ZN(n11155) );
  AOI211_X1 U13624 ( .C1(n13253), .C2(P2_REG2_REG_13__SCAN_IN), .A(n11156), 
        .B(n11155), .ZN(n11157) );
  OAI21_X1 U13625 ( .B1(n13197), .B2(n14340), .A(n11157), .ZN(n11158) );
  AOI21_X1 U13626 ( .B1(n14344), .B2(n13199), .A(n11158), .ZN(n11159) );
  OAI21_X1 U13627 ( .B1(n14342), .B2(n13248), .A(n11159), .ZN(P2_U3252) );
  NAND2_X1 U13628 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13687) );
  NAND2_X1 U13629 ( .A1(n13622), .A2(n14252), .ZN(n11161) );
  NAND2_X1 U13630 ( .A1(n13620), .A2(n14254), .ZN(n11160) );
  NAND2_X1 U13631 ( .A1(n11161), .A2(n11160), .ZN(n14567) );
  NAND2_X1 U13632 ( .A1(n14379), .A2(n14567), .ZN(n11162) );
  OAI211_X1 U13633 ( .C1(n14425), .C2(n15145), .A(n13687), .B(n11162), .ZN(
        n11172) );
  NOR2_X1 U13634 ( .A1(n13535), .A2(n11165), .ZN(n11166) );
  AOI21_X1 U13635 ( .B1(n15148), .B2(n13481), .A(n11166), .ZN(n11180) );
  NAND2_X1 U13636 ( .A1(n15148), .A2(n13491), .ZN(n11168) );
  NAND2_X1 U13637 ( .A1(n13481), .A2(n13621), .ZN(n11167) );
  NAND2_X1 U13638 ( .A1(n11168), .A2(n11167), .ZN(n11169) );
  XNOR2_X1 U13639 ( .A(n11169), .B(n13395), .ZN(n11179) );
  XOR2_X1 U13640 ( .A(n11180), .B(n11179), .Z(n11181) );
  XNOR2_X1 U13641 ( .A(n11182), .B(n11181), .ZN(n11170) );
  NOR2_X1 U13642 ( .A1(n11170), .A2(n14401), .ZN(n11171) );
  AOI211_X1 U13643 ( .C1(n14407), .C2(n15148), .A(n11172), .B(n11171), .ZN(
        n11173) );
  INV_X1 U13644 ( .A(n11173), .ZN(P1_U3213) );
  MUX2_X1 U13645 ( .A(n11175), .B(n11174), .S(n14865), .Z(n11178) );
  AOI22_X1 U13646 ( .A1(n14268), .A2(n9612), .B1(n14901), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U13647 ( .A1(n11178), .A2(n11177), .ZN(P3_U3233) );
  NAND2_X1 U13648 ( .A1(n11193), .A2(n13491), .ZN(n11184) );
  NAND2_X1 U13649 ( .A1(n13481), .A2(n13620), .ZN(n11183) );
  NAND2_X1 U13650 ( .A1(n11184), .A2(n11183), .ZN(n11185) );
  XNOR2_X1 U13651 ( .A(n11185), .B(n10689), .ZN(n11189) );
  NOR2_X1 U13652 ( .A1(n13535), .A2(n11186), .ZN(n11187) );
  AOI21_X1 U13653 ( .B1(n11193), .B2(n13481), .A(n11187), .ZN(n11188) );
  NAND2_X1 U13654 ( .A1(n11189), .A2(n11188), .ZN(n11282) );
  OAI21_X1 U13655 ( .B1(n11189), .B2(n11188), .A(n11282), .ZN(n11191) );
  INV_X1 U13656 ( .A(n11283), .ZN(n11190) );
  AOI21_X1 U13657 ( .B1(n11192), .B2(n11191), .A(n11190), .ZN(n11200) );
  AND2_X1 U13658 ( .A1(n11193), .A2(n14588), .ZN(n14580) );
  AOI21_X1 U13659 ( .B1(n14379), .B2(n11195), .A(n11194), .ZN(n11196) );
  OAI21_X1 U13660 ( .B1(n14425), .B2(n11197), .A(n11196), .ZN(n11198) );
  AOI21_X1 U13661 ( .B1(n14580), .B2(n14369), .A(n11198), .ZN(n11199) );
  OAI21_X1 U13662 ( .B1(n11200), .B2(n14401), .A(n11199), .ZN(P1_U3221) );
  AOI21_X1 U13663 ( .B1(n11202), .B2(n11201), .A(n12928), .ZN(n11204) );
  NAND2_X1 U13664 ( .A1(n11204), .A2(n11203), .ZN(n11210) );
  OAI21_X1 U13665 ( .B1(n12940), .B2(n11206), .A(n11205), .ZN(n11207) );
  AOI21_X1 U13666 ( .B1(n12942), .B2(n11208), .A(n11207), .ZN(n11209) );
  OAI211_X1 U13667 ( .C1(n14765), .C2(n12924), .A(n11210), .B(n11209), .ZN(
        P2_U3189) );
  NOR2_X2 U13668 ( .A1(n14238), .A2(n11211), .ZN(n14245) );
  AOI211_X1 U13669 ( .C1(n14238), .C2(n11211), .A(n14576), .B(n14245), .ZN(
        n14239) );
  INV_X1 U13670 ( .A(n14239), .ZN(n11227) );
  NAND2_X1 U13671 ( .A1(n11492), .A2(n11490), .ZN(n11212) );
  OR2_X1 U13672 ( .A1(n11492), .A2(n11490), .ZN(n11214) );
  NAND2_X1 U13673 ( .A1(n11215), .A2(n11214), .ZN(n11411) );
  XNOR2_X1 U13674 ( .A(n11411), .B(n11410), .ZN(n11222) );
  INV_X1 U13675 ( .A(n11410), .ZN(n11217) );
  OAI21_X1 U13676 ( .B1(n6576), .B2(n11217), .A(n11417), .ZN(n11220) );
  NAND2_X1 U13677 ( .A1(n13617), .A2(n14252), .ZN(n11219) );
  NAND2_X1 U13678 ( .A1(n14361), .A2(n14254), .ZN(n11218) );
  NAND2_X1 U13679 ( .A1(n11219), .A2(n11218), .ZN(n14378) );
  AOI21_X1 U13680 ( .B1(n11220), .B2(n14597), .A(n14378), .ZN(n11221) );
  OAI21_X1 U13681 ( .B1(n14571), .B2(n11222), .A(n11221), .ZN(n14240) );
  NAND2_X1 U13682 ( .A1(n14240), .A2(n15146), .ZN(n11226) );
  OAI22_X1 U13683 ( .A1(n15146), .A2(n11223), .B1(n14382), .B2(n15144), .ZN(
        n11224) );
  AOI21_X1 U13684 ( .B1(n14238), .B2(n15149), .A(n11224), .ZN(n11225) );
  OAI211_X1 U13685 ( .C1(n13998), .C2(n11227), .A(n11226), .B(n11225), .ZN(
        P1_U3281) );
  XNOR2_X1 U13686 ( .A(n11867), .B(n12964), .ZN(n12010) );
  NOR2_X1 U13687 ( .A1(n14339), .A2(n12965), .ZN(n11228) );
  NAND2_X1 U13688 ( .A1(n14339), .A2(n12965), .ZN(n11230) );
  XOR2_X1 U13689 ( .A(n12010), .B(n11381), .Z(n11375) );
  INV_X1 U13690 ( .A(n12965), .ZN(n11234) );
  NOR2_X1 U13691 ( .A1(n14339), .A2(n11234), .ZN(n11232) );
  NAND2_X1 U13692 ( .A1(n14339), .A2(n11234), .ZN(n11235) );
  XNOR2_X1 U13693 ( .A(n11396), .B(n12010), .ZN(n11372) );
  INV_X1 U13694 ( .A(n11867), .ZN(n11244) );
  AOI21_X1 U13695 ( .B1(n11867), .B2(n11236), .A(n13221), .ZN(n11237) );
  AND2_X1 U13696 ( .A1(n11237), .A2(n11389), .ZN(n11371) );
  NAND2_X1 U13697 ( .A1(n11371), .A2(n13251), .ZN(n11243) );
  NAND2_X1 U13698 ( .A1(n12963), .A2(n6433), .ZN(n11239) );
  NAND2_X1 U13699 ( .A1(n12906), .A2(n12965), .ZN(n11238) );
  NAND2_X1 U13700 ( .A1(n11239), .A2(n11238), .ZN(n11664) );
  INV_X1 U13701 ( .A(n11664), .ZN(n11240) );
  OAI22_X1 U13702 ( .A1(n13253), .A2(n11240), .B1(n11662), .B2(n14716), .ZN(
        n11241) );
  AOI21_X1 U13703 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n13253), .A(n11241), 
        .ZN(n11242) );
  OAI211_X1 U13704 ( .C1(n11244), .C2(n13242), .A(n11243), .B(n11242), .ZN(
        n11245) );
  AOI21_X1 U13705 ( .B1(n11372), .B2(n13199), .A(n11245), .ZN(n11246) );
  OAI21_X1 U13706 ( .B1(n11375), .B2(n13248), .A(n11246), .ZN(P2_U3251) );
  INV_X1 U13707 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11251) );
  MUX2_X1 U13708 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11251), .S(n13756), .Z(
        n13758) );
  INV_X1 U13709 ( .A(n11247), .ZN(n11248) );
  AOI21_X1 U13710 ( .B1(n11249), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11248), 
        .ZN(n11250) );
  XNOR2_X1 U13711 ( .A(n11250), .B(n14510), .ZN(n14507) );
  NOR2_X1 U13712 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14507), .ZN(n14506) );
  AOI21_X1 U13713 ( .B1(n11250), .B2(n14510), .A(n14506), .ZN(n13759) );
  NAND2_X1 U13714 ( .A1(n13758), .A2(n13759), .ZN(n13757) );
  OAI21_X1 U13715 ( .B1(n11252), .B2(n11251), .A(n13757), .ZN(n11256) );
  INV_X1 U13716 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11253) );
  MUX2_X1 U13717 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n11253), .S(n11254), .Z(
        n11255) );
  NAND2_X1 U13718 ( .A1(n11254), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13773) );
  OAI211_X1 U13719 ( .C1(n11254), .C2(P1_REG2_REG_17__SCAN_IN), .A(n11256), 
        .B(n13773), .ZN(n13772) );
  OAI211_X1 U13720 ( .C1(n11256), .C2(n11255), .A(n14492), .B(n13772), .ZN(
        n11267) );
  NAND2_X1 U13721 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13569)
         );
  XOR2_X1 U13722 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n13756), .Z(n13753) );
  AOI21_X1 U13723 ( .B1(n15088), .B2(n11258), .A(n11257), .ZN(n11260) );
  INV_X1 U13724 ( .A(n11260), .ZN(n11261) );
  XNOR2_X1 U13725 ( .A(n11260), .B(n11259), .ZN(n14505) );
  NOR2_X1 U13726 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14505), .ZN(n14504) );
  AOI21_X1 U13727 ( .B1(n11261), .B2(n14510), .A(n14504), .ZN(n13754) );
  NAND2_X1 U13728 ( .A1(n13753), .A2(n13754), .ZN(n13752) );
  INV_X1 U13729 ( .A(n13752), .ZN(n11262) );
  AOI21_X1 U13730 ( .B1(n13756), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11262), 
        .ZN(n13766) );
  XNOR2_X1 U13731 ( .A(n13764), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13763) );
  XNOR2_X1 U13732 ( .A(n13766), .B(n13763), .ZN(n11263) );
  NAND2_X1 U13733 ( .A1(n14486), .A2(n11263), .ZN(n11264) );
  NAND2_X1 U13734 ( .A1(n13569), .A2(n11264), .ZN(n11265) );
  AOI21_X1 U13735 ( .B1(n14497), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11265), 
        .ZN(n11266) );
  OAI211_X1 U13736 ( .C1(n14524), .C2(n13764), .A(n11267), .B(n11266), .ZN(
        P1_U3260) );
  INV_X1 U13737 ( .A(n11268), .ZN(n11270) );
  OAI222_X1 U13738 ( .A1(P3_U3151), .A2(n9602), .B1(n12821), .B2(n11270), .C1(
        n11269), .C2(n12817), .ZN(P3_U3271) );
  NAND2_X1 U13739 ( .A1(n11274), .A2(n13366), .ZN(n11272) );
  OR2_X1 U13740 ( .A1(n11271), .A2(P2_U3088), .ZN(n12043) );
  OAI211_X1 U13741 ( .C1(n11273), .C2(n13377), .A(n11272), .B(n12043), .ZN(
        P2_U3304) );
  NAND2_X1 U13742 ( .A1(n11274), .A2(n14184), .ZN(n11276) );
  OAI211_X1 U13743 ( .C1(n11277), .C2(n14195), .A(n11276), .B(n11275), .ZN(
        P1_U3332) );
  OAI22_X1 U13744 ( .A1(n11293), .A2(n11278), .B1(n11366), .B2(n13535), .ZN(
        n11350) );
  NAND2_X1 U13745 ( .A1(n14587), .A2(n13491), .ZN(n11280) );
  NAND2_X1 U13746 ( .A1(n13481), .A2(n13619), .ZN(n11279) );
  NAND2_X1 U13747 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  XNOR2_X1 U13748 ( .A(n11281), .B(n13537), .ZN(n11349) );
  XOR2_X1 U13749 ( .A(n11350), .B(n11349), .Z(n11285) );
  NAND2_X1 U13750 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  OAI21_X1 U13751 ( .B1(n11285), .B2(n11284), .A(n11361), .ZN(n11286) );
  NAND2_X1 U13752 ( .A1(n11286), .A2(n14421), .ZN(n11292) );
  INV_X1 U13753 ( .A(n11287), .ZN(n11290) );
  INV_X1 U13754 ( .A(n14425), .ZN(n13602) );
  INV_X1 U13755 ( .A(n14379), .ZN(n13604) );
  NAND2_X1 U13756 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13711) );
  OAI21_X1 U13757 ( .B1(n13604), .B2(n11288), .A(n13711), .ZN(n11289) );
  AOI21_X1 U13758 ( .B1(n11290), .B2(n13602), .A(n11289), .ZN(n11291) );
  OAI211_X1 U13759 ( .C1(n11293), .C2(n14419), .A(n11292), .B(n11291), .ZN(
        P1_U3231) );
  NAND2_X1 U13760 ( .A1(n11295), .A2(n11294), .ZN(n11297) );
  NAND2_X1 U13761 ( .A1(n14918), .A2(n10644), .ZN(n11296) );
  NAND2_X1 U13762 ( .A1(n11297), .A2(n11296), .ZN(n14912) );
  NAND2_X1 U13763 ( .A1(n14912), .A2(n14914), .ZN(n14913) );
  NAND2_X1 U13764 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  AND2_X1 U13765 ( .A1(n14913), .A2(n11300), .ZN(n14895) );
  NAND2_X1 U13766 ( .A1(n14895), .A2(n11301), .ZN(n14894) );
  NAND2_X1 U13767 ( .A1(n9611), .A2(n11302), .ZN(n11303) );
  NAND2_X1 U13768 ( .A1(n14894), .A2(n11303), .ZN(n14866) );
  NAND2_X1 U13769 ( .A1(n14866), .A2(n14867), .ZN(n11305) );
  NAND2_X1 U13770 ( .A1(n14890), .A2(n14864), .ZN(n11304) );
  NAND2_X1 U13771 ( .A1(n11305), .A2(n11304), .ZN(n14851) );
  INV_X1 U13772 ( .A(n14851), .ZN(n11307) );
  INV_X1 U13773 ( .A(n14859), .ZN(n11308) );
  NAND2_X1 U13774 ( .A1(n14873), .A2(n11308), .ZN(n11309) );
  NAND2_X1 U13775 ( .A1(n14855), .A2(n12218), .ZN(n11311) );
  XNOR2_X1 U13776 ( .A(n11312), .B(n11644), .ZN(n11318) );
  XNOR2_X1 U13777 ( .A(n11314), .B(n11313), .ZN(n11319) );
  INV_X1 U13778 ( .A(n14924), .ZN(n14875) );
  OAI22_X1 U13779 ( .A1(n11315), .A2(n14917), .B1(n11647), .B2(n14915), .ZN(
        n11316) );
  AOI21_X1 U13780 ( .B1(n11319), .B2(n14875), .A(n11316), .ZN(n11317) );
  OAI21_X1 U13781 ( .B1(n11318), .B2(n14877), .A(n11317), .ZN(n14958) );
  INV_X1 U13782 ( .A(n11319), .ZN(n14956) );
  INV_X1 U13783 ( .A(n12068), .ZN(n11320) );
  OAI22_X1 U13784 ( .A1(n14956), .A2(n14879), .B1(n11320), .B2(n14910), .ZN(
        n11321) );
  OAI21_X1 U13785 ( .B1(n14958), .B2(n11321), .A(n14927), .ZN(n11323) );
  NAND2_X1 U13786 ( .A1(n14268), .A2(n12067), .ZN(n11322) );
  OAI211_X1 U13787 ( .C1(n11324), .C2(n14927), .A(n11323), .B(n11322), .ZN(
        P3_U3226) );
  INV_X1 U13788 ( .A(n11325), .ZN(n11326) );
  OAI222_X1 U13789 ( .A1(n11328), .A2(P3_U3151), .B1(n12817), .B2(n11327), 
        .C1(n12821), .C2(n11326), .ZN(P3_U3270) );
  NAND2_X1 U13790 ( .A1(n11330), .A2(n11329), .ZN(n11332) );
  XOR2_X1 U13791 ( .A(n11332), .B(n11331), .Z(n11339) );
  INV_X1 U13792 ( .A(n11333), .ZN(n11334) );
  AOI22_X1 U13793 ( .A1(n12898), .A2(n11334), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11335) );
  OAI21_X1 U13794 ( .B1(n12908), .B2(n11336), .A(n11335), .ZN(n11337) );
  AOI21_X1 U13795 ( .B1(n11847), .B2(n12911), .A(n11337), .ZN(n11338) );
  OAI21_X1 U13796 ( .B1(n11339), .B2(n12928), .A(n11338), .ZN(P2_U3208) );
  INV_X1 U13797 ( .A(n14846), .ZN(n11348) );
  INV_X1 U13798 ( .A(n12248), .ZN(n11347) );
  OAI211_X1 U13799 ( .C1(n11342), .C2(n11341), .A(n11340), .B(n12229), .ZN(
        n11346) );
  NAND2_X1 U13800 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n14795) );
  INV_X1 U13801 ( .A(n14795), .ZN(n11344) );
  INV_X1 U13802 ( .A(n12242), .ZN(n12210) );
  OAI22_X1 U13803 ( .A1(n12210), .A2(n14840), .B1(n14839), .B2(n12244), .ZN(
        n11343) );
  AOI211_X1 U13804 ( .C1(n12219), .C2(n14845), .A(n11344), .B(n11343), .ZN(
        n11345) );
  OAI211_X1 U13805 ( .C1(n11348), .C2(n11347), .A(n11346), .B(n11345), .ZN(
        P3_U3161) );
  INV_X1 U13806 ( .A(n11349), .ZN(n11352) );
  INV_X1 U13807 ( .A(n11350), .ZN(n11351) );
  NAND2_X1 U13808 ( .A1(n11352), .A2(n11351), .ZN(n11359) );
  AND2_X1 U13809 ( .A1(n11361), .A2(n11359), .ZN(n11363) );
  NAND2_X1 U13810 ( .A1(n11358), .A2(n13491), .ZN(n11354) );
  NAND2_X1 U13811 ( .A1(n13481), .A2(n13618), .ZN(n11353) );
  NAND2_X1 U13812 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  XNOR2_X1 U13813 ( .A(n11355), .B(n13395), .ZN(n11495) );
  NOR2_X1 U13814 ( .A1(n13535), .A2(n11356), .ZN(n11357) );
  AOI21_X1 U13815 ( .B1(n11358), .B2(n13481), .A(n11357), .ZN(n11493) );
  XNOR2_X1 U13816 ( .A(n11495), .B(n11493), .ZN(n11362) );
  OAI211_X1 U13817 ( .C1(n11363), .C2(n11362), .A(n14421), .B(n11499), .ZN(
        n11370) );
  AOI21_X1 U13818 ( .B1(n14415), .B2(n13617), .A(n11364), .ZN(n11365) );
  OAI21_X1 U13819 ( .B1(n11366), .B2(n14394), .A(n11365), .ZN(n11367) );
  AOI21_X1 U13820 ( .B1(n11368), .B2(n13602), .A(n11367), .ZN(n11369) );
  OAI211_X1 U13821 ( .C1(n14593), .C2(n14419), .A(n11370), .B(n11369), .ZN(
        P1_U3217) );
  INV_X1 U13822 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11377) );
  AOI211_X1 U13823 ( .C1(n13261), .C2(n11867), .A(n11664), .B(n11371), .ZN(
        n11374) );
  NAND2_X1 U13824 ( .A1(n11372), .A2(n14753), .ZN(n11373) );
  OAI211_X1 U13825 ( .C1(n11375), .C2(n14749), .A(n11374), .B(n11373), .ZN(
        n11378) );
  NAND2_X1 U13826 ( .A1(n11378), .A2(n14754), .ZN(n11376) );
  OAI21_X1 U13827 ( .B1(n14754), .B2(n11377), .A(n11376), .ZN(P2_U3472) );
  NAND2_X1 U13828 ( .A1(n11378), .A2(n6436), .ZN(n11379) );
  OAI21_X1 U13829 ( .B1(n6436), .B2(n11450), .A(n11379), .ZN(P2_U3513) );
  INV_X1 U13830 ( .A(n12963), .ZN(n11569) );
  XNOR2_X1 U13831 ( .A(n14332), .B(n11569), .ZN(n12013) );
  AND2_X1 U13832 ( .A1(n11867), .A2(n12964), .ZN(n11380) );
  OR2_X1 U13833 ( .A1(n11867), .A2(n12964), .ZN(n11382) );
  XOR2_X1 U13834 ( .A(n12013), .B(n11578), .Z(n14335) );
  INV_X1 U13835 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U13836 ( .A1(n12962), .A2(n6433), .ZN(n11384) );
  NAND2_X1 U13837 ( .A1(n12906), .A2(n12964), .ZN(n11383) );
  NAND2_X1 U13838 ( .A1(n11384), .A2(n11383), .ZN(n14331) );
  AOI22_X1 U13839 ( .A1(n14714), .A2(n14331), .B1(n12938), .B2(n13239), .ZN(
        n11385) );
  OAI21_X1 U13840 ( .B1(n11386), .B2(n14714), .A(n11385), .ZN(n11392) );
  NAND2_X1 U13841 ( .A1(n14332), .A2(n11389), .ZN(n11390) );
  NAND3_X1 U13842 ( .A1(n11572), .A2(n13206), .A3(n11390), .ZN(n14333) );
  NOR2_X1 U13843 ( .A1(n14333), .A2(n13197), .ZN(n11391) );
  AOI211_X1 U13844 ( .C1(n13194), .C2(n14332), .A(n11392), .B(n11391), .ZN(
        n11398) );
  INV_X1 U13845 ( .A(n12964), .ZN(n11393) );
  AND2_X1 U13846 ( .A1(n11867), .A2(n11393), .ZN(n11395) );
  OR2_X1 U13847 ( .A1(n11867), .A2(n11393), .ZN(n11394) );
  XNOR2_X1 U13848 ( .A(n11568), .B(n12013), .ZN(n14337) );
  NAND2_X1 U13849 ( .A1(n14337), .A2(n13199), .ZN(n11397) );
  OAI211_X1 U13850 ( .C1(n14335), .C2(n13248), .A(n11398), .B(n11397), .ZN(
        P2_U3250) );
  NAND2_X1 U13851 ( .A1(n12218), .A2(n14907), .ZN(n14948) );
  INV_X1 U13852 ( .A(n14879), .ZN(n14926) );
  OAI21_X1 U13853 ( .B1(n11400), .B2(n11401), .A(n11399), .ZN(n14951) );
  INV_X1 U13854 ( .A(n14951), .ZN(n11405) );
  AOI22_X1 U13855 ( .A1(n12254), .A2(n14889), .B1(n14892), .B2(n12255), .ZN(
        n11404) );
  OAI211_X1 U13856 ( .C1(n6578), .C2(n11310), .A(n14920), .B(n11402), .ZN(
        n11403) );
  OAI211_X1 U13857 ( .C1(n11405), .C2(n14924), .A(n11404), .B(n11403), .ZN(
        n14949) );
  AOI21_X1 U13858 ( .B1(n14926), .B2(n14951), .A(n14949), .ZN(n11407) );
  MUX2_X1 U13859 ( .A(n11407), .B(n11406), .S(n14865), .Z(n11409) );
  NAND2_X1 U13860 ( .A1(n14901), .A2(n12221), .ZN(n11408) );
  OAI211_X1 U13861 ( .C1(n12466), .C2(n14948), .A(n11409), .B(n11408), .ZN(
        P3_U3227) );
  NAND2_X1 U13862 ( .A1(n11411), .A2(n11410), .ZN(n11413) );
  INV_X1 U13863 ( .A(n14253), .ZN(n14395) );
  OR2_X1 U13864 ( .A1(n14238), .A2(n14395), .ZN(n11412) );
  NAND2_X1 U13865 ( .A1(n11413), .A2(n11412), .ZN(n14250) );
  NAND2_X1 U13866 ( .A1(n14250), .A2(n11418), .ZN(n11415) );
  OR2_X1 U13867 ( .A1(n14406), .A2(n13397), .ZN(n11414) );
  NAND2_X1 U13868 ( .A1(n11415), .A2(n11414), .ZN(n11597) );
  XNOR2_X1 U13869 ( .A(n11597), .B(n11419), .ZN(n14432) );
  NAND2_X1 U13870 ( .A1(n11417), .A2(n11416), .ZN(n14243) );
  AOI21_X1 U13871 ( .B1(n14243), .B2(n14249), .A(n6492), .ZN(n11420) );
  OAI21_X1 U13872 ( .B1(n11420), .B2(n11419), .A(n11608), .ZN(n14430) );
  NOR2_X1 U13873 ( .A1(n14430), .A2(n14065), .ZN(n11428) );
  AOI211_X1 U13874 ( .C1(n14428), .C2(n14244), .A(n14576), .B(n11615), .ZN(
        n14426) );
  NAND2_X1 U13875 ( .A1(n14386), .A2(n14254), .ZN(n11422) );
  NAND2_X1 U13876 ( .A1(n14361), .A2(n14252), .ZN(n11421) );
  NAND2_X1 U13877 ( .A1(n11422), .A2(n11421), .ZN(n14427) );
  AOI21_X1 U13878 ( .B1(n14426), .B2(n13782), .A(n14427), .ZN(n11426) );
  AOI22_X1 U13879 ( .A1(n14042), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11423), 
        .B2(n14040), .ZN(n11425) );
  NAND2_X1 U13880 ( .A1(n14428), .A2(n15149), .ZN(n11424) );
  OAI211_X1 U13881 ( .C1(n11426), .C2(n14042), .A(n11425), .B(n11424), .ZN(
        n11427) );
  AOI211_X1 U13882 ( .C1(n13863), .C2(n14432), .A(n11428), .B(n11427), .ZN(
        n11429) );
  INV_X1 U13883 ( .A(n11429), .ZN(P1_U3279) );
  INV_X1 U13884 ( .A(n11430), .ZN(n11432) );
  OAI222_X1 U13885 ( .A1(P3_U3151), .A2(n11433), .B1(n12821), .B2(n11432), 
        .C1(n11431), .C2(n12817), .ZN(P3_U3269) );
  NOR2_X1 U13886 ( .A1(n11446), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n13019) );
  MUX2_X1 U13887 ( .A(n11081), .B(P2_REG2_REG_12__SCAN_IN), .S(n11447), .Z(
        n13020) );
  OAI21_X1 U13888 ( .B1(n13026), .B2(P2_REG2_REG_12__SCAN_IN), .A(n13018), 
        .ZN(n14664) );
  INV_X1 U13889 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11434) );
  MUX2_X1 U13890 ( .A(n11434), .B(P2_REG2_REG_13__SCAN_IN), .S(n11448), .Z(
        n14665) );
  NOR2_X1 U13891 ( .A1(n14664), .A2(n14665), .ZN(n14663) );
  AOI21_X1 U13892 ( .B1(n11448), .B2(P2_REG2_REG_13__SCAN_IN), .A(n14663), 
        .ZN(n11435) );
  OR2_X1 U13893 ( .A1(n11435), .A2(n11451), .ZN(n11436) );
  XNOR2_X1 U13894 ( .A(n11435), .B(n14672), .ZN(n14671) );
  NAND2_X1 U13895 ( .A1(n14671), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U13896 ( .A1(n11436), .A2(n14670), .ZN(n11437) );
  NAND2_X1 U13897 ( .A1(n14681), .A2(n11437), .ZN(n11438) );
  XNOR2_X1 U13898 ( .A(n11452), .B(n11437), .ZN(n14684) );
  NAND2_X1 U13899 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14684), .ZN(n14682) );
  NAND2_X1 U13900 ( .A1(n11444), .A2(n11439), .ZN(n11440) );
  OAI21_X1 U13901 ( .B1(n11444), .B2(n11439), .A(n11440), .ZN(n11441) );
  OAI211_X1 U13902 ( .C1(n11442), .C2(n11441), .A(n11584), .B(n14683), .ZN(
        n11460) );
  NAND2_X1 U13903 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n11695)
         );
  NOR2_X1 U13904 ( .A1(n11444), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11443) );
  AOI21_X1 U13905 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n11444), .A(n11443), 
        .ZN(n11456) );
  INV_X1 U13906 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14352) );
  AOI21_X1 U13907 ( .B1(n11446), .B2(P2_REG1_REG_11__SCAN_IN), .A(n11445), 
        .ZN(n13028) );
  MUX2_X1 U13908 ( .A(n14352), .B(P2_REG1_REG_12__SCAN_IN), .S(n11447), .Z(
        n13027) );
  AOI21_X1 U13909 ( .B1(n14352), .B2(n11447), .A(n13029), .ZN(n14662) );
  MUX2_X1 U13910 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11449), .S(n11448), .Z(
        n14661) );
  NAND2_X1 U13911 ( .A1(n14662), .A2(n14661), .ZN(n14660) );
  OAI21_X1 U13912 ( .B1(n11449), .B2(n14657), .A(n14660), .ZN(n14675) );
  MUX2_X1 U13913 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n11450), .S(n14672), .Z(
        n14674) );
  NAND2_X1 U13914 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  OAI21_X1 U13915 ( .B1(n11450), .B2(n11451), .A(n14673), .ZN(n11453) );
  NAND2_X1 U13916 ( .A1(n14681), .A2(n11453), .ZN(n11454) );
  XNOR2_X1 U13917 ( .A(n11453), .B(n11452), .ZN(n14686) );
  NAND2_X1 U13918 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14686), .ZN(n14685) );
  NAND2_X1 U13919 ( .A1(n11454), .A2(n14685), .ZN(n11455) );
  NAND2_X1 U13920 ( .A1(n11455), .A2(n11456), .ZN(n11587) );
  OAI211_X1 U13921 ( .C1(n11456), .C2(n11455), .A(n14696), .B(n11587), .ZN(
        n11457) );
  NAND2_X1 U13922 ( .A1(n11695), .A2(n11457), .ZN(n11458) );
  AOI21_X1 U13923 ( .B1(n14680), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11458), 
        .ZN(n11459) );
  OAI211_X1 U13924 ( .C1(n14658), .C2(n11588), .A(n11460), .B(n11459), .ZN(
        P2_U3230) );
  MUX2_X1 U13925 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n8117), .Z(n11464) );
  XNOR2_X1 U13926 ( .A(n11464), .B(n14800), .ZN(n14803) );
  OAI21_X1 U13927 ( .B1(n11464), .B2(n11475), .A(n14802), .ZN(n11466) );
  MUX2_X1 U13928 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n8117), .Z(n11537) );
  XNOR2_X1 U13929 ( .A(n11537), .B(n11526), .ZN(n11465) );
  NAND2_X1 U13930 ( .A1(n11466), .A2(n11465), .ZN(n11535) );
  OAI21_X1 U13931 ( .B1(n11466), .B2(n11465), .A(n11535), .ZN(n11485) );
  INV_X1 U13932 ( .A(n11526), .ZN(n11536) );
  NAND2_X1 U13933 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11475), .ZN(n11470) );
  INV_X1 U13934 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U13935 ( .A1(n14800), .A2(n14991), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11475), .ZN(n14807) );
  NAND2_X1 U13936 ( .A1(n11467), .A2(n11474), .ZN(n11469) );
  NAND2_X1 U13937 ( .A1(n11469), .A2(n11468), .ZN(n14806) );
  NAND2_X1 U13938 ( .A1(n14807), .A2(n14806), .ZN(n14805) );
  NAND2_X1 U13939 ( .A1(n11470), .A2(n14805), .ZN(n11524) );
  XNOR2_X1 U13940 ( .A(n11524), .B(n11526), .ZN(n11471) );
  NAND2_X1 U13941 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11471), .ZN(n11525) );
  OAI21_X1 U13942 ( .B1(n11471), .B2(P3_REG1_REG_11__SCAN_IN), .A(n11525), 
        .ZN(n11472) );
  NAND2_X1 U13943 ( .A1(n11472), .A2(n14809), .ZN(n11483) );
  AND2_X1 U13944 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12200) );
  NAND2_X1 U13945 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11475), .ZN(n11477) );
  OAI21_X1 U13946 ( .B1(n11475), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11477), 
        .ZN(n14813) );
  NOR2_X1 U13947 ( .A1(n14814), .A2(n14813), .ZN(n14812) );
  INV_X1 U13948 ( .A(n14812), .ZN(n11476) );
  NAND2_X1 U13949 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  INV_X1 U13950 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14295) );
  AOI21_X1 U13951 ( .B1(n11479), .B2(n14295), .A(n11521), .ZN(n11480) );
  NOR2_X1 U13952 ( .A1(n14815), .A2(n11480), .ZN(n11481) );
  AOI211_X1 U13953 ( .C1(n14799), .C2(P3_ADDR_REG_11__SCAN_IN), .A(n12200), 
        .B(n11481), .ZN(n11482) );
  OAI211_X1 U13954 ( .C1(n12393), .C2(n11536), .A(n11483), .B(n11482), .ZN(
        n11484) );
  AOI21_X1 U13955 ( .B1(n11485), .B2(n14810), .A(n11484), .ZN(n11486) );
  INV_X1 U13956 ( .A(n11486), .ZN(P3_U3193) );
  NAND2_X1 U13957 ( .A1(n11492), .A2(n13491), .ZN(n11488) );
  NAND2_X1 U13958 ( .A1(n10123), .A2(n13617), .ZN(n11487) );
  NAND2_X1 U13959 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  XNOR2_X1 U13960 ( .A(n11489), .B(n13395), .ZN(n13386) );
  NOR2_X1 U13961 ( .A1(n13535), .A2(n11490), .ZN(n11491) );
  AOI21_X1 U13962 ( .B1(n11492), .B2(n13481), .A(n11491), .ZN(n13384) );
  XNOR2_X1 U13963 ( .A(n13386), .B(n13384), .ZN(n11497) );
  INV_X1 U13964 ( .A(n11493), .ZN(n11494) );
  NAND2_X1 U13965 ( .A1(n11495), .A2(n11494), .ZN(n11498) );
  INV_X1 U13966 ( .A(n13387), .ZN(n11501) );
  AOI21_X1 U13967 ( .B1(n11499), .B2(n11498), .A(n11497), .ZN(n11500) );
  OAI21_X1 U13968 ( .B1(n11501), .B2(n11500), .A(n14421), .ZN(n11506) );
  INV_X1 U13969 ( .A(n11502), .ZN(n11504) );
  NAND2_X1 U13970 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13728)
         );
  OAI21_X1 U13971 ( .B1(n13604), .B2(n14438), .A(n13728), .ZN(n11503) );
  AOI21_X1 U13972 ( .B1(n11504), .B2(n13602), .A(n11503), .ZN(n11505) );
  OAI211_X1 U13973 ( .C1(n6870), .C2(n14419), .A(n11506), .B(n11505), .ZN(
        P1_U3236) );
  INV_X1 U13974 ( .A(n11507), .ZN(n11508) );
  AOI21_X1 U13975 ( .B1(n11510), .B2(n11509), .A(n11508), .ZN(n11516) );
  NAND2_X1 U13976 ( .A1(n12942), .A2(n11511), .ZN(n11512) );
  NAND2_X1 U13977 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n13024)
         );
  OAI211_X1 U13978 ( .C1(n12940), .C2(n11513), .A(n11512), .B(n13024), .ZN(
        n11514) );
  AOI21_X1 U13979 ( .B1(n14345), .B2(n12911), .A(n11514), .ZN(n11515) );
  OAI21_X1 U13980 ( .B1(n11516), .B2(n12928), .A(n11515), .ZN(P2_U3196) );
  INV_X1 U13981 ( .A(n11517), .ZN(n11519) );
  OAI222_X1 U13982 ( .A1(n8117), .A2(P3_U3151), .B1(n12821), .B2(n11519), .C1(
        n11518), .C2(n12817), .ZN(P3_U3268) );
  INV_X1 U13983 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U13984 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12267), .B1(n12263), 
        .B2(n15066), .ZN(n11523) );
  AOI21_X1 U13985 ( .B1(n6575), .B2(n11523), .A(n12260), .ZN(n11544) );
  INV_X1 U13986 ( .A(n11524), .ZN(n11527) );
  INV_X1 U13987 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11528) );
  MUX2_X1 U13988 ( .A(n11528), .B(P3_REG1_REG_12__SCAN_IN), .S(n12267), .Z(
        n11529) );
  OAI21_X1 U13989 ( .B1(n11530), .B2(n11529), .A(n12266), .ZN(n11542) );
  INV_X1 U13990 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U13991 ( .A1(n14801), .A2(n12267), .ZN(n11533) );
  INV_X1 U13992 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11531) );
  NOR2_X1 U13993 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11531), .ZN(n12122) );
  INV_X1 U13994 ( .A(n12122), .ZN(n11532) );
  OAI211_X1 U13995 ( .C1(n11534), .C2(n14797), .A(n11533), .B(n11532), .ZN(
        n11541) );
  MUX2_X1 U13996 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n8117), .Z(n12264) );
  XNOR2_X1 U13997 ( .A(n12264), .B(n12263), .ZN(n11539) );
  OAI21_X1 U13998 ( .B1(n11537), .B2(n11536), .A(n11535), .ZN(n11538) );
  AOI211_X1 U13999 ( .C1(n11539), .C2(n11538), .A(n14781), .B(n12262), .ZN(
        n11540) );
  AOI211_X1 U14000 ( .C1(n14809), .C2(n11542), .A(n11541), .B(n11540), .ZN(
        n11543) );
  OAI21_X1 U14001 ( .B1(n11544), .B2(n14815), .A(n11543), .ZN(P3_U3194) );
  INV_X1 U14002 ( .A(n11545), .ZN(n11546) );
  AOI21_X1 U14003 ( .B1(n11548), .B2(n11547), .A(n11546), .ZN(n11553) );
  OAI22_X1 U14004 ( .A1(n12210), .A2(n11647), .B1(n14290), .B2(n12244), .ZN(
        n11549) );
  AOI211_X1 U14005 ( .C1(n12219), .C2(n14830), .A(n11550), .B(n11549), .ZN(
        n11552) );
  NAND2_X1 U14006 ( .A1(n12248), .A2(n14831), .ZN(n11551) );
  OAI211_X1 U14007 ( .C1(n11553), .C2(n12237), .A(n11552), .B(n11551), .ZN(
        P3_U3171) );
  INV_X1 U14008 ( .A(n11554), .ZN(n11558) );
  OAI222_X1 U14009 ( .A1(n11556), .A2(P1_U3086), .B1(n14198), .B2(n11558), 
        .C1(n11555), .C2(n14195), .ZN(P1_U3331) );
  OAI222_X1 U14010 ( .A1(n13377), .A2(n11559), .B1(n13373), .B2(n11558), .C1(
        P2_U3088), .C2(n11557), .ZN(P2_U3303) );
  XNOR2_X1 U14011 ( .A(n11561), .B(n11560), .ZN(n11566) );
  NOR2_X1 U14012 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9332), .ZN(n14655) );
  NOR2_X1 U14013 ( .A1(n12940), .A2(n11562), .ZN(n11563) );
  AOI211_X1 U14014 ( .C1(n12942), .C2(n14338), .A(n14655), .B(n11563), .ZN(
        n11565) );
  NAND2_X1 U14015 ( .A1(n14339), .A2(n12911), .ZN(n11564) );
  OAI211_X1 U14016 ( .C1(n11566), .C2(n12928), .A(n11565), .B(n11564), .ZN(
        P2_U3206) );
  NOR2_X1 U14017 ( .A1(n14332), .A2(n11569), .ZN(n11567) );
  NAND2_X1 U14018 ( .A1(n14332), .A2(n11569), .ZN(n11570) );
  XNOR2_X1 U14019 ( .A(n14321), .B(n12962), .ZN(n12008) );
  OAI21_X1 U14020 ( .B1(n6565), .B2(n12008), .A(n11635), .ZN(n11571) );
  INV_X1 U14021 ( .A(n11571), .ZN(n14329) );
  AOI21_X1 U14022 ( .B1(n11572), .B2(n14321), .A(n13221), .ZN(n11573) );
  NAND2_X1 U14023 ( .A1(n11573), .A2(n11636), .ZN(n14323) );
  NOR2_X1 U14024 ( .A1(n14714), .A2(n11439), .ZN(n11576) );
  AND2_X1 U14025 ( .A1(n12963), .A2(n12906), .ZN(n11574) );
  AOI21_X1 U14026 ( .B1(n12961), .B2(n6433), .A(n11574), .ZN(n14322) );
  OAI22_X1 U14027 ( .A1(n13253), .A2(n14322), .B1(n11696), .B2(n14716), .ZN(
        n11575) );
  AOI211_X1 U14028 ( .C1(n14321), .C2(n13194), .A(n11576), .B(n11575), .ZN(
        n11577) );
  OAI21_X1 U14029 ( .B1(n14323), .B2(n13197), .A(n11577), .ZN(n11581) );
  NOR2_X1 U14030 ( .A1(n11579), .A2(n6923), .ZN(n14326) );
  NAND2_X1 U14031 ( .A1(n11579), .A2(n6923), .ZN(n11632) );
  INV_X1 U14032 ( .A(n11632), .ZN(n14325) );
  NOR3_X1 U14033 ( .A1(n14326), .A2(n14325), .A3(n13248), .ZN(n11580) );
  AOI211_X1 U14034 ( .C1(n14329), .C2(n13199), .A(n11581), .B(n11580), .ZN(
        n11582) );
  INV_X1 U14035 ( .A(n11582), .ZN(P2_U3249) );
  OR2_X1 U14036 ( .A1(n11589), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U14037 ( .A1(n11589), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U14038 ( .A1(n11583), .A2(n13038), .ZN(n13034) );
  XOR2_X1 U14039 ( .A(n13034), .B(n13036), .Z(n11594) );
  INV_X1 U14040 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14041 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12872)
         );
  OAI21_X1 U14042 ( .B1(n14705), .B2(n11585), .A(n12872), .ZN(n11586) );
  AOI21_X1 U14043 ( .B1(n11589), .B2(n14694), .A(n11586), .ZN(n11593) );
  INV_X1 U14044 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14330) );
  OAI21_X1 U14045 ( .B1(n14330), .B2(n11588), .A(n11587), .ZN(n11591) );
  INV_X1 U14046 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U14047 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n11589), .B1(n13044), 
        .B2(n13043), .ZN(n11590) );
  NAND2_X1 U14048 ( .A1(n11590), .A2(n11591), .ZN(n13042) );
  OAI211_X1 U14049 ( .C1(n11591), .C2(n11590), .A(n13042), .B(n14696), .ZN(
        n11592) );
  OAI211_X1 U14050 ( .C1(n11594), .C2(n14700), .A(n11593), .B(n11592), .ZN(
        P2_U3231) );
  NAND2_X1 U14051 ( .A1(n11626), .A2(n11625), .ZN(n11624) );
  NAND2_X1 U14052 ( .A1(n11624), .A2(n11598), .ZN(n11601) );
  INV_X1 U14053 ( .A(n11601), .ZN(n11600) );
  INV_X1 U14054 ( .A(n11612), .ZN(n11599) );
  NAND2_X1 U14055 ( .A1(n11601), .A2(n11612), .ZN(n11602) );
  NAND2_X1 U14056 ( .A1(n13822), .A2(n11602), .ZN(n11606) );
  NAND2_X1 U14057 ( .A1(n14385), .A2(n14254), .ZN(n11603) );
  OAI21_X1 U14058 ( .B1(n11604), .B2(n13949), .A(n11603), .ZN(n11605) );
  AOI21_X1 U14059 ( .B1(n11606), .B2(n14554), .A(n11605), .ZN(n14154) );
  NAND2_X1 U14060 ( .A1(n14428), .A2(n14416), .ZN(n11607) );
  INV_X1 U14061 ( .A(n11625), .ZN(n11609) );
  OR2_X1 U14062 ( .A1(n13412), .A2(n14386), .ZN(n11610) );
  NAND2_X1 U14063 ( .A1(n11611), .A2(n11610), .ZN(n11613) );
  NAND2_X1 U14064 ( .A1(n11613), .A2(n11612), .ZN(n13801) );
  OAI21_X1 U14065 ( .B1(n11613), .B2(n11612), .A(n13801), .ZN(n14152) );
  AOI21_X1 U14066 ( .B1(n11616), .B2(n14149), .A(n14576), .ZN(n11617) );
  NAND2_X1 U14067 ( .A1(n11617), .A2(n14054), .ZN(n14150) );
  OAI22_X1 U14068 ( .A1(n15146), .A2(n11251), .B1(n14393), .B2(n15144), .ZN(
        n11618) );
  AOI21_X1 U14069 ( .B1(n14149), .B2(n15149), .A(n11618), .ZN(n11619) );
  OAI21_X1 U14070 ( .B1(n14150), .B2(n13998), .A(n11619), .ZN(n11620) );
  AOI21_X1 U14071 ( .B1(n14152), .B2(n14248), .A(n11620), .ZN(n11621) );
  OAI21_X1 U14072 ( .B1(n14154), .B2(n14042), .A(n11621), .ZN(P1_U3277) );
  XOR2_X1 U14073 ( .A(n11622), .B(n11625), .Z(n14161) );
  XNOR2_X1 U14074 ( .A(n11614), .B(n6865), .ZN(n14159) );
  NAND2_X1 U14075 ( .A1(n14159), .A2(n14025), .ZN(n11623) );
  AOI22_X1 U14076 ( .A1(n14414), .A2(n14254), .B1(n14252), .B2(n14416), .ZN(
        n14155) );
  OAI211_X1 U14077 ( .C1(n15144), .C2(n14424), .A(n11623), .B(n14155), .ZN(
        n11629) );
  OAI21_X1 U14078 ( .B1(n11626), .B2(n11625), .A(n11624), .ZN(n14156) );
  AOI22_X1 U14079 ( .A1(n13412), .A2(n15149), .B1(n14258), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n11627) );
  OAI21_X1 U14080 ( .B1(n14156), .B2(n13978), .A(n11627), .ZN(n11628) );
  AOI21_X1 U14081 ( .B1(n15146), .B2(n11629), .A(n11628), .ZN(n11630) );
  OAI21_X1 U14082 ( .B1(n14065), .B2(n14161), .A(n11630), .ZN(P1_U3278) );
  NAND2_X1 U14083 ( .A1(n14321), .A2(n12962), .ZN(n11631) );
  NAND2_X1 U14084 ( .A1(n11632), .A2(n11631), .ZN(n11745) );
  XNOR2_X1 U14085 ( .A(n12876), .B(n12961), .ZN(n12011) );
  XNOR2_X1 U14086 ( .A(n11745), .B(n11744), .ZN(n13340) );
  INV_X1 U14087 ( .A(n12962), .ZN(n11633) );
  OR2_X1 U14088 ( .A1(n14321), .A2(n11633), .ZN(n11634) );
  XNOR2_X1 U14089 ( .A(n11706), .B(n11744), .ZN(n13338) );
  INV_X1 U14090 ( .A(n12876), .ZN(n13335) );
  AOI211_X1 U14091 ( .C1(n12876), .C2(n11636), .A(n13221), .B(n13235), .ZN(
        n13336) );
  NAND2_X1 U14092 ( .A1(n13336), .A2(n13251), .ZN(n11640) );
  AND2_X1 U14093 ( .A1(n12962), .A2(n12906), .ZN(n11637) );
  AOI21_X1 U14094 ( .B1(n12960), .B2(n6433), .A(n11637), .ZN(n13334) );
  OAI22_X1 U14095 ( .A1(n13253), .A2(n13334), .B1(n12873), .B2(n14716), .ZN(
        n11638) );
  AOI21_X1 U14096 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n10962), .A(n11638), 
        .ZN(n11639) );
  OAI211_X1 U14097 ( .C1(n13335), .C2(n13242), .A(n11640), .B(n11639), .ZN(
        n11641) );
  AOI21_X1 U14098 ( .B1(n13199), .B2(n13338), .A(n11641), .ZN(n11642) );
  OAI21_X1 U14099 ( .B1(n13340), .B2(n13248), .A(n11642), .ZN(P2_U3248) );
  AND2_X1 U14100 ( .A1(n12254), .A2(n12067), .ZN(n11643) );
  NAND2_X1 U14101 ( .A1(n14838), .A2(n14837), .ZN(n14836) );
  NAND2_X1 U14102 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  NAND2_X1 U14103 ( .A1(n12253), .A2(n14830), .ZN(n11650) );
  XNOR2_X1 U14104 ( .A(n11670), .B(n11669), .ZN(n11651) );
  OAI222_X1 U14105 ( .A1(n14917), .A2(n14839), .B1(n14915), .B2(n11672), .C1(
        n11651), .C2(n14877), .ZN(n14969) );
  INV_X1 U14106 ( .A(n14969), .ZN(n11657) );
  XNOR2_X1 U14107 ( .A(n11652), .B(n11669), .ZN(n14971) );
  INV_X1 U14108 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11654) );
  NOR2_X1 U14109 ( .A1(n12090), .A2(n14954), .ZN(n14970) );
  AOI22_X1 U14110 ( .A1(n14902), .A2(n14970), .B1(n14901), .B2(n12097), .ZN(
        n11653) );
  OAI21_X1 U14111 ( .B1(n11654), .B2(n14927), .A(n11653), .ZN(n11655) );
  AOI21_X1 U14112 ( .B1(n14971), .B2(n14281), .A(n11655), .ZN(n11656) );
  OAI21_X1 U14113 ( .B1(n11657), .B2(n14865), .A(n11656), .ZN(P3_U3223) );
  AOI21_X1 U14114 ( .B1(n11660), .B2(n11659), .A(n11658), .ZN(n11667) );
  OAI22_X1 U14115 ( .A1(n12940), .A2(n11662), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11661), .ZN(n11663) );
  AOI21_X1 U14116 ( .B1(n12942), .B2(n11664), .A(n11663), .ZN(n11666) );
  NAND2_X1 U14117 ( .A1(n11867), .A2(n12911), .ZN(n11665) );
  OAI211_X1 U14118 ( .C1(n11667), .C2(n12928), .A(n11666), .B(n11665), .ZN(
        P2_U3187) );
  XNOR2_X1 U14119 ( .A(n11668), .B(n11674), .ZN(n14306) );
  INV_X1 U14120 ( .A(n14286), .ZN(n11673) );
  INV_X1 U14121 ( .A(n12201), .ZN(n14292) );
  NAND2_X1 U14122 ( .A1(n11675), .A2(n11674), .ZN(n12412) );
  OAI211_X1 U14123 ( .C1(n11675), .C2(n11674), .A(n12412), .B(n14920), .ZN(
        n11677) );
  AOI22_X1 U14124 ( .A1(n14889), .A2(n12668), .B1(n12252), .B2(n14892), .ZN(
        n11676) );
  NAND2_X1 U14125 ( .A1(n11677), .A2(n11676), .ZN(n14308) );
  NAND2_X1 U14126 ( .A1(n14308), .A2(n14927), .ZN(n11681) );
  NAND2_X1 U14127 ( .A1(n12410), .A2(n14907), .ZN(n14304) );
  INV_X1 U14128 ( .A(n12123), .ZN(n11678) );
  OAI22_X1 U14129 ( .A1(n12466), .A2(n14304), .B1(n11678), .B2(n14910), .ZN(
        n11679) );
  AOI21_X1 U14130 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n14865), .A(n11679), 
        .ZN(n11680) );
  OAI211_X1 U14131 ( .C1(n14306), .C2(n12583), .A(n11681), .B(n11680), .ZN(
        P3_U3221) );
  XNOR2_X1 U14132 ( .A(n11682), .B(n12668), .ZN(n11683) );
  XNOR2_X1 U14133 ( .A(n11684), .B(n11683), .ZN(n11691) );
  INV_X1 U14134 ( .A(n12413), .ZN(n14280) );
  NOR2_X1 U14135 ( .A1(n12245), .A2(n14280), .ZN(n11688) );
  NAND2_X1 U14136 ( .A1(n12242), .A2(n14272), .ZN(n11686) );
  AND2_X1 U14137 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12270) );
  INV_X1 U14138 ( .A(n12270), .ZN(n11685) );
  OAI211_X1 U14139 ( .C1(n12652), .C2(n12244), .A(n11686), .B(n11685), .ZN(
        n11687) );
  AOI211_X1 U14140 ( .C1(n11689), .C2(n12248), .A(n11688), .B(n11687), .ZN(
        n11690) );
  OAI21_X1 U14141 ( .B1(n11691), .B2(n12237), .A(n11690), .ZN(P3_U3174) );
  AOI21_X1 U14142 ( .B1(n11694), .B2(n11693), .A(n11692), .ZN(n11700) );
  NOR2_X1 U14143 ( .A1(n12908), .A2(n14322), .ZN(n11698) );
  OAI21_X1 U14144 ( .B1(n12940), .B2(n11696), .A(n11695), .ZN(n11697) );
  AOI211_X1 U14145 ( .C1(n14321), .C2(n12943), .A(n11698), .B(n11697), .ZN(
        n11699) );
  OAI21_X1 U14146 ( .B1(n11700), .B2(n12928), .A(n11699), .ZN(P2_U3198) );
  INV_X1 U14147 ( .A(n13367), .ZN(n11702) );
  OAI222_X1 U14148 ( .A1(n8937), .A2(P1_U3086), .B1(n14198), .B2(n11702), .C1(
        n11701), .C2(n14195), .ZN(P1_U3327) );
  NAND2_X1 U14149 ( .A1(n13367), .A2(n11959), .ZN(n11704) );
  AND2_X2 U14150 ( .A1(n11704), .A2(n11703), .ZN(n13077) );
  INV_X2 U14151 ( .A(n13077), .ZN(n13266) );
  INV_X1 U14152 ( .A(n12961), .ZN(n11707) );
  NAND2_X1 U14153 ( .A1(n12876), .A2(n11707), .ZN(n11705) );
  OR2_X1 U14154 ( .A1(n12876), .A2(n11707), .ZN(n11708) );
  NAND2_X1 U14155 ( .A1(n11709), .A2(n11708), .ZN(n13231) );
  INV_X1 U14156 ( .A(n12960), .ZN(n11747) );
  NOR2_X1 U14157 ( .A1(n13330), .A2(n11747), .ZN(n11711) );
  NAND2_X1 U14158 ( .A1(n13330), .A2(n11747), .ZN(n11710) );
  INV_X1 U14159 ( .A(n12959), .ZN(n11712) );
  AND2_X1 U14160 ( .A1(n13326), .A2(n11712), .ZN(n11713) );
  INV_X1 U14161 ( .A(n12958), .ZN(n11714) );
  NAND2_X1 U14162 ( .A1(n13321), .A2(n11714), .ZN(n11716) );
  OR2_X1 U14163 ( .A1(n13321), .A2(n11714), .ZN(n11715) );
  NAND2_X1 U14164 ( .A1(n11716), .A2(n11715), .ZN(n13203) );
  INV_X1 U14165 ( .A(n12957), .ZN(n11717) );
  OR2_X1 U14166 ( .A1(n13195), .A2(n11717), .ZN(n11718) );
  XNOR2_X1 U14167 ( .A(n13307), .B(n12956), .ZN(n13173) );
  NAND2_X1 U14168 ( .A1(n13169), .A2(n13173), .ZN(n13168) );
  OR2_X1 U14169 ( .A1(n11719), .A2(n13307), .ZN(n11720) );
  NAND2_X1 U14170 ( .A1(n13168), .A2(n11720), .ZN(n13156) );
  INV_X1 U14171 ( .A(n12955), .ZN(n12882) );
  NAND2_X1 U14172 ( .A1(n13159), .A2(n12882), .ZN(n11721) );
  OR2_X1 U14173 ( .A1(n13159), .A2(n12882), .ZN(n11722) );
  INV_X1 U14174 ( .A(n12954), .ZN(n12859) );
  NAND2_X1 U14175 ( .A1(n13296), .A2(n12859), .ZN(n11725) );
  OR2_X1 U14176 ( .A1(n13296), .A2(n12859), .ZN(n11723) );
  NAND2_X1 U14177 ( .A1(n11725), .A2(n11723), .ZN(n13139) );
  XNOR2_X1 U14178 ( .A(n13131), .B(n12918), .ZN(n13122) );
  INV_X1 U14179 ( .A(n13122), .ZN(n13117) );
  NAND2_X1 U14180 ( .A1(n13118), .A2(n13117), .ZN(n13116) );
  INV_X1 U14181 ( .A(n12918), .ZN(n12953) );
  NAND2_X1 U14182 ( .A1(n13102), .A2(n11726), .ZN(n11727) );
  NAND2_X1 U14183 ( .A1(n13266), .A2(n12950), .ZN(n11760) );
  OR2_X1 U14184 ( .A1(n13266), .A2(n12950), .ZN(n11728) );
  NAND2_X1 U14185 ( .A1(n11760), .A2(n11728), .ZN(n13070) );
  NAND2_X1 U14186 ( .A1(n13071), .A2(n13070), .ZN(n13069) );
  OAI21_X1 U14187 ( .B1(n11933), .B2(n13266), .A(n13069), .ZN(n11736) );
  NAND2_X1 U14188 ( .A1(n9198), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11735) );
  INV_X1 U14189 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11765) );
  OR2_X1 U14190 ( .A1(n11730), .A2(n11765), .ZN(n11734) );
  OR2_X1 U14191 ( .A1(n11731), .A2(n11764), .ZN(n11733) );
  INV_X1 U14192 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15051) );
  OR2_X1 U14193 ( .A1(n11966), .A2(n15051), .ZN(n11732) );
  AND4_X1 U14194 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11951) );
  NAND2_X1 U14195 ( .A1(n12950), .A2(n12906), .ZN(n11743) );
  AOI21_X1 U14196 ( .B1(n11737), .B2(P2_B_REG_SCAN_IN), .A(n15177), .ZN(n13058) );
  INV_X1 U14197 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U14198 ( .A1(n11962), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11739) );
  NAND2_X1 U14199 ( .A1(n9530), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11738) );
  OAI211_X1 U14200 ( .C1(n11741), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        n12948) );
  NAND2_X1 U14201 ( .A1(n13058), .A2(n12948), .ZN(n11742) );
  NAND2_X1 U14202 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  NAND2_X1 U14203 ( .A1(n12876), .A2(n12961), .ZN(n11879) );
  XNOR2_X1 U14204 ( .A(n13330), .B(n11747), .ZN(n13230) );
  INV_X1 U14205 ( .A(n13230), .ZN(n13247) );
  OR2_X1 U14206 ( .A1(n13330), .A2(n12960), .ZN(n11748) );
  NAND2_X1 U14207 ( .A1(n13326), .A2(n12959), .ZN(n11749) );
  AND2_X1 U14208 ( .A1(n13321), .A2(n12958), .ZN(n11751) );
  OR2_X1 U14209 ( .A1(n13321), .A2(n12958), .ZN(n11752) );
  XNOR2_X1 U14210 ( .A(n13195), .B(n12957), .ZN(n13187) );
  INV_X1 U14211 ( .A(n13187), .ZN(n11753) );
  NAND2_X1 U14212 ( .A1(n13307), .A2(n12956), .ZN(n11754) );
  NAND2_X1 U14213 ( .A1(n13174), .A2(n11754), .ZN(n13154) );
  OR2_X1 U14214 ( .A1(n13159), .A2(n12955), .ZN(n11755) );
  NAND2_X1 U14215 ( .A1(n13154), .A2(n11755), .ZN(n11757) );
  NAND2_X1 U14216 ( .A1(n13159), .A2(n12955), .ZN(n11756) );
  NAND2_X1 U14217 ( .A1(n13290), .A2(n12918), .ZN(n11758) );
  OR2_X1 U14218 ( .A1(n13282), .A2(n11929), .ZN(n11759) );
  OR2_X2 U14219 ( .A1(n13098), .A2(n13097), .ZN(n13274) );
  INV_X1 U14220 ( .A(n13070), .ZN(n13075) );
  NAND2_X1 U14221 ( .A1(n13076), .A2(n13075), .ZN(n13074) );
  INV_X1 U14222 ( .A(n13330), .ZN(n13243) );
  INV_X1 U14223 ( .A(n13195), .ZN(n13314) );
  NAND2_X1 U14224 ( .A1(n13260), .A2(n13079), .ZN(n13062) );
  OAI211_X1 U14225 ( .C1(n13260), .C2(n13079), .A(n13206), .B(n13062), .ZN(
        n13263) );
  INV_X1 U14226 ( .A(n13260), .ZN(n11950) );
  OAI22_X1 U14227 ( .A1(n14714), .A2(n11765), .B1(n11764), .B2(n14716), .ZN(
        n11766) );
  AOI21_X1 U14228 ( .B1(n11950), .B2(n13194), .A(n11766), .ZN(n11767) );
  OAI21_X1 U14229 ( .B1(n13263), .B2(n13197), .A(n11767), .ZN(n11768) );
  AOI21_X1 U14230 ( .B1(n13259), .B2(n13183), .A(n11768), .ZN(n11769) );
  OAI21_X1 U14231 ( .B1(n6451), .B2(n13253), .A(n11769), .ZN(P2_U3236) );
  INV_X1 U14232 ( .A(n11770), .ZN(n11774) );
  OAI222_X1 U14233 ( .A1(P1_U3086), .A2(n8261), .B1(n14198), .B2(n11774), .C1(
        n11771), .C2(n14195), .ZN(P1_U3326) );
  OAI222_X1 U14234 ( .A1(n13373), .A2(n11774), .B1(n11773), .B2(P2_U3088), 
        .C1(n11772), .C2(n13377), .ZN(P2_U3298) );
  INV_X1 U14235 ( .A(n11775), .ZN(n14190) );
  OAI222_X1 U14236 ( .A1(n13373), .A2(n14190), .B1(n12039), .B2(P2_U3088), 
        .C1(n11776), .C2(n13377), .ZN(P2_U3300) );
  NOR2_X1 U14237 ( .A1(n11777), .A2(n12023), .ZN(n11778) );
  NAND2_X2 U14238 ( .A1(n11779), .A2(n11778), .ZN(n11797) );
  BUF_X8 U14239 ( .A(n7348), .Z(n11985) );
  MUX2_X1 U14240 ( .A(n12963), .B(n14332), .S(n11985), .Z(n11875) );
  NAND2_X1 U14241 ( .A1(n11780), .A2(n12028), .ZN(n11781) );
  OAI211_X1 U14242 ( .C1(n11783), .C2(n11797), .A(n11782), .B(n11781), .ZN(
        n11787) );
  MUX2_X1 U14243 ( .A(n11784), .B(n12978), .S(n11797), .Z(n11788) );
  NAND2_X1 U14244 ( .A1(n11787), .A2(n11788), .ZN(n11786) );
  MUX2_X1 U14245 ( .A(n11784), .B(n12978), .S(n7348), .Z(n11785) );
  NAND2_X1 U14246 ( .A1(n11786), .A2(n11785), .ZN(n11792) );
  INV_X1 U14247 ( .A(n11787), .ZN(n11790) );
  INV_X1 U14248 ( .A(n11788), .ZN(n11789) );
  NAND2_X1 U14249 ( .A1(n11790), .A2(n11789), .ZN(n11791) );
  MUX2_X1 U14250 ( .A(n12977), .B(n11793), .S(n11797), .Z(n11795) );
  MUX2_X1 U14251 ( .A(n12977), .B(n11793), .S(n7348), .Z(n11794) );
  INV_X1 U14252 ( .A(n11795), .ZN(n11796) );
  MUX2_X1 U14253 ( .A(n14730), .B(n12976), .S(n11797), .Z(n11801) );
  NAND2_X1 U14254 ( .A1(n11800), .A2(n11801), .ZN(n11799) );
  MUX2_X1 U14255 ( .A(n14730), .B(n12976), .S(n11985), .Z(n11798) );
  NAND2_X1 U14256 ( .A1(n11799), .A2(n11798), .ZN(n11805) );
  INV_X1 U14257 ( .A(n11800), .ZN(n11803) );
  INV_X1 U14258 ( .A(n11801), .ZN(n11802) );
  NAND2_X1 U14259 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  MUX2_X1 U14260 ( .A(n12975), .B(n11806), .S(n11985), .Z(n11807) );
  MUX2_X1 U14261 ( .A(n12974), .B(n11810), .S(n11985), .Z(n11814) );
  NAND2_X1 U14262 ( .A1(n11813), .A2(n11814), .ZN(n11812) );
  NAND2_X1 U14263 ( .A1(n11812), .A2(n11811), .ZN(n11818) );
  INV_X1 U14264 ( .A(n11813), .ZN(n11816) );
  INV_X1 U14265 ( .A(n11814), .ZN(n11815) );
  NAND2_X1 U14266 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  MUX2_X1 U14267 ( .A(n12973), .B(n11819), .S(n11967), .Z(n11821) );
  MUX2_X1 U14268 ( .A(n12973), .B(n11819), .S(n11985), .Z(n11820) );
  INV_X1 U14269 ( .A(n11821), .ZN(n11822) );
  MUX2_X1 U14270 ( .A(n12972), .B(n14746), .S(n11985), .Z(n11826) );
  NAND2_X1 U14271 ( .A1(n11825), .A2(n11826), .ZN(n11824) );
  NAND2_X1 U14272 ( .A1(n11824), .A2(n11823), .ZN(n11830) );
  INV_X1 U14273 ( .A(n11825), .ZN(n11828) );
  INV_X1 U14274 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U14275 ( .A1(n11828), .A2(n11827), .ZN(n11829) );
  MUX2_X1 U14276 ( .A(n12971), .B(n14755), .S(n11967), .Z(n11832) );
  MUX2_X1 U14277 ( .A(n12971), .B(n14755), .S(n11985), .Z(n11831) );
  MUX2_X1 U14278 ( .A(n12969), .B(n11834), .S(n11985), .Z(n11838) );
  NAND2_X1 U14279 ( .A1(n11837), .A2(n11838), .ZN(n11836) );
  NAND2_X1 U14280 ( .A1(n11836), .A2(n11835), .ZN(n11842) );
  INV_X1 U14281 ( .A(n11837), .ZN(n11840) );
  INV_X1 U14282 ( .A(n11838), .ZN(n11839) );
  NAND2_X1 U14283 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  MUX2_X1 U14284 ( .A(n12968), .B(n11843), .S(n11967), .Z(n11845) );
  MUX2_X1 U14285 ( .A(n12968), .B(n11843), .S(n11985), .Z(n11844) );
  INV_X1 U14286 ( .A(n11845), .ZN(n11846) );
  MUX2_X1 U14287 ( .A(n12967), .B(n11847), .S(n11985), .Z(n11851) );
  NAND2_X1 U14288 ( .A1(n11850), .A2(n11851), .ZN(n11849) );
  NAND2_X1 U14289 ( .A1(n11849), .A2(n11848), .ZN(n11855) );
  INV_X1 U14290 ( .A(n11850), .ZN(n11853) );
  INV_X1 U14291 ( .A(n11851), .ZN(n11852) );
  NAND2_X1 U14292 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  MUX2_X1 U14293 ( .A(n12966), .B(n14345), .S(n11967), .Z(n11857) );
  MUX2_X1 U14294 ( .A(n12966), .B(n14345), .S(n11985), .Z(n11856) );
  MUX2_X1 U14295 ( .A(n12965), .B(n14339), .S(n11985), .Z(n11862) );
  NAND2_X1 U14296 ( .A1(n11861), .A2(n11862), .ZN(n11860) );
  NAND2_X1 U14297 ( .A1(n11860), .A2(n11859), .ZN(n11866) );
  INV_X1 U14298 ( .A(n11861), .ZN(n11864) );
  INV_X1 U14299 ( .A(n11862), .ZN(n11863) );
  NAND2_X1 U14300 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  NAND2_X1 U14301 ( .A1(n11866), .A2(n11865), .ZN(n11870) );
  MUX2_X1 U14302 ( .A(n12964), .B(n11867), .S(n11967), .Z(n11871) );
  NAND2_X1 U14303 ( .A1(n11870), .A2(n11871), .ZN(n11869) );
  MUX2_X1 U14304 ( .A(n12964), .B(n11867), .S(n11985), .Z(n11868) );
  INV_X1 U14305 ( .A(n11870), .ZN(n11873) );
  INV_X1 U14306 ( .A(n11871), .ZN(n11872) );
  MUX2_X1 U14307 ( .A(n12961), .B(n12876), .S(n11985), .Z(n11883) );
  AND2_X1 U14308 ( .A1(n12962), .A2(n11967), .ZN(n11877) );
  NOR2_X1 U14309 ( .A1(n12962), .A2(n11967), .ZN(n11876) );
  MUX2_X1 U14310 ( .A(n11877), .B(n11876), .S(n14321), .Z(n11878) );
  AOI21_X1 U14311 ( .B1(n11883), .B2(n11879), .A(n11878), .ZN(n11880) );
  NAND2_X1 U14312 ( .A1(n11881), .A2(n11880), .ZN(n11885) );
  NOR2_X1 U14313 ( .A1(n12876), .A2(n12961), .ZN(n11882) );
  OR2_X1 U14314 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  NAND2_X1 U14315 ( .A1(n11885), .A2(n11884), .ZN(n11888) );
  MUX2_X1 U14316 ( .A(n12960), .B(n13330), .S(n11967), .Z(n11889) );
  NAND2_X1 U14317 ( .A1(n11888), .A2(n11889), .ZN(n11887) );
  MUX2_X1 U14318 ( .A(n12960), .B(n13330), .S(n11985), .Z(n11886) );
  NAND2_X1 U14319 ( .A1(n11887), .A2(n11886), .ZN(n11893) );
  INV_X1 U14320 ( .A(n11888), .ZN(n11891) );
  INV_X1 U14321 ( .A(n11889), .ZN(n11890) );
  NAND2_X1 U14322 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  MUX2_X1 U14323 ( .A(n12959), .B(n13326), .S(n11985), .Z(n11897) );
  NAND2_X1 U14324 ( .A1(n11896), .A2(n11897), .ZN(n11895) );
  MUX2_X1 U14325 ( .A(n12959), .B(n13326), .S(n11967), .Z(n11894) );
  NAND2_X1 U14326 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  INV_X1 U14327 ( .A(n11896), .ZN(n11899) );
  INV_X1 U14328 ( .A(n11897), .ZN(n11898) );
  NAND2_X1 U14329 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  MUX2_X1 U14330 ( .A(n12958), .B(n13321), .S(n11967), .Z(n11903) );
  MUX2_X1 U14331 ( .A(n12958), .B(n13321), .S(n11985), .Z(n11902) );
  INV_X1 U14332 ( .A(n11903), .ZN(n11904) );
  MUX2_X1 U14333 ( .A(n12957), .B(n13195), .S(n11985), .Z(n11908) );
  NAND2_X1 U14334 ( .A1(n11907), .A2(n11908), .ZN(n11906) );
  NAND2_X1 U14335 ( .A1(n11906), .A2(n11905), .ZN(n11912) );
  INV_X1 U14336 ( .A(n11907), .ZN(n11910) );
  INV_X1 U14337 ( .A(n11908), .ZN(n11909) );
  NAND2_X1 U14338 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  MUX2_X1 U14339 ( .A(n12956), .B(n13307), .S(n11967), .Z(n11914) );
  MUX2_X1 U14340 ( .A(n12956), .B(n13307), .S(n11985), .Z(n11913) );
  MUX2_X1 U14341 ( .A(n12955), .B(n13159), .S(n11985), .Z(n11918) );
  NAND2_X1 U14342 ( .A1(n11917), .A2(n11918), .ZN(n11916) );
  NAND2_X1 U14343 ( .A1(n11916), .A2(n11915), .ZN(n11922) );
  INV_X1 U14344 ( .A(n11917), .ZN(n11920) );
  INV_X1 U14345 ( .A(n11918), .ZN(n11919) );
  NAND2_X1 U14346 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  NAND2_X1 U14347 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  MUX2_X1 U14348 ( .A(n12954), .B(n13296), .S(n11967), .Z(n11924) );
  NAND2_X1 U14349 ( .A1(n11923), .A2(n11924), .ZN(n11928) );
  MUX2_X1 U14350 ( .A(n12954), .B(n13296), .S(n11985), .Z(n11927) );
  INV_X1 U14351 ( .A(n11923), .ZN(n11926) );
  INV_X1 U14352 ( .A(n11924), .ZN(n11925) );
  MUX2_X1 U14353 ( .A(n12918), .B(n13290), .S(n11985), .Z(n11931) );
  MUX2_X1 U14354 ( .A(n11929), .B(n13282), .S(n11985), .Z(n11939) );
  MUX2_X1 U14355 ( .A(n12016), .B(n12952), .S(n11985), .Z(n11938) );
  AOI22_X1 U14356 ( .A1(n11932), .A2(n11931), .B1(n11939), .B2(n11938), .ZN(
        n11945) );
  MUX2_X1 U14357 ( .A(n13131), .B(n12953), .S(n11985), .Z(n11930) );
  OAI21_X1 U14358 ( .B1(n11932), .B2(n11931), .A(n11930), .ZN(n11944) );
  MUX2_X1 U14359 ( .A(n12951), .B(n13272), .S(n11967), .Z(n11947) );
  MUX2_X1 U14360 ( .A(n11934), .B(n13092), .S(n11985), .Z(n11948) );
  INV_X1 U14361 ( .A(n11938), .ZN(n11941) );
  INV_X1 U14362 ( .A(n11939), .ZN(n11940) );
  AOI21_X1 U14363 ( .B1(n11945), .B2(n11944), .A(n11943), .ZN(n11958) );
  INV_X1 U14364 ( .A(n11946), .ZN(n11949) );
  NOR3_X1 U14365 ( .A1(n11949), .A2(n11936), .A3(n11935), .ZN(n11957) );
  MUX2_X1 U14366 ( .A(n12949), .B(n11950), .S(n11967), .Z(n11972) );
  MUX2_X1 U14367 ( .A(n11951), .B(n13260), .S(n11985), .Z(n11973) );
  AOI21_X1 U14368 ( .B1(n11972), .B2(n11973), .A(n11954), .ZN(n11955) );
  INV_X1 U14369 ( .A(n11955), .ZN(n11956) );
  NAND2_X1 U14370 ( .A1(n13363), .A2(n11959), .ZN(n11961) );
  MUX2_X1 U14371 ( .A(n12948), .B(n13055), .S(n11967), .Z(n11980) );
  INV_X1 U14372 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n11965) );
  NAND2_X1 U14373 ( .A1(n9198), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U14374 ( .A1(n11962), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n11963) );
  OAI211_X1 U14375 ( .C1(n11966), .C2(n11965), .A(n11964), .B(n11963), .ZN(
        n13057) );
  NAND2_X1 U14376 ( .A1(n11967), .A2(n13057), .ZN(n11981) );
  OAI211_X1 U14377 ( .C1(n11969), .C2(n12031), .A(n11981), .B(n11968), .ZN(
        n11970) );
  AND2_X1 U14378 ( .A1(n11970), .A2(n12948), .ZN(n11971) );
  AOI21_X1 U14379 ( .B1(n13055), .B2(n11985), .A(n11971), .ZN(n11979) );
  OAI22_X1 U14380 ( .A1(n11980), .A2(n11979), .B1(n11973), .B2(n11972), .ZN(
        n11978) );
  NAND2_X1 U14381 ( .A1(n14185), .A2(n11974), .ZN(n11976) );
  INV_X1 U14382 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U14383 ( .A1(n13059), .A2(n13057), .ZN(n11977) );
  NAND2_X1 U14384 ( .A1(n11982), .A2(n11977), .ZN(n11989) );
  INV_X1 U14385 ( .A(n11981), .ZN(n11984) );
  INV_X1 U14386 ( .A(n11982), .ZN(n11983) );
  AOI211_X1 U14387 ( .C1(n11985), .C2(n13059), .A(n11984), .B(n11983), .ZN(
        n11986) );
  OAI21_X2 U14388 ( .B1(n11988), .B2(n7384), .A(n11987), .ZN(n12035) );
  NOR2_X1 U14389 ( .A1(n12035), .A2(n14709), .ZN(n12025) );
  INV_X1 U14390 ( .A(n11989), .ZN(n12021) );
  XNOR2_X1 U14391 ( .A(n13258), .B(n12948), .ZN(n12020) );
  XNOR2_X1 U14392 ( .A(n13159), .B(n12882), .ZN(n13155) );
  NOR4_X1 U14393 ( .A1(n14708), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11995) );
  NAND4_X1 U14394 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11997) );
  NOR4_X1 U14395 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12003) );
  NAND4_X1 U14396 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  NOR3_X1 U14397 ( .A1(n12007), .A2(n12006), .A3(n12005), .ZN(n12009) );
  NAND4_X1 U14398 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12012) );
  NOR4_X1 U14399 ( .A1(n13203), .A2(n13230), .A3(n12013), .A4(n12012), .ZN(
        n12014) );
  XNOR2_X1 U14400 ( .A(n13326), .B(n12959), .ZN(n13217) );
  NAND4_X1 U14401 ( .A1(n13173), .A2(n12014), .A3(n13187), .A4(n13217), .ZN(
        n12015) );
  NOR4_X1 U14402 ( .A1(n13122), .A2(n13155), .A3(n13139), .A4(n12015), .ZN(
        n12017) );
  XNOR2_X1 U14403 ( .A(n12016), .B(n12952), .ZN(n13112) );
  NAND4_X1 U14404 ( .A1(n13070), .A2(n12017), .A3(n13098), .A4(n13112), .ZN(
        n12018) );
  NAND2_X1 U14405 ( .A1(n6479), .A2(n12023), .ZN(n12024) );
  NOR2_X1 U14406 ( .A1(n12025), .A2(n12024), .ZN(n12037) );
  OAI22_X1 U14407 ( .A1(n12040), .A2(n12028), .B1(n12027), .B2(n12026), .ZN(
        n12029) );
  INV_X1 U14408 ( .A(n12029), .ZN(n12034) );
  INV_X1 U14409 ( .A(n11779), .ZN(n14709) );
  OAI22_X1 U14410 ( .A1(n14709), .A2(n12031), .B1(n13053), .B2(n12030), .ZN(
        n12032) );
  NAND2_X1 U14411 ( .A1(n12035), .A2(n12032), .ZN(n12033) );
  OAI21_X1 U14412 ( .B1(n12035), .B2(n12034), .A(n12033), .ZN(n12036) );
  NOR2_X1 U14413 ( .A1(n12037), .A2(n12036), .ZN(n12044) );
  INV_X1 U14414 ( .A(n14723), .ZN(n14725) );
  NOR4_X1 U14415 ( .A1(n14725), .A2(n12919), .A3(n12039), .A4(n12038), .ZN(
        n12042) );
  OAI21_X1 U14416 ( .B1(n12040), .B2(n12043), .A(P2_B_REG_SCAN_IN), .ZN(n12041) );
  OAI22_X1 U14417 ( .A1(n12044), .A2(n12043), .B1(n12042), .B2(n12041), .ZN(
        P2_U3328) );
  XNOR2_X1 U14418 ( .A(n12477), .B(n12045), .ZN(n12052) );
  INV_X1 U14419 ( .A(n12052), .ZN(n12046) );
  NAND2_X1 U14420 ( .A1(n12046), .A2(n12229), .ZN(n12058) );
  INV_X1 U14421 ( .A(n12047), .ZN(n12048) );
  NAND4_X1 U14422 ( .A1(n12057), .A2(n12229), .A3(n12048), .A4(n12052), .ZN(
        n12056) );
  AOI22_X1 U14423 ( .A1(n12452), .A2(n12242), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12050) );
  NAND2_X1 U14424 ( .A1(n12480), .A2(n12248), .ZN(n12049) );
  OAI211_X1 U14425 ( .C1(n12473), .C2(n12244), .A(n12050), .B(n12049), .ZN(
        n12054) );
  NOR4_X1 U14426 ( .A1(n12052), .A2(n12051), .A3(n12452), .A4(n12237), .ZN(
        n12053) );
  AOI211_X1 U14427 ( .C1(n12219), .C2(n12479), .A(n12054), .B(n12053), .ZN(
        n12055) );
  OAI211_X1 U14428 ( .C1(n12058), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        P3_U3160) );
  INV_X1 U14429 ( .A(n12059), .ZN(n12061) );
  OAI222_X1 U14430 ( .A1(n12062), .A2(P3_U3151), .B1(n12821), .B2(n12061), 
        .C1(n12060), .C2(n12817), .ZN(P3_U3265) );
  OAI211_X1 U14431 ( .C1(n12065), .C2(n12064), .A(n12063), .B(n12229), .ZN(
        n12072) );
  AOI21_X1 U14432 ( .B1(n12219), .B2(n12067), .A(n12066), .ZN(n12071) );
  AOI22_X1 U14433 ( .A1(n12220), .A2(n14826), .B1(n12242), .B2(n14855), .ZN(
        n12070) );
  NAND2_X1 U14434 ( .A1(n12248), .A2(n12068), .ZN(n12069) );
  NAND4_X1 U14435 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        P3_U3153) );
  INV_X1 U14436 ( .A(n12236), .ZN(n12073) );
  AOI21_X1 U14437 ( .B1(n12075), .B2(n12074), .A(n12073), .ZN(n12082) );
  NOR2_X1 U14438 ( .A1(n12801), .A2(n12245), .ZN(n12080) );
  NAND2_X1 U14439 ( .A1(n12242), .A2(n12668), .ZN(n12078) );
  INV_X1 U14440 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12076) );
  NOR2_X1 U14441 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12076), .ZN(n12284) );
  INV_X1 U14442 ( .A(n12284), .ZN(n12077) );
  OAI211_X1 U14443 ( .C1(n12638), .C2(n12244), .A(n12078), .B(n12077), .ZN(
        n12079) );
  AOI211_X1 U14444 ( .C1(n12675), .C2(n12248), .A(n12080), .B(n12079), .ZN(
        n12081) );
  OAI21_X1 U14445 ( .B1(n12082), .B2(n12237), .A(n12081), .ZN(P3_U3155) );
  AOI21_X1 U14446 ( .B1(n12547), .B2(n12083), .A(n6438), .ZN(n12088) );
  AOI22_X1 U14447 ( .A1(n12220), .A2(n12536), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12085) );
  NAND2_X1 U14448 ( .A1(n12248), .A2(n12539), .ZN(n12084) );
  OAI211_X1 U14449 ( .C1(n12558), .C2(n12210), .A(n12085), .B(n12084), .ZN(
        n12086) );
  AOI21_X1 U14450 ( .B1(n12709), .B2(n12219), .A(n12086), .ZN(n12087) );
  OAI21_X1 U14451 ( .B1(n12088), .B2(n12237), .A(n12087), .ZN(P3_U3156) );
  AOI22_X1 U14452 ( .A1(n12220), .A2(n12252), .B1(n12242), .B2(n12253), .ZN(
        n12089) );
  NAND2_X1 U14453 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n14818)
         );
  OAI211_X1 U14454 ( .C1(n12090), .C2(n12245), .A(n12089), .B(n14818), .ZN(
        n12096) );
  INV_X1 U14455 ( .A(n12091), .ZN(n12092) );
  AOI211_X1 U14456 ( .C1(n12094), .C2(n12093), .A(n12237), .B(n12092), .ZN(
        n12095) );
  AOI211_X1 U14457 ( .C1(n12097), .C2(n12248), .A(n12096), .B(n12095), .ZN(
        n12098) );
  INV_X1 U14458 ( .A(n12098), .ZN(P3_U3157) );
  XNOR2_X1 U14459 ( .A(n12099), .B(n12100), .ZN(n12105) );
  NAND2_X1 U14460 ( .A1(n12242), .A2(n12589), .ZN(n12101) );
  NAND2_X1 U14461 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12397)
         );
  OAI211_X1 U14462 ( .C1(n12559), .C2(n12244), .A(n12101), .B(n12397), .ZN(
        n12103) );
  NOR2_X1 U14463 ( .A1(n12782), .A2(n12245), .ZN(n12102) );
  AOI211_X1 U14464 ( .C1(n12594), .C2(n12248), .A(n12103), .B(n12102), .ZN(
        n12104) );
  OAI21_X1 U14465 ( .B1(n12105), .B2(n12237), .A(n12104), .ZN(P3_U3159) );
  INV_X1 U14466 ( .A(n12107), .ZN(n12108) );
  AOI21_X1 U14467 ( .B1(n12109), .B2(n12106), .A(n12108), .ZN(n12114) );
  AOI22_X1 U14468 ( .A1(n12220), .A2(n12535), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12111) );
  NAND2_X1 U14469 ( .A1(n12248), .A2(n12563), .ZN(n12110) );
  OAI211_X1 U14470 ( .C1(n12559), .C2(n12210), .A(n12111), .B(n12110), .ZN(
        n12112) );
  AOI21_X1 U14471 ( .B1(n12562), .B2(n12219), .A(n12112), .ZN(n12113) );
  OAI21_X1 U14472 ( .B1(n12114), .B2(n12237), .A(n12113), .ZN(P3_U3163) );
  NAND2_X1 U14473 ( .A1(n12116), .A2(n12115), .ZN(n12120) );
  XNOR2_X1 U14474 ( .A(n12117), .B(n12118), .ZN(n12198) );
  OAI22_X1 U14475 ( .A1(n12198), .A2(n12252), .B1(n12117), .B2(n12118), .ZN(
        n12119) );
  XOR2_X1 U14476 ( .A(n12120), .B(n12119), .Z(n12121) );
  NAND2_X1 U14477 ( .A1(n12121), .A2(n12229), .ZN(n12127) );
  AOI21_X1 U14478 ( .B1(n12219), .B2(n12410), .A(n12122), .ZN(n12126) );
  AOI22_X1 U14479 ( .A1(n12220), .A2(n12668), .B1(n12242), .B2(n12252), .ZN(
        n12125) );
  NAND2_X1 U14480 ( .A1(n12248), .A2(n12123), .ZN(n12124) );
  NAND4_X1 U14481 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        P3_U3164) );
  INV_X1 U14482 ( .A(n12699), .ZN(n12518) );
  INV_X1 U14483 ( .A(n12128), .ZN(n12167) );
  INV_X1 U14484 ( .A(n12129), .ZN(n12131) );
  NOR3_X1 U14485 ( .A1(n12167), .A2(n12131), .A3(n12130), .ZN(n12134) );
  INV_X1 U14486 ( .A(n12132), .ZN(n12133) );
  OAI21_X1 U14487 ( .B1(n12134), .B2(n12133), .A(n12229), .ZN(n12139) );
  AOI22_X1 U14488 ( .A1(n12512), .A2(n12220), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12135) );
  OAI21_X1 U14489 ( .B1(n12136), .B2(n12210), .A(n12135), .ZN(n12137) );
  AOI21_X1 U14490 ( .B1(n12516), .B2(n12248), .A(n12137), .ZN(n12138) );
  OAI211_X1 U14491 ( .C1(n12518), .C2(n12245), .A(n12139), .B(n12138), .ZN(
        P3_U3165) );
  NAND2_X1 U14492 ( .A1(n12236), .A2(n12140), .ZN(n12240) );
  NAND2_X1 U14493 ( .A1(n12240), .A2(n12141), .ZN(n12143) );
  XNOR2_X1 U14494 ( .A(n12143), .B(n12142), .ZN(n12148) );
  NAND2_X1 U14495 ( .A1(n12242), .A2(n12667), .ZN(n12144) );
  NAND2_X1 U14496 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12326)
         );
  OAI211_X1 U14497 ( .C1(n12637), .C2(n12244), .A(n12144), .B(n12326), .ZN(
        n12146) );
  NOR2_X1 U14498 ( .A1(n12794), .A2(n12245), .ZN(n12145) );
  AOI211_X1 U14499 ( .C1(n12643), .C2(n12248), .A(n12146), .B(n12145), .ZN(
        n12147) );
  OAI21_X1 U14500 ( .B1(n12148), .B2(n12237), .A(n12147), .ZN(P3_U3166) );
  XNOR2_X1 U14501 ( .A(n12150), .B(n12149), .ZN(n12151) );
  NAND2_X1 U14502 ( .A1(n12151), .A2(n12229), .ZN(n12156) );
  AOI21_X1 U14503 ( .B1(n12219), .B2(n14859), .A(n12152), .ZN(n12155) );
  AOI22_X1 U14504 ( .A1(n12220), .A2(n14855), .B1(n12242), .B2(n14890), .ZN(
        n12154) );
  NAND2_X1 U14505 ( .A1(n12248), .A2(n14860), .ZN(n12153) );
  NAND4_X1 U14506 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        P3_U3167) );
  XNOR2_X1 U14507 ( .A(n12157), .B(n12158), .ZN(n12163) );
  NAND2_X1 U14508 ( .A1(n12242), .A2(n12416), .ZN(n12159) );
  NAND2_X1 U14509 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12347)
         );
  OAI211_X1 U14510 ( .C1(n12622), .C2(n12244), .A(n12159), .B(n12347), .ZN(
        n12161) );
  INV_X1 U14511 ( .A(n12430), .ZN(n12790) );
  NOR2_X1 U14512 ( .A1(n12790), .A2(n12245), .ZN(n12160) );
  AOI211_X1 U14513 ( .C1(n12626), .C2(n12248), .A(n12161), .B(n12160), .ZN(
        n12162) );
  OAI21_X1 U14514 ( .B1(n12163), .B2(n12237), .A(n12162), .ZN(P3_U3168) );
  INV_X1 U14515 ( .A(n12443), .ZN(n12771) );
  INV_X1 U14516 ( .A(n12164), .ZN(n12166) );
  NOR3_X1 U14517 ( .A1(n6438), .A2(n12166), .A3(n12165), .ZN(n12168) );
  OAI21_X1 U14518 ( .B1(n12168), .B2(n12167), .A(n12229), .ZN(n12172) );
  AOI22_X1 U14519 ( .A1(n12220), .A2(n12447), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12169) );
  OAI21_X1 U14520 ( .B1(n12525), .B2(n12210), .A(n12169), .ZN(n12170) );
  AOI21_X1 U14521 ( .B1(n12528), .B2(n12248), .A(n12170), .ZN(n12171) );
  OAI211_X1 U14522 ( .C1(n12771), .C2(n12245), .A(n12172), .B(n12171), .ZN(
        P3_U3169) );
  OAI21_X1 U14523 ( .B1(n12175), .B2(n12174), .A(n12173), .ZN(n12176) );
  NAND2_X1 U14524 ( .A1(n12176), .A2(n12229), .ZN(n12182) );
  AOI21_X1 U14525 ( .B1(n12219), .B2(n14864), .A(n12177), .ZN(n12181) );
  AOI22_X1 U14526 ( .A1(n12220), .A2(n12255), .B1(n12242), .B2(n9611), .ZN(
        n12180) );
  NAND2_X1 U14527 ( .A1(n12248), .A2(n12178), .ZN(n12179) );
  NAND4_X1 U14528 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        P3_U3170) );
  XNOR2_X1 U14529 ( .A(n12183), .B(n12184), .ZN(n12189) );
  AOI22_X1 U14530 ( .A1(n12220), .A2(n12575), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12186) );
  NAND2_X1 U14531 ( .A1(n12248), .A2(n12577), .ZN(n12185) );
  OAI211_X1 U14532 ( .C1(n12604), .C2(n12210), .A(n12186), .B(n12185), .ZN(
        n12187) );
  AOI21_X1 U14533 ( .B1(n12721), .B2(n12219), .A(n12187), .ZN(n12188) );
  OAI21_X1 U14534 ( .B1(n12189), .B2(n12237), .A(n12188), .ZN(P3_U3173) );
  INV_X1 U14535 ( .A(n12191), .ZN(n12192) );
  AOI21_X1 U14536 ( .B1(n12535), .B2(n12190), .A(n12192), .ZN(n12197) );
  AOI22_X1 U14537 ( .A1(n12242), .A2(n12575), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12194) );
  NAND2_X1 U14538 ( .A1(n12248), .A2(n12551), .ZN(n12193) );
  OAI211_X1 U14539 ( .C1(n12525), .C2(n12244), .A(n12194), .B(n12193), .ZN(
        n12195) );
  AOI21_X1 U14540 ( .B1(n12714), .B2(n12219), .A(n12195), .ZN(n12196) );
  OAI21_X1 U14541 ( .B1(n12197), .B2(n12237), .A(n12196), .ZN(P3_U3175) );
  XNOR2_X1 U14542 ( .A(n12198), .B(n12252), .ZN(n12199) );
  NAND2_X1 U14543 ( .A1(n12199), .A2(n12229), .ZN(n12205) );
  AOI21_X1 U14544 ( .B1(n12219), .B2(n12201), .A(n12200), .ZN(n12204) );
  AOI22_X1 U14545 ( .A1(n12220), .A2(n14272), .B1(n12242), .B2(n14825), .ZN(
        n12203) );
  NAND2_X1 U14546 ( .A1(n12248), .A2(n14293), .ZN(n12202) );
  NAND4_X1 U14547 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        P3_U3176) );
  XNOR2_X1 U14548 ( .A(n12206), .B(n12207), .ZN(n12213) );
  AND2_X1 U14549 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12377) );
  AOI21_X1 U14550 ( .B1(n12220), .B2(n12574), .A(n12377), .ZN(n12209) );
  NAND2_X1 U14551 ( .A1(n12248), .A2(n12610), .ZN(n12208) );
  OAI211_X1 U14552 ( .C1(n12637), .C2(n12210), .A(n12209), .B(n12208), .ZN(
        n12211) );
  AOI21_X1 U14553 ( .B1(n12609), .B2(n12219), .A(n12211), .ZN(n12212) );
  OAI21_X1 U14554 ( .B1(n12213), .B2(n12237), .A(n12212), .ZN(P3_U3178) );
  OAI211_X1 U14555 ( .C1(n12216), .C2(n12215), .A(n12214), .B(n12229), .ZN(
        n12225) );
  AOI21_X1 U14556 ( .B1(n12219), .B2(n12218), .A(n12217), .ZN(n12224) );
  AOI22_X1 U14557 ( .A1(n12220), .A2(n12254), .B1(n12242), .B2(n12255), .ZN(
        n12223) );
  NAND2_X1 U14558 ( .A1(n12248), .A2(n12221), .ZN(n12222) );
  NAND4_X1 U14559 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        P3_U3179) );
  INV_X1 U14560 ( .A(n12507), .ZN(n12766) );
  OAI21_X1 U14561 ( .B1(n12228), .B2(n12226), .A(n12227), .ZN(n12230) );
  NAND2_X1 U14562 ( .A1(n12230), .A2(n12229), .ZN(n12234) );
  AOI22_X1 U14563 ( .A1(n12447), .A2(n12242), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12231) );
  OAI21_X1 U14564 ( .B1(n12502), .B2(n12244), .A(n12231), .ZN(n12232) );
  AOI21_X1 U14565 ( .B1(n12506), .B2(n12248), .A(n12232), .ZN(n12233) );
  OAI211_X1 U14566 ( .C1(n12766), .C2(n12245), .A(n12234), .B(n12233), .ZN(
        P3_U3180) );
  NAND2_X1 U14567 ( .A1(n12236), .A2(n12235), .ZN(n12239) );
  AOI21_X1 U14568 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12241) );
  NAND2_X1 U14569 ( .A1(n12241), .A2(n12240), .ZN(n12250) );
  NAND2_X1 U14570 ( .A1(n12242), .A2(n14273), .ZN(n12243) );
  NAND2_X1 U14571 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12304)
         );
  OAI211_X1 U14572 ( .C1(n12651), .C2(n12244), .A(n12243), .B(n12304), .ZN(
        n12247) );
  INV_X1 U14573 ( .A(n12424), .ZN(n12797) );
  NOR2_X1 U14574 ( .A1(n12797), .A2(n12245), .ZN(n12246) );
  AOI211_X1 U14575 ( .C1(n12659), .C2(n12248), .A(n12247), .B(n12246), .ZN(
        n12249) );
  NAND2_X1 U14576 ( .A1(n12250), .A2(n12249), .ZN(P3_U3181) );
  MUX2_X1 U14577 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12251), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14578 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12461), .S(P3_U3897), .Z(
        P3_U3521) );
  INV_X1 U14579 ( .A(n12485), .ZN(n12460) );
  MUX2_X1 U14580 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12460), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14581 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12452), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14582 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12512), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14583 ( .A(n12447), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12258), .Z(
        P3_U3516) );
  MUX2_X1 U14584 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12536), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14585 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12547), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14586 ( .A(n12535), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12258), .Z(
        P3_U3513) );
  MUX2_X1 U14587 ( .A(n12575), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12258), .Z(
        P3_U3512) );
  MUX2_X1 U14588 ( .A(n12588), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12258), .Z(
        P3_U3511) );
  MUX2_X1 U14589 ( .A(n12574), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12258), .Z(
        P3_U3510) );
  MUX2_X1 U14590 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12589), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14591 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12429), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14592 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12416), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14593 ( .A(n12667), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12258), .Z(
        P3_U3506) );
  MUX2_X1 U14594 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14273), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14595 ( .A(n12668), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12258), .Z(
        P3_U3504) );
  MUX2_X1 U14596 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14272), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14597 ( .A(n12252), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12258), .Z(
        P3_U3502) );
  MUX2_X1 U14598 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14825), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14599 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12253), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14600 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n14826), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14601 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12254), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14602 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n14855), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14603 ( .A(n12255), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12258), .Z(
        P3_U3496) );
  MUX2_X1 U14604 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n14890), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14605 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n9611), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14606 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n14891), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14607 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12257), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14608 ( .A(n12259), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12258), .Z(
        P3_U3491) );
  INV_X1 U14609 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14276) );
  AOI21_X1 U14610 ( .B1(n14276), .B2(n12261), .A(n12279), .ZN(n12276) );
  MUX2_X1 U14611 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n8117), .Z(n12289) );
  XNOR2_X1 U14612 ( .A(n12289), .B(n12278), .ZN(n12265) );
  OAI21_X1 U14613 ( .B1(n6571), .B2(n12265), .A(n12288), .ZN(n12274) );
  NAND2_X1 U14614 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12268), .ZN(n12282) );
  OAI21_X1 U14615 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12268), .A(n12282), 
        .ZN(n12269) );
  NAND2_X1 U14616 ( .A1(n12269), .A2(n14809), .ZN(n12272) );
  AOI21_X1 U14617 ( .B1(n14799), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12270), 
        .ZN(n12271) );
  OAI211_X1 U14618 ( .C1(n12393), .C2(n14216), .A(n12272), .B(n12271), .ZN(
        n12273) );
  AOI21_X1 U14619 ( .B1(n12274), .B2(n14810), .A(n12273), .ZN(n12275) );
  OAI21_X1 U14620 ( .B1(n12276), .B2(n14815), .A(n12275), .ZN(P3_U3195) );
  NAND2_X1 U14621 ( .A1(n12309), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12298) );
  OAI21_X1 U14622 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12309), .A(n12298), 
        .ZN(n12287) );
  NOR2_X1 U14623 ( .A1(n12280), .A2(n12287), .ZN(n12297) );
  AOI21_X1 U14624 ( .B1(n12280), .B2(n12287), .A(n12297), .ZN(n12296) );
  NAND2_X1 U14625 ( .A1(n14216), .A2(n12281), .ZN(n12283) );
  NAND2_X1 U14626 ( .A1(n12283), .A2(n12282), .ZN(n12303) );
  XNOR2_X1 U14627 ( .A(n12309), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n12286) );
  INV_X1 U14628 ( .A(n12286), .ZN(n12302) );
  XNOR2_X1 U14629 ( .A(n12303), .B(n12302), .ZN(n12294) );
  AOI21_X1 U14630 ( .B1(n14799), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12284), 
        .ZN(n12285) );
  OAI21_X1 U14631 ( .B1(n12393), .B2(n12309), .A(n12285), .ZN(n12293) );
  MUX2_X1 U14632 ( .A(n12287), .B(n12286), .S(n8117), .Z(n12291) );
  NOR2_X1 U14633 ( .A1(n12290), .A2(n12291), .ZN(n12307) );
  AOI211_X1 U14634 ( .C1(n12291), .C2(n12290), .A(n14781), .B(n12307), .ZN(
        n12292) );
  AOI211_X1 U14635 ( .C1(n14809), .C2(n12294), .A(n12293), .B(n12292), .ZN(
        n12295) );
  OAI21_X1 U14636 ( .B1(n12296), .B2(n14815), .A(n12295), .ZN(P3_U3196) );
  INV_X1 U14637 ( .A(n12297), .ZN(n12299) );
  NAND2_X1 U14638 ( .A1(n12300), .A2(n12332), .ZN(n12317) );
  INV_X1 U14639 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15036) );
  AOI21_X1 U14640 ( .B1(n12301), .B2(n15036), .A(n12319), .ZN(n12316) );
  INV_X1 U14641 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12744) );
  XNOR2_X1 U14642 ( .A(n12323), .B(n12744), .ZN(n12314) );
  NAND2_X1 U14643 ( .A1(n14801), .A2(n6851), .ZN(n12305) );
  OAI211_X1 U14644 ( .C1(n12306), .C2(n14797), .A(n12305), .B(n12304), .ZN(
        n12313) );
  MUX2_X1 U14645 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n8117), .Z(n12308) );
  MUX2_X1 U14646 ( .A(n15036), .B(n12744), .S(n8117), .Z(n12310) );
  AOI211_X1 U14647 ( .C1(n12311), .C2(n12310), .A(n14781), .B(n12330), .ZN(
        n12312) );
  AOI211_X1 U14648 ( .C1(n14809), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12315) );
  OAI21_X1 U14649 ( .B1(n12316), .B2(n14815), .A(n12315), .ZN(P3_U3197) );
  INV_X1 U14650 ( .A(n12317), .ZN(n12318) );
  INV_X1 U14651 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U14652 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12344), .B1(n14222), 
        .B2(n12320), .ZN(n12321) );
  AOI21_X1 U14653 ( .B1(n6491), .B2(n12321), .A(n12340), .ZN(n12339) );
  XNOR2_X1 U14654 ( .A(n12344), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12324) );
  OAI21_X1 U14655 ( .B1(n12325), .B2(n12324), .A(n12343), .ZN(n12337) );
  NAND2_X1 U14656 ( .A1(n14801), .A2(n12344), .ZN(n12327) );
  OAI211_X1 U14657 ( .C1(n12328), .C2(n14797), .A(n12327), .B(n12326), .ZN(
        n12336) );
  INV_X1 U14658 ( .A(n12329), .ZN(n12331) );
  MUX2_X1 U14659 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n8117), .Z(n12351) );
  XNOR2_X1 U14660 ( .A(n12351), .B(n14222), .ZN(n12333) );
  NOR2_X1 U14661 ( .A1(n12334), .A2(n12333), .ZN(n12350) );
  AOI211_X1 U14662 ( .C1(n12334), .C2(n12333), .A(n14781), .B(n12350), .ZN(
        n12335) );
  AOI211_X1 U14663 ( .C1(n14809), .C2(n12337), .A(n12336), .B(n12335), .ZN(
        n12338) );
  OAI21_X1 U14664 ( .B1(n12339), .B2(n14815), .A(n12338), .ZN(P3_U3198) );
  INV_X1 U14665 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12342) );
  AOI21_X1 U14666 ( .B1(n12342), .B2(n12341), .A(n12358), .ZN(n12357) );
  INV_X1 U14667 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12740) );
  OAI21_X1 U14668 ( .B1(n12345), .B2(P3_REG1_REG_17__SCAN_IN), .A(n12372), 
        .ZN(n12346) );
  NAND2_X1 U14669 ( .A1(n14809), .A2(n12346), .ZN(n12348) );
  OAI211_X1 U14670 ( .C1(n12349), .C2(n14797), .A(n12348), .B(n12347), .ZN(
        n12355) );
  AOI21_X1 U14671 ( .B1(n12351), .B2(n14222), .A(n12350), .ZN(n12353) );
  MUX2_X1 U14672 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n8117), .Z(n12366) );
  XNOR2_X1 U14673 ( .A(n12366), .B(n14210), .ZN(n12352) );
  NOR2_X1 U14674 ( .A1(n12353), .A2(n12352), .ZN(n12365) );
  AOI211_X1 U14675 ( .C1(n12353), .C2(n12352), .A(n14781), .B(n12365), .ZN(
        n12354) );
  AOI211_X1 U14676 ( .C1(n14801), .C2(n12359), .A(n12355), .B(n12354), .ZN(
        n12356) );
  OAI21_X1 U14677 ( .B1(n12357), .B2(n14815), .A(n12356), .ZN(P3_U3199) );
  INV_X1 U14678 ( .A(n12358), .ZN(n12363) );
  OR2_X1 U14679 ( .A1(n12360), .A2(n12359), .ZN(n12362) );
  NAND2_X1 U14680 ( .A1(n14230), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12383) );
  OAI21_X1 U14681 ( .B1(n14230), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12383), 
        .ZN(n12361) );
  AND3_X1 U14682 ( .A1(n12363), .A2(n12362), .A3(n12361), .ZN(n12364) );
  NOR2_X1 U14683 ( .A1(n12385), .A2(n12364), .ZN(n12382) );
  INV_X1 U14684 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12367) );
  INV_X1 U14685 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12732) );
  MUX2_X1 U14686 ( .A(n12367), .B(n12732), .S(n8117), .Z(n12368) );
  OAI21_X1 U14687 ( .B1(n12369), .B2(n12368), .A(n12388), .ZN(n12380) );
  NAND2_X1 U14688 ( .A1(n14210), .A2(n12370), .ZN(n12373) );
  XNOR2_X1 U14689 ( .A(n14230), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12371) );
  AOI21_X1 U14690 ( .B1(n12373), .B2(n12372), .A(n12371), .ZN(n12394) );
  INV_X1 U14691 ( .A(n12394), .ZN(n12375) );
  NAND3_X1 U14692 ( .A1(n12373), .A2(n12372), .A3(n12371), .ZN(n12374) );
  AOI21_X1 U14693 ( .B1(n12375), .B2(n12374), .A(n12399), .ZN(n12376) );
  OAI21_X1 U14694 ( .B1(n14230), .B2(n12393), .A(n12378), .ZN(n12379) );
  AOI21_X1 U14695 ( .B1(n12380), .B2(n14810), .A(n12379), .ZN(n12381) );
  OAI21_X1 U14696 ( .B1(n12382), .B2(n14815), .A(n12381), .ZN(P3_U3200) );
  XNOR2_X1 U14697 ( .A(n12392), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12389) );
  INV_X1 U14698 ( .A(n12383), .ZN(n12384) );
  INV_X1 U14699 ( .A(n12386), .ZN(n12387) );
  XNOR2_X1 U14700 ( .A(n12392), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12395) );
  MUX2_X1 U14701 ( .A(n12389), .B(n12395), .S(n8117), .Z(n12390) );
  NOR2_X1 U14702 ( .A1(n12393), .A2(n12392), .ZN(n12400) );
  INV_X1 U14703 ( .A(n12395), .ZN(n12396) );
  NAND2_X1 U14704 ( .A1(n14799), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12398) );
  INV_X1 U14705 ( .A(P3_B_REG_SCAN_IN), .ZN(n12403) );
  NOR2_X1 U14706 ( .A1(n8119), .A2(n12403), .ZN(n12404) );
  NOR2_X1 U14707 ( .A1(n14915), .A2(n12404), .ZN(n12462) );
  INV_X1 U14708 ( .A(n12462), .ZN(n12405) );
  NOR2_X1 U14709 ( .A1(n12406), .A2(n12405), .ZN(n14297) );
  NOR2_X1 U14710 ( .A1(n12407), .A2(n14910), .ZN(n12468) );
  AOI21_X1 U14711 ( .B1(n14297), .B2(n14927), .A(n12468), .ZN(n14270) );
  NAND2_X1 U14712 ( .A1(n14865), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12408) );
  OAI211_X1 U14713 ( .C1(n12754), .C2(n12677), .A(n14270), .B(n12408), .ZN(
        P3_U3202) );
  XNOR2_X1 U14714 ( .A(n12409), .B(n12457), .ZN(n12687) );
  NAND2_X1 U14715 ( .A1(n14272), .A2(n12410), .ZN(n12411) );
  AND2_X1 U14716 ( .A1(n12413), .A2(n12668), .ZN(n12414) );
  NAND2_X1 U14717 ( .A1(n12415), .A2(n14273), .ZN(n12615) );
  NAND2_X1 U14718 ( .A1(n12417), .A2(n12416), .ZN(n12419) );
  INV_X1 U14719 ( .A(n12419), .ZN(n12418) );
  OR2_X1 U14720 ( .A1(n12418), .A2(n12634), .ZN(n12425) );
  INV_X1 U14721 ( .A(n12425), .ZN(n12421) );
  NAND2_X1 U14722 ( .A1(n12424), .A2(n12667), .ZN(n12632) );
  AND2_X1 U14723 ( .A1(n12632), .A2(n12419), .ZN(n12420) );
  AND2_X1 U14724 ( .A1(n12615), .A2(n12423), .ZN(n12422) );
  INV_X1 U14725 ( .A(n12423), .ZN(n12427) );
  OR2_X1 U14726 ( .A1(n12424), .A2(n12667), .ZN(n12631) );
  AND2_X1 U14727 ( .A1(n12631), .A2(n12425), .ZN(n12616) );
  AND2_X1 U14728 ( .A1(n12616), .A2(n12619), .ZN(n12426) );
  NAND2_X1 U14729 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  INV_X1 U14730 ( .A(n12598), .ZN(n12432) );
  OR2_X1 U14731 ( .A1(n12609), .A2(n12589), .ZN(n12433) );
  OR2_X1 U14732 ( .A1(n12782), .A2(n12604), .ZN(n12434) );
  NAND2_X1 U14733 ( .A1(n12587), .A2(n12434), .ZN(n12573) );
  NAND2_X1 U14734 ( .A1(n12721), .A2(n12588), .ZN(n12435) );
  OR2_X1 U14735 ( .A1(n12562), .A2(n12575), .ZN(n12436) );
  NAND2_X1 U14736 ( .A1(n12437), .A2(n12436), .ZN(n12546) );
  NOR2_X1 U14737 ( .A1(n12714), .A2(n12535), .ZN(n12438) );
  INV_X1 U14738 ( .A(n12714), .ZN(n12553) );
  NAND2_X1 U14739 ( .A1(n12533), .A2(n12439), .ZN(n12441) );
  NAND2_X1 U14740 ( .A1(n12709), .A2(n12547), .ZN(n12440) );
  NAND2_X1 U14741 ( .A1(n12441), .A2(n12440), .ZN(n12521) );
  OR2_X1 U14742 ( .A1(n12443), .A2(n12536), .ZN(n12442) );
  NAND2_X1 U14743 ( .A1(n12521), .A2(n12442), .ZN(n12445) );
  NAND2_X1 U14744 ( .A1(n12443), .A2(n12536), .ZN(n12444) );
  NAND2_X1 U14745 ( .A1(n12445), .A2(n12444), .ZN(n12511) );
  NAND2_X1 U14746 ( .A1(n12511), .A2(n12446), .ZN(n12449) );
  NAND2_X1 U14747 ( .A1(n12699), .A2(n12447), .ZN(n12448) );
  NAND2_X1 U14748 ( .A1(n12449), .A2(n12448), .ZN(n12500) );
  OR2_X1 U14749 ( .A1(n12507), .A2(n12512), .ZN(n12450) );
  NAND2_X1 U14750 ( .A1(n12484), .A2(n12451), .ZN(n12455) );
  OR2_X1 U14751 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  NAND2_X1 U14752 ( .A1(n12479), .A2(n12460), .ZN(n12456) );
  XNOR2_X1 U14753 ( .A(n12458), .B(n12457), .ZN(n12459) );
  NAND2_X1 U14754 ( .A1(n12459), .A2(n14920), .ZN(n12464) );
  NAND2_X1 U14755 ( .A1(n12683), .A2(n14927), .ZN(n12470) );
  NAND2_X1 U14756 ( .A1(n12465), .A2(n14907), .ZN(n12686) );
  NOR2_X1 U14757 ( .A1(n12686), .A2(n12466), .ZN(n12467) );
  AOI211_X1 U14758 ( .C1(n14865), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12468), 
        .B(n12467), .ZN(n12469) );
  OAI211_X1 U14759 ( .C1(n12687), .C2(n12583), .A(n12470), .B(n12469), .ZN(
        P3_U3204) );
  AOI21_X1 U14760 ( .B1(n12471), .B2(n12477), .A(n14877), .ZN(n12475) );
  OAI22_X1 U14761 ( .A1(n12473), .A2(n14915), .B1(n12502), .B2(n14917), .ZN(
        n12474) );
  AOI21_X1 U14762 ( .B1(n12475), .B2(n12472), .A(n12474), .ZN(n12689) );
  NAND2_X1 U14763 ( .A1(n12491), .A2(n12476), .ZN(n12478) );
  XNOR2_X1 U14764 ( .A(n12478), .B(n12477), .ZN(n12688) );
  INV_X1 U14765 ( .A(n12479), .ZN(n12758) );
  AOI22_X1 U14766 ( .A1(n14865), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n12480), 
        .B2(n14901), .ZN(n12481) );
  OAI21_X1 U14767 ( .B1(n12758), .B2(n12677), .A(n12481), .ZN(n12482) );
  AOI21_X1 U14768 ( .B1(n12688), .B2(n14281), .A(n12482), .ZN(n12483) );
  OAI21_X1 U14769 ( .B1(n12689), .B2(n14865), .A(n12483), .ZN(P3_U3205) );
  XNOR2_X1 U14770 ( .A(n12484), .B(n12492), .ZN(n12490) );
  NOR2_X1 U14771 ( .A1(n12486), .A2(n14917), .ZN(n12487) );
  INV_X1 U14772 ( .A(n12693), .ZN(n12498) );
  OAI21_X1 U14773 ( .B1(n12493), .B2(n12492), .A(n12491), .ZN(n12692) );
  AOI22_X1 U14774 ( .A1(n14865), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n14901), 
        .B2(n12494), .ZN(n12495) );
  OAI21_X1 U14775 ( .B1(n12762), .B2(n12677), .A(n12495), .ZN(n12496) );
  AOI21_X1 U14776 ( .B1(n12692), .B2(n14281), .A(n12496), .ZN(n12497) );
  OAI21_X1 U14777 ( .B1(n12498), .B2(n14865), .A(n12497), .ZN(P3_U3206) );
  XNOR2_X1 U14778 ( .A(n12499), .B(n12501), .ZN(n12696) );
  XOR2_X1 U14779 ( .A(n12501), .B(n12500), .Z(n12505) );
  OAI22_X1 U14780 ( .A1(n12502), .A2(n14915), .B1(n12526), .B2(n14917), .ZN(
        n12503) );
  AOI21_X1 U14781 ( .B1(n12696), .B2(n14875), .A(n12503), .ZN(n12504) );
  OAI21_X1 U14782 ( .B1(n12505), .B2(n14877), .A(n12504), .ZN(n12695) );
  AOI21_X1 U14783 ( .B1(n14926), .B2(n12696), .A(n12695), .ZN(n12510) );
  AOI22_X1 U14784 ( .A1(n14865), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n14901), 
        .B2(n12506), .ZN(n12509) );
  NAND2_X1 U14785 ( .A1(n12507), .A2(n14268), .ZN(n12508) );
  OAI211_X1 U14786 ( .C1(n12510), .C2(n14865), .A(n12509), .B(n12508), .ZN(
        P3_U3207) );
  XNOR2_X1 U14787 ( .A(n12511), .B(n12514), .ZN(n12513) );
  AOI222_X1 U14788 ( .A1(n14920), .A2(n12513), .B1(n12512), .B2(n14889), .C1(
        n12536), .C2(n14892), .ZN(n12702) );
  XNOR2_X1 U14789 ( .A(n12515), .B(n12514), .ZN(n12700) );
  AOI22_X1 U14790 ( .A1(n14865), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n14901), 
        .B2(n12516), .ZN(n12517) );
  OAI21_X1 U14791 ( .B1(n12518), .B2(n12677), .A(n12517), .ZN(n12519) );
  AOI21_X1 U14792 ( .B1(n12700), .B2(n14281), .A(n12519), .ZN(n12520) );
  OAI21_X1 U14793 ( .B1(n12702), .B2(n14865), .A(n12520), .ZN(P3_U3208) );
  XNOR2_X1 U14794 ( .A(n12522), .B(n12523), .ZN(n12524) );
  OAI222_X1 U14795 ( .A1(n14915), .A2(n12526), .B1(n14917), .B2(n12525), .C1(
        n12524), .C2(n14877), .ZN(n12703) );
  INV_X1 U14796 ( .A(n12703), .ZN(n12532) );
  OAI21_X1 U14797 ( .B1(n6528), .B2(n7823), .A(n12527), .ZN(n12704) );
  AOI22_X1 U14798 ( .A1(n14865), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n14901), 
        .B2(n12528), .ZN(n12529) );
  OAI21_X1 U14799 ( .B1(n12771), .B2(n12677), .A(n12529), .ZN(n12530) );
  AOI21_X1 U14800 ( .B1(n12704), .B2(n14281), .A(n12530), .ZN(n12531) );
  OAI21_X1 U14801 ( .B1(n12532), .B2(n14865), .A(n12531), .ZN(P3_U3209) );
  XNOR2_X1 U14802 ( .A(n12533), .B(n12540), .ZN(n12534) );
  NAND2_X1 U14803 ( .A1(n12534), .A2(n14920), .ZN(n12538) );
  AOI22_X1 U14804 ( .A1(n12536), .A2(n14889), .B1(n14892), .B2(n12535), .ZN(
        n12537) );
  NAND2_X1 U14805 ( .A1(n12538), .A2(n12537), .ZN(n12713) );
  NAND2_X1 U14806 ( .A1(n12713), .A2(n14927), .ZN(n12545) );
  AOI22_X1 U14807 ( .A1(n14865), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n14901), 
        .B2(n12539), .ZN(n12544) );
  OR2_X1 U14808 ( .A1(n12541), .A2(n12540), .ZN(n12708) );
  NAND3_X1 U14809 ( .A1(n12708), .A2(n12707), .A3(n14281), .ZN(n12543) );
  NAND2_X1 U14810 ( .A1(n12709), .A2(n14268), .ZN(n12542) );
  NAND4_X1 U14811 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        P3_U3210) );
  XOR2_X1 U14812 ( .A(n12546), .B(n12549), .Z(n12548) );
  AOI222_X1 U14813 ( .A1(n14920), .A2(n12548), .B1(n12575), .B2(n14892), .C1(
        n12547), .C2(n14889), .ZN(n12717) );
  XOR2_X1 U14814 ( .A(n12550), .B(n12549), .Z(n12715) );
  AOI22_X1 U14815 ( .A1(n14865), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14901), 
        .B2(n12551), .ZN(n12552) );
  OAI21_X1 U14816 ( .B1(n12553), .B2(n12677), .A(n12552), .ZN(n12554) );
  AOI21_X1 U14817 ( .B1(n12715), .B2(n14281), .A(n12554), .ZN(n12555) );
  OAI21_X1 U14818 ( .B1(n12717), .B2(n14865), .A(n12555), .ZN(P3_U3211) );
  XOR2_X1 U14819 ( .A(n12560), .B(n12556), .Z(n12557) );
  OAI222_X1 U14820 ( .A1(n14917), .A2(n12559), .B1(n14915), .B2(n12558), .C1(
        n14877), .C2(n12557), .ZN(n12718) );
  INV_X1 U14821 ( .A(n12718), .ZN(n12567) );
  XOR2_X1 U14822 ( .A(n12561), .B(n12560), .Z(n12719) );
  INV_X1 U14823 ( .A(n12562), .ZN(n12777) );
  AOI22_X1 U14824 ( .A1(n14865), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14901), 
        .B2(n12563), .ZN(n12564) );
  OAI21_X1 U14825 ( .B1(n12777), .B2(n12677), .A(n12564), .ZN(n12565) );
  AOI21_X1 U14826 ( .B1(n12719), .B2(n14281), .A(n12565), .ZN(n12566) );
  OAI21_X1 U14827 ( .B1(n12567), .B2(n14865), .A(n12566), .ZN(P3_U3212) );
  NAND2_X1 U14828 ( .A1(n12569), .A2(n12568), .ZN(n12570) );
  NAND2_X1 U14829 ( .A1(n12571), .A2(n12570), .ZN(n12724) );
  XNOR2_X1 U14830 ( .A(n12573), .B(n12572), .ZN(n12576) );
  AOI222_X1 U14831 ( .A1(n14920), .A2(n12576), .B1(n12575), .B2(n14889), .C1(
        n12574), .C2(n14892), .ZN(n12723) );
  OR2_X1 U14832 ( .A1(n12723), .A2(n14865), .ZN(n12582) );
  INV_X1 U14833 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12579) );
  INV_X1 U14834 ( .A(n12577), .ZN(n12578) );
  OAI22_X1 U14835 ( .A1(n14927), .A2(n12579), .B1(n12578), .B2(n14910), .ZN(
        n12580) );
  AOI21_X1 U14836 ( .B1(n12721), .B2(n14268), .A(n12580), .ZN(n12581) );
  OAI211_X1 U14837 ( .C1(n12724), .C2(n12583), .A(n12582), .B(n12581), .ZN(
        P3_U3213) );
  NAND2_X1 U14838 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  NAND3_X1 U14839 ( .A1(n12587), .A2(n14920), .A3(n12586), .ZN(n12591) );
  AOI22_X1 U14840 ( .A1(n12589), .A2(n14892), .B1(n14889), .B2(n12588), .ZN(
        n12590) );
  XNOR2_X1 U14841 ( .A(n12593), .B(n12592), .ZN(n12725) );
  AOI22_X1 U14842 ( .A1(n14865), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14901), 
        .B2(n12594), .ZN(n12595) );
  OAI21_X1 U14843 ( .B1(n12782), .B2(n12677), .A(n12595), .ZN(n12596) );
  AOI21_X1 U14844 ( .B1(n12725), .B2(n14281), .A(n12596), .ZN(n12597) );
  OAI21_X1 U14845 ( .B1(n12727), .B2(n14865), .A(n12597), .ZN(P3_U3214) );
  INV_X1 U14846 ( .A(n12599), .ZN(n12600) );
  AOI21_X1 U14847 ( .B1(n12602), .B2(n12601), .A(n12600), .ZN(n12603) );
  OAI222_X1 U14848 ( .A1(n14917), .A2(n12637), .B1(n14915), .B2(n12604), .C1(
        n14877), .C2(n12603), .ZN(n12730) );
  INV_X1 U14849 ( .A(n12730), .ZN(n12614) );
  INV_X1 U14850 ( .A(n12605), .ZN(n12606) );
  AOI21_X1 U14851 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12731) );
  INV_X1 U14852 ( .A(n12609), .ZN(n12786) );
  AOI22_X1 U14853 ( .A1(n14865), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14901), 
        .B2(n12610), .ZN(n12611) );
  OAI21_X1 U14854 ( .B1(n12786), .B2(n12677), .A(n12611), .ZN(n12612) );
  AOI21_X1 U14855 ( .B1(n12731), .B2(n14281), .A(n12612), .ZN(n12613) );
  OAI21_X1 U14856 ( .B1(n12614), .B2(n14865), .A(n12613), .ZN(P3_U3215) );
  NAND2_X1 U14857 ( .A1(n6462), .A2(n12615), .ZN(n12648) );
  NAND2_X1 U14858 ( .A1(n12648), .A2(n12616), .ZN(n12618) );
  NAND2_X1 U14859 ( .A1(n12618), .A2(n12617), .ZN(n12620) );
  XNOR2_X1 U14860 ( .A(n12620), .B(n12619), .ZN(n12621) );
  OAI222_X1 U14861 ( .A1(n14917), .A2(n12651), .B1(n14915), .B2(n12622), .C1(
        n12621), .C2(n14877), .ZN(n12734) );
  INV_X1 U14862 ( .A(n12734), .ZN(n12630) );
  OAI21_X1 U14863 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n12735) );
  AOI22_X1 U14864 ( .A1(n14865), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14901), 
        .B2(n12626), .ZN(n12627) );
  OAI21_X1 U14865 ( .B1(n12790), .B2(n12677), .A(n12627), .ZN(n12628) );
  AOI21_X1 U14866 ( .B1(n12735), .B2(n14281), .A(n12628), .ZN(n12629) );
  OAI21_X1 U14867 ( .B1(n12630), .B2(n14865), .A(n12629), .ZN(P3_U3216) );
  NAND2_X1 U14868 ( .A1(n12648), .A2(n12631), .ZN(n12633) );
  NAND2_X1 U14869 ( .A1(n12633), .A2(n12632), .ZN(n12635) );
  XNOR2_X1 U14870 ( .A(n12635), .B(n12634), .ZN(n12636) );
  OAI222_X1 U14871 ( .A1(n14917), .A2(n12638), .B1(n14915), .B2(n12637), .C1(
        n12636), .C2(n14877), .ZN(n12738) );
  INV_X1 U14872 ( .A(n12738), .ZN(n12647) );
  OR2_X1 U14873 ( .A1(n12672), .A2(n12639), .ZN(n12654) );
  NAND2_X1 U14874 ( .A1(n12654), .A2(n12640), .ZN(n12642) );
  XNOR2_X1 U14875 ( .A(n12642), .B(n12641), .ZN(n12739) );
  AOI22_X1 U14876 ( .A1(n14865), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14901), 
        .B2(n12643), .ZN(n12644) );
  OAI21_X1 U14877 ( .B1(n12794), .B2(n12677), .A(n12644), .ZN(n12645) );
  AOI21_X1 U14878 ( .B1(n12739), .B2(n14281), .A(n12645), .ZN(n12646) );
  OAI21_X1 U14879 ( .B1(n12647), .B2(n14865), .A(n12646), .ZN(P3_U3217) );
  XOR2_X1 U14880 ( .A(n12649), .B(n12648), .Z(n12650) );
  OAI222_X1 U14881 ( .A1(n14917), .A2(n12652), .B1(n14915), .B2(n12651), .C1(
        n14877), .C2(n12650), .ZN(n12742) );
  INV_X1 U14882 ( .A(n12742), .ZN(n12663) );
  AND2_X1 U14883 ( .A1(n12654), .A2(n12653), .ZN(n12658) );
  OR2_X1 U14884 ( .A1(n12672), .A2(n12671), .ZN(n12674) );
  NAND3_X1 U14885 ( .A1(n12674), .A2(n12656), .A3(n12655), .ZN(n12657) );
  NAND2_X1 U14886 ( .A1(n12658), .A2(n12657), .ZN(n12743) );
  AOI22_X1 U14887 ( .A1(n14865), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14901), 
        .B2(n12659), .ZN(n12660) );
  OAI21_X1 U14888 ( .B1(n12677), .B2(n12797), .A(n12660), .ZN(n12661) );
  AOI21_X1 U14889 ( .B1(n12743), .B2(n14281), .A(n12661), .ZN(n12662) );
  OAI21_X1 U14890 ( .B1(n12663), .B2(n14865), .A(n12662), .ZN(P3_U3218) );
  NAND2_X1 U14891 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  NAND3_X1 U14892 ( .A1(n6462), .A2(n14920), .A3(n12666), .ZN(n12670) );
  AOI22_X1 U14893 ( .A1(n14892), .A2(n12668), .B1(n12667), .B2(n14889), .ZN(
        n12669) );
  NAND2_X1 U14894 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  NAND2_X1 U14895 ( .A1(n12674), .A2(n12673), .ZN(n12746) );
  AOI22_X1 U14896 ( .A1(n14865), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14901), 
        .B2(n12675), .ZN(n12676) );
  OAI21_X1 U14897 ( .B1(n12677), .B2(n12801), .A(n12676), .ZN(n12678) );
  AOI21_X1 U14898 ( .B1(n12746), .B2(n14281), .A(n12678), .ZN(n12679) );
  OAI21_X1 U14899 ( .B1(n12748), .B2(n14865), .A(n12679), .ZN(P3_U3219) );
  INV_X1 U14900 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12680) );
  NOR2_X1 U14901 ( .A1(n14993), .A2(n12680), .ZN(n12681) );
  AOI21_X1 U14902 ( .B1(n14297), .B2(n14993), .A(n12681), .ZN(n12682) );
  OAI21_X1 U14903 ( .B1(n12754), .B2(n12751), .A(n12682), .ZN(P3_U3490) );
  NAND2_X1 U14904 ( .A1(n12685), .A2(n12684), .ZN(n14955) );
  MUX2_X1 U14905 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n12755), .S(n14993), .Z(
        P3_U3488) );
  NAND2_X1 U14906 ( .A1(n12688), .A2(n14972), .ZN(n12690) );
  AND2_X1 U14907 ( .A1(n12690), .A2(n12689), .ZN(n12756) );
  MUX2_X1 U14908 ( .A(n15058), .B(n12759), .S(n14993), .Z(n12694) );
  OAI21_X1 U14909 ( .B1(n12762), .B2(n12751), .A(n12694), .ZN(P3_U3486) );
  AOI21_X1 U14910 ( .B1(n14966), .B2(n12696), .A(n12695), .ZN(n12763) );
  MUX2_X1 U14911 ( .A(n12697), .B(n12763), .S(n14993), .Z(n12698) );
  OAI21_X1 U14912 ( .B1(n12766), .B2(n12751), .A(n12698), .ZN(P3_U3485) );
  AOI22_X1 U14913 ( .A1(n12700), .A2(n14972), .B1(n14907), .B2(n12699), .ZN(
        n12701) );
  NAND2_X1 U14914 ( .A1(n12702), .A2(n12701), .ZN(n12767) );
  MUX2_X1 U14915 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12767), .S(n14993), .Z(
        P3_U3484) );
  AOI21_X1 U14916 ( .B1(n14972), .B2(n12704), .A(n12703), .ZN(n12768) );
  MUX2_X1 U14917 ( .A(n12705), .B(n12768), .S(n14993), .Z(n12706) );
  OAI21_X1 U14918 ( .B1(n12771), .B2(n12751), .A(n12706), .ZN(P3_U3483) );
  NAND3_X1 U14919 ( .A1(n12708), .A2(n12707), .A3(n14972), .ZN(n12711) );
  NAND2_X1 U14920 ( .A1(n12709), .A2(n14907), .ZN(n12710) );
  NAND2_X1 U14921 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  MUX2_X1 U14922 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12772), .S(n14993), .Z(
        P3_U3482) );
  AOI22_X1 U14923 ( .A1(n12715), .A2(n14972), .B1(n14907), .B2(n12714), .ZN(
        n12716) );
  NAND2_X1 U14924 ( .A1(n12717), .A2(n12716), .ZN(n12773) );
  MUX2_X1 U14925 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12773), .S(n14993), .Z(
        P3_U3481) );
  INV_X1 U14926 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n15069) );
  AOI21_X1 U14927 ( .B1(n12719), .B2(n14972), .A(n12718), .ZN(n12774) );
  MUX2_X1 U14928 ( .A(n15069), .B(n12774), .S(n14993), .Z(n12720) );
  OAI21_X1 U14929 ( .B1(n12777), .B2(n12751), .A(n12720), .ZN(P3_U3480) );
  NAND2_X1 U14930 ( .A1(n12721), .A2(n14907), .ZN(n12722) );
  OAI211_X1 U14931 ( .C1(n14305), .C2(n12724), .A(n12723), .B(n12722), .ZN(
        n12778) );
  MUX2_X1 U14932 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12778), .S(n14993), .Z(
        P3_U3479) );
  NAND2_X1 U14933 ( .A1(n12725), .A2(n14972), .ZN(n12726) );
  NAND2_X1 U14934 ( .A1(n12727), .A2(n12726), .ZN(n12779) );
  MUX2_X1 U14935 ( .A(n12779), .B(P3_REG1_REG_19__SCAN_IN), .S(n14990), .Z(
        n12728) );
  INV_X1 U14936 ( .A(n12728), .ZN(n12729) );
  OAI21_X1 U14937 ( .B1(n12751), .B2(n12782), .A(n12729), .ZN(P3_U3478) );
  AOI21_X1 U14938 ( .B1(n12731), .B2(n14972), .A(n12730), .ZN(n12783) );
  MUX2_X1 U14939 ( .A(n12732), .B(n12783), .S(n14993), .Z(n12733) );
  OAI21_X1 U14940 ( .B1(n12786), .B2(n12751), .A(n12733), .ZN(P3_U3477) );
  INV_X1 U14941 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12736) );
  AOI21_X1 U14942 ( .B1(n14972), .B2(n12735), .A(n12734), .ZN(n12787) );
  MUX2_X1 U14943 ( .A(n12736), .B(n12787), .S(n14993), .Z(n12737) );
  OAI21_X1 U14944 ( .B1(n12790), .B2(n12751), .A(n12737), .ZN(P3_U3476) );
  AOI21_X1 U14945 ( .B1(n12739), .B2(n14972), .A(n12738), .ZN(n12791) );
  MUX2_X1 U14946 ( .A(n12740), .B(n12791), .S(n14993), .Z(n12741) );
  OAI21_X1 U14947 ( .B1(n12794), .B2(n12751), .A(n12741), .ZN(P3_U3475) );
  AOI21_X1 U14948 ( .B1(n14972), .B2(n12743), .A(n12742), .ZN(n12795) );
  MUX2_X1 U14949 ( .A(n12744), .B(n12795), .S(n14993), .Z(n12745) );
  OAI21_X1 U14950 ( .B1(n12797), .B2(n12751), .A(n12745), .ZN(P3_U3474) );
  NAND2_X1 U14951 ( .A1(n12746), .A2(n14972), .ZN(n12747) );
  INV_X1 U14952 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12749) );
  MUX2_X1 U14953 ( .A(n12799), .B(n12749), .S(n14990), .Z(n12750) );
  OAI21_X1 U14954 ( .B1(n12751), .B2(n12801), .A(n12750), .ZN(P3_U3473) );
  NAND2_X1 U14955 ( .A1(n14973), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U14956 ( .A1(n14297), .A2(n14975), .ZN(n12752) );
  OAI211_X1 U14957 ( .C1(n12754), .C2(n12802), .A(n12753), .B(n12752), .ZN(
        P3_U3458) );
  INV_X1 U14958 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12757) );
  INV_X1 U14959 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12760) );
  MUX2_X1 U14960 ( .A(n12760), .B(n12759), .S(n14975), .Z(n12761) );
  OAI21_X1 U14961 ( .B1(n12762), .B2(n12802), .A(n12761), .ZN(P3_U3454) );
  INV_X1 U14962 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12764) );
  MUX2_X1 U14963 ( .A(n12764), .B(n12763), .S(n14975), .Z(n12765) );
  OAI21_X1 U14964 ( .B1(n12766), .B2(n12802), .A(n12765), .ZN(P3_U3453) );
  MUX2_X1 U14965 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12767), .S(n14975), .Z(
        P3_U3452) );
  INV_X1 U14966 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12769) );
  MUX2_X1 U14967 ( .A(n12769), .B(n12768), .S(n14975), .Z(n12770) );
  OAI21_X1 U14968 ( .B1(n12771), .B2(n12802), .A(n12770), .ZN(P3_U3451) );
  MUX2_X1 U14969 ( .A(n12772), .B(P3_REG0_REG_23__SCAN_IN), .S(n14973), .Z(
        P3_U3450) );
  MUX2_X1 U14970 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12773), .S(n14975), .Z(
        P3_U3449) );
  INV_X1 U14971 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12775) );
  MUX2_X1 U14972 ( .A(n12775), .B(n12774), .S(n14975), .Z(n12776) );
  OAI21_X1 U14973 ( .B1(n12777), .B2(n12802), .A(n12776), .ZN(P3_U3448) );
  MUX2_X1 U14974 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12778), .S(n14975), .Z(
        P3_U3447) );
  MUX2_X1 U14975 ( .A(n12779), .B(P3_REG0_REG_19__SCAN_IN), .S(n14973), .Z(
        n12780) );
  INV_X1 U14976 ( .A(n12780), .ZN(n12781) );
  OAI21_X1 U14977 ( .B1(n12802), .B2(n12782), .A(n12781), .ZN(P3_U3446) );
  INV_X1 U14978 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12784) );
  MUX2_X1 U14979 ( .A(n12784), .B(n12783), .S(n14975), .Z(n12785) );
  OAI21_X1 U14980 ( .B1(n12786), .B2(n12802), .A(n12785), .ZN(P3_U3444) );
  INV_X1 U14981 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12788) );
  MUX2_X1 U14982 ( .A(n12788), .B(n12787), .S(n14975), .Z(n12789) );
  OAI21_X1 U14983 ( .B1(n12790), .B2(n12802), .A(n12789), .ZN(P3_U3441) );
  INV_X1 U14984 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12792) );
  MUX2_X1 U14985 ( .A(n12792), .B(n12791), .S(n14975), .Z(n12793) );
  OAI21_X1 U14986 ( .B1(n12794), .B2(n12802), .A(n12793), .ZN(P3_U3438) );
  INV_X1 U14987 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n15041) );
  MUX2_X1 U14988 ( .A(n15041), .B(n12795), .S(n14975), .Z(n12796) );
  OAI21_X1 U14989 ( .B1(n12797), .B2(n12802), .A(n12796), .ZN(P3_U3435) );
  INV_X1 U14990 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U14991 ( .A(n12799), .B(n12798), .S(n14973), .Z(n12800) );
  OAI21_X1 U14992 ( .B1(n12802), .B2(n12801), .A(n12800), .ZN(P3_U3432) );
  MUX2_X1 U14993 ( .A(n12804), .B(P3_D_REG_1__SCAN_IN), .S(n12803), .Z(
        P3_U3377) );
  MUX2_X1 U14994 ( .A(P3_D_REG_0__SCAN_IN), .B(n12806), .S(n12805), .Z(
        P3_U3376) );
  NAND3_X1 U14995 ( .A1(n12807), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12809) );
  OAI22_X1 U14996 ( .A1(n12810), .A2(n12809), .B1(n12808), .B2(n12817), .ZN(
        n12811) );
  AOI21_X1 U14997 ( .B1(n12812), .B2(n14227), .A(n12811), .ZN(n12813) );
  INV_X1 U14998 ( .A(n12813), .ZN(P3_U3264) );
  INV_X1 U14999 ( .A(n12814), .ZN(n12815) );
  OAI222_X1 U15000 ( .A1(n12817), .A2(n12816), .B1(n12821), .B2(n12815), .C1(
        P3_U3151), .C2(n7420), .ZN(P3_U3266) );
  INV_X1 U15001 ( .A(n12818), .ZN(n12820) );
  OAI222_X1 U15002 ( .A1(n12821), .A2(n12820), .B1(n8119), .B2(P3_U3151), .C1(
        n12819), .C2(n12817), .ZN(P3_U3267) );
  INV_X1 U15003 ( .A(n12822), .ZN(n12828) );
  AOI22_X1 U15004 ( .A1(n12823), .A2(n6591), .B1(n12934), .B2(n12955), .ZN(
        n12827) );
  AOI22_X1 U15005 ( .A1(n12956), .A2(n12906), .B1(n6433), .B2(n12954), .ZN(
        n13300) );
  AOI22_X1 U15006 ( .A1(n13160), .A2(n12898), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12824) );
  OAI21_X1 U15007 ( .B1(n13300), .B2(n12908), .A(n12824), .ZN(n12825) );
  AOI21_X1 U15008 ( .B1(n13159), .B2(n12943), .A(n12825), .ZN(n12826) );
  OAI21_X1 U15009 ( .B1(n12828), .B2(n12827), .A(n12826), .ZN(P2_U3188) );
  INV_X1 U15010 ( .A(n13326), .ZN(n13227) );
  OAI21_X1 U15011 ( .B1(n12831), .B2(n12830), .A(n12829), .ZN(n12832) );
  NAND2_X1 U15012 ( .A1(n12832), .A2(n6591), .ZN(n12836) );
  NAND2_X1 U15013 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13054)
         );
  INV_X1 U15014 ( .A(n13054), .ZN(n12834) );
  AOI22_X1 U15015 ( .A1(n12958), .A2(n6433), .B1(n12906), .B2(n12960), .ZN(
        n13219) );
  NOR2_X1 U15016 ( .A1(n13219), .A2(n12908), .ZN(n12833) );
  AOI211_X1 U15017 ( .C1(n12898), .C2(n13224), .A(n12834), .B(n12833), .ZN(
        n12835) );
  OAI211_X1 U15018 ( .C1(n13227), .C2(n12924), .A(n12836), .B(n12835), .ZN(
        P2_U3191) );
  INV_X1 U15019 ( .A(n12837), .ZN(n12838) );
  NAND2_X1 U15020 ( .A1(n12950), .A2(n13221), .ZN(n12839) );
  XNOR2_X1 U15021 ( .A(n12840), .B(n12839), .ZN(n12841) );
  XNOR2_X1 U15022 ( .A(n13077), .B(n12841), .ZN(n12842) );
  XNOR2_X1 U15023 ( .A(n12843), .B(n12842), .ZN(n12848) );
  AOI22_X1 U15024 ( .A1(n12906), .A2(n12951), .B1(n12949), .B2(n6433), .ZN(
        n13072) );
  INV_X1 U15025 ( .A(n13080), .ZN(n12844) );
  AOI22_X1 U15026 ( .A1(n12898), .A2(n12844), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12845) );
  OAI21_X1 U15027 ( .B1(n12908), .B2(n13072), .A(n12845), .ZN(n12846) );
  AOI21_X1 U15028 ( .B1(n13266), .B2(n12943), .A(n12846), .ZN(n12847) );
  OAI21_X1 U15029 ( .B1(n12848), .B2(n12928), .A(n12847), .ZN(P2_U3192) );
  OAI211_X1 U15030 ( .C1(n12851), .C2(n12850), .A(n12849), .B(n6591), .ZN(
        n12857) );
  NAND2_X1 U15031 ( .A1(n12956), .A2(n6433), .ZN(n12853) );
  NAND2_X1 U15032 ( .A1(n12958), .A2(n12906), .ZN(n12852) );
  NAND2_X1 U15033 ( .A1(n12853), .A2(n12852), .ZN(n13311) );
  OAI22_X1 U15034 ( .A1(n12940), .A2(n13192), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12854), .ZN(n12855) );
  AOI21_X1 U15035 ( .B1(n13311), .B2(n12942), .A(n12855), .ZN(n12856) );
  OAI211_X1 U15036 ( .C1(n13314), .C2(n12924), .A(n12857), .B(n12856), .ZN(
        P2_U3195) );
  NOR3_X1 U15037 ( .A1(n12860), .A2(n12859), .A3(n12858), .ZN(n12865) );
  AOI21_X1 U15038 ( .B1(n12861), .B2(n12862), .A(n12928), .ZN(n12864) );
  OAI21_X1 U15039 ( .B1(n12865), .B2(n12864), .A(n12863), .ZN(n12869) );
  NOR2_X1 U15040 ( .A1(n12940), .A2(n13128), .ZN(n12867) );
  AOI22_X1 U15041 ( .A1(n12952), .A2(n6433), .B1(n12906), .B2(n12954), .ZN(
        n13120) );
  NOR2_X1 U15042 ( .A1(n12908), .A2(n13120), .ZN(n12866) );
  AOI211_X1 U15043 ( .C1(P2_REG3_REG_25__SCAN_IN), .C2(P2_U3088), .A(n12867), 
        .B(n12866), .ZN(n12868) );
  OAI211_X1 U15044 ( .C1(n13290), .C2(n12924), .A(n12869), .B(n12868), .ZN(
        P2_U3197) );
  AOI21_X1 U15045 ( .B1(n6559), .B2(n12871), .A(n12870), .ZN(n12878) );
  NOR2_X1 U15046 ( .A1(n12908), .A2(n13334), .ZN(n12875) );
  OAI21_X1 U15047 ( .B1(n12940), .B2(n12873), .A(n12872), .ZN(n12874) );
  AOI211_X1 U15048 ( .C1(n12876), .C2(n12943), .A(n12875), .B(n12874), .ZN(
        n12877) );
  OAI21_X1 U15049 ( .B1(n12878), .B2(n12928), .A(n12877), .ZN(P2_U3200) );
  INV_X1 U15050 ( .A(n13296), .ZN(n13146) );
  OAI211_X1 U15051 ( .C1(n12880), .C2(n12879), .A(n12861), .B(n6591), .ZN(
        n12886) );
  OAI22_X1 U15052 ( .A1(n12882), .A2(n12919), .B1(n12918), .B2(n15177), .ZN(
        n13143) );
  INV_X1 U15053 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12883) );
  OAI22_X1 U15054 ( .A1(n12940), .A2(n13147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12883), .ZN(n12884) );
  AOI21_X1 U15055 ( .B1(n13143), .B2(n12942), .A(n12884), .ZN(n12885) );
  OAI211_X1 U15056 ( .C1(n13146), .C2(n12924), .A(n12886), .B(n12885), .ZN(
        P2_U3201) );
  INV_X1 U15057 ( .A(n12887), .ZN(n12889) );
  NAND2_X1 U15058 ( .A1(n12889), .A2(n12888), .ZN(n12890) );
  XNOR2_X1 U15059 ( .A(n12891), .B(n12890), .ZN(n12895) );
  AOI22_X1 U15060 ( .A1(n12957), .A2(n6433), .B1(n12906), .B2(n12959), .ZN(
        n13204) );
  AOI22_X1 U15061 ( .A1(n12898), .A2(n13210), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12892) );
  OAI21_X1 U15062 ( .B1(n13204), .B2(n12908), .A(n12892), .ZN(n12893) );
  AOI21_X1 U15063 ( .B1(n13321), .B2(n12943), .A(n12893), .ZN(n12894) );
  OAI21_X1 U15064 ( .B1(n12895), .B2(n12928), .A(n12894), .ZN(P2_U3205) );
  AOI22_X1 U15065 ( .A1(n6486), .A2(n6591), .B1(n12934), .B2(n12956), .ZN(
        n12902) );
  AND2_X1 U15066 ( .A1(n12957), .A2(n12906), .ZN(n12896) );
  AOI21_X1 U15067 ( .B1(n12955), .B2(n6433), .A(n12896), .ZN(n13170) );
  INV_X1 U15068 ( .A(n12897), .ZN(n13178) );
  AOI22_X1 U15069 ( .A1(n13178), .A2(n12898), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12899) );
  OAI21_X1 U15070 ( .B1(n13170), .B2(n12908), .A(n12899), .ZN(n12900) );
  AOI21_X1 U15071 ( .B1(n13307), .B2(n12911), .A(n12900), .ZN(n12901) );
  OAI21_X1 U15072 ( .B1(n12903), .B2(n12902), .A(n12901), .ZN(P2_U3207) );
  XNOR2_X1 U15073 ( .A(n12905), .B(n12904), .ZN(n12913) );
  AND2_X1 U15074 ( .A1(n12961), .A2(n12906), .ZN(n12907) );
  AOI21_X1 U15075 ( .B1(n12959), .B2(n6433), .A(n12907), .ZN(n13232) );
  NOR2_X1 U15076 ( .A1(n12908), .A2(n13232), .ZN(n12910) );
  NAND2_X1 U15077 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14703)
         );
  OAI21_X1 U15078 ( .B1(n12940), .B2(n13238), .A(n14703), .ZN(n12909) );
  AOI211_X1 U15079 ( .C1(n13330), .C2(n12911), .A(n12910), .B(n12909), .ZN(
        n12912) );
  OAI21_X1 U15080 ( .B1(n12913), .B2(n12928), .A(n12912), .ZN(P2_U3210) );
  NAND3_X1 U15081 ( .A1(n12914), .A2(n12934), .A3(n12953), .ZN(n12915) );
  OAI21_X1 U15082 ( .B1(n12863), .B2(n12928), .A(n12915), .ZN(n12927) );
  INV_X1 U15083 ( .A(n12916), .ZN(n12926) );
  NAND2_X1 U15084 ( .A1(n12951), .A2(n6433), .ZN(n12921) );
  OR2_X1 U15085 ( .A1(n12919), .A2(n12918), .ZN(n12920) );
  NAND2_X1 U15086 ( .A1(n12921), .A2(n12920), .ZN(n13279) );
  OAI22_X1 U15087 ( .A1(n12940), .A2(n13105), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15039), .ZN(n12922) );
  AOI21_X1 U15088 ( .B1(n12942), .B2(n13279), .A(n12922), .ZN(n12923) );
  OAI21_X1 U15089 ( .B1(n13282), .B2(n12924), .A(n12923), .ZN(n12925) );
  NAND2_X1 U15090 ( .A1(n12931), .A2(n12930), .ZN(n12933) );
  XNOR2_X1 U15091 ( .A(n12933), .B(n12932), .ZN(n12935) );
  NAND3_X1 U15092 ( .A1(n12935), .A2(n12934), .A3(n12963), .ZN(n12947) );
  INV_X1 U15093 ( .A(n12935), .ZN(n12937) );
  NAND3_X1 U15094 ( .A1(n12937), .A2(n6591), .A3(n12936), .ZN(n12946) );
  INV_X1 U15095 ( .A(n12938), .ZN(n12939) );
  OAI22_X1 U15096 ( .A1(n12940), .A2(n12939), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9384), .ZN(n12941) );
  AOI21_X1 U15097 ( .B1(n12942), .B2(n14331), .A(n12941), .ZN(n12945) );
  NAND2_X1 U15098 ( .A1(n14332), .A2(n12943), .ZN(n12944) );
  NAND4_X1 U15099 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        P2_U3213) );
  INV_X2 U15100 ( .A(P2_U3947), .ZN(n12970) );
  MUX2_X1 U15101 ( .A(n13057), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12970), .Z(
        P2_U3562) );
  MUX2_X1 U15102 ( .A(n12948), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12970), .Z(
        P2_U3561) );
  MUX2_X1 U15103 ( .A(n12949), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12970), .Z(
        P2_U3560) );
  MUX2_X1 U15104 ( .A(n12950), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12970), .Z(
        P2_U3559) );
  MUX2_X1 U15105 ( .A(n12951), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12970), .Z(
        P2_U3558) );
  MUX2_X1 U15106 ( .A(n12952), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12970), .Z(
        P2_U3557) );
  MUX2_X1 U15107 ( .A(n12953), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12970), .Z(
        P2_U3556) );
  MUX2_X1 U15108 ( .A(n12954), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12970), .Z(
        P2_U3555) );
  MUX2_X1 U15109 ( .A(n12955), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12970), .Z(
        P2_U3554) );
  MUX2_X1 U15110 ( .A(n12956), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12970), .Z(
        P2_U3553) );
  MUX2_X1 U15111 ( .A(n12957), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12970), .Z(
        P2_U3552) );
  MUX2_X1 U15112 ( .A(n12958), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12970), .Z(
        P2_U3551) );
  MUX2_X1 U15113 ( .A(n12959), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12970), .Z(
        P2_U3550) );
  MUX2_X1 U15114 ( .A(n12960), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12970), .Z(
        P2_U3549) );
  MUX2_X1 U15115 ( .A(n12961), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12970), .Z(
        P2_U3548) );
  MUX2_X1 U15116 ( .A(n12962), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12970), .Z(
        P2_U3547) );
  MUX2_X1 U15117 ( .A(n12963), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12970), .Z(
        P2_U3546) );
  MUX2_X1 U15118 ( .A(n12964), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12970), .Z(
        P2_U3545) );
  MUX2_X1 U15119 ( .A(n12965), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12970), .Z(
        P2_U3544) );
  MUX2_X1 U15120 ( .A(n12966), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12970), .Z(
        P2_U3543) );
  MUX2_X1 U15121 ( .A(n12967), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12970), .Z(
        P2_U3542) );
  MUX2_X1 U15122 ( .A(n12968), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12970), .Z(
        P2_U3541) );
  MUX2_X1 U15123 ( .A(n12969), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12970), .Z(
        P2_U3540) );
  MUX2_X1 U15124 ( .A(n12971), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12970), .Z(
        P2_U3539) );
  MUX2_X1 U15125 ( .A(n12972), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12970), .Z(
        P2_U3538) );
  MUX2_X1 U15126 ( .A(n12973), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12970), .Z(
        P2_U3537) );
  MUX2_X1 U15127 ( .A(n12974), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12970), .Z(
        P2_U3536) );
  MUX2_X1 U15128 ( .A(n12975), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12970), .Z(
        P2_U3535) );
  MUX2_X1 U15129 ( .A(n12976), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12970), .Z(
        P2_U3534) );
  MUX2_X1 U15130 ( .A(n12977), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12970), .Z(
        P2_U3533) );
  MUX2_X1 U15131 ( .A(n12978), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12970), .Z(
        P2_U3532) );
  MUX2_X1 U15132 ( .A(n12979), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12970), .Z(
        P2_U3531) );
  NAND2_X1 U15133 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n12981) );
  AOI211_X1 U15134 ( .C1(n12982), .C2(n12981), .A(n12980), .B(n14700), .ZN(
        n12983) );
  AOI21_X1 U15135 ( .B1(n14694), .B2(n12984), .A(n12983), .ZN(n12993) );
  AOI22_X1 U15136 ( .A1(n14680), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n12992) );
  AND2_X1 U15137 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n12990) );
  MUX2_X1 U15138 ( .A(n12986), .B(P2_REG1_REG_1__SCAN_IN), .S(n12985), .Z(
        n12989) );
  INV_X1 U15139 ( .A(n12987), .ZN(n12988) );
  OAI211_X1 U15140 ( .C1(n12990), .C2(n12989), .A(n14696), .B(n12988), .ZN(
        n12991) );
  NAND3_X1 U15141 ( .A1(n12993), .A2(n12992), .A3(n12991), .ZN(P2_U3215) );
  XOR2_X1 U15142 ( .A(n12995), .B(n12994), .Z(n12996) );
  AOI22_X1 U15143 ( .A1(n12997), .A2(n14694), .B1(n14696), .B2(n12996), .ZN(
        n13003) );
  AOI22_X1 U15144 ( .A1(n14680), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n13002) );
  NAND2_X1 U15145 ( .A1(n12999), .A2(n12998), .ZN(n13000) );
  NAND3_X1 U15146 ( .A1(n14683), .A2(n13006), .A3(n13000), .ZN(n13001) );
  NAND3_X1 U15147 ( .A1(n13003), .A2(n13002), .A3(n13001), .ZN(P2_U3216) );
  AND3_X1 U15148 ( .A1(n13006), .A2(n13005), .A3(n13004), .ZN(n13007) );
  NOR3_X1 U15149 ( .A1(n14700), .A2(n13008), .A3(n13007), .ZN(n13009) );
  AOI21_X1 U15150 ( .B1(n14694), .B2(n13010), .A(n13009), .ZN(n13017) );
  AOI22_X1 U15151 ( .A1(n14680), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(P2_U3088), 
        .B2(P2_REG3_REG_3__SCAN_IN), .ZN(n13016) );
  OAI211_X1 U15152 ( .C1(n13014), .C2(n13013), .A(n14696), .B(n13012), .ZN(
        n13015) );
  NAND3_X1 U15153 ( .A1(n13017), .A2(n13016), .A3(n13015), .ZN(P2_U3217) );
  INV_X1 U15154 ( .A(n13018), .ZN(n13023) );
  NOR3_X1 U15155 ( .A1(n13021), .A2(n13020), .A3(n13019), .ZN(n13022) );
  OAI21_X1 U15156 ( .B1(n13023), .B2(n13022), .A(n14683), .ZN(n13033) );
  OAI21_X1 U15157 ( .B1(n14705), .B2(n14458), .A(n13024), .ZN(n13025) );
  AOI21_X1 U15158 ( .B1(n13026), .B2(n14694), .A(n13025), .ZN(n13032) );
  NOR2_X1 U15159 ( .A1(n13028), .A2(n13027), .ZN(n13030) );
  OAI21_X1 U15160 ( .B1(n13030), .B2(n13029), .A(n14696), .ZN(n13031) );
  NAND3_X1 U15161 ( .A1(n13033), .A2(n13032), .A3(n13031), .ZN(P2_U3226) );
  INV_X1 U15162 ( .A(n13034), .ZN(n13035) );
  NAND2_X1 U15163 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NOR2_X1 U15164 ( .A1(n14691), .A2(n13040), .ZN(n13041) );
  XNOR2_X1 U15165 ( .A(n13041), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13052) );
  INV_X1 U15166 ( .A(n13052), .ZN(n13049) );
  OAI21_X1 U15167 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(n13045) );
  XOR2_X1 U15168 ( .A(n14693), .B(n13045), .Z(n14697) );
  NAND2_X1 U15169 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14697), .ZN(n14695) );
  NAND2_X1 U15170 ( .A1(n13045), .A2(n14693), .ZN(n13046) );
  NAND2_X1 U15171 ( .A1(n14695), .A2(n13046), .ZN(n13047) );
  XNOR2_X1 U15172 ( .A(n13047), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13051) );
  AOI21_X1 U15173 ( .B1(n13051), .B2(n14696), .A(n14694), .ZN(n13048) );
  XNOR2_X1 U15174 ( .A(n13063), .B(n13059), .ZN(n13056) );
  NAND2_X1 U15175 ( .A1(n13056), .A2(n13206), .ZN(n13254) );
  NAND2_X1 U15176 ( .A1(n13058), .A2(n13057), .ZN(n13256) );
  NOR2_X1 U15177 ( .A1(n10962), .A2(n13256), .ZN(n13067) );
  INV_X1 U15178 ( .A(n13059), .ZN(n13255) );
  NOR2_X1 U15179 ( .A1(n13255), .A2(n13242), .ZN(n13060) );
  AOI211_X1 U15180 ( .C1(n13253), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13067), 
        .B(n13060), .ZN(n13061) );
  OAI21_X1 U15181 ( .B1(n13254), .B2(n13197), .A(n13061), .ZN(P2_U3234) );
  INV_X1 U15182 ( .A(n13062), .ZN(n13065) );
  INV_X1 U15183 ( .A(n13063), .ZN(n13064) );
  OAI211_X1 U15184 ( .C1(n13258), .C2(n13065), .A(n13064), .B(n13206), .ZN(
        n13257) );
  NOR2_X1 U15185 ( .A1(n13258), .A2(n13242), .ZN(n13066) );
  AOI211_X1 U15186 ( .C1(n13253), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13067), 
        .B(n13066), .ZN(n13068) );
  OAI21_X1 U15187 ( .B1(n13197), .B2(n13257), .A(n13068), .ZN(P2_U3235) );
  OAI211_X1 U15188 ( .C1(n13071), .C2(n13070), .A(n13069), .B(n14753), .ZN(
        n13073) );
  OAI21_X1 U15189 ( .B1(n13076), .B2(n13075), .A(n13074), .ZN(n13269) );
  INV_X1 U15190 ( .A(n13269), .ZN(n13085) );
  NOR2_X1 U15191 ( .A1(n13077), .A2(n13094), .ZN(n13078) );
  OAI22_X1 U15192 ( .A1(n14714), .A2(n13081), .B1(n13080), .B2(n14716), .ZN(
        n13082) );
  AOI21_X1 U15193 ( .B1(n13266), .B2(n13194), .A(n13082), .ZN(n13083) );
  OAI21_X1 U15194 ( .B1(n13264), .B2(n13197), .A(n13083), .ZN(n13084) );
  AOI21_X1 U15195 ( .B1(n13085), .B2(n13183), .A(n13084), .ZN(n13086) );
  OAI21_X1 U15196 ( .B1(n13268), .B2(n13253), .A(n13086), .ZN(P2_U3237) );
  XNOR2_X1 U15197 ( .A(n13087), .B(n13098), .ZN(n13270) );
  INV_X1 U15198 ( .A(n13270), .ZN(n13101) );
  INV_X1 U15199 ( .A(n13088), .ZN(n13089) );
  AOI22_X1 U15200 ( .A1(n14714), .A2(n13271), .B1(n13089), .B2(n13239), .ZN(
        n13090) );
  OAI21_X1 U15201 ( .B1(n13091), .B2(n14714), .A(n13090), .ZN(n13096) );
  NOR2_X1 U15202 ( .A1(n13092), .A2(n13104), .ZN(n13093) );
  NOR2_X1 U15203 ( .A1(n13275), .A2(n13197), .ZN(n13095) );
  AOI211_X1 U15204 ( .C1(n13194), .C2(n13272), .A(n13096), .B(n13095), .ZN(
        n13100) );
  NAND2_X1 U15205 ( .A1(n13098), .A2(n13097), .ZN(n13273) );
  NAND3_X1 U15206 ( .A1(n13274), .A2(n13273), .A3(n13183), .ZN(n13099) );
  OAI211_X1 U15207 ( .C1(n13101), .C2(n13115), .A(n13100), .B(n13099), .ZN(
        P2_U3238) );
  XOR2_X1 U15208 ( .A(n13102), .B(n13112), .Z(n13286) );
  NOR2_X1 U15209 ( .A1(n13282), .A2(n13126), .ZN(n13103) );
  INV_X1 U15210 ( .A(n13281), .ZN(n13110) );
  NOR2_X1 U15211 ( .A1(n14716), .A2(n13105), .ZN(n13106) );
  AOI21_X1 U15212 ( .B1(n14714), .B2(n13279), .A(n13106), .ZN(n13108) );
  NAND2_X1 U15213 ( .A1(n10962), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13107) );
  OAI211_X1 U15214 ( .C1(n13282), .C2(n13242), .A(n13108), .B(n13107), .ZN(
        n13109) );
  AOI21_X1 U15215 ( .B1(n13110), .B2(n13251), .A(n13109), .ZN(n13114) );
  XOR2_X1 U15216 ( .A(n13112), .B(n13111), .Z(n13284) );
  NAND2_X1 U15217 ( .A1(n13284), .A2(n13183), .ZN(n13113) );
  OAI211_X1 U15218 ( .C1(n13286), .C2(n13115), .A(n13114), .B(n13113), .ZN(
        P2_U3239) );
  OAI21_X1 U15219 ( .B1(n13118), .B2(n13117), .A(n13116), .ZN(n13119) );
  NAND2_X1 U15220 ( .A1(n13119), .A2(n14753), .ZN(n13121) );
  NAND2_X1 U15221 ( .A1(n13121), .A2(n13120), .ZN(n13293) );
  INV_X1 U15222 ( .A(n13293), .ZN(n13135) );
  OR2_X1 U15223 ( .A1(n13123), .A2(n13122), .ZN(n13124) );
  NAND2_X1 U15224 ( .A1(n13125), .A2(n13124), .ZN(n13288) );
  NOR2_X1 U15225 ( .A1(n13145), .A2(n13290), .ZN(n13127) );
  OAI22_X1 U15226 ( .A1(n14714), .A2(n13129), .B1(n13128), .B2(n14716), .ZN(
        n13130) );
  AOI21_X1 U15227 ( .B1(n13131), .B2(n13194), .A(n13130), .ZN(n13132) );
  OAI21_X1 U15228 ( .B1(n13289), .B2(n13197), .A(n13132), .ZN(n13133) );
  AOI21_X1 U15229 ( .B1(n13183), .B2(n13288), .A(n13133), .ZN(n13134) );
  OAI21_X1 U15230 ( .B1(n13135), .B2(n13253), .A(n13134), .ZN(P2_U3240) );
  INV_X1 U15231 ( .A(n13136), .ZN(n13137) );
  XNOR2_X1 U15232 ( .A(n13137), .B(n13139), .ZN(n13294) );
  NAND2_X1 U15233 ( .A1(n13138), .A2(n13139), .ZN(n13140) );
  AOI21_X1 U15234 ( .B1(n13141), .B2(n13140), .A(n7052), .ZN(n13142) );
  AOI211_X1 U15235 ( .C1(n13294), .C2(n13144), .A(n13143), .B(n13142), .ZN(
        n13298) );
  AOI211_X1 U15236 ( .C1(n13296), .C2(n13157), .A(n13221), .B(n13145), .ZN(
        n13295) );
  NOR2_X1 U15237 ( .A1(n13146), .A2(n13242), .ZN(n13150) );
  OAI22_X1 U15238 ( .A1(n14714), .A2(n13148), .B1(n13147), .B2(n14716), .ZN(
        n13149) );
  AOI211_X1 U15239 ( .C1(n13295), .C2(n13251), .A(n13150), .B(n13149), .ZN(
        n13153) );
  NAND2_X1 U15240 ( .A1(n13294), .A2(n13151), .ZN(n13152) );
  OAI211_X1 U15241 ( .C1(n13298), .C2(n10962), .A(n13153), .B(n13152), .ZN(
        P2_U3241) );
  XNOR2_X1 U15242 ( .A(n13154), .B(n13155), .ZN(n13305) );
  XNOR2_X1 U15243 ( .A(n13156), .B(n13155), .ZN(n13303) );
  NAND2_X1 U15244 ( .A1(n13303), .A2(n13199), .ZN(n13167) );
  AOI21_X1 U15245 ( .B1(n13159), .B2(n6558), .A(n13221), .ZN(n13158) );
  NAND2_X1 U15246 ( .A1(n13158), .A2(n13157), .ZN(n13301) );
  INV_X1 U15247 ( .A(n13301), .ZN(n13165) );
  INV_X1 U15248 ( .A(n13160), .ZN(n13161) );
  OAI22_X1 U15249 ( .A1(n13300), .A2(n13253), .B1(n13161), .B2(n14716), .ZN(
        n13162) );
  AOI21_X1 U15250 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(n13253), .A(n13162), 
        .ZN(n13163) );
  OAI21_X1 U15251 ( .B1(n11763), .B2(n13242), .A(n13163), .ZN(n13164) );
  AOI21_X1 U15252 ( .B1(n13165), .B2(n13251), .A(n13164), .ZN(n13166) );
  OAI211_X1 U15253 ( .C1(n13305), .C2(n13248), .A(n13167), .B(n13166), .ZN(
        P2_U3242) );
  OAI211_X1 U15254 ( .C1(n13169), .C2(n13173), .A(n13168), .B(n14753), .ZN(
        n13171) );
  INV_X1 U15255 ( .A(n13172), .ZN(n13176) );
  INV_X1 U15256 ( .A(n13173), .ZN(n13175) );
  OAI21_X1 U15257 ( .B1(n13176), .B2(n13175), .A(n13174), .ZN(n13310) );
  INV_X1 U15258 ( .A(n13310), .ZN(n13184) );
  INV_X1 U15259 ( .A(n13307), .ZN(n13181) );
  AOI21_X1 U15260 ( .B1(n13307), .B2(n13189), .A(n13221), .ZN(n13177) );
  AND2_X1 U15261 ( .A1(n13177), .A2(n6558), .ZN(n13306) );
  NAND2_X1 U15262 ( .A1(n13306), .A2(n13251), .ZN(n13180) );
  AOI22_X1 U15263 ( .A1(n10962), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13178), 
        .B2(n13239), .ZN(n13179) );
  OAI211_X1 U15264 ( .C1(n13181), .C2(n13242), .A(n13180), .B(n13179), .ZN(
        n13182) );
  AOI21_X1 U15265 ( .B1(n13184), .B2(n13183), .A(n13182), .ZN(n13185) );
  OAI21_X1 U15266 ( .B1(n13309), .B2(n13253), .A(n13185), .ZN(P2_U3243) );
  XNOR2_X1 U15267 ( .A(n13186), .B(n13187), .ZN(n13318) );
  XNOR2_X1 U15268 ( .A(n13188), .B(n13187), .ZN(n13316) );
  OAI211_X1 U15269 ( .C1(n13209), .C2(n13314), .A(n13206), .B(n13189), .ZN(
        n13313) );
  NAND2_X1 U15270 ( .A1(n13311), .A2(n14714), .ZN(n13191) );
  NAND2_X1 U15271 ( .A1(n10962), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13190) );
  OAI211_X1 U15272 ( .C1(n14716), .C2(n13192), .A(n13191), .B(n13190), .ZN(
        n13193) );
  AOI21_X1 U15273 ( .B1(n13195), .B2(n13194), .A(n13193), .ZN(n13196) );
  OAI21_X1 U15274 ( .B1(n13313), .B2(n13197), .A(n13196), .ZN(n13198) );
  AOI21_X1 U15275 ( .B1(n13316), .B2(n13199), .A(n13198), .ZN(n13200) );
  OAI21_X1 U15276 ( .B1(n13248), .B2(n13318), .A(n13200), .ZN(P2_U3244) );
  XNOR2_X1 U15277 ( .A(n13201), .B(n13203), .ZN(n13323) );
  AOI21_X1 U15278 ( .B1(n13203), .B2(n13202), .A(n6504), .ZN(n13205) );
  OAI21_X1 U15279 ( .B1(n13205), .B2(n7052), .A(n13204), .ZN(n13319) );
  INV_X1 U15280 ( .A(n13321), .ZN(n13213) );
  NAND2_X1 U15281 ( .A1(n13222), .A2(n13321), .ZN(n13207) );
  NAND2_X1 U15282 ( .A1(n13207), .A2(n13206), .ZN(n13208) );
  NOR2_X1 U15283 ( .A1(n13209), .A2(n13208), .ZN(n13320) );
  NAND2_X1 U15284 ( .A1(n13320), .A2(n13251), .ZN(n13212) );
  AOI22_X1 U15285 ( .A1(n10962), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13210), 
        .B2(n13239), .ZN(n13211) );
  OAI211_X1 U15286 ( .C1(n13213), .C2(n13242), .A(n13212), .B(n13211), .ZN(
        n13214) );
  AOI21_X1 U15287 ( .B1(n13319), .B2(n14714), .A(n13214), .ZN(n13215) );
  OAI21_X1 U15288 ( .B1(n13248), .B2(n13323), .A(n13215), .ZN(P2_U3245) );
  XNOR2_X1 U15289 ( .A(n13216), .B(n13217), .ZN(n13328) );
  XOR2_X1 U15290 ( .A(n13218), .B(n13217), .Z(n13220) );
  OAI21_X1 U15291 ( .B1(n13220), .B2(n7052), .A(n13219), .ZN(n13324) );
  AOI21_X1 U15292 ( .B1(n13236), .B2(n13326), .A(n13221), .ZN(n13223) );
  AND2_X1 U15293 ( .A1(n13223), .A2(n13222), .ZN(n13325) );
  NAND2_X1 U15294 ( .A1(n13325), .A2(n13251), .ZN(n13226) );
  AOI22_X1 U15295 ( .A1(n10962), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13224), 
        .B2(n13239), .ZN(n13225) );
  OAI211_X1 U15296 ( .C1(n13227), .C2(n13242), .A(n13226), .B(n13225), .ZN(
        n13228) );
  AOI21_X1 U15297 ( .B1(n13324), .B2(n14714), .A(n13228), .ZN(n13229) );
  OAI21_X1 U15298 ( .B1(n13248), .B2(n13328), .A(n13229), .ZN(P2_U3246) );
  XNOR2_X1 U15299 ( .A(n13231), .B(n13230), .ZN(n13234) );
  INV_X1 U15300 ( .A(n13232), .ZN(n13233) );
  AOI21_X1 U15301 ( .B1(n13234), .B2(n14753), .A(n13233), .ZN(n13332) );
  INV_X1 U15302 ( .A(n13236), .ZN(n13237) );
  AOI211_X1 U15303 ( .C1(n13330), .C2(n6776), .A(n13221), .B(n13237), .ZN(
        n13329) );
  INV_X1 U15304 ( .A(n13238), .ZN(n13240) );
  AOI22_X1 U15305 ( .A1(n10962), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13240), 
        .B2(n13239), .ZN(n13241) );
  OAI21_X1 U15306 ( .B1(n13243), .B2(n13242), .A(n13241), .ZN(n13250) );
  INV_X1 U15307 ( .A(n13244), .ZN(n13245) );
  AOI21_X1 U15308 ( .B1(n13247), .B2(n13246), .A(n13245), .ZN(n13333) );
  NOR2_X1 U15309 ( .A1(n13333), .A2(n13248), .ZN(n13249) );
  AOI211_X1 U15310 ( .C1(n13329), .C2(n13251), .A(n13250), .B(n13249), .ZN(
        n13252) );
  OAI21_X1 U15311 ( .B1(n13253), .B2(n13332), .A(n13252), .ZN(P2_U3247) );
  OAI211_X1 U15312 ( .C1(n13255), .C2(n14764), .A(n13254), .B(n13256), .ZN(
        n13342) );
  MUX2_X1 U15313 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13342), .S(n6436), .Z(
        P2_U3530) );
  OAI211_X1 U15314 ( .C1(n13258), .C2(n14764), .A(n13257), .B(n13256), .ZN(
        n13343) );
  MUX2_X1 U15315 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13343), .S(n6436), .Z(
        P2_U3529) );
  NAND2_X1 U15316 ( .A1(n11950), .A2(n13261), .ZN(n13262) );
  INV_X1 U15317 ( .A(n13264), .ZN(n13265) );
  AOI21_X1 U15318 ( .B1(n13261), .B2(n13266), .A(n13265), .ZN(n13267) );
  OAI211_X1 U15319 ( .C1(n14749), .C2(n13269), .A(n13268), .B(n13267), .ZN(
        n13345) );
  MUX2_X1 U15320 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13345), .S(n6436), .Z(
        P2_U3527) );
  NAND2_X1 U15321 ( .A1(n13270), .A2(n14753), .ZN(n13278) );
  AOI21_X1 U15322 ( .B1(n13272), .B2(n13261), .A(n13271), .ZN(n13277) );
  NAND3_X1 U15323 ( .A1(n13274), .A2(n13273), .A3(n13287), .ZN(n13276) );
  NAND4_X1 U15324 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13346) );
  MUX2_X1 U15325 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13346), .S(n6436), .Z(
        P2_U3526) );
  INV_X1 U15326 ( .A(n13279), .ZN(n13280) );
  OAI211_X1 U15327 ( .C1(n13282), .C2(n14764), .A(n13281), .B(n13280), .ZN(
        n13283) );
  AOI21_X1 U15328 ( .B1(n13284), .B2(n13287), .A(n13283), .ZN(n13285) );
  OAI21_X1 U15329 ( .B1(n13286), .B2(n7052), .A(n13285), .ZN(n13347) );
  MUX2_X1 U15330 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13347), .S(n6436), .Z(
        P2_U3525) );
  AND2_X1 U15331 ( .A1(n13288), .A2(n13287), .ZN(n13292) );
  OAI21_X1 U15332 ( .B1(n13290), .B2(n14764), .A(n13289), .ZN(n13291) );
  MUX2_X1 U15333 ( .A(n13348), .B(P2_REG1_REG_25__SCAN_IN), .S(n14776), .Z(
        P2_U3524) );
  INV_X1 U15334 ( .A(n13294), .ZN(n13299) );
  AOI21_X1 U15335 ( .B1(n13261), .B2(n13296), .A(n13295), .ZN(n13297) );
  OAI211_X1 U15336 ( .C1(n14761), .C2(n13299), .A(n13298), .B(n13297), .ZN(
        n13349) );
  MUX2_X1 U15337 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13349), .S(n6436), .Z(
        P2_U3523) );
  OAI211_X1 U15338 ( .C1(n11763), .C2(n14764), .A(n13301), .B(n13300), .ZN(
        n13302) );
  AOI21_X1 U15339 ( .B1(n13303), .B2(n14753), .A(n13302), .ZN(n13304) );
  OAI21_X1 U15340 ( .B1(n14749), .B2(n13305), .A(n13304), .ZN(n13350) );
  MUX2_X1 U15341 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13350), .S(n6436), .Z(
        P2_U3522) );
  AOI21_X1 U15342 ( .B1(n13261), .B2(n13307), .A(n13306), .ZN(n13308) );
  OAI211_X1 U15343 ( .C1(n14749), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        n13351) );
  MUX2_X1 U15344 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13351), .S(n6436), .Z(
        P2_U3521) );
  INV_X1 U15345 ( .A(n13311), .ZN(n13312) );
  OAI211_X1 U15346 ( .C1(n13314), .C2(n14764), .A(n13313), .B(n13312), .ZN(
        n13315) );
  AOI21_X1 U15347 ( .B1(n13316), .B2(n14753), .A(n13315), .ZN(n13317) );
  OAI21_X1 U15348 ( .B1(n14749), .B2(n13318), .A(n13317), .ZN(n13352) );
  MUX2_X1 U15349 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13352), .S(n6436), .Z(
        P2_U3520) );
  AOI211_X1 U15350 ( .C1(n13261), .C2(n13321), .A(n13320), .B(n13319), .ZN(
        n13322) );
  OAI21_X1 U15351 ( .B1(n14749), .B2(n13323), .A(n13322), .ZN(n13353) );
  MUX2_X1 U15352 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13353), .S(n6436), .Z(
        P2_U3519) );
  AOI211_X1 U15353 ( .C1(n13261), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        n13327) );
  OAI21_X1 U15354 ( .B1(n14749), .B2(n13328), .A(n13327), .ZN(n13354) );
  MUX2_X1 U15355 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13354), .S(n6436), .Z(
        P2_U3518) );
  AOI21_X1 U15356 ( .B1(n13261), .B2(n13330), .A(n13329), .ZN(n13331) );
  OAI211_X1 U15357 ( .C1(n13333), .C2(n14749), .A(n13332), .B(n13331), .ZN(
        n13355) );
  MUX2_X1 U15358 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13355), .S(n6436), .Z(
        P2_U3517) );
  OAI21_X1 U15359 ( .B1(n13335), .B2(n14764), .A(n13334), .ZN(n13337) );
  AOI211_X1 U15360 ( .C1(n13338), .C2(n14753), .A(n13337), .B(n13336), .ZN(
        n13339) );
  OAI21_X1 U15361 ( .B1(n14749), .B2(n13340), .A(n13339), .ZN(n13356) );
  MUX2_X1 U15362 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13356), .S(n6436), .Z(
        P2_U3516) );
  MUX2_X1 U15363 ( .A(n13341), .B(P2_REG1_REG_2__SCAN_IN), .S(n14776), .Z(
        P2_U3501) );
  MUX2_X1 U15364 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13342), .S(n14754), .Z(
        P2_U3498) );
  MUX2_X1 U15365 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13343), .S(n14754), .Z(
        P2_U3497) );
  MUX2_X1 U15366 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13345), .S(n14754), .Z(
        P2_U3495) );
  MUX2_X1 U15367 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13346), .S(n14754), .Z(
        P2_U3494) );
  MUX2_X1 U15368 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13347), .S(n14754), .Z(
        P2_U3493) );
  MUX2_X1 U15369 ( .A(n13348), .B(P2_REG0_REG_25__SCAN_IN), .S(n14769), .Z(
        P2_U3492) );
  MUX2_X1 U15370 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13349), .S(n14754), .Z(
        P2_U3491) );
  MUX2_X1 U15371 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13350), .S(n14754), .Z(
        P2_U3490) );
  MUX2_X1 U15372 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13351), .S(n14754), .Z(
        P2_U3489) );
  MUX2_X1 U15373 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13352), .S(n14754), .Z(
        P2_U3488) );
  MUX2_X1 U15374 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13353), .S(n14754), .Z(
        P2_U3487) );
  MUX2_X1 U15375 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13354), .S(n14754), .Z(
        P2_U3486) );
  MUX2_X1 U15376 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13355), .S(n14754), .Z(
        P2_U3484) );
  MUX2_X1 U15377 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13356), .S(n14754), .Z(
        P2_U3481) );
  NAND3_X1 U15378 ( .A1(n13357), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13359) );
  OAI22_X1 U15379 ( .A1(n13360), .A2(n13359), .B1(n13358), .B2(n13377), .ZN(
        n13361) );
  AOI21_X1 U15380 ( .B1(n14185), .B2(n13366), .A(n13361), .ZN(n13362) );
  INV_X1 U15381 ( .A(n13362), .ZN(P2_U3296) );
  INV_X1 U15382 ( .A(n13363), .ZN(n14188) );
  OAI222_X1 U15383 ( .A1(n13373), .A2(n14188), .B1(n13365), .B2(P2_U3088), 
        .C1(n13364), .C2(n13377), .ZN(P2_U3297) );
  NAND2_X1 U15384 ( .A1(n13367), .A2(n13366), .ZN(n13369) );
  OAI211_X1 U15385 ( .C1(n13377), .C2(n13370), .A(n13369), .B(n13368), .ZN(
        P2_U3299) );
  INV_X1 U15386 ( .A(n13371), .ZN(n14193) );
  OAI222_X1 U15387 ( .A1(n13373), .A2(n14193), .B1(n13372), .B2(P2_U3088), 
        .C1(n15097), .C2(n13377), .ZN(P2_U3301) );
  INV_X1 U15388 ( .A(n13374), .ZN(n14197) );
  OAI222_X1 U15389 ( .A1(n13377), .A2(n13376), .B1(n13373), .B2(n14197), .C1(
        P2_U3088), .C2(n13375), .ZN(P2_U3302) );
  INV_X1 U15390 ( .A(n13378), .ZN(n13379) );
  MUX2_X1 U15391 ( .A(n13379), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15392 ( .A1(n14093), .A2(n13491), .ZN(n13381) );
  NAND2_X1 U15393 ( .A1(n10123), .A2(n13817), .ZN(n13380) );
  NAND2_X1 U15394 ( .A1(n13381), .A2(n13380), .ZN(n13382) );
  XNOR2_X1 U15395 ( .A(n13382), .B(n13537), .ZN(n13530) );
  AOI22_X1 U15396 ( .A1(n14093), .A2(n13481), .B1(n13485), .B2(n13817), .ZN(
        n13531) );
  XNOR2_X1 U15397 ( .A(n13530), .B(n13531), .ZN(n13533) );
  AOI22_X1 U15398 ( .A1(n14428), .A2(n13491), .B1(n10123), .B2(n14416), .ZN(
        n13383) );
  XNOR2_X1 U15399 ( .A(n13383), .B(n13395), .ZN(n13408) );
  AOI22_X1 U15400 ( .A1(n14428), .A2(n13481), .B1(n13485), .B2(n14416), .ZN(
        n13407) );
  INV_X1 U15401 ( .A(n13384), .ZN(n13385) );
  NAND2_X1 U15402 ( .A1(n14238), .A2(n13491), .ZN(n13389) );
  NAND2_X1 U15403 ( .A1(n13481), .A2(n14253), .ZN(n13388) );
  NAND2_X1 U15404 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  XNOR2_X1 U15405 ( .A(n13390), .B(n13537), .ZN(n13399) );
  NAND2_X1 U15406 ( .A1(n14238), .A2(n10123), .ZN(n13392) );
  NAND2_X1 U15407 ( .A1(n13485), .A2(n14253), .ZN(n13391) );
  NAND2_X1 U15408 ( .A1(n13392), .A2(n13391), .ZN(n13400) );
  NAND2_X1 U15409 ( .A1(n13399), .A2(n13400), .ZN(n14371) );
  NAND2_X1 U15410 ( .A1(n14406), .A2(n13491), .ZN(n13394) );
  NAND2_X1 U15411 ( .A1(n10123), .A2(n14361), .ZN(n13393) );
  NAND2_X1 U15412 ( .A1(n13394), .A2(n13393), .ZN(n13396) );
  XNOR2_X1 U15413 ( .A(n13396), .B(n13395), .ZN(n13404) );
  NOR2_X1 U15414 ( .A1(n13535), .A2(n13397), .ZN(n13398) );
  AOI21_X1 U15415 ( .B1(n14406), .B2(n13481), .A(n13398), .ZN(n13405) );
  XNOR2_X1 U15416 ( .A(n13404), .B(n13405), .ZN(n14399) );
  INV_X1 U15417 ( .A(n13399), .ZN(n13402) );
  INV_X1 U15418 ( .A(n13400), .ZN(n13401) );
  NAND2_X1 U15419 ( .A1(n13402), .A2(n13401), .ZN(n14400) );
  INV_X1 U15420 ( .A(n13404), .ZN(n13406) );
  XNOR2_X1 U15421 ( .A(n13408), .B(n13407), .ZN(n14360) );
  NAND2_X1 U15422 ( .A1(n13412), .A2(n13491), .ZN(n13410) );
  NAND2_X1 U15423 ( .A1(n10123), .A2(n14386), .ZN(n13409) );
  NAND2_X1 U15424 ( .A1(n13410), .A2(n13409), .ZN(n13411) );
  XNOR2_X1 U15425 ( .A(n13411), .B(n10689), .ZN(n13413) );
  XNOR2_X1 U15426 ( .A(n13415), .B(n13413), .ZN(n14412) );
  AOI22_X1 U15427 ( .A1(n13412), .A2(n13481), .B1(n13485), .B2(n14386), .ZN(
        n14413) );
  NAND2_X1 U15428 ( .A1(n14412), .A2(n14413), .ZN(n14411) );
  INV_X1 U15429 ( .A(n13413), .ZN(n13414) );
  NAND2_X1 U15430 ( .A1(n14149), .A2(n13491), .ZN(n13418) );
  NAND2_X1 U15431 ( .A1(n14414), .A2(n10123), .ZN(n13417) );
  NAND2_X1 U15432 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  XNOR2_X1 U15433 ( .A(n13419), .B(n13537), .ZN(n13420) );
  AOI22_X1 U15434 ( .A1(n14149), .A2(n13481), .B1(n13485), .B2(n14414), .ZN(
        n13421) );
  XNOR2_X1 U15435 ( .A(n13420), .B(n13421), .ZN(n14384) );
  INV_X1 U15436 ( .A(n13420), .ZN(n13422) );
  AOI22_X1 U15437 ( .A1(n14146), .A2(n13481), .B1(n13485), .B2(n14385), .ZN(
        n13426) );
  NAND2_X1 U15438 ( .A1(n14146), .A2(n13491), .ZN(n13424) );
  NAND2_X1 U15439 ( .A1(n14385), .A2(n13481), .ZN(n13423) );
  NAND2_X1 U15440 ( .A1(n13424), .A2(n13423), .ZN(n13425) );
  XNOR2_X1 U15441 ( .A(n13425), .B(n13537), .ZN(n13428) );
  XOR2_X1 U15442 ( .A(n13426), .B(n13428), .Z(n13567) );
  INV_X1 U15443 ( .A(n13426), .ZN(n13427) );
  OAI22_X1 U15444 ( .A1(n14045), .A2(n13536), .B1(n13568), .B2(n13535), .ZN(
        n13433) );
  NAND2_X1 U15445 ( .A1(n14141), .A2(n13491), .ZN(n13430) );
  NAND2_X1 U15446 ( .A1(n14021), .A2(n10123), .ZN(n13429) );
  NAND2_X1 U15447 ( .A1(n13430), .A2(n13429), .ZN(n13431) );
  XNOR2_X1 U15448 ( .A(n13431), .B(n13537), .ZN(n13432) );
  XOR2_X1 U15449 ( .A(n13433), .B(n13432), .Z(n13601) );
  INV_X1 U15450 ( .A(n13432), .ZN(n13435) );
  INV_X1 U15451 ( .A(n13433), .ZN(n13434) );
  NAND2_X1 U15452 ( .A1(n13435), .A2(n13434), .ZN(n13436) );
  NAND2_X1 U15453 ( .A1(n13437), .A2(n13436), .ZN(n13522) );
  INV_X1 U15454 ( .A(n13522), .ZN(n13443) );
  AND2_X1 U15455 ( .A1(n14001), .A2(n13485), .ZN(n13438) );
  AOI21_X1 U15456 ( .B1(n14134), .B2(n13481), .A(n13438), .ZN(n13444) );
  NAND2_X1 U15457 ( .A1(n14134), .A2(n13491), .ZN(n13440) );
  NAND2_X1 U15458 ( .A1(n14001), .A2(n13481), .ZN(n13439) );
  NAND2_X1 U15459 ( .A1(n13440), .A2(n13439), .ZN(n13441) );
  XNOR2_X1 U15460 ( .A(n13441), .B(n13537), .ZN(n13446) );
  XOR2_X1 U15461 ( .A(n13444), .B(n13446), .Z(n13521) );
  NAND2_X1 U15462 ( .A1(n13443), .A2(n13442), .ZN(n13523) );
  INV_X1 U15463 ( .A(n13444), .ZN(n13445) );
  NAND2_X1 U15464 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NAND2_X1 U15465 ( .A1(n13523), .A2(n13447), .ZN(n13583) );
  AND2_X1 U15466 ( .A1(n14022), .A2(n13485), .ZN(n13448) );
  AOI21_X1 U15467 ( .B1(n14130), .B2(n13481), .A(n13448), .ZN(n13451) );
  AOI22_X1 U15468 ( .A1(n14130), .A2(n13491), .B1(n10123), .B2(n14022), .ZN(
        n13449) );
  XNOR2_X1 U15469 ( .A(n13449), .B(n13537), .ZN(n13450) );
  XOR2_X1 U15470 ( .A(n13451), .B(n13450), .Z(n13582) );
  INV_X1 U15471 ( .A(n13450), .ZN(n13453) );
  INV_X1 U15472 ( .A(n13451), .ZN(n13452) );
  NAND2_X1 U15473 ( .A1(n13453), .A2(n13452), .ZN(n13454) );
  AOI22_X1 U15474 ( .A1(n14125), .A2(n13491), .B1(n10123), .B2(n14002), .ZN(
        n13455) );
  XNOR2_X1 U15475 ( .A(n13455), .B(n13537), .ZN(n13458) );
  AOI22_X1 U15476 ( .A1(n14125), .A2(n10123), .B1(n13485), .B2(n14002), .ZN(
        n13457) );
  XNOR2_X1 U15477 ( .A(n13458), .B(n13457), .ZN(n13552) );
  NAND2_X1 U15478 ( .A1(n13458), .A2(n13457), .ZN(n13459) );
  NAND2_X1 U15479 ( .A1(n13549), .A2(n13459), .ZN(n13590) );
  INV_X1 U15480 ( .A(n13984), .ZN(n13950) );
  OAI22_X1 U15481 ( .A1(n13599), .A2(n13536), .B1(n13950), .B2(n13535), .ZN(
        n13464) );
  NAND2_X1 U15482 ( .A1(n14120), .A2(n13491), .ZN(n13461) );
  NAND2_X1 U15483 ( .A1(n13481), .A2(n13984), .ZN(n13460) );
  NAND2_X1 U15484 ( .A1(n13461), .A2(n13460), .ZN(n13462) );
  XNOR2_X1 U15485 ( .A(n13462), .B(n13537), .ZN(n13463) );
  XOR2_X1 U15486 ( .A(n13464), .B(n13463), .Z(n13591) );
  NAND2_X1 U15487 ( .A1(n13590), .A2(n13591), .ZN(n13589) );
  INV_X1 U15488 ( .A(n13463), .ZN(n13466) );
  INV_X1 U15489 ( .A(n13464), .ZN(n13465) );
  NAND2_X1 U15490 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  NAND2_X1 U15491 ( .A1(n13589), .A2(n13467), .ZN(n13506) );
  NAND2_X1 U15492 ( .A1(n14112), .A2(n13491), .ZN(n13469) );
  NAND2_X1 U15493 ( .A1(n10123), .A2(n13934), .ZN(n13468) );
  NAND2_X1 U15494 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  XNOR2_X1 U15495 ( .A(n13470), .B(n13537), .ZN(n13471) );
  AOI22_X1 U15496 ( .A1(n14112), .A2(n13481), .B1(n13485), .B2(n13934), .ZN(
        n13472) );
  XNOR2_X1 U15497 ( .A(n13471), .B(n13472), .ZN(n13507) );
  INV_X1 U15498 ( .A(n13471), .ZN(n13473) );
  NAND2_X1 U15499 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U15500 ( .A1(n14106), .A2(n13491), .ZN(n13476) );
  NAND2_X1 U15501 ( .A1(n13481), .A2(n13837), .ZN(n13475) );
  NAND2_X1 U15502 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  XNOR2_X1 U15503 ( .A(n13477), .B(n13537), .ZN(n13478) );
  AOI22_X1 U15504 ( .A1(n14106), .A2(n13481), .B1(n13485), .B2(n13837), .ZN(
        n13479) );
  XNOR2_X1 U15505 ( .A(n13478), .B(n13479), .ZN(n13575) );
  INV_X1 U15506 ( .A(n13478), .ZN(n13480) );
  NAND2_X1 U15507 ( .A1(n13924), .A2(n13491), .ZN(n13483) );
  NAND2_X1 U15508 ( .A1(n13481), .A2(n13933), .ZN(n13482) );
  NAND2_X1 U15509 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  XNOR2_X1 U15510 ( .A(n13484), .B(n13537), .ZN(n13486) );
  AOI22_X1 U15511 ( .A1(n13924), .A2(n10123), .B1(n13485), .B2(n13933), .ZN(
        n13487) );
  XNOR2_X1 U15512 ( .A(n13486), .B(n13487), .ZN(n13559) );
  NAND2_X1 U15513 ( .A1(n13558), .A2(n13559), .ZN(n13490) );
  INV_X1 U15514 ( .A(n13486), .ZN(n13488) );
  NAND2_X1 U15515 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  NAND2_X1 U15516 ( .A1(n13490), .A2(n13489), .ZN(n13608) );
  OAI22_X1 U15517 ( .A1(n7250), .A2(n13536), .B1(n13881), .B2(n13535), .ZN(
        n13496) );
  NAND2_X1 U15518 ( .A1(n14098), .A2(n13491), .ZN(n13493) );
  NAND2_X1 U15519 ( .A1(n10123), .A2(n13839), .ZN(n13492) );
  NAND2_X1 U15520 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  XNOR2_X1 U15521 ( .A(n13494), .B(n13537), .ZN(n13495) );
  XOR2_X1 U15522 ( .A(n13496), .B(n13495), .Z(n13609) );
  NAND2_X1 U15523 ( .A1(n13608), .A2(n13609), .ZN(n13500) );
  INV_X1 U15524 ( .A(n13495), .ZN(n13498) );
  INV_X1 U15525 ( .A(n13496), .ZN(n13497) );
  NAND2_X1 U15526 ( .A1(n13498), .A2(n13497), .ZN(n13499) );
  NAND2_X1 U15527 ( .A1(n13500), .A2(n13499), .ZN(n13534) );
  XOR2_X1 U15528 ( .A(n13533), .B(n13534), .Z(n13505) );
  OAI22_X1 U15529 ( .A1(n14394), .A2(n13881), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15068), .ZN(n13501) );
  AOI21_X1 U15530 ( .B1(n14415), .B2(n13851), .A(n13501), .ZN(n13502) );
  OAI21_X1 U15531 ( .B1(n13889), .B2(n14425), .A(n13502), .ZN(n13503) );
  AOI21_X1 U15532 ( .B1(n14093), .B2(n14407), .A(n13503), .ZN(n13504) );
  OAI21_X1 U15533 ( .B1(n13505), .B2(n14401), .A(n13504), .ZN(P1_U3214) );
  XOR2_X1 U15534 ( .A(n13507), .B(n13506), .Z(n13512) );
  NOR2_X1 U15535 ( .A1(n14425), .A2(n13953), .ZN(n13510) );
  AOI22_X1 U15536 ( .A1(n14415), .A2(n13837), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13508) );
  OAI21_X1 U15537 ( .B1(n13950), .B2(n14394), .A(n13508), .ZN(n13509) );
  AOI211_X1 U15538 ( .C1(n14112), .C2(n14407), .A(n13510), .B(n13509), .ZN(
        n13511) );
  OAI21_X1 U15539 ( .B1(n13512), .B2(n14401), .A(n13511), .ZN(P1_U3216) );
  OAI211_X1 U15540 ( .C1(n13515), .C2(n13514), .A(n13513), .B(n14421), .ZN(
        n13520) );
  AOI22_X1 U15541 ( .A1(n14417), .A2(n13626), .B1(n14415), .B2(n13624), .ZN(
        n13519) );
  MUX2_X1 U15542 ( .A(n14425), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13518) );
  NAND2_X1 U15543 ( .A1(n14407), .A2(n13516), .ZN(n13517) );
  NAND4_X1 U15544 ( .A1(n13520), .A2(n13519), .A3(n13518), .A4(n13517), .ZN(
        P1_U3218) );
  INV_X1 U15545 ( .A(n14134), .ZN(n13529) );
  AOI21_X1 U15546 ( .B1(n13522), .B2(n13521), .A(n14401), .ZN(n13524) );
  NAND2_X1 U15547 ( .A1(n13524), .A2(n13523), .ZN(n13528) );
  NOR2_X1 U15548 ( .A1(n14425), .A2(n14026), .ZN(n13526) );
  NAND2_X1 U15549 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13785)
         );
  OAI21_X1 U15550 ( .B1(n13828), .B2(n14397), .A(n13785), .ZN(n13525) );
  AOI211_X1 U15551 ( .C1(n14417), .C2(n14021), .A(n13526), .B(n13525), .ZN(
        n13527) );
  OAI211_X1 U15552 ( .C1(n13529), .C2(n14419), .A(n13528), .B(n13527), .ZN(
        P1_U3219) );
  INV_X1 U15553 ( .A(n13530), .ZN(n13532) );
  AOI22_X1 U15554 ( .A1(n13534), .A2(n13533), .B1(n13532), .B2(n13531), .ZN(
        n13542) );
  OAI22_X1 U15555 ( .A1(n13869), .A2(n10124), .B1(n13880), .B2(n13536), .ZN(
        n13540) );
  OAI22_X1 U15556 ( .A1(n13869), .A2(n13536), .B1(n13880), .B2(n13535), .ZN(
        n13538) );
  XNOR2_X1 U15557 ( .A(n13538), .B(n13537), .ZN(n13539) );
  XOR2_X1 U15558 ( .A(n13540), .B(n13539), .Z(n13541) );
  XNOR2_X1 U15559 ( .A(n13542), .B(n13541), .ZN(n13548) );
  NAND2_X1 U15560 ( .A1(n13616), .A2(n14254), .ZN(n13544) );
  NAND2_X1 U15561 ( .A1(n13817), .A2(n14252), .ZN(n13543) );
  NAND2_X1 U15562 ( .A1(n13544), .A2(n13543), .ZN(n14084) );
  AOI22_X1 U15563 ( .A1(n14379), .A2(n14084), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13545) );
  OAI21_X1 U15564 ( .B1(n13864), .B2(n14425), .A(n13545), .ZN(n13546) );
  AOI21_X1 U15565 ( .B1(n14085), .B2(n14407), .A(n13546), .ZN(n13547) );
  OAI21_X1 U15566 ( .B1(n13548), .B2(n14401), .A(n13547), .ZN(P1_U3220) );
  INV_X1 U15567 ( .A(n13549), .ZN(n13550) );
  AOI21_X1 U15568 ( .B1(n13552), .B2(n13551), .A(n13550), .ZN(n13557) );
  NOR2_X1 U15569 ( .A1(n14425), .A2(n13994), .ZN(n13555) );
  AOI22_X1 U15570 ( .A1(n14415), .A2(n13984), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13553) );
  OAI21_X1 U15571 ( .B1(n13828), .B2(n14394), .A(n13553), .ZN(n13554) );
  AOI211_X1 U15572 ( .C1(n14125), .C2(n14407), .A(n13555), .B(n13554), .ZN(
        n13556) );
  OAI21_X1 U15573 ( .B1(n13557), .B2(n14401), .A(n13556), .ZN(P1_U3223) );
  XOR2_X1 U15574 ( .A(n13559), .B(n13558), .Z(n13565) );
  NAND2_X1 U15575 ( .A1(n13837), .A2(n14252), .ZN(n13561) );
  NAND2_X1 U15576 ( .A1(n13839), .A2(n14254), .ZN(n13560) );
  NAND2_X1 U15577 ( .A1(n13561), .A2(n13560), .ZN(n13916) );
  AOI22_X1 U15578 ( .A1(n14379), .A2(n13916), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13562) );
  OAI21_X1 U15579 ( .B1(n13921), .B2(n14425), .A(n13562), .ZN(n13563) );
  AOI21_X1 U15580 ( .B1(n13924), .B2(n14407), .A(n13563), .ZN(n13564) );
  OAI21_X1 U15581 ( .B1(n13565), .B2(n14401), .A(n13564), .ZN(P1_U3225) );
  XOR2_X1 U15582 ( .A(n13567), .B(n13566), .Z(n13573) );
  OAI22_X1 U15583 ( .A1(n13568), .A2(n13951), .B1(n13820), .B2(n13949), .ZN(
        n14051) );
  NAND2_X1 U15584 ( .A1(n14051), .A2(n14379), .ZN(n13570) );
  OAI211_X1 U15585 ( .C1(n14425), .C2(n14059), .A(n13570), .B(n13569), .ZN(
        n13571) );
  AOI21_X1 U15586 ( .B1(n14146), .B2(n14407), .A(n13571), .ZN(n13572) );
  OAI21_X1 U15587 ( .B1(n13573), .B2(n14401), .A(n13572), .ZN(P1_U3228) );
  XOR2_X1 U15588 ( .A(n13575), .B(n13574), .Z(n13580) );
  NOR2_X1 U15589 ( .A1(n14425), .A2(n13940), .ZN(n13578) );
  INV_X1 U15590 ( .A(n13934), .ZN(n13835) );
  AOI22_X1 U15591 ( .A1(n14415), .A2(n13933), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13576) );
  OAI21_X1 U15592 ( .B1(n13835), .B2(n14394), .A(n13576), .ZN(n13577) );
  AOI211_X1 U15593 ( .C1(n14106), .C2(n14407), .A(n13578), .B(n13577), .ZN(
        n13579) );
  OAI21_X1 U15594 ( .B1(n13580), .B2(n14401), .A(n13579), .ZN(P1_U3229) );
  INV_X1 U15595 ( .A(n14130), .ZN(n14011) );
  OAI211_X1 U15596 ( .C1(n13583), .C2(n13582), .A(n13581), .B(n14421), .ZN(
        n13588) );
  NOR2_X1 U15597 ( .A1(n14425), .A2(n14008), .ZN(n13586) );
  OAI22_X1 U15598 ( .A1(n13830), .A2(n14397), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13584), .ZN(n13585) );
  AOI211_X1 U15599 ( .C1(n14417), .C2(n14001), .A(n13586), .B(n13585), .ZN(
        n13587) );
  OAI211_X1 U15600 ( .C1(n14011), .C2(n14419), .A(n13588), .B(n13587), .ZN(
        P1_U3233) );
  OAI21_X1 U15601 ( .B1(n13591), .B2(n13590), .A(n13589), .ZN(n13592) );
  NAND2_X1 U15602 ( .A1(n13592), .A2(n14421), .ZN(n13598) );
  INV_X1 U15603 ( .A(n13593), .ZN(n13969) );
  AND2_X1 U15604 ( .A1(n13934), .A2(n14254), .ZN(n13594) );
  AOI21_X1 U15605 ( .B1(n14002), .B2(n14252), .A(n13594), .ZN(n14117) );
  INV_X1 U15606 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13595) );
  OAI22_X1 U15607 ( .A1(n14117), .A2(n13604), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13595), .ZN(n13596) );
  AOI21_X1 U15608 ( .B1(n13969), .B2(n13602), .A(n13596), .ZN(n13597) );
  OAI211_X1 U15609 ( .C1(n14419), .C2(n13599), .A(n13598), .B(n13597), .ZN(
        P1_U3235) );
  XOR2_X1 U15610 ( .A(n13601), .B(n13600), .Z(n13607) );
  AOI22_X1 U15611 ( .A1(n14001), .A2(n14254), .B1(n14252), .B2(n14385), .ZN(
        n14036) );
  NAND2_X1 U15612 ( .A1(n13602), .A2(n14041), .ZN(n13603) );
  NAND2_X1 U15613 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14526)
         );
  OAI211_X1 U15614 ( .C1(n14036), .C2(n13604), .A(n13603), .B(n14526), .ZN(
        n13605) );
  AOI21_X1 U15615 ( .B1(n14141), .B2(n14407), .A(n13605), .ZN(n13606) );
  OAI21_X1 U15616 ( .B1(n13607), .B2(n14401), .A(n13606), .ZN(P1_U3238) );
  XOR2_X1 U15617 ( .A(n13609), .B(n13608), .Z(n13615) );
  NAND2_X1 U15618 ( .A1(n13933), .A2(n14252), .ZN(n13611) );
  NAND2_X1 U15619 ( .A1(n13817), .A2(n14254), .ZN(n13610) );
  NAND2_X1 U15620 ( .A1(n13611), .A2(n13610), .ZN(n14097) );
  AOI22_X1 U15621 ( .A1(n14379), .A2(n14097), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13612) );
  OAI21_X1 U15622 ( .B1(n13898), .B2(n14425), .A(n13612), .ZN(n13613) );
  AOI21_X1 U15623 ( .B1(n14098), .B2(n14407), .A(n13613), .ZN(n13614) );
  OAI21_X1 U15624 ( .B1(n13615), .B2(n14401), .A(n13614), .ZN(P1_U3240) );
  MUX2_X1 U15625 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13793), .S(n13644), .Z(
        P1_U3591) );
  MUX2_X1 U15626 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13847), .S(n13644), .Z(
        P1_U3590) );
  MUX2_X1 U15627 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13616), .S(n13644), .Z(
        P1_U3589) );
  MUX2_X1 U15628 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13851), .S(n13644), .Z(
        P1_U3588) );
  MUX2_X1 U15629 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13817), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15630 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13839), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15631 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13933), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15632 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13837), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15633 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13934), .S(n13644), .Z(
        P1_U3583) );
  MUX2_X1 U15634 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13984), .S(n13644), .Z(
        P1_U3582) );
  MUX2_X1 U15635 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14002), .S(n13644), .Z(
        P1_U3581) );
  MUX2_X1 U15636 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14022), .S(n13644), .Z(
        P1_U3580) );
  MUX2_X1 U15637 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14001), .S(n13644), .Z(
        P1_U3579) );
  MUX2_X1 U15638 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14021), .S(n13644), .Z(
        P1_U3578) );
  MUX2_X1 U15639 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14385), .S(n13644), .Z(
        P1_U3577) );
  MUX2_X1 U15640 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14414), .S(n13644), .Z(
        P1_U3576) );
  MUX2_X1 U15641 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14386), .S(n13644), .Z(
        P1_U3575) );
  MUX2_X1 U15642 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14416), .S(n13644), .Z(
        P1_U3574) );
  MUX2_X1 U15643 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14361), .S(n13644), .Z(
        P1_U3573) );
  MUX2_X1 U15644 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14253), .S(n13644), .Z(
        P1_U3572) );
  MUX2_X1 U15645 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13617), .S(n13644), .Z(
        P1_U3571) );
  MUX2_X1 U15646 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13618), .S(n13644), .Z(
        P1_U3570) );
  MUX2_X1 U15647 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13619), .S(n13644), .Z(
        P1_U3569) );
  MUX2_X1 U15648 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13620), .S(n13644), .Z(
        P1_U3568) );
  MUX2_X1 U15649 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13621), .S(n13644), .Z(
        P1_U3567) );
  MUX2_X1 U15650 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13622), .S(n13644), .Z(
        P1_U3566) );
  MUX2_X1 U15651 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13623), .S(n13644), .Z(
        P1_U3565) );
  MUX2_X1 U15652 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13624), .S(n13644), .Z(
        P1_U3564) );
  MUX2_X1 U15653 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13625), .S(n13644), .Z(
        P1_U3563) );
  MUX2_X1 U15654 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13626), .S(n13644), .Z(
        P1_U3562) );
  MUX2_X1 U15655 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13627), .S(n13644), .Z(
        P1_U3561) );
  MUX2_X1 U15656 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13628), .S(n13644), .Z(
        P1_U3560) );
  OAI211_X1 U15657 ( .C1(n13641), .C2(n13630), .A(n14492), .B(n13629), .ZN(
        n13638) );
  MUX2_X1 U15658 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9827), .S(n13631), .Z(
        n13632) );
  OAI21_X1 U15659 ( .B1(n8543), .B2(n14476), .A(n13632), .ZN(n13633) );
  NAND3_X1 U15660 ( .A1(n14486), .A2(n13653), .A3(n13633), .ZN(n13637) );
  NAND2_X1 U15661 ( .A1(n14494), .A2(n13634), .ZN(n13636) );
  AOI22_X1 U15662 ( .A1(n14497), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13635) );
  NAND4_X1 U15663 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        P1_U3244) );
  NOR2_X1 U15664 ( .A1(n14191), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13639) );
  MUX2_X1 U15665 ( .A(n13641), .B(n13640), .S(n14191), .Z(n13643) );
  NAND2_X1 U15666 ( .A1(n13643), .A2(n13642), .ZN(n13645) );
  OAI211_X1 U15667 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6587), .A(n13645), .B(
        n13644), .ZN(n14502) );
  AOI22_X1 U15668 ( .A1(n14497), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13657) );
  XNOR2_X1 U15669 ( .A(n13647), .B(n13646), .ZN(n13648) );
  OAI22_X1 U15670 ( .A1(n13648), .A2(n14520), .B1(n14524), .B2(n13650), .ZN(
        n13649) );
  INV_X1 U15671 ( .A(n13649), .ZN(n13656) );
  MUX2_X1 U15672 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9830), .S(n13650), .Z(
        n13651) );
  NAND3_X1 U15673 ( .A1(n13653), .A2(n13652), .A3(n13651), .ZN(n13654) );
  NAND3_X1 U15674 ( .A1(n14486), .A2(n13666), .A3(n13654), .ZN(n13655) );
  NAND4_X1 U15675 ( .A1(n14502), .A2(n13657), .A3(n13656), .A4(n13655), .ZN(
        P1_U3245) );
  INV_X1 U15676 ( .A(n14497), .ZN(n14528) );
  OAI22_X1 U15677 ( .A1(n14528), .A2(n13659), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13658), .ZN(n13660) );
  AOI21_X1 U15678 ( .B1(n13663), .B2(n14494), .A(n13660), .ZN(n13670) );
  OAI211_X1 U15679 ( .C1(n13662), .C2(n13661), .A(n14492), .B(n14488), .ZN(
        n13669) );
  MUX2_X1 U15680 ( .A(n9833), .B(P1_REG1_REG_3__SCAN_IN), .S(n13663), .Z(
        n13664) );
  NAND3_X1 U15681 ( .A1(n13666), .A2(n13665), .A3(n13664), .ZN(n13667) );
  NAND3_X1 U15682 ( .A1(n14486), .A2(n14482), .A3(n13667), .ZN(n13668) );
  NAND3_X1 U15683 ( .A1(n13670), .A2(n13669), .A3(n13668), .ZN(P1_U3246) );
  OAI21_X1 U15684 ( .B1(n14528), .B2(n13672), .A(n13671), .ZN(n13673) );
  AOI21_X1 U15685 ( .B1(n13674), .B2(n14494), .A(n13673), .ZN(n13686) );
  OAI21_X1 U15686 ( .B1(n13677), .B2(n13676), .A(n13675), .ZN(n13678) );
  NAND2_X1 U15687 ( .A1(n14486), .A2(n13678), .ZN(n13685) );
  MUX2_X1 U15688 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9853), .S(n13679), .Z(
        n13681) );
  NAND3_X1 U15689 ( .A1(n13681), .A2(n14491), .A3(n13680), .ZN(n13682) );
  NAND3_X1 U15690 ( .A1(n14492), .A2(n13683), .A3(n13682), .ZN(n13684) );
  NAND3_X1 U15691 ( .A1(n13686), .A2(n13685), .A3(n13684), .ZN(P1_U3248) );
  INV_X1 U15692 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13688) );
  OAI21_X1 U15693 ( .B1(n14528), .B2(n13688), .A(n13687), .ZN(n13689) );
  AOI21_X1 U15694 ( .B1(n13696), .B2(n14494), .A(n13689), .ZN(n13704) );
  MUX2_X1 U15695 ( .A(n9858), .B(P1_REG2_REG_7__SCAN_IN), .S(n13696), .Z(
        n13690) );
  NAND3_X1 U15696 ( .A1(n13692), .A2(n13691), .A3(n13690), .ZN(n13693) );
  NAND3_X1 U15697 ( .A1(n14492), .A2(n13694), .A3(n13693), .ZN(n13703) );
  INV_X1 U15698 ( .A(n13695), .ZN(n13698) );
  MUX2_X1 U15699 ( .A(n14609), .B(P1_REG1_REG_7__SCAN_IN), .S(n13696), .Z(
        n13697) );
  NAND2_X1 U15700 ( .A1(n13698), .A2(n13697), .ZN(n13700) );
  OAI211_X1 U15701 ( .C1(n13701), .C2(n13700), .A(n14486), .B(n13699), .ZN(
        n13702) );
  NAND3_X1 U15702 ( .A1(n13704), .A2(n13703), .A3(n13702), .ZN(P1_U3250) );
  INV_X1 U15703 ( .A(n13705), .ZN(n13710) );
  NOR3_X1 U15704 ( .A1(n13708), .A2(n13707), .A3(n13706), .ZN(n13709) );
  OAI21_X1 U15705 ( .B1(n13710), .B2(n13709), .A(n14486), .ZN(n13723) );
  OAI21_X1 U15706 ( .B1(n14528), .B2(n13712), .A(n13711), .ZN(n13713) );
  AOI21_X1 U15707 ( .B1(n13714), .B2(n14494), .A(n13713), .ZN(n13722) );
  MUX2_X1 U15708 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9873), .S(n13715), .Z(
        n13716) );
  NAND3_X1 U15709 ( .A1(n13718), .A2(n13717), .A3(n13716), .ZN(n13719) );
  NAND3_X1 U15710 ( .A1(n14492), .A2(n13720), .A3(n13719), .ZN(n13721) );
  NAND3_X1 U15711 ( .A1(n13723), .A2(n13722), .A3(n13721), .ZN(P1_U3252) );
  OAI21_X1 U15712 ( .B1(n13726), .B2(n13725), .A(n13724), .ZN(n13727) );
  NAND2_X1 U15713 ( .A1(n13727), .A2(n14486), .ZN(n13739) );
  OAI21_X1 U15714 ( .B1(n14528), .B2(n13729), .A(n13728), .ZN(n13730) );
  AOI21_X1 U15715 ( .B1(n13731), .B2(n14494), .A(n13730), .ZN(n13738) );
  MUX2_X1 U15716 ( .A(n10004), .B(P1_REG2_REG_11__SCAN_IN), .S(n13731), .Z(
        n13732) );
  NAND3_X1 U15717 ( .A1(n13734), .A2(n13733), .A3(n13732), .ZN(n13735) );
  NAND3_X1 U15718 ( .A1(n13736), .A2(n14492), .A3(n13735), .ZN(n13737) );
  NAND3_X1 U15719 ( .A1(n13739), .A2(n13738), .A3(n13737), .ZN(P1_U3254) );
  OAI211_X1 U15720 ( .C1(n13742), .C2(n13741), .A(n14486), .B(n13740), .ZN(
        n13751) );
  INV_X1 U15721 ( .A(n13743), .ZN(n13744) );
  AOI22_X1 U15722 ( .A1(n14494), .A2(n13744), .B1(n14497), .B2(
        P1_ADDR_REG_13__SCAN_IN), .ZN(n13750) );
  NAND2_X1 U15723 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14408)
         );
  OAI211_X1 U15724 ( .C1(n13747), .C2(n13746), .A(n13745), .B(n14492), .ZN(
        n13748) );
  AND2_X1 U15725 ( .A1(n14408), .A2(n13748), .ZN(n13749) );
  NAND3_X1 U15726 ( .A1(n13751), .A2(n13750), .A3(n13749), .ZN(P1_U3256) );
  NAND2_X1 U15727 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14391)
         );
  OAI211_X1 U15728 ( .C1(n13754), .C2(n13753), .A(n14486), .B(n13752), .ZN(
        n13755) );
  AND2_X1 U15729 ( .A1(n14391), .A2(n13755), .ZN(n13762) );
  AOI22_X1 U15730 ( .A1(n14494), .A2(n13756), .B1(n14497), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n13761) );
  OAI211_X1 U15731 ( .C1(n13759), .C2(n13758), .A(n14492), .B(n13757), .ZN(
        n13760) );
  NAND3_X1 U15732 ( .A1(n13762), .A2(n13761), .A3(n13760), .ZN(P1_U3259) );
  INV_X1 U15733 ( .A(n13763), .ZN(n13767) );
  INV_X1 U15734 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13765) );
  OAI22_X1 U15735 ( .A1(n13767), .A2(n13766), .B1(n13765), .B2(n13764), .ZN(
        n13768) );
  XNOR2_X1 U15736 ( .A(n14523), .B(n13768), .ZN(n14516) );
  NAND2_X1 U15737 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14516), .ZN(n14515) );
  NAND2_X1 U15738 ( .A1(n13775), .A2(n13768), .ZN(n13769) );
  NAND2_X1 U15739 ( .A1(n14515), .A2(n13769), .ZN(n13771) );
  XNOR2_X1 U15740 ( .A(n13771), .B(n13770), .ZN(n13781) );
  INV_X1 U15741 ( .A(n13781), .ZN(n13779) );
  NAND2_X1 U15742 ( .A1(n13773), .A2(n13772), .ZN(n13774) );
  XNOR2_X1 U15743 ( .A(n14523), .B(n13774), .ZN(n14518) );
  NAND2_X1 U15744 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14518), .ZN(n14517) );
  NAND2_X1 U15745 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  NAND2_X1 U15746 ( .A1(n14517), .A2(n13776), .ZN(n13777) );
  XOR2_X1 U15747 ( .A(n13777), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13780) );
  OAI21_X1 U15748 ( .B1(n13780), .B2(n14520), .A(n14524), .ZN(n13778) );
  AOI21_X1 U15749 ( .B1(n14486), .B2(n13779), .A(n13778), .ZN(n13784) );
  AOI22_X1 U15750 ( .A1(n13781), .A2(n14486), .B1(n13780), .B2(n14492), .ZN(
        n13783) );
  MUX2_X1 U15751 ( .A(n13784), .B(n13783), .S(n13782), .Z(n13786) );
  OAI211_X1 U15752 ( .C1(n13787), .C2(n14528), .A(n13786), .B(n13785), .ZN(
        P1_U3262) );
  NAND2_X1 U15753 ( .A1(n14045), .A2(n14057), .ZN(n14039) );
  NOR2_X1 U15754 ( .A1(n13789), .A2(n13845), .ZN(n13791) );
  XNOR2_X1 U15755 ( .A(n13791), .B(n13790), .ZN(n14066) );
  NAND2_X1 U15756 ( .A1(n14066), .A2(n13792), .ZN(n13795) );
  AOI21_X1 U15757 ( .B1(n14475), .B2(P1_B_REG_SCAN_IN), .A(n13951), .ZN(n13848) );
  NAND2_X1 U15758 ( .A1(n13848), .A2(n13793), .ZN(n14069) );
  NOR2_X1 U15759 ( .A1(n14042), .A2(n14069), .ZN(n13798) );
  AOI21_X1 U15760 ( .B1(n14258), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13798), 
        .ZN(n13794) );
  OAI211_X1 U15761 ( .C1(n14068), .C2(n14260), .A(n13795), .B(n13794), .ZN(
        P1_U3263) );
  XNOR2_X1 U15762 ( .A(n13845), .B(n14071), .ZN(n13796) );
  NAND2_X1 U15763 ( .A1(n13796), .A2(n14548), .ZN(n14070) );
  NOR2_X1 U15764 ( .A1(n14071), .A2(n14260), .ZN(n13797) );
  AOI211_X1 U15765 ( .C1(n14258), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13798), 
        .B(n13797), .ZN(n13799) );
  OAI21_X1 U15766 ( .B1(n13998), .B2(n14070), .A(n13799), .ZN(P1_U3264) );
  OR2_X1 U15767 ( .A1(n14149), .A2(n14414), .ZN(n13800) );
  NAND2_X1 U15768 ( .A1(n13801), .A2(n13800), .ZN(n14048) );
  NAND2_X1 U15769 ( .A1(n14146), .A2(n14385), .ZN(n13802) );
  NAND2_X1 U15770 ( .A1(n14048), .A2(n13802), .ZN(n13804) );
  OR2_X1 U15771 ( .A1(n14146), .A2(n14385), .ZN(n13803) );
  NAND2_X1 U15772 ( .A1(n13804), .A2(n13803), .ZN(n14033) );
  NOR2_X1 U15773 ( .A1(n14141), .A2(n14021), .ZN(n13805) );
  NAND2_X1 U15774 ( .A1(n14141), .A2(n14021), .ZN(n13806) );
  INV_X1 U15775 ( .A(n14013), .ZN(n14000) );
  NAND2_X1 U15776 ( .A1(n14130), .A2(n14022), .ZN(n13987) );
  AND2_X1 U15777 ( .A1(n13986), .A2(n13987), .ZN(n13808) );
  OR2_X1 U15778 ( .A1(n14125), .A2(n14002), .ZN(n13809) );
  NAND2_X1 U15779 ( .A1(n13975), .A2(n13974), .ZN(n13973) );
  OR2_X1 U15780 ( .A1(n14120), .A2(n13984), .ZN(n13810) );
  NAND2_X1 U15781 ( .A1(n13973), .A2(n13810), .ZN(n13960) );
  INV_X1 U15782 ( .A(n13931), .ZN(n13929) );
  OR2_X1 U15783 ( .A1(n14106), .A2(n13837), .ZN(n13811) );
  NAND2_X1 U15784 ( .A1(n13924), .A2(n13933), .ZN(n13813) );
  NAND2_X1 U15785 ( .A1(n13913), .A2(n13813), .ZN(n13905) );
  NAND2_X1 U15786 ( .A1(n13905), .A2(n13904), .ZN(n13815) );
  NAND2_X1 U15787 ( .A1(n14098), .A2(n13839), .ZN(n13814) );
  INV_X1 U15788 ( .A(n13876), .ZN(n13816) );
  OR2_X1 U15789 ( .A1(n14093), .A2(n13817), .ZN(n13818) );
  INV_X1 U15790 ( .A(n13862), .ZN(n13858) );
  NOR2_X1 U15791 ( .A1(n13859), .A2(n13858), .ZN(n13861) );
  AOI21_X1 U15792 ( .B1(n14085), .B2(n13851), .A(n13861), .ZN(n13819) );
  XNOR2_X1 U15793 ( .A(n13819), .B(n13842), .ZN(n14082) );
  NAND2_X1 U15794 ( .A1(n14149), .A2(n13820), .ZN(n13821) );
  NAND2_X1 U15795 ( .A1(n14134), .A2(n13826), .ZN(n13827) );
  OR2_X1 U15796 ( .A1(n14130), .A2(n13828), .ZN(n13829) );
  INV_X1 U15797 ( .A(n13986), .ZN(n13982) );
  OR2_X1 U15798 ( .A1(n14125), .A2(n13830), .ZN(n13831) );
  NAND2_X1 U15799 ( .A1(n13981), .A2(n13831), .ZN(n13966) );
  NAND2_X1 U15800 ( .A1(n14120), .A2(n13950), .ZN(n13834) );
  AND2_X1 U15801 ( .A1(n14112), .A2(n13835), .ZN(n13836) );
  INV_X1 U15802 ( .A(n13837), .ZN(n13952) );
  OR2_X1 U15803 ( .A1(n14106), .A2(n13952), .ZN(n13838) );
  NOR2_X1 U15805 ( .A1(n14085), .A2(n13880), .ZN(n13841) );
  OAI22_X1 U15806 ( .A1(n6475), .A2(n13841), .B1(n13869), .B2(n13851), .ZN(
        n13843) );
  XNOR2_X1 U15807 ( .A(n13843), .B(n13842), .ZN(n14080) );
  INV_X1 U15808 ( .A(n13844), .ZN(n14075) );
  AOI21_X1 U15809 ( .B1(n13868), .B2(n13844), .A(n14576), .ZN(n13846) );
  NAND2_X1 U15810 ( .A1(n14072), .A2(n14247), .ZN(n13855) );
  NAND2_X1 U15811 ( .A1(n13848), .A2(n13847), .ZN(n14074) );
  OAI22_X1 U15812 ( .A1(n13850), .A2(n14074), .B1(n13849), .B2(n15144), .ZN(
        n13853) );
  NAND2_X1 U15813 ( .A1(n13851), .A2(n14252), .ZN(n14073) );
  NOR2_X1 U15814 ( .A1(n14042), .A2(n14073), .ZN(n13852) );
  AOI211_X1 U15815 ( .C1(n14258), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13853), 
        .B(n13852), .ZN(n13854) );
  OAI211_X1 U15816 ( .C1(n14075), .C2(n14260), .A(n13855), .B(n13854), .ZN(
        n13856) );
  AOI21_X1 U15817 ( .B1(n14080), .B2(n13863), .A(n13856), .ZN(n13857) );
  OAI21_X1 U15818 ( .B1(n14082), .B2(n14065), .A(n13857), .ZN(P1_U3356) );
  AND2_X1 U15819 ( .A1(n13859), .A2(n13858), .ZN(n13860) );
  NOR2_X1 U15820 ( .A1(n13861), .A2(n13860), .ZN(n14086) );
  INV_X1 U15821 ( .A(n14086), .ZN(n13874) );
  XNOR2_X1 U15822 ( .A(n6475), .B(n13862), .ZN(n14083) );
  NAND2_X1 U15823 ( .A1(n14083), .A2(n13863), .ZN(n13873) );
  INV_X1 U15824 ( .A(n13864), .ZN(n13865) );
  AOI22_X1 U15825 ( .A1(n15146), .A2(n14084), .B1(n13865), .B2(n14040), .ZN(
        n13866) );
  OAI21_X1 U15826 ( .B1(n13867), .B2(n15146), .A(n13866), .ZN(n13871) );
  OAI211_X1 U15827 ( .C1(n13869), .C2(n13887), .A(n14548), .B(n13868), .ZN(
        n14087) );
  NOR2_X1 U15828 ( .A1(n14087), .A2(n13998), .ZN(n13870) );
  AOI211_X1 U15829 ( .C1(n15149), .C2(n14085), .A(n13871), .B(n13870), .ZN(
        n13872) );
  OAI211_X1 U15830 ( .C1(n14065), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        P1_U3265) );
  XNOR2_X1 U15831 ( .A(n13875), .B(n13876), .ZN(n14095) );
  OAI21_X2 U15832 ( .B1(n13879), .B2(n6505), .A(n13878), .ZN(n13884) );
  AOI21_X1 U15833 ( .B1(n13851), .B2(n14254), .A(n13882), .ZN(n13883) );
  NAND2_X1 U15834 ( .A1(n14093), .A2(n13897), .ZN(n13885) );
  NAND2_X1 U15835 ( .A1(n13885), .A2(n14548), .ZN(n13886) );
  NOR2_X1 U15836 ( .A1(n13887), .A2(n13886), .ZN(n14092) );
  NAND2_X1 U15837 ( .A1(n14092), .A2(n14247), .ZN(n13892) );
  NAND2_X1 U15838 ( .A1(n14042), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n13888) );
  OAI21_X1 U15839 ( .B1(n15144), .B2(n13889), .A(n13888), .ZN(n13890) );
  AOI21_X1 U15840 ( .B1(n14093), .B2(n15149), .A(n13890), .ZN(n13891) );
  NAND2_X1 U15841 ( .A1(n13892), .A2(n13891), .ZN(n13893) );
  AOI21_X1 U15842 ( .B1(n14091), .B2(n15146), .A(n13893), .ZN(n13894) );
  OAI21_X1 U15843 ( .B1(n14095), .B2(n14065), .A(n13894), .ZN(P1_U3266) );
  XNOR2_X1 U15844 ( .A(n13895), .B(n13904), .ZN(n14102) );
  AOI21_X1 U15845 ( .B1(n14098), .B2(n13909), .A(n14576), .ZN(n13896) );
  AND2_X1 U15846 ( .A1(n13897), .A2(n13896), .ZN(n14096) );
  INV_X1 U15847 ( .A(n13898), .ZN(n13899) );
  AOI21_X1 U15848 ( .B1(n14040), .B2(n13899), .A(n14097), .ZN(n13902) );
  NAND2_X1 U15849 ( .A1(n14098), .A2(n15149), .ZN(n13901) );
  NAND2_X1 U15850 ( .A1(n14042), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n13900) );
  OAI211_X1 U15851 ( .C1(n14258), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        n13903) );
  AOI21_X1 U15852 ( .B1(n14096), .B2(n14247), .A(n13903), .ZN(n13907) );
  XOR2_X1 U15853 ( .A(n13905), .B(n13904), .Z(n14099) );
  NAND2_X1 U15854 ( .A1(n14099), .A2(n14248), .ZN(n13906) );
  OAI211_X1 U15855 ( .C1(n14102), .C2(n13978), .A(n13907), .B(n13906), .ZN(
        P1_U3267) );
  AOI21_X1 U15856 ( .B1(n13924), .B2(n13942), .A(n14576), .ZN(n13910) );
  NAND2_X1 U15857 ( .A1(n13910), .A2(n13909), .ZN(n14103) );
  XNOR2_X1 U15858 ( .A(n13911), .B(n13914), .ZN(n13912) );
  NAND2_X1 U15859 ( .A1(n13912), .A2(n14554), .ZN(n13920) );
  OAI211_X1 U15860 ( .C1(n13915), .C2(n13914), .A(n13913), .B(n14597), .ZN(
        n13918) );
  INV_X1 U15861 ( .A(n13916), .ZN(n13917) );
  AND2_X1 U15862 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  NAND2_X1 U15863 ( .A1(n13920), .A2(n13919), .ZN(n14105) );
  NAND2_X1 U15864 ( .A1(n14105), .A2(n15146), .ZN(n13926) );
  OAI22_X1 U15865 ( .A1(n15146), .A2(n13922), .B1(n13921), .B2(n15144), .ZN(
        n13923) );
  AOI21_X1 U15866 ( .B1(n13924), .B2(n15149), .A(n13923), .ZN(n13925) );
  OAI211_X1 U15867 ( .C1(n14103), .C2(n13998), .A(n13926), .B(n13925), .ZN(
        P1_U3268) );
  OAI21_X1 U15868 ( .B1(n13929), .B2(n13928), .A(n13927), .ZN(n13938) );
  OAI211_X1 U15869 ( .C1(n13932), .C2(n13931), .A(n13930), .B(n14554), .ZN(
        n13936) );
  AOI22_X1 U15870 ( .A1(n14252), .A2(n13934), .B1(n13933), .B2(n14254), .ZN(
        n13935) );
  NAND2_X1 U15871 ( .A1(n13936), .A2(n13935), .ZN(n13937) );
  AOI21_X1 U15872 ( .B1(n14597), .B2(n13938), .A(n13937), .ZN(n14108) );
  NAND2_X1 U15873 ( .A1(n14042), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n13939) );
  OAI21_X1 U15874 ( .B1(n15144), .B2(n13940), .A(n13939), .ZN(n13941) );
  AOI21_X1 U15875 ( .B1(n14106), .B2(n15149), .A(n13941), .ZN(n13945) );
  AOI21_X1 U15876 ( .B1(n14106), .B2(n13947), .A(n14576), .ZN(n13943) );
  NAND2_X1 U15877 ( .A1(n13943), .A2(n13942), .ZN(n14107) );
  OR2_X1 U15878 ( .A1(n14107), .A2(n13998), .ZN(n13944) );
  OAI211_X1 U15879 ( .C1(n14108), .C2(n14042), .A(n13945), .B(n13944), .ZN(
        P1_U3269) );
  XOR2_X1 U15880 ( .A(n13946), .B(n13961), .Z(n14116) );
  INV_X1 U15881 ( .A(n13947), .ZN(n13948) );
  AOI211_X1 U15882 ( .C1(n14112), .C2(n13967), .A(n14576), .B(n13948), .ZN(
        n14110) );
  NAND2_X1 U15883 ( .A1(n14112), .A2(n15149), .ZN(n13956) );
  OAI22_X1 U15884 ( .A1(n13952), .A2(n13951), .B1(n13950), .B2(n13949), .ZN(
        n14111) );
  INV_X1 U15885 ( .A(n13953), .ZN(n13954) );
  AOI22_X1 U15886 ( .A1(n15146), .A2(n14111), .B1(n13954), .B2(n14040), .ZN(
        n13955) );
  OAI211_X1 U15887 ( .C1(n15146), .C2(n13957), .A(n13956), .B(n13955), .ZN(
        n13958) );
  AOI21_X1 U15888 ( .B1(n14110), .B2(n14247), .A(n13958), .ZN(n13963) );
  AOI21_X1 U15889 ( .B1(n13961), .B2(n13960), .A(n13959), .ZN(n14113) );
  NAND2_X1 U15890 ( .A1(n14113), .A2(n14248), .ZN(n13962) );
  OAI211_X1 U15891 ( .C1(n14116), .C2(n13978), .A(n13963), .B(n13962), .ZN(
        P1_U3270) );
  INV_X1 U15892 ( .A(n13964), .ZN(n13965) );
  AOI21_X1 U15893 ( .B1(n13974), .B2(n13966), .A(n13965), .ZN(n14124) );
  AOI21_X1 U15894 ( .B1(n14120), .B2(n13979), .A(n14576), .ZN(n13968) );
  AND2_X1 U15895 ( .A1(n13968), .A2(n13967), .ZN(n14118) );
  NAND2_X1 U15896 ( .A1(n14120), .A2(n15149), .ZN(n13971) );
  AOI22_X1 U15897 ( .A1(n14042), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n13969), 
        .B2(n14040), .ZN(n13970) );
  OAI211_X1 U15898 ( .C1(n14258), .C2(n14117), .A(n13971), .B(n13970), .ZN(
        n13972) );
  AOI21_X1 U15899 ( .B1(n14118), .B2(n14247), .A(n13972), .ZN(n13977) );
  OAI21_X1 U15900 ( .B1(n13975), .B2(n13974), .A(n13973), .ZN(n14121) );
  NAND2_X1 U15901 ( .A1(n14121), .A2(n14248), .ZN(n13976) );
  OAI211_X1 U15902 ( .C1(n14124), .C2(n13978), .A(n13977), .B(n13976), .ZN(
        P1_U3271) );
  AOI21_X1 U15903 ( .B1(n14006), .B2(n14125), .A(n14576), .ZN(n13980) );
  NAND2_X1 U15904 ( .A1(n13980), .A2(n13979), .ZN(n14126) );
  OAI211_X1 U15905 ( .C1(n13983), .C2(n13982), .A(n13981), .B(n14554), .ZN(
        n13992) );
  AOI22_X1 U15906 ( .A1(n14022), .A2(n14252), .B1(n14254), .B2(n13984), .ZN(
        n13991) );
  INV_X1 U15907 ( .A(n13985), .ZN(n13989) );
  AOI21_X1 U15908 ( .B1(n14012), .B2(n13987), .A(n13986), .ZN(n13988) );
  OAI21_X1 U15909 ( .B1(n13989), .B2(n13988), .A(n14597), .ZN(n13990) );
  OR2_X1 U15910 ( .A1(n14127), .A2(n14042), .ZN(n13997) );
  NAND2_X1 U15911 ( .A1(n14042), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n13993) );
  OAI21_X1 U15912 ( .B1(n15144), .B2(n13994), .A(n13993), .ZN(n13995) );
  AOI21_X1 U15913 ( .B1(n14125), .B2(n15149), .A(n13995), .ZN(n13996) );
  OAI211_X1 U15914 ( .C1(n14126), .C2(n13998), .A(n13997), .B(n13996), .ZN(
        P1_U3272) );
  OAI211_X1 U15915 ( .C1(n6538), .C2(n14000), .A(n13999), .B(n14554), .ZN(
        n14004) );
  AOI22_X1 U15916 ( .A1(n14002), .A2(n14254), .B1(n14252), .B2(n14001), .ZN(
        n14003) );
  AND2_X1 U15917 ( .A1(n14004), .A2(n14003), .ZN(n14132) );
  INV_X1 U15918 ( .A(n14006), .ZN(n14007) );
  AOI211_X1 U15919 ( .C1(n14130), .C2(n14017), .A(n14576), .B(n14007), .ZN(
        n14129) );
  INV_X1 U15920 ( .A(n14008), .ZN(n14009) );
  AOI22_X1 U15921 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n14042), .B1(n14009), 
        .B2(n14040), .ZN(n14010) );
  OAI21_X1 U15922 ( .B1(n14011), .B2(n14260), .A(n14010), .ZN(n14015) );
  OAI21_X1 U15923 ( .B1(n6561), .B2(n14013), .A(n14012), .ZN(n14133) );
  NOR2_X1 U15924 ( .A1(n14133), .A2(n14065), .ZN(n14014) );
  AOI211_X1 U15925 ( .C1(n14129), .C2(n14247), .A(n14015), .B(n14014), .ZN(
        n14016) );
  OAI21_X1 U15926 ( .B1(n14258), .B2(n14132), .A(n14016), .ZN(P1_U3273) );
  AOI21_X1 U15927 ( .B1(n14134), .B2(n14039), .A(n14005), .ZN(n14135) );
  OAI21_X1 U15928 ( .B1(n14020), .B2(n14019), .A(n14018), .ZN(n14023) );
  INV_X1 U15929 ( .A(n14137), .ZN(n14024) );
  AOI21_X1 U15930 ( .B1(n14025), .B2(n14135), .A(n14024), .ZN(n14032) );
  INV_X1 U15931 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14027) );
  OAI22_X1 U15932 ( .A1(n15146), .A2(n14027), .B1(n14026), .B2(n15144), .ZN(
        n14030) );
  XNOR2_X1 U15933 ( .A(n14028), .B(n7130), .ZN(n14138) );
  NOR2_X1 U15934 ( .A1(n14138), .A2(n14065), .ZN(n14029) );
  AOI211_X1 U15935 ( .C1(n15149), .C2(n14134), .A(n14030), .B(n14029), .ZN(
        n14031) );
  OAI21_X1 U15936 ( .B1(n14032), .B2(n14042), .A(n14031), .ZN(P1_U3274) );
  XNOR2_X1 U15937 ( .A(n14033), .B(n6521), .ZN(n14143) );
  OAI211_X1 U15938 ( .C1(n14035), .C2(n6521), .A(n14034), .B(n14554), .ZN(
        n14037) );
  NAND2_X1 U15939 ( .A1(n14037), .A2(n14036), .ZN(n14139) );
  OR2_X1 U15940 ( .A1(n14045), .A2(n14057), .ZN(n14038) );
  AND3_X1 U15941 ( .A1(n14039), .A2(n14038), .A3(n14548), .ZN(n14140) );
  NAND2_X1 U15942 ( .A1(n14140), .A2(n14247), .ZN(n14044) );
  AOI22_X1 U15943 ( .A1(n14042), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14041), 
        .B2(n14040), .ZN(n14043) );
  OAI211_X1 U15944 ( .C1(n14045), .C2(n14260), .A(n14044), .B(n14043), .ZN(
        n14046) );
  AOI21_X1 U15945 ( .B1(n14139), .B2(n15146), .A(n14046), .ZN(n14047) );
  OAI21_X1 U15946 ( .B1(n14143), .B2(n14065), .A(n14047), .ZN(P1_U3275) );
  XNOR2_X1 U15947 ( .A(n14048), .B(n14050), .ZN(n14148) );
  OAI211_X1 U15948 ( .C1(n14050), .C2(n6567), .A(n14049), .B(n14554), .ZN(
        n14053) );
  INV_X1 U15949 ( .A(n14051), .ZN(n14052) );
  NAND2_X1 U15950 ( .A1(n14053), .A2(n14052), .ZN(n14144) );
  NAND2_X1 U15951 ( .A1(n14054), .A2(n14146), .ZN(n14055) );
  NAND2_X1 U15952 ( .A1(n14055), .A2(n14548), .ZN(n14056) );
  NOR2_X1 U15953 ( .A1(n14057), .A2(n14056), .ZN(n14145) );
  NAND2_X1 U15954 ( .A1(n14145), .A2(n14247), .ZN(n14062) );
  NAND2_X1 U15955 ( .A1(n14258), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14058) );
  OAI21_X1 U15956 ( .B1(n15144), .B2(n14059), .A(n14058), .ZN(n14060) );
  AOI21_X1 U15957 ( .B1(n14146), .B2(n15149), .A(n14060), .ZN(n14061) );
  NAND2_X1 U15958 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  AOI21_X1 U15959 ( .B1(n14144), .B2(n15146), .A(n14063), .ZN(n14064) );
  OAI21_X1 U15960 ( .B1(n14148), .B2(n14065), .A(n14064), .ZN(P1_U3276) );
  NAND2_X1 U15961 ( .A1(n14066), .A2(n14548), .ZN(n14067) );
  OAI211_X1 U15962 ( .C1(n14068), .C2(n14592), .A(n14067), .B(n14069), .ZN(
        n14162) );
  MUX2_X1 U15963 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14162), .S(n14615), .Z(
        P1_U3559) );
  OAI211_X1 U15964 ( .C1(n14071), .C2(n14592), .A(n14070), .B(n14069), .ZN(
        n14163) );
  MUX2_X1 U15965 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14163), .S(n14615), .Z(
        P1_U3558) );
  OAI211_X1 U15966 ( .C1(n14075), .C2(n14592), .A(n14074), .B(n14073), .ZN(
        n14076) );
  INV_X1 U15967 ( .A(n14076), .ZN(n14077) );
  OAI21_X1 U15968 ( .B1(n14082), .B2(n14578), .A(n14081), .ZN(n14164) );
  MUX2_X1 U15969 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14164), .S(n14615), .Z(
        P1_U3557) );
  NAND2_X1 U15970 ( .A1(n14083), .A2(n14554), .ZN(n14090) );
  AOI21_X1 U15971 ( .B1(n14085), .B2(n14588), .A(n14084), .ZN(n14089) );
  NAND2_X1 U15972 ( .A1(n14086), .A2(n14597), .ZN(n14088) );
  NAND4_X1 U15973 ( .A1(n14090), .A2(n14089), .A3(n14088), .A4(n14087), .ZN(
        n14165) );
  MUX2_X1 U15974 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14165), .S(n14615), .Z(
        P1_U3556) );
  OAI21_X1 U15975 ( .B1(n14095), .B2(n14578), .A(n14094), .ZN(n14166) );
  MUX2_X1 U15976 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14166), .S(n14615), .Z(
        P1_U3555) );
  AOI211_X1 U15977 ( .C1(n14588), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        n14101) );
  NAND2_X1 U15978 ( .A1(n14099), .A2(n14597), .ZN(n14100) );
  OAI211_X1 U15979 ( .C1(n14102), .C2(n14571), .A(n14101), .B(n14100), .ZN(
        n14167) );
  MUX2_X1 U15980 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14167), .S(n14615), .Z(
        P1_U3554) );
  OAI21_X1 U15981 ( .B1(n13788), .B2(n14592), .A(n14103), .ZN(n14104) );
  MUX2_X1 U15982 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14168), .S(n14615), .Z(
        P1_U3553) );
  INV_X1 U15983 ( .A(n14106), .ZN(n14109) );
  OAI211_X1 U15984 ( .C1(n14109), .C2(n14592), .A(n14108), .B(n14107), .ZN(
        n14169) );
  MUX2_X1 U15985 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14169), .S(n14615), .Z(
        P1_U3552) );
  AOI211_X1 U15986 ( .C1(n14588), .C2(n14112), .A(n14111), .B(n14110), .ZN(
        n14115) );
  NAND2_X1 U15987 ( .A1(n14113), .A2(n14597), .ZN(n14114) );
  OAI211_X1 U15988 ( .C1(n14116), .C2(n14571), .A(n14115), .B(n14114), .ZN(
        n14170) );
  MUX2_X1 U15989 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14170), .S(n14615), .Z(
        P1_U3551) );
  INV_X1 U15990 ( .A(n14117), .ZN(n14119) );
  AOI211_X1 U15991 ( .C1(n14588), .C2(n14120), .A(n14119), .B(n14118), .ZN(
        n14123) );
  NAND2_X1 U15992 ( .A1(n14121), .A2(n14597), .ZN(n14122) );
  OAI211_X1 U15993 ( .C1(n14124), .C2(n14571), .A(n14123), .B(n14122), .ZN(
        n14171) );
  MUX2_X1 U15994 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14171), .S(n14615), .Z(
        P1_U3550) );
  INV_X1 U15995 ( .A(n14125), .ZN(n14128) );
  OAI211_X1 U15996 ( .C1(n14128), .C2(n14592), .A(n14127), .B(n14126), .ZN(
        n14172) );
  MUX2_X1 U15997 ( .A(n14172), .B(P1_REG1_REG_21__SCAN_IN), .S(n14613), .Z(
        P1_U3549) );
  AOI21_X1 U15998 ( .B1(n14588), .B2(n14130), .A(n14129), .ZN(n14131) );
  OAI211_X1 U15999 ( .C1(n14578), .C2(n14133), .A(n14132), .B(n14131), .ZN(
        n14173) );
  MUX2_X1 U16000 ( .A(n14173), .B(P1_REG1_REG_20__SCAN_IN), .S(n14613), .Z(
        P1_U3548) );
  AOI22_X1 U16001 ( .A1(n14135), .A2(n14548), .B1(n14588), .B2(n14134), .ZN(
        n14136) );
  OAI211_X1 U16002 ( .C1(n14138), .C2(n14578), .A(n14137), .B(n14136), .ZN(
        n14174) );
  MUX2_X1 U16003 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14174), .S(n14615), .Z(
        P1_U3547) );
  AOI211_X1 U16004 ( .C1(n14588), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14142) );
  OAI21_X1 U16005 ( .B1(n14143), .B2(n14578), .A(n14142), .ZN(n14175) );
  MUX2_X1 U16006 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14175), .S(n14615), .Z(
        P1_U3546) );
  AOI211_X1 U16007 ( .C1(n14588), .C2(n14146), .A(n14145), .B(n14144), .ZN(
        n14147) );
  OAI21_X1 U16008 ( .B1(n14148), .B2(n14578), .A(n14147), .ZN(n14176) );
  MUX2_X1 U16009 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14176), .S(n14615), .Z(
        P1_U3545) );
  INV_X1 U16010 ( .A(n14149), .ZN(n14388) );
  OAI21_X1 U16011 ( .B1(n14388), .B2(n14592), .A(n14150), .ZN(n14151) );
  AOI21_X1 U16012 ( .B1(n14152), .B2(n14597), .A(n14151), .ZN(n14153) );
  NAND2_X1 U16013 ( .A1(n14154), .A2(n14153), .ZN(n14177) );
  MUX2_X1 U16014 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14177), .S(n14615), .Z(
        P1_U3544) );
  OAI21_X1 U16015 ( .B1(n11614), .B2(n14592), .A(n14155), .ZN(n14158) );
  NOR2_X1 U16016 ( .A1(n14156), .A2(n14571), .ZN(n14157) );
  AOI211_X1 U16017 ( .C1(n14548), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        n14160) );
  OAI21_X1 U16018 ( .B1(n14578), .B2(n14161), .A(n14160), .ZN(n14178) );
  MUX2_X1 U16019 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14178), .S(n14615), .Z(
        P1_U3543) );
  MUX2_X1 U16020 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14162), .S(n14601), .Z(
        P1_U3527) );
  MUX2_X1 U16021 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14163), .S(n14601), .Z(
        P1_U3526) );
  MUX2_X1 U16022 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14164), .S(n14601), .Z(
        P1_U3525) );
  MUX2_X1 U16023 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14165), .S(n14601), .Z(
        P1_U3524) );
  MUX2_X1 U16024 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14166), .S(n14601), .Z(
        P1_U3523) );
  MUX2_X1 U16025 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14167), .S(n14601), .Z(
        P1_U3522) );
  MUX2_X1 U16026 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14168), .S(n14601), .Z(
        P1_U3521) );
  MUX2_X1 U16027 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14169), .S(n14601), .Z(
        P1_U3520) );
  MUX2_X1 U16028 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14170), .S(n14601), .Z(
        P1_U3519) );
  MUX2_X1 U16029 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14171), .S(n14601), .Z(
        P1_U3518) );
  MUX2_X1 U16030 ( .A(n14172), .B(P1_REG0_REG_21__SCAN_IN), .S(n14599), .Z(
        P1_U3517) );
  MUX2_X1 U16031 ( .A(n14173), .B(P1_REG0_REG_20__SCAN_IN), .S(n14599), .Z(
        P1_U3516) );
  MUX2_X1 U16032 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14174), .S(n14601), .Z(
        P1_U3515) );
  MUX2_X1 U16033 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14175), .S(n14601), .Z(
        P1_U3513) );
  MUX2_X1 U16034 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14176), .S(n14601), .Z(
        P1_U3510) );
  MUX2_X1 U16035 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14177), .S(n14601), .Z(
        P1_U3507) );
  MUX2_X1 U16036 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14178), .S(n14601), .Z(
        P1_U3504) );
  NAND3_X1 U16037 ( .A1(n14179), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14181) );
  OAI22_X1 U16038 ( .A1(n14182), .A2(n14181), .B1(n14180), .B2(n14195), .ZN(
        n14183) );
  AOI21_X1 U16039 ( .B1(n14185), .B2(n14184), .A(n14183), .ZN(n14186) );
  INV_X1 U16040 ( .A(n14186), .ZN(P1_U3324) );
  OAI222_X1 U16041 ( .A1(P1_U3086), .A2(n8260), .B1(n14198), .B2(n14188), .C1(
        n14187), .C2(n14195), .ZN(P1_U3325) );
  OAI222_X1 U16042 ( .A1(P1_U3086), .A2(n14191), .B1(n14198), .B2(n14190), 
        .C1(n14189), .C2(n14195), .ZN(P1_U3328) );
  OAI222_X1 U16043 ( .A1(P1_U3086), .A2(n14194), .B1(n14198), .B2(n14193), 
        .C1(n14192), .C2(n14195), .ZN(P1_U3329) );
  OAI222_X1 U16044 ( .A1(n9793), .A2(P1_U3086), .B1(n14198), .B2(n14197), .C1(
        n14196), .C2(n14195), .ZN(P1_U3330) );
  MUX2_X1 U16045 ( .A(n14200), .B(n14199), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16046 ( .A(n14201), .ZN(n14202) );
  MUX2_X1 U16047 ( .A(n14202), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16048 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14206) );
  OAI21_X1 U16049 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14206), 
        .ZN(U28) );
  AOI21_X1 U16050 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14207) );
  OAI21_X1 U16051 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14207), 
        .ZN(U29) );
  AOI22_X1 U16052 ( .A1(n14208), .A2(n14227), .B1(SI_17_), .B2(n14226), .ZN(
        n14209) );
  OAI21_X1 U16053 ( .B1(P3_U3151), .B2(n14210), .A(n14209), .ZN(P3_U3278) );
  AOI21_X1 U16054 ( .B1(n14213), .B2(n14212), .A(n14211), .ZN(SUB_1596_U61) );
  AOI22_X1 U16055 ( .A1(n14214), .A2(n14227), .B1(SI_13_), .B2(n14226), .ZN(
        n14215) );
  OAI21_X1 U16056 ( .B1(P3_U3151), .B2(n14216), .A(n14215), .ZN(P3_U3282) );
  AOI21_X1 U16057 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(SUB_1596_U57) );
  AOI22_X1 U16058 ( .A1(n14220), .A2(n14227), .B1(SI_16_), .B2(n14226), .ZN(
        n14221) );
  OAI21_X1 U16059 ( .B1(P3_U3151), .B2(n14222), .A(n14221), .ZN(P3_U3279) );
  OAI21_X1 U16060 ( .B1(n14225), .B2(n14224), .A(n14223), .ZN(SUB_1596_U55) );
  AOI22_X1 U16061 ( .A1(n14228), .A2(n14227), .B1(SI_18_), .B2(n14226), .ZN(
        n14229) );
  OAI21_X1 U16062 ( .B1(P3_U3151), .B2(n14230), .A(n14229), .ZN(P3_U3277) );
  AOI21_X1 U16063 ( .B1(n14654), .B2(n14233), .A(n14232), .ZN(SUB_1596_U54) );
  OAI21_X1 U16064 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14237) );
  XNOR2_X1 U16065 ( .A(n14237), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  AND2_X1 U16066 ( .A1(n14238), .A2(n14588), .ZN(n14370) );
  NOR3_X1 U16067 ( .A1(n14240), .A2(n14239), .A3(n14370), .ZN(n14242) );
  INV_X1 U16068 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U16069 ( .A1(n14601), .A2(n14242), .B1(n14241), .B2(n14599), .ZN(
        P1_U3495) );
  AOI22_X1 U16070 ( .A1(n14615), .A2(n14242), .B1(n10012), .B2(n14613), .ZN(
        P1_U3540) );
  XNOR2_X1 U16071 ( .A(n14243), .B(n14249), .ZN(n14437) );
  OAI211_X1 U16072 ( .C1(n14434), .C2(n14245), .A(n14548), .B(n14244), .ZN(
        n14433) );
  INV_X1 U16073 ( .A(n14433), .ZN(n14246) );
  AOI22_X1 U16074 ( .A1(n14437), .A2(n14248), .B1(n14247), .B2(n14246), .ZN(
        n14263) );
  XNOR2_X1 U16075 ( .A(n14250), .B(n14249), .ZN(n14251) );
  NAND2_X1 U16076 ( .A1(n14251), .A2(n14554), .ZN(n14256) );
  AOI22_X1 U16077 ( .A1(n14254), .A2(n14416), .B1(n14253), .B2(n14252), .ZN(
        n14255) );
  NAND2_X1 U16078 ( .A1(n14256), .A2(n14255), .ZN(n14435) );
  NOR2_X1 U16079 ( .A1(n15144), .A2(n14410), .ZN(n14257) );
  AOI21_X1 U16080 ( .B1(n14258), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14257), 
        .ZN(n14259) );
  OAI21_X1 U16081 ( .B1(n14434), .B2(n14260), .A(n14259), .ZN(n14261) );
  AOI21_X1 U16082 ( .B1(n14435), .B2(n15146), .A(n14261), .ZN(n14262) );
  NAND2_X1 U16083 ( .A1(n14263), .A2(n14262), .ZN(P1_U3280) );
  AOI21_X1 U16084 ( .B1(n14266), .B2(n14265), .A(n14264), .ZN(n14267) );
  XOR2_X1 U16085 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14267), .Z(SUB_1596_U63)
         );
  AOI22_X1 U16086 ( .A1(n14298), .A2(n14268), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14865), .ZN(n14269) );
  NAND2_X1 U16087 ( .A1(n14270), .A2(n14269), .ZN(P3_U3203) );
  XOR2_X1 U16088 ( .A(n14279), .B(n14271), .Z(n14274) );
  AOI222_X1 U16089 ( .A1(n14920), .A2(n14274), .B1(n14273), .B2(n14889), .C1(
        n14272), .C2(n14892), .ZN(n14299) );
  OAI22_X1 U16090 ( .A1(n14927), .A2(n14276), .B1(n14910), .B2(n14275), .ZN(
        n14277) );
  INV_X1 U16091 ( .A(n14277), .ZN(n14283) );
  XOR2_X1 U16092 ( .A(n14279), .B(n14278), .Z(n14302) );
  NOR2_X1 U16093 ( .A1(n14280), .A2(n14954), .ZN(n14301) );
  AOI22_X1 U16094 ( .A1(n14302), .A2(n14281), .B1(n14902), .B2(n14301), .ZN(
        n14282) );
  OAI211_X1 U16095 ( .C1(n14865), .C2(n14299), .A(n14283), .B(n14282), .ZN(
        P3_U3220) );
  XNOR2_X1 U16096 ( .A(n14285), .B(n14284), .ZN(n14311) );
  XNOR2_X1 U16097 ( .A(n14286), .B(n14287), .ZN(n14288) );
  OAI222_X1 U16098 ( .A1(n14917), .A2(n14290), .B1(n14915), .B2(n14289), .C1(
        n14288), .C2(n14877), .ZN(n14309) );
  AOI21_X1 U16099 ( .B1(n14311), .B2(n14291), .A(n14309), .ZN(n14296) );
  NOR2_X1 U16100 ( .A1(n14292), .A2(n14954), .ZN(n14310) );
  AOI22_X1 U16101 ( .A1(n14902), .A2(n14310), .B1(n14901), .B2(n14293), .ZN(
        n14294) );
  OAI221_X1 U16102 ( .B1(n14865), .B2(n14296), .C1(n14927), .C2(n14295), .A(
        n14294), .ZN(P3_U3222) );
  AOI21_X1 U16103 ( .B1(n14298), .B2(n14907), .A(n14297), .ZN(n14314) );
  INV_X1 U16104 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16105 ( .A1(n14993), .A2(n14314), .B1(n15115), .B2(n14990), .ZN(
        P3_U3489) );
  INV_X1 U16106 ( .A(n14299), .ZN(n14300) );
  AOI211_X1 U16107 ( .C1(n14302), .C2(n14972), .A(n14301), .B(n14300), .ZN(
        n14316) );
  INV_X1 U16108 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U16109 ( .A1(n14993), .A2(n14316), .B1(n14303), .B2(n14990), .ZN(
        P3_U3472) );
  OAI21_X1 U16110 ( .B1(n14306), .B2(n14305), .A(n14304), .ZN(n14307) );
  NOR2_X1 U16111 ( .A1(n14308), .A2(n14307), .ZN(n14318) );
  AOI22_X1 U16112 ( .A1(n14993), .A2(n14318), .B1(n11528), .B2(n14990), .ZN(
        P3_U3471) );
  AOI211_X1 U16113 ( .C1(n14311), .C2(n14972), .A(n14310), .B(n14309), .ZN(
        n14320) );
  INV_X1 U16114 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U16115 ( .A1(n14993), .A2(n14320), .B1(n14312), .B2(n14990), .ZN(
        P3_U3470) );
  INV_X1 U16116 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U16117 ( .A1(n14975), .A2(n14314), .B1(n14313), .B2(n14973), .ZN(
        P3_U3457) );
  INV_X1 U16118 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U16119 ( .A1(n14975), .A2(n14316), .B1(n14315), .B2(n14973), .ZN(
        P3_U3429) );
  INV_X1 U16120 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U16121 ( .A1(n14975), .A2(n14318), .B1(n14317), .B2(n14973), .ZN(
        P3_U3426) );
  INV_X1 U16122 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U16123 ( .A1(n14975), .A2(n14320), .B1(n14319), .B2(n14973), .ZN(
        P3_U3423) );
  INV_X1 U16124 ( .A(n14321), .ZN(n14324) );
  OAI211_X1 U16125 ( .C1(n14324), .C2(n14764), .A(n14323), .B(n14322), .ZN(
        n14328) );
  NOR3_X1 U16126 ( .A1(n14326), .A2(n14325), .A3(n14749), .ZN(n14327) );
  AOI211_X1 U16127 ( .C1(n14329), .C2(n14753), .A(n14328), .B(n14327), .ZN(
        n14354) );
  AOI22_X1 U16128 ( .A1(n6436), .A2(n14354), .B1(n14330), .B2(n14776), .ZN(
        P2_U3515) );
  AOI21_X1 U16129 ( .B1(n14332), .B2(n13261), .A(n14331), .ZN(n14334) );
  OAI211_X1 U16130 ( .C1(n14335), .C2(n14749), .A(n14334), .B(n14333), .ZN(
        n14336) );
  AOI21_X1 U16131 ( .B1(n14337), .B2(n14753), .A(n14336), .ZN(n14356) );
  AOI22_X1 U16132 ( .A1(n6436), .A2(n14356), .B1(n9369), .B2(n14776), .ZN(
        P2_U3514) );
  AOI21_X1 U16133 ( .B1(n14339), .B2(n13261), .A(n14338), .ZN(n14341) );
  OAI211_X1 U16134 ( .C1(n14342), .C2(n14749), .A(n14341), .B(n14340), .ZN(
        n14343) );
  AOI21_X1 U16135 ( .B1(n14344), .B2(n14753), .A(n14343), .ZN(n14357) );
  AOI22_X1 U16136 ( .A1(n6436), .A2(n14357), .B1(n11449), .B2(n14776), .ZN(
        P2_U3512) );
  INV_X1 U16137 ( .A(n14345), .ZN(n14347) );
  OAI21_X1 U16138 ( .B1(n14347), .B2(n14764), .A(n14346), .ZN(n14348) );
  AOI21_X1 U16139 ( .B1(n14349), .B2(n14736), .A(n14348), .ZN(n14350) );
  AND2_X1 U16140 ( .A1(n14351), .A2(n14350), .ZN(n14358) );
  AOI22_X1 U16141 ( .A1(n6436), .A2(n14358), .B1(n14352), .B2(n14776), .ZN(
        P2_U3511) );
  INV_X1 U16142 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U16143 ( .A1(n14754), .A2(n14354), .B1(n14353), .B2(n14769), .ZN(
        P2_U3478) );
  INV_X1 U16144 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16145 ( .A1(n14754), .A2(n14356), .B1(n14355), .B2(n14769), .ZN(
        P2_U3475) );
  AOI22_X1 U16146 ( .A1(n14754), .A2(n14357), .B1(n9335), .B2(n14769), .ZN(
        P2_U3469) );
  AOI22_X1 U16147 ( .A1(n14754), .A2(n14358), .B1(n9315), .B2(n14769), .ZN(
        P2_U3466) );
  AOI21_X1 U16148 ( .B1(n14360), .B2(n14359), .A(n6562), .ZN(n14364) );
  AOI22_X1 U16149 ( .A1(n14417), .A2(n14361), .B1(n14415), .B2(n14386), .ZN(
        n14363) );
  NAND2_X1 U16150 ( .A1(n14428), .A2(n14407), .ZN(n14362) );
  OAI211_X1 U16151 ( .C1(n14364), .C2(n14401), .A(n14363), .B(n14362), .ZN(
        n14365) );
  INV_X1 U16152 ( .A(n14365), .ZN(n14367) );
  OAI211_X1 U16153 ( .C1(n14425), .C2(n14368), .A(n14367), .B(n14366), .ZN(
        P1_U3215) );
  AOI22_X1 U16154 ( .A1(n14370), .A2(n14369), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14381) );
  INV_X1 U16155 ( .A(n14400), .ZN(n14376) );
  AOI21_X1 U16156 ( .B1(n14371), .B2(n14400), .A(n14375), .ZN(n14373) );
  NOR2_X1 U16157 ( .A1(n14373), .A2(n7032), .ZN(n14374) );
  AOI211_X1 U16158 ( .C1(n14376), .C2(n14375), .A(n14401), .B(n14374), .ZN(
        n14377) );
  AOI21_X1 U16159 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14380) );
  OAI211_X1 U16160 ( .C1(n14382), .C2(n14425), .A(n14381), .B(n14380), .ZN(
        P1_U3224) );
  XNOR2_X1 U16161 ( .A(n14383), .B(n14384), .ZN(n14390) );
  AOI22_X1 U16162 ( .A1(n14417), .A2(n14386), .B1(n14415), .B2(n14385), .ZN(
        n14387) );
  OAI21_X1 U16163 ( .B1(n14388), .B2(n14419), .A(n14387), .ZN(n14389) );
  AOI21_X1 U16164 ( .B1(n14390), .B2(n14421), .A(n14389), .ZN(n14392) );
  OAI211_X1 U16165 ( .C1(n14425), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U3226) );
  OAI22_X1 U16166 ( .A1(n14397), .A2(n14396), .B1(n14395), .B2(n14394), .ZN(
        n14405) );
  INV_X1 U16167 ( .A(n14398), .ZN(n14403) );
  AOI21_X1 U16168 ( .B1(n14372), .B2(n14400), .A(n14399), .ZN(n14402) );
  NOR3_X1 U16169 ( .A1(n14403), .A2(n14402), .A3(n14401), .ZN(n14404) );
  AOI211_X1 U16170 ( .C1(n14407), .C2(n14406), .A(n14405), .B(n14404), .ZN(
        n14409) );
  OAI211_X1 U16171 ( .C1(n14425), .C2(n14410), .A(n14409), .B(n14408), .ZN(
        P1_U3234) );
  OAI21_X1 U16172 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14422) );
  AOI22_X1 U16173 ( .A1(n14417), .A2(n14416), .B1(n14415), .B2(n14414), .ZN(
        n14418) );
  OAI21_X1 U16174 ( .B1(n11614), .B2(n14419), .A(n14418), .ZN(n14420) );
  AOI21_X1 U16175 ( .B1(n14422), .B2(n14421), .A(n14420), .ZN(n14423) );
  NAND2_X1 U16176 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14512)
         );
  OAI211_X1 U16177 ( .C1(n14425), .C2(n14424), .A(n14423), .B(n14512), .ZN(
        P1_U3241) );
  AOI211_X1 U16178 ( .C1(n14588), .C2(n14428), .A(n14427), .B(n14426), .ZN(
        n14429) );
  OAI21_X1 U16179 ( .B1(n14578), .B2(n14430), .A(n14429), .ZN(n14431) );
  AOI21_X1 U16180 ( .B1(n14554), .B2(n14432), .A(n14431), .ZN(n14445) );
  AOI22_X1 U16181 ( .A1(n14615), .A2(n14445), .B1(n15088), .B2(n14613), .ZN(
        P1_U3542) );
  OAI21_X1 U16182 ( .B1(n14434), .B2(n14592), .A(n14433), .ZN(n14436) );
  AOI211_X1 U16183 ( .C1(n14597), .C2(n14437), .A(n14436), .B(n14435), .ZN(
        n14447) );
  AOI22_X1 U16184 ( .A1(n14615), .A2(n14447), .B1(n10221), .B2(n14613), .ZN(
        P1_U3541) );
  OAI211_X1 U16185 ( .C1(n6870), .C2(n14592), .A(n14439), .B(n14438), .ZN(
        n14442) );
  NOR2_X1 U16186 ( .A1(n14440), .A2(n14578), .ZN(n14441) );
  AOI211_X1 U16187 ( .C1(n14443), .C2(n14554), .A(n14442), .B(n14441), .ZN(
        n14449) );
  AOI22_X1 U16188 ( .A1(n14615), .A2(n14449), .B1(n8443), .B2(n14613), .ZN(
        P1_U3539) );
  INV_X1 U16189 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U16190 ( .A1(n14601), .A2(n14445), .B1(n14444), .B2(n14599), .ZN(
        P1_U3501) );
  INV_X1 U16191 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U16192 ( .A1(n14601), .A2(n14447), .B1(n14446), .B2(n14599), .ZN(
        P1_U3498) );
  INV_X1 U16193 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16194 ( .A1(n14601), .A2(n14449), .B1(n14448), .B2(n14599), .ZN(
        P1_U3492) );
  OAI21_X1 U16195 ( .B1(n14452), .B2(n14451), .A(n14450), .ZN(n14453) );
  XNOR2_X1 U16196 ( .A(n14453), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16197 ( .A1(n14458), .A2(n14457), .B1(n14458), .B2(n14456), .C1(
        n14455), .C2(n14454), .ZN(SUB_1596_U68) );
  OAI21_X1 U16198 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(SUB_1596_U67) );
  OAI21_X1 U16199 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14465) );
  XNOR2_X1 U16200 ( .A(n14465), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16201 ( .B1(n14468), .B2(n14467), .A(n14466), .ZN(n14469) );
  XOR2_X1 U16202 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14469), .Z(SUB_1596_U65)
         );
  INV_X1 U16203 ( .A(n14472), .ZN(n14471) );
  OAI222_X1 U16204 ( .A1(n14474), .A2(n14473), .B1(n14474), .B2(n14472), .C1(
        n14471), .C2(n14470), .ZN(SUB_1596_U64) );
  OAI21_X1 U16205 ( .B1(n14475), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6587), .ZN(
        n14477) );
  XNOR2_X1 U16206 ( .A(n14477), .B(n14476), .ZN(n14480) );
  AOI22_X1 U16207 ( .A1(n14497), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14478) );
  OAI21_X1 U16208 ( .B1(n14480), .B2(n14479), .A(n14478), .ZN(P1_U3243) );
  MUX2_X1 U16209 ( .A(n9826), .B(P1_REG1_REG_4__SCAN_IN), .S(n14493), .Z(
        n14483) );
  NAND3_X1 U16210 ( .A1(n14483), .A2(n14482), .A3(n14481), .ZN(n14484) );
  NAND3_X1 U16211 ( .A1(n14486), .A2(n14485), .A3(n14484), .ZN(n14501) );
  MUX2_X1 U16212 ( .A(n10612), .B(P1_REG2_REG_4__SCAN_IN), .S(n14493), .Z(
        n14489) );
  NAND3_X1 U16213 ( .A1(n14489), .A2(n14488), .A3(n14487), .ZN(n14490) );
  NAND3_X1 U16214 ( .A1(n14492), .A2(n14491), .A3(n14490), .ZN(n14500) );
  NAND2_X1 U16215 ( .A1(n14494), .A2(n14493), .ZN(n14499) );
  INV_X1 U16216 ( .A(n14495), .ZN(n14496) );
  AOI21_X1 U16217 ( .B1(n14497), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14496), .ZN(
        n14498) );
  AND4_X1 U16218 ( .A1(n14501), .A2(n14500), .A3(n14499), .A4(n14498), .ZN(
        n14503) );
  NAND2_X1 U16219 ( .A1(n14503), .A2(n14502), .ZN(P1_U3247) );
  AOI21_X1 U16220 ( .B1(n14505), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14504), 
        .ZN(n14509) );
  AOI21_X1 U16221 ( .B1(n14507), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14506), 
        .ZN(n14508) );
  OAI222_X1 U16222 ( .A1(n14524), .A2(n14510), .B1(n14522), .B2(n14509), .C1(
        n14520), .C2(n14508), .ZN(n14511) );
  INV_X1 U16223 ( .A(n14511), .ZN(n14513) );
  OAI211_X1 U16224 ( .C1(n14514), .C2(n14528), .A(n14513), .B(n14512), .ZN(
        P1_U3258) );
  OAI21_X1 U16225 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n14516), .A(n14515), 
        .ZN(n14521) );
  OAI21_X1 U16226 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n14518), .A(n14517), 
        .ZN(n14519) );
  OAI222_X1 U16227 ( .A1(n14524), .A2(n14523), .B1(n14522), .B2(n14521), .C1(
        n14520), .C2(n14519), .ZN(n14525) );
  INV_X1 U16228 ( .A(n14525), .ZN(n14527) );
  OAI211_X1 U16229 ( .C1(n14529), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        P1_U3261) );
  NOR2_X1 U16230 ( .A1(n14530), .A2(n15108), .ZN(P1_U3294) );
  AND2_X1 U16231 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14531), .ZN(P1_U3295) );
  AND2_X1 U16232 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14531), .ZN(P1_U3296) );
  AND2_X1 U16233 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14531), .ZN(P1_U3297) );
  AND2_X1 U16234 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14531), .ZN(P1_U3298) );
  AND2_X1 U16235 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14531), .ZN(P1_U3299) );
  AND2_X1 U16236 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14531), .ZN(P1_U3300) );
  AND2_X1 U16237 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14531), .ZN(P1_U3301) );
  AND2_X1 U16238 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14531), .ZN(P1_U3302) );
  AND2_X1 U16239 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14531), .ZN(P1_U3303) );
  AND2_X1 U16240 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14531), .ZN(P1_U3304) );
  AND2_X1 U16241 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14531), .ZN(P1_U3305) );
  AND2_X1 U16242 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14531), .ZN(P1_U3306) );
  AND2_X1 U16243 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14531), .ZN(P1_U3307) );
  AND2_X1 U16244 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14531), .ZN(P1_U3308) );
  AND2_X1 U16245 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14531), .ZN(P1_U3309) );
  AND2_X1 U16246 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14531), .ZN(P1_U3310) );
  AND2_X1 U16247 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14531), .ZN(P1_U3311) );
  AND2_X1 U16248 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14531), .ZN(P1_U3312) );
  AND2_X1 U16249 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14531), .ZN(P1_U3313) );
  NOR2_X1 U16250 ( .A1(n14530), .A2(n15131), .ZN(P1_U3314) );
  NOR2_X1 U16251 ( .A1(n14530), .A2(n15085), .ZN(P1_U3315) );
  AND2_X1 U16252 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14531), .ZN(P1_U3316) );
  AND2_X1 U16253 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14531), .ZN(P1_U3317) );
  AND2_X1 U16254 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14531), .ZN(P1_U3318) );
  AND2_X1 U16255 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14531), .ZN(P1_U3319) );
  AND2_X1 U16256 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14531), .ZN(P1_U3320) );
  NOR2_X1 U16257 ( .A1(n14530), .A2(n15123), .ZN(P1_U3321) );
  AND2_X1 U16258 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14531), .ZN(P1_U3322) );
  AND2_X1 U16259 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14531), .ZN(P1_U3323) );
  OAI22_X1 U16260 ( .A1(n14533), .A2(n14576), .B1(n14532), .B2(n14592), .ZN(
        n14536) );
  INV_X1 U16261 ( .A(n14534), .ZN(n14535) );
  AOI211_X1 U16262 ( .C1(n14597), .C2(n14537), .A(n14536), .B(n14535), .ZN(
        n14602) );
  INV_X1 U16263 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16264 ( .A1(n14601), .A2(n14602), .B1(n14538), .B2(n14599), .ZN(
        P1_U3462) );
  AOI211_X1 U16265 ( .C1(n14588), .C2(n8525), .A(n6579), .B(n14539), .ZN(
        n14603) );
  INV_X1 U16266 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U16267 ( .A1(n14601), .A2(n14603), .B1(n14540), .B2(n14599), .ZN(
        P1_U3465) );
  INV_X1 U16268 ( .A(n14541), .ZN(n14544) );
  OAI22_X1 U16269 ( .A1(n14542), .A2(n14576), .B1(n8735), .B2(n14592), .ZN(
        n14543) );
  NOR2_X1 U16270 ( .A1(n14544), .A2(n14543), .ZN(n14604) );
  INV_X1 U16271 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U16272 ( .A1(n14601), .A2(n14604), .B1(n14545), .B2(n14599), .ZN(
        P1_U3468) );
  AOI211_X1 U16273 ( .C1(n14549), .C2(n14548), .A(n14547), .B(n14546), .ZN(
        n14550) );
  OAI21_X1 U16274 ( .B1(n14551), .B2(n14578), .A(n14550), .ZN(n14552) );
  AOI21_X1 U16275 ( .B1(n13878), .B2(n14553), .A(n14552), .ZN(n14605) );
  INV_X1 U16276 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U16277 ( .A1(n14601), .A2(n14605), .B1(n15026), .B2(n14599), .ZN(
        P1_U3471) );
  AOI211_X1 U16278 ( .C1(n14588), .C2(n14557), .A(n14556), .B(n14555), .ZN(
        n14606) );
  INV_X1 U16279 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U16280 ( .A1(n14601), .A2(n14606), .B1(n14558), .B2(n14599), .ZN(
        P1_U3474) );
  OAI211_X1 U16281 ( .C1(n14561), .C2(n14592), .A(n14560), .B(n14559), .ZN(
        n14562) );
  INV_X1 U16282 ( .A(n14562), .ZN(n14608) );
  AOI22_X1 U16283 ( .A1(n14601), .A2(n14608), .B1(n8560), .B2(n14599), .ZN(
        P1_U3477) );
  XNOR2_X1 U16284 ( .A(n14563), .B(n14564), .ZN(n14570) );
  XNOR2_X1 U16285 ( .A(n14566), .B(n14565), .ZN(n14568) );
  AOI21_X1 U16286 ( .B1(n14568), .B2(n14597), .A(n14567), .ZN(n14569) );
  OAI21_X1 U16287 ( .B1(n14571), .B2(n14570), .A(n14569), .ZN(n15154) );
  INV_X1 U16288 ( .A(n14572), .ZN(n14574) );
  OAI21_X1 U16289 ( .B1(n14574), .B2(n14575), .A(n14573), .ZN(n15151) );
  OAI22_X1 U16290 ( .A1(n15151), .A2(n14576), .B1(n14575), .B2(n14592), .ZN(
        n14577) );
  NOR2_X1 U16291 ( .A1(n15154), .A2(n14577), .ZN(n14610) );
  AOI22_X1 U16292 ( .A1(n14601), .A2(n14610), .B1(n8484), .B2(n14599), .ZN(
        P1_U3480) );
  NOR2_X1 U16293 ( .A1(n14579), .A2(n14578), .ZN(n14583) );
  NOR4_X1 U16294 ( .A1(n14583), .A2(n14582), .A3(n14581), .A4(n14580), .ZN(
        n14611) );
  INV_X1 U16295 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U16296 ( .A1(n14601), .A2(n14611), .B1(n14584), .B2(n14599), .ZN(
        P1_U3483) );
  AOI211_X1 U16297 ( .C1(n14588), .C2(n14587), .A(n14586), .B(n14585), .ZN(
        n14612) );
  INV_X1 U16298 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14589) );
  AOI22_X1 U16299 ( .A1(n14601), .A2(n14612), .B1(n14589), .B2(n14599), .ZN(
        P1_U3486) );
  OAI211_X1 U16300 ( .C1(n14593), .C2(n14592), .A(n14591), .B(n14590), .ZN(
        n14596) );
  INV_X1 U16301 ( .A(n14594), .ZN(n14595) );
  AOI211_X1 U16302 ( .C1(n14598), .C2(n14597), .A(n14596), .B(n14595), .ZN(
        n14614) );
  INV_X1 U16303 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U16304 ( .A1(n14601), .A2(n14614), .B1(n14600), .B2(n14599), .ZN(
        P1_U3489) );
  AOI22_X1 U16305 ( .A1(n14615), .A2(n14602), .B1(n9827), .B2(n14613), .ZN(
        P1_U3529) );
  AOI22_X1 U16306 ( .A1(n14615), .A2(n14603), .B1(n9830), .B2(n14613), .ZN(
        P1_U3530) );
  AOI22_X1 U16307 ( .A1(n14615), .A2(n14604), .B1(n9833), .B2(n14613), .ZN(
        P1_U3531) );
  AOI22_X1 U16308 ( .A1(n14615), .A2(n14605), .B1(n9826), .B2(n14613), .ZN(
        P1_U3532) );
  AOI22_X1 U16309 ( .A1(n14615), .A2(n14606), .B1(n8575), .B2(n14613), .ZN(
        P1_U3533) );
  AOI22_X1 U16310 ( .A1(n14615), .A2(n14608), .B1(n14607), .B2(n14613), .ZN(
        P1_U3534) );
  AOI22_X1 U16311 ( .A1(n14615), .A2(n14610), .B1(n14609), .B2(n14613), .ZN(
        P1_U3535) );
  AOI22_X1 U16312 ( .A1(n14615), .A2(n14611), .B1(n9825), .B2(n14613), .ZN(
        P1_U3536) );
  AOI22_X1 U16313 ( .A1(n14615), .A2(n14612), .B1(n8457), .B2(n14613), .ZN(
        P1_U3537) );
  AOI22_X1 U16314 ( .A1(n14615), .A2(n14614), .B1(n8606), .B2(n14613), .ZN(
        P1_U3538) );
  NOR2_X1 U16315 ( .A1(n14680), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16316 ( .A(n14616), .ZN(n14618) );
  OAI21_X1 U16317 ( .B1(n14618), .B2(n14617), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14619) );
  OAI21_X1 U16318 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n14619), .ZN(n14630) );
  AOI211_X1 U16319 ( .C1(n14622), .C2(n14621), .A(n14620), .B(n14700), .ZN(
        n14623) );
  INV_X1 U16320 ( .A(n14623), .ZN(n14629) );
  OAI211_X1 U16321 ( .C1(n14626), .C2(n14625), .A(n14696), .B(n14624), .ZN(
        n14628) );
  NAND2_X1 U16322 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14680), .ZN(n14627) );
  NAND4_X1 U16323 ( .A1(n14630), .A2(n14629), .A3(n14628), .A4(n14627), .ZN(
        P2_U3218) );
  OAI21_X1 U16324 ( .B1(n14705), .B2(n9016), .A(n14631), .ZN(n14632) );
  AOI21_X1 U16325 ( .B1(n14633), .B2(n14694), .A(n14632), .ZN(n14642) );
  AOI211_X1 U16326 ( .C1(n6583), .C2(n14635), .A(n14700), .B(n14634), .ZN(
        n14636) );
  INV_X1 U16327 ( .A(n14636), .ZN(n14641) );
  OAI211_X1 U16328 ( .C1(n14639), .C2(n14638), .A(n14637), .B(n14696), .ZN(
        n14640) );
  NAND3_X1 U16329 ( .A1(n14642), .A2(n14641), .A3(n14640), .ZN(P2_U3221) );
  OAI21_X1 U16330 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14651) );
  OAI21_X1 U16331 ( .B1(n14648), .B2(n14647), .A(n14646), .ZN(n14649) );
  AOI222_X1 U16332 ( .A1(n14651), .A2(n14696), .B1(n14650), .B2(n14694), .C1(
        n14649), .C2(n14683), .ZN(n14653) );
  OAI211_X1 U16333 ( .C1(n14654), .C2(n14705), .A(n14653), .B(n14652), .ZN(
        P2_U3223) );
  INV_X1 U16334 ( .A(n14655), .ZN(n14656) );
  OAI21_X1 U16335 ( .B1(n14658), .B2(n14657), .A(n14656), .ZN(n14659) );
  AOI21_X1 U16336 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14680), .A(n14659), 
        .ZN(n14669) );
  OAI211_X1 U16337 ( .C1(n14662), .C2(n14661), .A(n14660), .B(n14696), .ZN(
        n14668) );
  AOI211_X1 U16338 ( .C1(n14665), .C2(n14664), .A(n14700), .B(n14663), .ZN(
        n14666) );
  INV_X1 U16339 ( .A(n14666), .ZN(n14667) );
  NAND3_X1 U16340 ( .A1(n14669), .A2(n14668), .A3(n14667), .ZN(P2_U3227) );
  AOI22_X1 U16341 ( .A1(n14680), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14679) );
  OAI211_X1 U16342 ( .C1(n14671), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14670), 
        .B(n14683), .ZN(n14678) );
  NAND2_X1 U16343 ( .A1(n14694), .A2(n14672), .ZN(n14677) );
  OAI211_X1 U16344 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14696), .ZN(
        n14676) );
  NAND4_X1 U16345 ( .A1(n14679), .A2(n14678), .A3(n14677), .A4(n14676), .ZN(
        P2_U3228) );
  AOI22_X1 U16346 ( .A1(n14680), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14690) );
  NAND2_X1 U16347 ( .A1(n14681), .A2(n14694), .ZN(n14689) );
  OAI211_X1 U16348 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14684), .A(n14683), 
        .B(n14682), .ZN(n14688) );
  OAI211_X1 U16349 ( .C1(n14686), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14696), 
        .B(n14685), .ZN(n14687) );
  NAND4_X1 U16350 ( .A1(n14690), .A2(n14689), .A3(n14688), .A4(n14687), .ZN(
        P2_U3229) );
  INV_X1 U16351 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14706) );
  AOI21_X1 U16352 ( .B1(n14692), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14691), 
        .ZN(n14701) );
  NAND2_X1 U16353 ( .A1(n14694), .A2(n14693), .ZN(n14699) );
  OAI211_X1 U16354 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14697), .A(n14696), 
        .B(n14695), .ZN(n14698) );
  OAI211_X1 U16355 ( .C1(n14701), .C2(n14700), .A(n14699), .B(n14698), .ZN(
        n14702) );
  INV_X1 U16356 ( .A(n14702), .ZN(n14704) );
  OAI211_X1 U16357 ( .C1(n14706), .C2(n14705), .A(n14704), .B(n14703), .ZN(
        P2_U3232) );
  AOI22_X1 U16358 ( .A1(n14710), .A2(n14709), .B1(n14708), .B2(n14707), .ZN(
        n14711) );
  NAND3_X1 U16359 ( .A1(n14714), .A2(n14712), .A3(n14711), .ZN(n14713) );
  OAI21_X1 U16360 ( .B1(n14714), .B2(P2_REG2_REG_0__SCAN_IN), .A(n14713), .ZN(
        n14715) );
  OAI21_X1 U16361 ( .B1(n10292), .B2(n14716), .A(n14715), .ZN(P2_U3265) );
  INV_X1 U16362 ( .A(n14717), .ZN(n14718) );
  AND2_X1 U16363 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14720), .ZN(P2_U3266) );
  AND2_X1 U16364 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14720), .ZN(P2_U3267) );
  AND2_X1 U16365 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14720), .ZN(P2_U3268) );
  INV_X1 U16366 ( .A(n14720), .ZN(n14719) );
  INV_X1 U16367 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15110) );
  NOR2_X1 U16368 ( .A1(n14719), .A2(n15110), .ZN(P2_U3269) );
  AND2_X1 U16369 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14720), .ZN(P2_U3270) );
  AND2_X1 U16370 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14720), .ZN(P2_U3271) );
  AND2_X1 U16371 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14720), .ZN(P2_U3272) );
  AND2_X1 U16372 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14720), .ZN(P2_U3273) );
  AND2_X1 U16373 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14720), .ZN(P2_U3274) );
  AND2_X1 U16374 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14720), .ZN(P2_U3275) );
  AND2_X1 U16375 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14720), .ZN(P2_U3276) );
  AND2_X1 U16376 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14720), .ZN(P2_U3277) );
  AND2_X1 U16377 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14720), .ZN(P2_U3278) );
  AND2_X1 U16378 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14720), .ZN(P2_U3279) );
  AND2_X1 U16379 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14720), .ZN(P2_U3280) );
  AND2_X1 U16380 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14720), .ZN(P2_U3281) );
  AND2_X1 U16381 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14720), .ZN(P2_U3282) );
  AND2_X1 U16382 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14720), .ZN(P2_U3283) );
  AND2_X1 U16383 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14720), .ZN(P2_U3284) );
  AND2_X1 U16384 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14720), .ZN(P2_U3285) );
  INV_X1 U16385 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15053) );
  NOR2_X1 U16386 ( .A1(n14719), .A2(n15053), .ZN(P2_U3286) );
  AND2_X1 U16387 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14720), .ZN(P2_U3287) );
  AND2_X1 U16388 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14720), .ZN(P2_U3288) );
  AND2_X1 U16389 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14720), .ZN(P2_U3289) );
  AND2_X1 U16390 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14720), .ZN(P2_U3290) );
  AND2_X1 U16391 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14720), .ZN(P2_U3291) );
  AND2_X1 U16392 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14720), .ZN(P2_U3292) );
  AND2_X1 U16393 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14720), .ZN(P2_U3293) );
  AND2_X1 U16394 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14720), .ZN(P2_U3294) );
  AND2_X1 U16395 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14720), .ZN(P2_U3295) );
  OAI21_X1 U16396 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(P2_U3416) );
  AOI21_X1 U16397 ( .B1(n14725), .B2(P2_D_REG_1__SCAN_IN), .A(n14724), .ZN(
        n14726) );
  INV_X1 U16398 ( .A(n14726), .ZN(P2_U3417) );
  INV_X1 U16399 ( .A(n14727), .ZN(n14729) );
  AOI211_X1 U16400 ( .C1(n13261), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        n14732) );
  OAI211_X1 U16401 ( .C1(n14749), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        n14734) );
  INV_X1 U16402 ( .A(n14734), .ZN(n14771) );
  INV_X1 U16403 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U16404 ( .A1(n14754), .A2(n14771), .B1(n14735), .B2(n14769), .ZN(
        P2_U3439) );
  NAND2_X1 U16405 ( .A1(n14737), .A2(n14736), .ZN(n14740) );
  INV_X1 U16406 ( .A(n14738), .ZN(n14739) );
  OAI211_X1 U16407 ( .C1(n14741), .C2(n14764), .A(n14740), .B(n14739), .ZN(
        n14742) );
  NOR2_X1 U16408 ( .A1(n14743), .A2(n14742), .ZN(n14772) );
  INV_X1 U16409 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U16410 ( .A1(n14754), .A2(n14772), .B1(n14744), .B2(n14769), .ZN(
        P2_U3442) );
  AOI21_X1 U16411 ( .B1(n14746), .B2(n13261), .A(n14745), .ZN(n14748) );
  OAI211_X1 U16412 ( .C1(n14750), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        n14751) );
  AOI21_X1 U16413 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14773) );
  AOI22_X1 U16414 ( .A1(n14754), .A2(n14773), .B1(n9220), .B2(n14769), .ZN(
        P2_U3451) );
  NAND2_X1 U16415 ( .A1(n14755), .A2(n13261), .ZN(n14756) );
  OAI211_X1 U16416 ( .C1(n14758), .C2(n14761), .A(n14757), .B(n14756), .ZN(
        n14759) );
  NOR2_X1 U16417 ( .A1(n14760), .A2(n14759), .ZN(n14775) );
  AOI22_X1 U16418 ( .A1(n14754), .A2(n14775), .B1(n9237), .B2(n14769), .ZN(
        P2_U3454) );
  NOR2_X1 U16419 ( .A1(n14762), .A2(n14761), .ZN(n14767) );
  OAI21_X1 U16420 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14766) );
  NOR3_X1 U16421 ( .A1(n14768), .A2(n14767), .A3(n14766), .ZN(n14777) );
  INV_X1 U16422 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14770) );
  AOI22_X1 U16423 ( .A1(n14754), .A2(n14777), .B1(n14770), .B2(n14769), .ZN(
        P2_U3460) );
  AOI22_X1 U16424 ( .A1(n6436), .A2(n14771), .B1(n9960), .B2(n14776), .ZN(
        P2_U3502) );
  AOI22_X1 U16425 ( .A1(n6436), .A2(n14772), .B1(n9962), .B2(n14776), .ZN(
        P2_U3503) );
  AOI22_X1 U16426 ( .A1(n6436), .A2(n14773), .B1(n9966), .B2(n14776), .ZN(
        P2_U3506) );
  AOI22_X1 U16427 ( .A1(n6436), .A2(n14775), .B1(n14774), .B2(n14776), .ZN(
        P2_U3507) );
  AOI22_X1 U16428 ( .A1(n6436), .A2(n14777), .B1(n9272), .B2(n14776), .ZN(
        P2_U3509) );
  NOR2_X1 U16429 ( .A1(P3_U3897), .A2(n14799), .ZN(P3_U3150) );
  INV_X1 U16430 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14798) );
  AOI21_X1 U16431 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14782) );
  NOR2_X1 U16432 ( .A1(n14782), .A2(n14781), .ZN(n14794) );
  AOI21_X1 U16433 ( .B1(n14785), .B2(n14784), .A(n14783), .ZN(n14792) );
  OAI21_X1 U16434 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14790) );
  AOI22_X1 U16435 ( .A1(n14790), .A2(n14809), .B1(n14789), .B2(n14801), .ZN(
        n14791) );
  OAI21_X1 U16436 ( .B1(n14792), .B2(n14815), .A(n14791), .ZN(n14793) );
  NOR2_X1 U16437 ( .A1(n14794), .A2(n14793), .ZN(n14796) );
  OAI211_X1 U16438 ( .C1(n14798), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        P3_U3190) );
  AOI22_X1 U16439 ( .A1(n14801), .A2(n14800), .B1(n14799), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n14820) );
  OAI21_X1 U16440 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14811) );
  OAI21_X1 U16441 ( .B1(n14807), .B2(n14806), .A(n14805), .ZN(n14808) );
  AOI22_X1 U16442 ( .A1(n14811), .A2(n14810), .B1(n14809), .B2(n14808), .ZN(
        n14819) );
  AOI21_X1 U16443 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n14816) );
  OR2_X1 U16444 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  NAND4_X1 U16445 ( .A1(n14820), .A2(n14819), .A3(n14818), .A4(n14817), .ZN(
        P3_U3192) );
  XNOR2_X1 U16446 ( .A(n14822), .B(n11649), .ZN(n14829) );
  INV_X1 U16447 ( .A(n14829), .ZN(n14967) );
  OAI211_X1 U16448 ( .C1(n14824), .C2(n11649), .A(n14920), .B(n14823), .ZN(
        n14828) );
  AOI22_X1 U16449 ( .A1(n14892), .A2(n14826), .B1(n14825), .B2(n14889), .ZN(
        n14827) );
  OAI211_X1 U16450 ( .C1(n14924), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14964) );
  AOI21_X1 U16451 ( .B1(n14926), .B2(n14967), .A(n14964), .ZN(n14834) );
  AND2_X1 U16452 ( .A1(n14830), .A2(n14907), .ZN(n14965) );
  AOI22_X1 U16453 ( .A1(n14902), .A2(n14965), .B1(n14831), .B2(n14901), .ZN(
        n14832) );
  OAI221_X1 U16454 ( .B1(n14865), .B2(n14834), .C1(n14927), .C2(n14833), .A(
        n14832), .ZN(P3_U3224) );
  XNOR2_X1 U16455 ( .A(n14835), .B(n14837), .ZN(n14844) );
  INV_X1 U16456 ( .A(n14844), .ZN(n14962) );
  OAI21_X1 U16457 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14842) );
  OAI22_X1 U16458 ( .A1(n14840), .A2(n14917), .B1(n14839), .B2(n14915), .ZN(
        n14841) );
  AOI21_X1 U16459 ( .B1(n14842), .B2(n14920), .A(n14841), .ZN(n14843) );
  OAI21_X1 U16460 ( .B1(n14924), .B2(n14844), .A(n14843), .ZN(n14960) );
  AOI21_X1 U16461 ( .B1(n14926), .B2(n14962), .A(n14960), .ZN(n14849) );
  AND2_X1 U16462 ( .A1(n14845), .A2(n14907), .ZN(n14961) );
  AOI22_X1 U16463 ( .A1(n14902), .A2(n14961), .B1(n14901), .B2(n14846), .ZN(
        n14847) );
  OAI221_X1 U16464 ( .B1(n14865), .B2(n14849), .C1(n14927), .C2(n14848), .A(
        n14847), .ZN(P3_U3225) );
  XNOR2_X1 U16465 ( .A(n14850), .B(n14854), .ZN(n14946) );
  INV_X1 U16466 ( .A(n14852), .ZN(n14853) );
  AOI21_X1 U16467 ( .B1(n14854), .B2(n14851), .A(n14853), .ZN(n14858) );
  AOI22_X1 U16468 ( .A1(n14892), .A2(n14890), .B1(n14855), .B2(n14889), .ZN(
        n14857) );
  NAND2_X1 U16469 ( .A1(n14946), .A2(n14875), .ZN(n14856) );
  OAI211_X1 U16470 ( .C1(n14858), .C2(n14877), .A(n14857), .B(n14856), .ZN(
        n14944) );
  AOI21_X1 U16471 ( .B1(n14926), .B2(n14946), .A(n14944), .ZN(n14863) );
  AND2_X1 U16472 ( .A1(n14859), .A2(n14907), .ZN(n14945) );
  AOI22_X1 U16473 ( .A1(n14902), .A2(n14945), .B1(n14901), .B2(n14860), .ZN(
        n14861) );
  OAI221_X1 U16474 ( .B1(n14865), .B2(n14863), .C1(n14927), .C2(n14862), .A(
        n14861), .ZN(P3_U3228) );
  AND2_X1 U16475 ( .A1(n14864), .A2(n14907), .ZN(n14941) );
  AOI22_X1 U16476 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n14865), .B1(n14902), 
        .B2(n14941), .ZN(n14883) );
  XNOR2_X1 U16477 ( .A(n14868), .B(n14867), .ZN(n14878) );
  AND2_X1 U16478 ( .A1(n14870), .A2(n14869), .ZN(n14872) );
  XNOR2_X1 U16479 ( .A(n14872), .B(n14871), .ZN(n14942) );
  OAI22_X1 U16480 ( .A1(n14873), .A2(n14915), .B1(n14916), .B2(n14917), .ZN(
        n14874) );
  AOI21_X1 U16481 ( .B1(n14942), .B2(n14875), .A(n14874), .ZN(n14876) );
  OAI21_X1 U16482 ( .B1(n14878), .B2(n14877), .A(n14876), .ZN(n14940) );
  INV_X1 U16483 ( .A(n14942), .ZN(n14880) );
  NOR2_X1 U16484 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  OAI21_X1 U16485 ( .B1(n14940), .B2(n14881), .A(n14927), .ZN(n14882) );
  OAI211_X1 U16486 ( .C1(n14884), .C2(n14910), .A(n14883), .B(n14882), .ZN(
        P3_U3229) );
  NAND2_X1 U16487 ( .A1(n14886), .A2(n14885), .ZN(n14888) );
  NAND2_X1 U16488 ( .A1(n14888), .A2(n14893), .ZN(n14887) );
  OAI21_X1 U16489 ( .B1(n14888), .B2(n14893), .A(n14887), .ZN(n14938) );
  INV_X1 U16490 ( .A(n14938), .ZN(n14898) );
  AOI22_X1 U16491 ( .A1(n14892), .A2(n14891), .B1(n14890), .B2(n14889), .ZN(
        n14897) );
  OAI211_X1 U16492 ( .C1(n14895), .C2(n11301), .A(n14920), .B(n14894), .ZN(
        n14896) );
  OAI211_X1 U16493 ( .C1(n14898), .C2(n14924), .A(n14897), .B(n14896), .ZN(
        n14936) );
  AOI21_X1 U16494 ( .B1(n14926), .B2(n14938), .A(n14936), .ZN(n14905) );
  NOR2_X1 U16495 ( .A1(n14899), .A2(n14954), .ZN(n14937) );
  AOI22_X1 U16496 ( .A1(n14902), .A2(n14937), .B1(n14901), .B2(n14900), .ZN(
        n14903) );
  OAI221_X1 U16497 ( .B1(n14865), .B2(n14905), .C1(n14927), .C2(n14904), .A(
        n14903), .ZN(P3_U3230) );
  XNOR2_X1 U16498 ( .A(n14914), .B(n14906), .ZN(n14923) );
  INV_X1 U16499 ( .A(n14923), .ZN(n14934) );
  NAND2_X1 U16500 ( .A1(n14933), .A2(n14908), .ZN(n14909) );
  OAI21_X1 U16501 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14925) );
  OAI21_X1 U16502 ( .B1(n14912), .B2(n14914), .A(n14913), .ZN(n14921) );
  OAI22_X1 U16503 ( .A1(n14918), .A2(n14917), .B1(n14916), .B2(n14915), .ZN(
        n14919) );
  AOI21_X1 U16504 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14922) );
  OAI21_X1 U16505 ( .B1(n14924), .B2(n14923), .A(n14922), .ZN(n14932) );
  AOI211_X1 U16506 ( .C1(n14926), .C2(n14934), .A(n14925), .B(n14932), .ZN(
        n14928) );
  AOI22_X1 U16507 ( .A1(n14865), .A2(n15096), .B1(n14928), .B2(n14927), .ZN(
        P3_U3231) );
  AOI211_X1 U16508 ( .C1(n14972), .C2(n14931), .A(n14930), .B(n14929), .ZN(
        n14976) );
  INV_X1 U16509 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15070) );
  AOI22_X1 U16510 ( .A1(n14975), .A2(n14976), .B1(n15070), .B2(n14973), .ZN(
        P3_U3393) );
  AOI211_X1 U16511 ( .C1(n14934), .C2(n14966), .A(n14933), .B(n14932), .ZN(
        n14977) );
  INV_X1 U16512 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14935) );
  AOI22_X1 U16513 ( .A1(n14975), .A2(n14977), .B1(n14935), .B2(n14973), .ZN(
        P3_U3396) );
  AOI211_X1 U16514 ( .C1(n14966), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14979) );
  INV_X1 U16515 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U16516 ( .A1(n14975), .A2(n14979), .B1(n14939), .B2(n14973), .ZN(
        P3_U3399) );
  AOI211_X1 U16517 ( .C1(n14942), .C2(n14966), .A(n14941), .B(n14940), .ZN(
        n14981) );
  INV_X1 U16518 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U16519 ( .A1(n14975), .A2(n14981), .B1(n14943), .B2(n14973), .ZN(
        P3_U3402) );
  AOI211_X1 U16520 ( .C1(n14946), .C2(n14966), .A(n14945), .B(n14944), .ZN(
        n14983) );
  INV_X1 U16521 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14947) );
  AOI22_X1 U16522 ( .A1(n14975), .A2(n14983), .B1(n14947), .B2(n14973), .ZN(
        P3_U3405) );
  INV_X1 U16523 ( .A(n14948), .ZN(n14950) );
  AOI211_X1 U16524 ( .C1(n14966), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14984) );
  INV_X1 U16525 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U16526 ( .A1(n14975), .A2(n14984), .B1(n14952), .B2(n14973), .ZN(
        P3_U3408) );
  OAI22_X1 U16527 ( .A1(n14956), .A2(n14955), .B1(n14954), .B2(n14953), .ZN(
        n14957) );
  NOR2_X1 U16528 ( .A1(n14958), .A2(n14957), .ZN(n14985) );
  INV_X1 U16529 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U16530 ( .A1(n14975), .A2(n14985), .B1(n14959), .B2(n14973), .ZN(
        P3_U3411) );
  AOI211_X1 U16531 ( .C1(n14962), .C2(n14966), .A(n14961), .B(n14960), .ZN(
        n14987) );
  INV_X1 U16532 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16533 ( .A1(n14975), .A2(n14987), .B1(n14963), .B2(n14973), .ZN(
        P3_U3414) );
  AOI211_X1 U16534 ( .C1(n14967), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14989) );
  INV_X1 U16535 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U16536 ( .A1(n14975), .A2(n14989), .B1(n14968), .B2(n14973), .ZN(
        P3_U3417) );
  AOI211_X1 U16537 ( .C1(n14972), .C2(n14971), .A(n14970), .B(n14969), .ZN(
        n14992) );
  INV_X1 U16538 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U16539 ( .A1(n14975), .A2(n14992), .B1(n14974), .B2(n14973), .ZN(
        P3_U3420) );
  AOI22_X1 U16540 ( .A1(n14993), .A2(n14976), .B1(n10510), .B2(n14990), .ZN(
        P3_U3460) );
  AOI22_X1 U16541 ( .A1(n14993), .A2(n14977), .B1(n10440), .B2(n14990), .ZN(
        P3_U3461) );
  INV_X1 U16542 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16543 ( .A1(n14993), .A2(n14979), .B1(n14978), .B2(n14990), .ZN(
        P3_U3462) );
  AOI22_X1 U16544 ( .A1(n14993), .A2(n14981), .B1(n14980), .B2(n14990), .ZN(
        P3_U3463) );
  AOI22_X1 U16545 ( .A1(n14993), .A2(n14983), .B1(n14982), .B2(n14990), .ZN(
        P3_U3464) );
  AOI22_X1 U16546 ( .A1(n14993), .A2(n14984), .B1(n10414), .B2(n14990), .ZN(
        P3_U3465) );
  AOI22_X1 U16547 ( .A1(n14993), .A2(n14985), .B1(n10479), .B2(n14990), .ZN(
        P3_U3466) );
  AOI22_X1 U16548 ( .A1(n14993), .A2(n14987), .B1(n14986), .B2(n14990), .ZN(
        P3_U3467) );
  INV_X1 U16549 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n14988) );
  AOI22_X1 U16550 ( .A1(n14993), .A2(n14989), .B1(n14988), .B2(n14990), .ZN(
        P3_U3468) );
  AOI22_X1 U16551 ( .A1(n14993), .A2(n14992), .B1(n14991), .B2(n14990), .ZN(
        P3_U3469) );
  NOR2_X1 U16552 ( .A1(keyinput12), .A2(keyinput28), .ZN(n14994) );
  NAND3_X1 U16553 ( .A1(keyinput7), .A2(keyinput55), .A3(n14994), .ZN(n15000)
         );
  NAND3_X1 U16554 ( .A1(keyinput34), .A2(keyinput32), .A3(keyinput51), .ZN(
        n14999) );
  NOR3_X1 U16555 ( .A1(keyinput23), .A2(keyinput10), .A3(keyinput57), .ZN(
        n14997) );
  INV_X1 U16556 ( .A(keyinput15), .ZN(n14995) );
  NOR3_X1 U16557 ( .A1(keyinput20), .A2(keyinput62), .A3(n14995), .ZN(n14996)
         );
  NAND4_X1 U16558 ( .A1(keyinput26), .A2(n14997), .A3(keyinput60), .A4(n14996), 
        .ZN(n14998) );
  NOR4_X1 U16559 ( .A1(keyinput46), .A2(n15000), .A3(n14999), .A4(n14998), 
        .ZN(n15143) );
  NAND3_X1 U16560 ( .A1(keyinput33), .A2(keyinput19), .A3(keyinput41), .ZN(
        n15022) );
  NOR3_X1 U16561 ( .A1(keyinput13), .A2(keyinput3), .A3(keyinput25), .ZN(
        n15005) );
  INV_X1 U16562 ( .A(keyinput29), .ZN(n15001) );
  NOR4_X1 U16563 ( .A1(keyinput24), .A2(keyinput11), .A3(keyinput4), .A4(
        n15001), .ZN(n15004) );
  INV_X1 U16564 ( .A(keyinput6), .ZN(n15002) );
  NOR4_X1 U16565 ( .A1(keyinput37), .A2(keyinput50), .A3(keyinput43), .A4(
        n15002), .ZN(n15003) );
  NAND4_X1 U16566 ( .A1(keyinput38), .A2(n15005), .A3(n15004), .A4(n15003), 
        .ZN(n15021) );
  NOR3_X1 U16567 ( .A1(keyinput54), .A2(keyinput40), .A3(keyinput61), .ZN(
        n15019) );
  NAND2_X1 U16568 ( .A1(keyinput44), .A2(keyinput31), .ZN(n15009) );
  NOR2_X1 U16569 ( .A1(keyinput1), .A2(keyinput8), .ZN(n15007) );
  NOR4_X1 U16570 ( .A1(keyinput14), .A2(keyinput2), .A3(keyinput18), .A4(
        keyinput5), .ZN(n15006) );
  NAND4_X1 U16571 ( .A1(keyinput36), .A2(keyinput63), .A3(n15007), .A4(n15006), 
        .ZN(n15008) );
  NOR4_X1 U16572 ( .A1(keyinput53), .A2(keyinput9), .A3(n15009), .A4(n15008), 
        .ZN(n15018) );
  NOR2_X1 U16573 ( .A1(keyinput17), .A2(keyinput0), .ZN(n15010) );
  NAND3_X1 U16574 ( .A1(keyinput22), .A2(keyinput16), .A3(n15010), .ZN(n15016)
         );
  NAND3_X1 U16575 ( .A1(keyinput56), .A2(keyinput49), .A3(keyinput39), .ZN(
        n15015) );
  NOR2_X1 U16576 ( .A1(keyinput47), .A2(keyinput59), .ZN(n15013) );
  INV_X1 U16577 ( .A(keyinput52), .ZN(n15011) );
  NOR4_X1 U16578 ( .A1(keyinput42), .A2(keyinput27), .A3(keyinput35), .A4(
        n15011), .ZN(n15012) );
  NAND4_X1 U16579 ( .A1(keyinput30), .A2(keyinput58), .A3(n15013), .A4(n15012), 
        .ZN(n15014) );
  NOR4_X1 U16580 ( .A1(keyinput48), .A2(n15016), .A3(n15015), .A4(n15014), 
        .ZN(n15017) );
  NAND4_X1 U16581 ( .A1(keyinput21), .A2(n15019), .A3(n15018), .A4(n15017), 
        .ZN(n15020) );
  NOR4_X1 U16582 ( .A1(keyinput45), .A2(n15022), .A3(n15021), .A4(n15020), 
        .ZN(n15142) );
  AOI22_X1 U16583 ( .A1(n6649), .A2(keyinput57), .B1(keyinput26), .B2(n15024), 
        .ZN(n15023) );
  OAI221_X1 U16584 ( .B1(n6649), .B2(keyinput57), .C1(n15024), .C2(keyinput26), 
        .A(n15023), .ZN(n15034) );
  INV_X1 U16585 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15027) );
  AOI22_X1 U16586 ( .A1(n15027), .A2(keyinput7), .B1(keyinput55), .B2(n15026), 
        .ZN(n15025) );
  OAI221_X1 U16587 ( .B1(n15027), .B2(keyinput7), .C1(n15026), .C2(keyinput55), 
        .A(n15025), .ZN(n15033) );
  XNOR2_X1 U16588 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput28), .ZN(n15031) );
  XNOR2_X1 U16589 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput12), .ZN(n15030)
         );
  XNOR2_X1 U16590 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput10), .ZN(n15029) );
  XNOR2_X1 U16591 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput23), .ZN(n15028)
         );
  NAND4_X1 U16592 ( .A1(n15031), .A2(n15030), .A3(n15029), .A4(n15028), .ZN(
        n15032) );
  NOR3_X1 U16593 ( .A1(n15034), .A2(n15033), .A3(n15032), .ZN(n15081) );
  AOI22_X1 U16594 ( .A1(n15037), .A2(keyinput34), .B1(keyinput32), .B2(n15036), 
        .ZN(n15035) );
  OAI221_X1 U16595 ( .B1(n15037), .B2(keyinput34), .C1(n15036), .C2(keyinput32), .A(n15035), .ZN(n15048) );
  AOI22_X1 U16596 ( .A1(n9047), .A2(keyinput15), .B1(keyinput62), .B2(n15039), 
        .ZN(n15038) );
  OAI221_X1 U16597 ( .B1(n9047), .B2(keyinput15), .C1(n15039), .C2(keyinput62), 
        .A(n15038), .ZN(n15047) );
  AOI22_X1 U16598 ( .A1(n15042), .A2(keyinput60), .B1(n15041), .B2(keyinput20), 
        .ZN(n15040) );
  OAI221_X1 U16599 ( .B1(n15042), .B2(keyinput60), .C1(n15041), .C2(keyinput20), .A(n15040), .ZN(n15046) );
  XNOR2_X1 U16600 ( .A(P3_REG0_REG_14__SCAN_IN), .B(keyinput51), .ZN(n15044)
         );
  XNOR2_X1 U16601 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput46), .ZN(n15043) );
  NAND2_X1 U16602 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  NOR4_X1 U16603 ( .A1(n15048), .A2(n15047), .A3(n15046), .A4(n15045), .ZN(
        n15080) );
  AOI22_X1 U16604 ( .A1(n15051), .A2(keyinput44), .B1(n15050), .B2(keyinput53), 
        .ZN(n15049) );
  OAI221_X1 U16605 ( .B1(n15051), .B2(keyinput44), .C1(n15050), .C2(keyinput53), .A(n15049), .ZN(n15063) );
  AOI22_X1 U16606 ( .A1(n15053), .A2(keyinput9), .B1(n11406), .B2(keyinput31), 
        .ZN(n15052) );
  OAI221_X1 U16607 ( .B1(n15053), .B2(keyinput9), .C1(n11406), .C2(keyinput31), 
        .A(n15052), .ZN(n15062) );
  AOI22_X1 U16608 ( .A1(n15056), .A2(keyinput36), .B1(n15055), .B2(keyinput1), 
        .ZN(n15054) );
  OAI221_X1 U16609 ( .B1(n15056), .B2(keyinput36), .C1(n15055), .C2(keyinput1), 
        .A(n15054), .ZN(n15061) );
  INV_X1 U16610 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U16611 ( .A1(n15059), .A2(keyinput63), .B1(n15058), .B2(keyinput8), 
        .ZN(n15057) );
  OAI221_X1 U16612 ( .B1(n15059), .B2(keyinput63), .C1(n15058), .C2(keyinput8), 
        .A(n15057), .ZN(n15060) );
  NOR4_X1 U16613 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15079) );
  AOI22_X1 U16614 ( .A1(n15066), .A2(keyinput54), .B1(n15065), .B2(keyinput40), 
        .ZN(n15064) );
  OAI221_X1 U16615 ( .B1(n15066), .B2(keyinput54), .C1(n15065), .C2(keyinput40), .A(n15064), .ZN(n15077) );
  AOI22_X1 U16616 ( .A1(n15069), .A2(keyinput61), .B1(keyinput21), .B2(n15068), 
        .ZN(n15067) );
  OAI221_X1 U16617 ( .B1(n15069), .B2(keyinput61), .C1(n15068), .C2(keyinput21), .A(n15067), .ZN(n15076) );
  XOR2_X1 U16618 ( .A(n15070), .B(keyinput18), .Z(n15074) );
  XNOR2_X1 U16619 ( .A(P1_REG3_REG_12__SCAN_IN), .B(keyinput2), .ZN(n15073) );
  XNOR2_X1 U16620 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput14), .ZN(n15072) );
  XNOR2_X1 U16621 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput5), .ZN(n15071) );
  NAND4_X1 U16622 ( .A1(n15074), .A2(n15073), .A3(n15072), .A4(n15071), .ZN(
        n15075) );
  NOR3_X1 U16623 ( .A1(n15077), .A2(n15076), .A3(n15075), .ZN(n15078) );
  NAND4_X1 U16624 ( .A1(n15081), .A2(n15080), .A3(n15079), .A4(n15078), .ZN(
        n15141) );
  AOI22_X1 U16625 ( .A1(n15083), .A2(keyinput29), .B1(n9876), .B2(keyinput11), 
        .ZN(n15082) );
  OAI221_X1 U16626 ( .B1(n15083), .B2(keyinput29), .C1(n9876), .C2(keyinput11), 
        .A(n15082), .ZN(n15094) );
  AOI22_X1 U16627 ( .A1(n9833), .A2(keyinput24), .B1(n15085), .B2(keyinput4), 
        .ZN(n15084) );
  OAI221_X1 U16628 ( .B1(n9833), .B2(keyinput24), .C1(n15085), .C2(keyinput4), 
        .A(n15084), .ZN(n15093) );
  AOI22_X1 U16629 ( .A1(n15088), .A2(keyinput37), .B1(n15087), .B2(keyinput6), 
        .ZN(n15086) );
  OAI221_X1 U16630 ( .B1(n15088), .B2(keyinput37), .C1(n15087), .C2(keyinput6), 
        .A(n15086), .ZN(n15092) );
  XNOR2_X1 U16631 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput50), .ZN(n15090) );
  XNOR2_X1 U16632 ( .A(keyinput43), .B(P1_REG2_REG_0__SCAN_IN), .ZN(n15089) );
  NAND2_X1 U16633 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  NOR4_X1 U16634 ( .A1(n15094), .A2(n15093), .A3(n15092), .A4(n15091), .ZN(
        n15139) );
  AOI22_X1 U16635 ( .A1(n15097), .A2(keyinput19), .B1(keyinput41), .B2(n15096), 
        .ZN(n15095) );
  OAI221_X1 U16636 ( .B1(n15097), .B2(keyinput19), .C1(n15096), .C2(keyinput41), .A(n15095), .ZN(n15106) );
  AOI22_X1 U16637 ( .A1(n10004), .A2(keyinput38), .B1(n15099), .B2(keyinput25), 
        .ZN(n15098) );
  OAI221_X1 U16638 ( .B1(n10004), .B2(keyinput38), .C1(n15099), .C2(keyinput25), .A(n15098), .ZN(n15105) );
  XNOR2_X1 U16639 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput33), .ZN(n15103)
         );
  XNOR2_X1 U16640 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput45), .ZN(n15102) );
  XNOR2_X1 U16641 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput13), .ZN(n15101) );
  XNOR2_X1 U16642 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput3), .ZN(n15100)
         );
  NAND4_X1 U16643 ( .A1(n15103), .A2(n15102), .A3(n15101), .A4(n15100), .ZN(
        n15104) );
  NOR3_X1 U16644 ( .A1(n15106), .A2(n15105), .A3(n15104), .ZN(n15138) );
  AOI22_X1 U16645 ( .A1(n9975), .A2(keyinput59), .B1(keyinput58), .B2(n15108), 
        .ZN(n15107) );
  OAI221_X1 U16646 ( .B1(n9975), .B2(keyinput59), .C1(n15108), .C2(keyinput58), 
        .A(n15107), .ZN(n15120) );
  AOI22_X1 U16647 ( .A1(n15110), .A2(keyinput30), .B1(keyinput47), .B2(n9960), 
        .ZN(n15109) );
  OAI221_X1 U16648 ( .B1(n15110), .B2(keyinput30), .C1(n9960), .C2(keyinput47), 
        .A(n15109), .ZN(n15119) );
  AOI22_X1 U16649 ( .A1(n15113), .A2(keyinput52), .B1(n15112), .B2(keyinput35), 
        .ZN(n15111) );
  OAI221_X1 U16650 ( .B1(n15113), .B2(keyinput52), .C1(n15112), .C2(keyinput35), .A(n15111), .ZN(n15118) );
  AOI22_X1 U16651 ( .A1(n15116), .A2(keyinput42), .B1(keyinput27), .B2(n15115), 
        .ZN(n15114) );
  OAI221_X1 U16652 ( .B1(n15116), .B2(keyinput42), .C1(n15115), .C2(keyinput27), .A(n15114), .ZN(n15117) );
  NOR4_X1 U16653 ( .A1(n15120), .A2(n15119), .A3(n15118), .A4(n15117), .ZN(
        n15137) );
  AOI22_X1 U16654 ( .A1(n7481), .A2(keyinput49), .B1(keyinput39), .B2(n15122), 
        .ZN(n15121) );
  OAI221_X1 U16655 ( .B1(n7481), .B2(keyinput49), .C1(n15122), .C2(keyinput39), 
        .A(n15121), .ZN(n15128) );
  XNOR2_X1 U16656 ( .A(n15123), .B(keyinput16), .ZN(n15127) );
  XOR2_X1 U16657 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput22), .Z(n15126) );
  XNOR2_X1 U16658 ( .A(n15124), .B(keyinput0), .ZN(n15125) );
  OR4_X1 U16659 ( .A1(n15128), .A2(n15127), .A3(n15126), .A4(n15125), .ZN(
        n15135) );
  AOI22_X1 U16660 ( .A1(n15131), .A2(keyinput56), .B1(n15130), .B2(keyinput48), 
        .ZN(n15129) );
  OAI221_X1 U16661 ( .B1(n15131), .B2(keyinput56), .C1(n15130), .C2(keyinput48), .A(n15129), .ZN(n15134) );
  XNOR2_X1 U16662 ( .A(n15132), .B(keyinput17), .ZN(n15133) );
  NOR3_X1 U16663 ( .A1(n15135), .A2(n15134), .A3(n15133), .ZN(n15136) );
  NAND4_X1 U16664 ( .A1(n15139), .A2(n15138), .A3(n15137), .A4(n15136), .ZN(
        n15140) );
  AOI211_X1 U16665 ( .C1(n15143), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        n15156) );
  OAI22_X1 U16666 ( .A1(n15146), .A2(n9858), .B1(n15145), .B2(n15144), .ZN(
        n15147) );
  AOI21_X1 U16667 ( .B1(n15149), .B2(n15148), .A(n15147), .ZN(n15150) );
  OAI21_X1 U16668 ( .B1(n15152), .B2(n15151), .A(n15150), .ZN(n15153) );
  AOI21_X1 U16669 ( .B1(n15154), .B2(n15146), .A(n15153), .ZN(n15155) );
  XNOR2_X1 U16670 ( .A(n15156), .B(n15155), .ZN(P1_U3286) );
  OAI21_X1 U16671 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(SUB_1596_U59) );
  OAI21_X1 U16672 ( .B1(n15162), .B2(n15161), .A(n15160), .ZN(SUB_1596_U58) );
  XOR2_X1 U16673 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15163), .Z(SUB_1596_U53) );
  AOI21_X1 U16674 ( .B1(n15166), .B2(n15165), .A(n15164), .ZN(SUB_1596_U56) );
  OAI21_X1 U16675 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(SUB_1596_U60) );
  AOI21_X1 U16676 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(SUB_1596_U5) );
  NAND2_X1 U7248 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  CLKBUF_X1 U7199 ( .A(n9191), .Z(n11974) );
  NAND2_X1 U7205 ( .A1(n13930), .A2(n13838), .ZN(n13911) );
  CLKBUF_X2 U7220 ( .A(n9138), .Z(n9530) );
  NAND2_X1 U7228 ( .A1(n6943), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8253) );
  CLKBUF_X1 U7236 ( .A(n9107), .Z(n12023) );
  NAND2_X1 U7347 ( .A1(n9954), .A2(n9967), .ZN(n15177) );
endmodule

