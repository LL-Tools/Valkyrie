

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540;

  INV_X4 U4953 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  OR2_X1 U4954 ( .A1(n9690), .A2(n9438), .ZN(n8262) );
  XNOR2_X1 U4955 ( .A(n6836), .B(n5764), .ZN(n8367) );
  AOI21_X1 U4956 ( .B1(n5747), .B2(n5746), .A(n5745), .ZN(n5759) );
  NOR2_X1 U4957 ( .A1(n5114), .A2(n7508), .ZN(n7705) );
  AOI21_X1 U4958 ( .B1(n7751), .B2(n6486), .A(n6612), .ZN(n8472) );
  OR2_X1 U4959 ( .A1(n8815), .A2(n8814), .ZN(n8832) );
  XNOR2_X1 U4960 ( .A(n5625), .B(n5601), .ZN(n8363) );
  CLKBUF_X3 U4961 ( .A(n6333), .Z(n4455) );
  NAND2_X2 U4962 ( .A1(n6904), .A2(n6121), .ZN(n6317) );
  OR2_X1 U4963 ( .A1(n8791), .A2(n10157), .ZN(n8637) );
  INV_X1 U4964 ( .A(n6430), .ZN(n6672) );
  INV_X2 U4965 ( .A(n7928), .ZN(n6677) );
  CLKBUF_X1 U4966 ( .A(n8444), .Z(n4588) );
  CLKBUF_X1 U4967 ( .A(n6422), .Z(n7927) );
  INV_X1 U4968 ( .A(n8376), .ZN(n7460) );
  NAND2_X1 U4969 ( .A1(n4568), .A2(n4567), .ZN(n8632) );
  NAND2_X2 U4970 ( .A1(n4454), .A2(n6873), .ZN(n6430) );
  MUX2_X1 U4971 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10030), .S(n4462), .Z(n7452)
         );
  NAND2_X1 U4972 ( .A1(n4454), .A2(n6390), .ZN(n6453) );
  XNOR2_X1 U4973 ( .A(n5223), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U4974 ( .A(n5910), .B(n5909), .ZN(n6002) );
  NOR2_X1 U4975 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4675) );
  CLKBUF_X1 U4977 ( .A(n7509), .Z(n4448) );
  INV_X1 U4978 ( .A(n5181), .ZN(n4449) );
  XNOR2_X1 U4979 ( .A(n5173), .B(n5172), .ZN(n5175) );
  AOI21_X2 U4980 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8560) );
  NAND2_X2 U4981 ( .A1(n8106), .A2(n8105), .ZN(n8384) );
  NAND2_X2 U4982 ( .A1(n4919), .A2(n6556), .ZN(n4918) );
  XNOR2_X2 U4983 ( .A(n9652), .B(n9650), .ZN(n9646) );
  NOR2_X2 U4984 ( .A1(n8017), .A2(n9886), .ZN(n5833) );
  NAND2_X1 U4985 ( .A1(n7412), .A2(n8596), .ZN(n4450) );
  INV_X1 U4986 ( .A(n6690), .ZN(n4451) );
  AND2_X1 U4987 ( .A1(n5814), .A2(n8268), .ZN(n5107) );
  OR2_X1 U4988 ( .A1(n9357), .A2(n6305), .ZN(n9698) );
  NOR2_X1 U4989 ( .A1(n7323), .A2(n7321), .ZN(n7326) );
  BUF_X1 U4990 ( .A(n5588), .Z(n4459) );
  INV_X1 U4991 ( .A(n4469), .ZN(n5589) );
  XNOR2_X1 U4992 ( .A(n8444), .B(n6124), .ZN(n8235) );
  NAND2_X1 U4993 ( .A1(n6020), .A2(n6019), .ZN(n7279) );
  INV_X1 U4994 ( .A(n6695), .ZN(n8766) );
  OR2_X1 U4996 ( .A1(n5700), .A2(n5699), .ZN(n5719) );
  INV_X1 U4997 ( .A(n6326), .ZN(n6307) );
  OAI21_X1 U4998 ( .B1(n9296), .B2(n9294), .A(n9292), .ZN(n9387) );
  CLKBUF_X2 U4999 ( .A(n5350), .Z(n4456) );
  CLKBUF_X2 U5000 ( .A(n5350), .Z(n4457) );
  AND2_X1 U5001 ( .A1(n5175), .A2(n5176), .ZN(n5326) );
  INV_X1 U5002 ( .A(n9498), .ZN(n5320) );
  AND2_X1 U5003 ( .A1(n5247), .A2(n5246), .ZN(n7650) );
  CLKBUF_X3 U5004 ( .A(n7650), .Z(n4466) );
  INV_X1 U5005 ( .A(n7496), .ZN(n5280) );
  INV_X1 U5006 ( .A(n5748), .ZN(n6390) );
  NAND2_X1 U5007 ( .A1(n6002), .A2(n6004), .ZN(n6816) );
  OAI211_X1 U5008 ( .C1(n6816), .C2(n6868), .A(n6455), .B(n6454), .ZN(n6739)
         );
  NAND2_X1 U5009 ( .A1(n6527), .A2(n6526), .ZN(n7875) );
  NAND2_X1 U5010 ( .A1(n5660), .A2(n5659), .ZN(n9752) );
  NAND2_X1 U5011 ( .A1(n5446), .A2(n5445), .ZN(n9338) );
  NAND2_X1 U5012 ( .A1(n5401), .A2(n5400), .ZN(n7968) );
  NAND3_X1 U5013 ( .A1(n5168), .A2(n4554), .A3(n5119), .ZN(n4809) );
  INV_X4 U5014 ( .A(n6390), .ZN(n6873) );
  AND2_X2 U5015 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7777) );
  INV_X1 U5016 ( .A(n9791), .ZN(n10003) );
  OR2_X1 U5017 ( .A1(n5215), .A2(n5276), .ZN(n4452) );
  AND2_X1 U5018 ( .A1(n5120), .A2(n5170), .ZN(n4453) );
  NAND2_X2 U5019 ( .A1(n5396), .A2(n5395), .ZN(n5412) );
  NAND2_X2 U5020 ( .A1(n5394), .A2(n5393), .ZN(n5396) );
  NOR2_X2 U5021 ( .A1(n5616), .A2(n9333), .ZN(n4624) );
  NAND2_X2 U5022 ( .A1(n8010), .A2(n5806), .ZN(n9876) );
  NAND2_X2 U5023 ( .A1(n8009), .A2(n8149), .ZN(n8010) );
  INV_X2 U5024 ( .A(n7301), .ZN(n10046) );
  NAND2_X1 U5025 ( .A1(n6002), .A2(n6004), .ZN(n4454) );
  OAI21_X2 U5026 ( .B1(n8409), .B2(n5030), .A(n5028), .ZN(n8478) );
  AOI22_X2 U5027 ( .A1(n7279), .A2(n7278), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7281), .ZN(n6021) );
  AOI21_X2 U5028 ( .B1(n4611), .B2(n4515), .A(n8583), .ZN(n8585) );
  NAND2_X2 U5029 ( .A1(n9876), .A2(n8154), .ZN(n9854) );
  INV_X1 U5030 ( .A(n10150), .ZN(n4567) );
  NAND2_X2 U5031 ( .A1(n7777), .A2(n5187), .ZN(n4706) );
  AND2_X2 U5032 ( .A1(n6411), .A2(n5877), .ZN(n4482) );
  NAND2_X1 U5033 ( .A1(n6904), .A2(n7457), .ZN(n6333) );
  INV_X2 U5034 ( .A(n7452), .ZN(n7321) );
  AND2_X1 U5035 ( .A1(n5175), .A2(n10027), .ZN(n5350) );
  NAND2_X2 U5036 ( .A1(n9245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4864) );
  BUF_X4 U5037 ( .A(n5326), .Z(n4458) );
  NOR2_X2 U5038 ( .A1(n8950), .A2(n6821), .ZN(n6826) );
  AOI21_X2 U5039 ( .B1(n8270), .B2(n8266), .A(n8265), .ZN(n8334) );
  OAI21_X2 U5040 ( .B1(n5600), .B2(n5599), .A(n5598), .ZN(n5625) );
  INV_X1 U5041 ( .A(n7084), .ZN(n10157) );
  AND2_X4 U5042 ( .A1(n5181), .A2(n10027), .ZN(n5325) );
  XNOR2_X2 U5043 ( .A(n6382), .B(n6381), .ZN(n8369) );
  NAND2_X4 U5044 ( .A1(n4707), .A2(n4706), .ZN(n5748) );
  AND3_X2 U5045 ( .A1(n5294), .A2(n5292), .A3(n5293), .ZN(n8444) );
  AOI21_X1 U5046 ( .B1(n4719), .B2(n4873), .A(n4718), .ZN(n8741) );
  AND2_X1 U5047 ( .A1(n6851), .A2(n6850), .ZN(n9650) );
  NAND2_X1 U5048 ( .A1(n8169), .A2(n8168), .ZN(n9749) );
  AOI21_X1 U5049 ( .B1(n5453), .B2(n5153), .A(n5152), .ZN(n8079) );
  NAND2_X1 U5050 ( .A1(n9024), .A2(n8710), .ZN(n9041) );
  NAND2_X1 U5051 ( .A1(n8661), .A2(n8645), .ZN(n8599) );
  NAND2_X1 U5052 ( .A1(n7817), .A2(n7317), .ZN(n10071) );
  INV_X1 U5053 ( .A(n8786), .ZN(n7805) );
  CLKBUF_X2 U5054 ( .A(n7085), .Z(n10126) );
  CLKBUF_X1 U5055 ( .A(n6736), .Z(n7404) );
  INV_X4 U5056 ( .A(n4455), .ZN(n6141) );
  CLKBUF_X2 U5057 ( .A(n5349), .Z(n5767) );
  INV_X2 U5058 ( .A(n6697), .ZN(n4889) );
  AND4_X1 U5059 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n7383)
         );
  INV_X1 U5060 ( .A(n7363), .ZN(n8638) );
  CLKBUF_X2 U5061 ( .A(n6849), .Z(n4469) );
  NAND2_X1 U5062 ( .A1(n5873), .A2(n5867), .ZN(n6904) );
  BUF_X1 U5064 ( .A(n5588), .Z(n4465) );
  INV_X1 U5065 ( .A(n5316), .ZN(n5588) );
  INV_X1 U5066 ( .A(n6412), .ZN(n6690) );
  NAND2_X1 U5067 ( .A1(n8433), .A2(n6383), .ZN(n6401) );
  INV_X1 U5068 ( .A(n8369), .ZN(n6383) );
  INV_X2 U5069 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U5070 ( .A1(n9658), .A2(n4513), .ZN(n6102) );
  NOR2_X1 U5071 ( .A1(n8954), .A2(n4571), .ZN(n6798) );
  AOI21_X1 U5072 ( .B1(n9673), .B2(n10071), .A(n6113), .ZN(n6830) );
  AND2_X1 U5073 ( .A1(n4657), .A2(n4656), .ZN(n9973) );
  AND2_X1 U5074 ( .A1(n6110), .A2(n6357), .ZN(n9682) );
  NOR2_X1 U5075 ( .A1(n9899), .A2(n9900), .ZN(n4656) );
  NAND2_X1 U5076 ( .A1(n4750), .A2(n9685), .ZN(n9899) );
  NAND2_X1 U5077 ( .A1(n8917), .A2(n4564), .ZN(n5994) );
  NAND2_X1 U5078 ( .A1(n5993), .A2(n8906), .ZN(n8917) );
  NAND2_X1 U5079 ( .A1(n4861), .A2(n4493), .ZN(n9662) );
  OAI21_X1 U5080 ( .B1(n6776), .B2(n4871), .A(n8734), .ZN(n6802) );
  NAND2_X1 U5081 ( .A1(n8889), .A2(n8890), .ZN(n8888) );
  NAND2_X1 U5082 ( .A1(n9697), .A2(n5819), .ZN(n5820) );
  NAND2_X1 U5083 ( .A1(n9713), .A2(n9717), .ZN(n9697) );
  NAND2_X1 U5084 ( .A1(n8462), .A2(n8399), .ZN(n8515) );
  OAI21_X1 U5085 ( .B1(n9750), .B2(n5671), .A(n5670), .ZN(n9734) );
  NAND2_X1 U5086 ( .A1(n8536), .A2(n5020), .ZN(n8462) );
  AOI21_X1 U5087 ( .B1(n9387), .B2(n4682), .A(n4680), .ZN(n4679) );
  AOI21_X1 U5088 ( .B1(n5093), .B2(n5145), .A(n4532), .ZN(n5092) );
  NAND2_X1 U5089 ( .A1(n9009), .A2(n6628), .ZN(n8999) );
  NAND2_X1 U5090 ( .A1(n9650), .A2(n8290), .ZN(n8208) );
  AOI21_X1 U5091 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8342) );
  AND2_X1 U5092 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  OR2_X1 U5093 ( .A1(n8733), .A2(n6805), .ZN(n8752) );
  NAND2_X1 U5094 ( .A1(n4595), .A2(n8693), .ZN(n9063) );
  AND2_X1 U5095 ( .A1(n8734), .A2(n8735), .ZN(n8731) );
  NAND2_X1 U5096 ( .A1(n4958), .A2(n5765), .ZN(n9665) );
  NAND2_X1 U5097 ( .A1(n5000), .A2(n4998), .ZN(n9074) );
  NAND2_X1 U5098 ( .A1(n8367), .A2(n6847), .ZN(n4958) );
  CLKBUF_X1 U5099 ( .A(n8560), .Z(n4599) );
  AOI21_X1 U5100 ( .B1(n9364), .B2(n9366), .A(n9365), .ZN(n9380) );
  NAND2_X1 U5101 ( .A1(n5737), .A2(n5736), .ZN(n9690) );
  NAND2_X1 U5102 ( .A1(n5751), .A2(n5750), .ZN(n6359) );
  NAND2_X1 U5103 ( .A1(n6573), .A2(n6572), .ZN(n9080) );
  NAND2_X1 U5104 ( .A1(n6662), .A2(n6661), .ZN(n8451) );
  AOI21_X2 U5105 ( .B1(n5816), .B2(n5106), .A(n5105), .ZN(n5103) );
  NAND2_X1 U5106 ( .A1(n5696), .A2(n5695), .ZN(n9357) );
  NAND2_X1 U5107 ( .A1(n6640), .A2(n6639), .ZN(n9180) );
  NOR3_X1 U5108 ( .A1(n4473), .A2(n9752), .A3(n5121), .ZN(n5834) );
  NAND2_X1 U5109 ( .A1(n6651), .A2(n6650), .ZN(n8970) );
  NAND2_X1 U5110 ( .A1(n5716), .A2(n5715), .ZN(n9706) );
  NOR2_X2 U5111 ( .A1(n9749), .A2(n8116), .ZN(n5816) );
  NAND2_X1 U5112 ( .A1(n5680), .A2(n5679), .ZN(n9736) );
  NAND2_X1 U5113 ( .A1(n4967), .A2(n6191), .ZN(n7946) );
  NAND2_X1 U5114 ( .A1(n5640), .A2(n5639), .ZN(n9418) );
  OR2_X1 U5115 ( .A1(n6610), .A2(n8401), .ZN(n9024) );
  NAND2_X1 U5116 ( .A1(n5717), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5117 ( .A1(n5968), .A2(n4771), .ZN(n8830) );
  NAND2_X1 U5118 ( .A1(n5603), .A2(n5602), .ZN(n9791) );
  XNOR2_X1 U5119 ( .A(n5673), .B(n5672), .ZN(n7843) );
  NOR2_X1 U5120 ( .A1(n7391), .A2(n4499), .ZN(n7394) );
  INV_X1 U5121 ( .A(n5719), .ZN(n5717) );
  NAND2_X1 U5122 ( .A1(n5540), .A2(n5539), .ZN(n9842) );
  AND2_X1 U5123 ( .A1(n7269), .A2(n7271), .ZN(n7391) );
  NAND2_X1 U5124 ( .A1(n5591), .A2(n5590), .ZN(n10006) );
  NAND2_X1 U5125 ( .A1(n6601), .A2(n6600), .ZN(n9060) );
  NAND2_X1 U5126 ( .A1(n6576), .A2(n6575), .ZN(n9225) );
  NAND2_X1 U5127 ( .A1(n7509), .A2(n5111), .ZN(n5110) );
  NAND2_X1 U5128 ( .A1(n6567), .A2(n6566), .ZN(n9231) );
  NAND2_X1 U5129 ( .A1(n4717), .A2(n6557), .ZN(n9149) );
  NAND2_X1 U5130 ( .A1(n5500), .A2(n5499), .ZN(n9886) );
  NAND2_X1 U5131 ( .A1(n5962), .A2(n4768), .ZN(n5963) );
  NAND2_X1 U5132 ( .A1(n4790), .A2(n8305), .ZN(n7509) );
  OR2_X1 U5133 ( .A1(n9963), .A2(n5803), .ZN(n9874) );
  NOR2_X1 U5134 ( .A1(n6534), .A2(n5076), .ZN(n5075) );
  NAND2_X1 U5135 ( .A1(n6547), .A2(n6546), .ZN(n9239) );
  NAND2_X1 U5136 ( .A1(n5461), .A2(n5460), .ZN(n8082) );
  AND3_X1 U5137 ( .A1(n7636), .A2(n6510), .A3(n4607), .ZN(n6511) );
  XNOR2_X1 U5138 ( .A(n6021), .B(n6478), .ZN(n7520) );
  NAND2_X1 U5139 ( .A1(n6537), .A2(n6536), .ZN(n8065) );
  AND2_X1 U5140 ( .A1(n7160), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7284) );
  XNOR2_X1 U5141 ( .A(n7993), .B(n8783), .ZN(n7870) );
  CLKBUF_X1 U5142 ( .A(n7993), .Z(n4615) );
  INV_X2 U5143 ( .A(n9814), .ZN(n10057) );
  AND2_X1 U5144 ( .A1(n8660), .A2(n8644), .ZN(n8598) );
  NAND2_X1 U5145 ( .A1(n6506), .A2(n6505), .ZN(n7909) );
  INV_X4 U5146 ( .A(n9850), .ZN(n10063) );
  NAND2_X1 U5147 ( .A1(n5101), .A2(n5791), .ZN(n7297) );
  OR2_X1 U5148 ( .A1(n7559), .A2(n7862), .ZN(n8662) );
  NAND2_X1 U5149 ( .A1(n5370), .A2(n4762), .ZN(n9325) );
  NOR2_X1 U5150 ( .A1(n10041), .A2(n9514), .ZN(n9636) );
  NAND2_X1 U5151 ( .A1(n4761), .A2(n5238), .ZN(n9493) );
  NAND2_X1 U5152 ( .A1(n6488), .A2(n6489), .ZN(n7541) );
  INV_X1 U5153 ( .A(n10117), .ZN(n8623) );
  NAND2_X1 U5154 ( .A1(n6737), .A2(n4678), .ZN(n10117) );
  INV_X1 U5155 ( .A(n8785), .ZN(n7862) );
  INV_X2 U5156 ( .A(n6329), .ZN(n6318) );
  AND3_X1 U5157 ( .A1(n5264), .A2(n5263), .A3(n5262), .ZN(n10067) );
  NAND4_X2 U5158 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n8791)
         );
  NAND4_X2 U5159 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n8785)
         );
  AND3_X2 U5160 ( .A1(n5309), .A2(n4549), .A3(n5308), .ZN(n8376) );
  BUF_X2 U5161 ( .A(n7111), .Z(n4460) );
  INV_X1 U5162 ( .A(n7383), .ZN(n8792) );
  CLKBUF_X3 U5163 ( .A(n7111), .Z(n8107) );
  AND2_X1 U5164 ( .A1(n6399), .A2(n6398), .ZN(n7085) );
  NOR2_X1 U5165 ( .A1(n8803), .A2(n5945), .ZN(n5949) );
  OR2_X2 U5166 ( .A1(n6904), .A2(n6865), .ZN(n9469) );
  NOR2_X2 U5167 ( .A1(n7017), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U5168 ( .A1(n6690), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6427) );
  OAI211_X1 U5169 ( .C1(n6816), .C2(n8798), .A(n6443), .B(n6444), .ZN(n7363)
         );
  AND3_X1 U5170 ( .A1(n6403), .A2(n6404), .A3(n6405), .ZN(n6407) );
  AOI21_X1 U5171 ( .B1(n5941), .B2(n8801), .A(n8800), .ZN(n8803) );
  CLKBUF_X2 U5172 ( .A(n6849), .Z(n4470) );
  NAND2_X2 U5173 ( .A1(n7011), .A2(n8771), .ZN(n6697) );
  CLKBUF_X3 U5174 ( .A(n6401), .Z(n7928) );
  NAND2_X1 U5175 ( .A1(n5824), .A2(n5825), .ZN(n5316) );
  NAND2_X1 U5176 ( .A1(n6384), .A2(n8369), .ZN(n6412) );
  XNOR2_X1 U5177 ( .A(n5900), .B(n5899), .ZN(n7810) );
  XNOR2_X1 U5178 ( .A(n6728), .B(n10304), .ZN(n8365) );
  NAND2_X1 U5179 ( .A1(n5174), .A2(n4527), .ZN(n4658) );
  NAND2_X1 U5180 ( .A1(n5849), .A2(n5848), .ZN(n8090) );
  NAND2_X1 U5181 ( .A1(n6686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6728) );
  XNOR2_X1 U5182 ( .A(n6685), .B(n6684), .ZN(n8612) );
  XNOR2_X1 U5183 ( .A(n5786), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8300) );
  OR2_X2 U5184 ( .A1(n5218), .A2(n10022), .ZN(n5220) );
  NAND2_X1 U5185 ( .A1(n4809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5173) );
  NAND3_X1 U5186 ( .A1(n5913), .A2(n5914), .A3(n5140), .ZN(n6004) );
  XNOR2_X1 U5187 ( .A(n5778), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U5188 ( .A1(n5221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U5189 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5910) );
  NOR2_X1 U5190 ( .A1(n7187), .A2(n7188), .ZN(n7186) );
  AND3_X1 U5191 ( .A1(n4453), .A2(n5167), .A3(n5171), .ZN(n5119) );
  OR2_X1 U5192 ( .A1(n6380), .A2(n5055), .ZN(n6382) );
  NOR2_X1 U5193 ( .A1(n7173), .A2(n5935), .ZN(n7187) );
  OAI21_X1 U5194 ( .B1(n5908), .B2(P2_IR_REG_26__SCAN_IN), .A(n5912), .ZN(
        n5914) );
  XNOR2_X1 U5195 ( .A(n5944), .B(n5943), .ZN(n8798) );
  INV_X1 U5196 ( .A(n4672), .ZN(n5916) );
  XNOR2_X1 U5197 ( .A(n5242), .B(SI_6_), .ZN(n5240) );
  BUF_X1 U5198 ( .A(n5888), .Z(n5881) );
  AND2_X1 U5199 ( .A1(n5165), .A2(n5164), .ZN(n4751) );
  NOR2_X1 U5200 ( .A1(n4597), .A2(n5907), .ZN(n5100) );
  AND2_X1 U5201 ( .A1(n5164), .A2(n5167), .ZN(n5113) );
  OAI211_X2 U5202 ( .C1(n5936), .C2(n4900), .A(n4899), .B(n4898), .ZN(n7185)
         );
  NOR2_X1 U5203 ( .A1(n4674), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5204 ( .A1(n5868), .A2(n5871), .ZN(n5169) );
  AND3_X1 U5205 ( .A1(n5161), .A2(n5160), .A3(n5159), .ZN(n5781) );
  AND2_X1 U5206 ( .A1(n5158), .A2(n5157), .ZN(n5518) );
  AND2_X1 U5207 ( .A1(n5163), .A2(n5224), .ZN(n5164) );
  AND2_X1 U5208 ( .A1(n5156), .A2(n5155), .ZN(n5517) );
  INV_X1 U5209 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5937) );
  NOR2_X1 U5210 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5155) );
  NOR2_X1 U5211 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5158) );
  NOR2_X1 U5212 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5156) );
  INV_X1 U5213 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5885) );
  NOR2_X1 U5214 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4965) );
  NOR2_X1 U5215 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5895) );
  NOR2_X1 U5216 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5893) );
  NOR2_X2 U5217 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5984) );
  NOR2_X1 U5218 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4676) );
  INV_X1 U5219 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4865) );
  INV_X1 U5220 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5877) );
  INV_X1 U5221 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5056) );
  INV_X4 U5222 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5223 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5886) );
  OAI21_X2 U5224 ( .B1(n7635), .B2(n7639), .A(n8666), .ZN(n7581) );
  AOI211_X2 U5225 ( .C1(n8351), .C2(n8350), .A(n8349), .B(n8348), .ZN(n8352)
         );
  OAI21_X1 U5226 ( .B1(n9020), .B2(n8700), .A(n5149), .ZN(n6750) );
  NAND2_X1 U5227 ( .A1(n5824), .A2(n5825), .ZN(n4461) );
  NAND2_X1 U5228 ( .A1(n5824), .A2(n5825), .ZN(n4462) );
  OAI21_X2 U5229 ( .B1(n7235), .B2(n5088), .A(n5086), .ZN(n10105) );
  NAND2_X2 U5230 ( .A1(n6435), .A2(n6434), .ZN(n7235) );
  NAND3_X2 U5231 ( .A1(n8310), .A2(n8245), .A3(n5110), .ZN(n7699) );
  AND2_X1 U5232 ( .A1(n5781), .A2(n5165), .ZN(n5112) );
  INV_X1 U5233 ( .A(n6430), .ZN(n4463) );
  XNOR2_X1 U5234 ( .A(n8576), .B(n6807), .ZN(n8948) );
  OAI211_X2 U5235 ( .C1(n6453), .C2(n5061), .A(n5060), .B(n5059), .ZN(n7016)
         );
  NAND2_X1 U5236 ( .A1(n4707), .A2(n4706), .ZN(n4464) );
  NAND2_X1 U5237 ( .A1(n9802), .A2(n8330), .ZN(n9770) );
  NAND2_X2 U5238 ( .A1(n7971), .A2(n5102), .ZN(n8009) );
  AOI21_X2 U5239 ( .B1(n8999), .B2(n6638), .A(n6637), .ZN(n8982) );
  NAND2_X2 U5240 ( .A1(n7972), .A2(n8247), .ZN(n7971) );
  NAND2_X2 U5241 ( .A1(n4764), .A2(n8144), .ZN(n7972) );
  NOR2_X4 U5242 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5303) );
  BUF_X4 U5243 ( .A(n6690), .Z(n4467) );
  CLKBUF_X1 U5244 ( .A(n6849), .Z(n4468) );
  NAND2_X1 U5245 ( .A1(n4461), .A2(n6390), .ZN(n6849) );
  OAI21_X2 U5246 ( .B1(n7297), .B2(n5794), .A(n5793), .ZN(n7550) );
  NOR2_X1 U5247 ( .A1(n8648), .A2(n6476), .ZN(n8659) );
  NOR2_X1 U5248 ( .A1(n8718), .A2(n8719), .ZN(n4987) );
  NAND2_X1 U5249 ( .A1(n7511), .A2(n7653), .ZN(n4760) );
  AND2_X1 U5250 ( .A1(n8358), .A2(n8223), .ZN(n8292) );
  INV_X1 U5251 ( .A(n8300), .ZN(n8260) );
  NAND2_X1 U5252 ( .A1(n7428), .A2(n8260), .ZN(n8356) );
  INV_X1 U5253 ( .A(n4458), .ZN(n5771) );
  NAND2_X1 U5254 ( .A1(n4888), .A2(n4887), .ZN(n8648) );
  NAND2_X1 U5255 ( .A1(n8665), .A2(n6697), .ZN(n4887) );
  NAND2_X1 U5256 ( .A1(n8641), .A2(n4889), .ZN(n4888) );
  AND2_X1 U5257 ( .A1(n4891), .A2(n4890), .ZN(n8698) );
  NOR2_X1 U5258 ( .A1(n9077), .A2(n8689), .ZN(n4890) );
  OR2_X1 U5259 ( .A1(n8216), .A2(n8209), .ZN(n8210) );
  INV_X1 U5260 ( .A(n5598), .ZN(n4963) );
  INV_X1 U5261 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5157) );
  INV_X1 U5262 ( .A(n5494), .ZN(n4942) );
  AND2_X1 U5263 ( .A1(n5049), .A2(n4548), .ZN(n5048) );
  NAND2_X1 U5264 ( .A1(n8446), .A2(n5050), .ZN(n5049) );
  NAND2_X1 U5265 ( .A1(n7189), .A2(n6009), .ZN(n6010) );
  INV_X1 U5266 ( .A(n7071), .ZN(n6038) );
  NAND2_X1 U5267 ( .A1(n5950), .A2(n6868), .ZN(n4909) );
  AND3_X1 U5268 ( .A1(n4906), .A2(n4903), .A3(n4553), .ZN(n5953) );
  NAND2_X1 U5269 ( .A1(n4785), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U5270 ( .A1(n8888), .A2(n5990), .ZN(n5993) );
  AOI21_X1 U5271 ( .B1(n8903), .B2(n8904), .A(n6088), .ZN(n6093) );
  AND2_X1 U5272 ( .A1(n9041), .A2(n4543), .ZN(n5099) );
  NAND2_X1 U5273 ( .A1(n4717), .A2(n4715), .ZN(n9073) );
  NOR2_X1 U5274 ( .A1(n8489), .A2(n4716), .ZN(n4715) );
  INV_X1 U5275 ( .A(n6557), .ZN(n4716) );
  AND2_X1 U5276 ( .A1(n6884), .A2(n6794), .ZN(n6992) );
  AND2_X1 U5277 ( .A1(n6167), .A2(n6168), .ZN(n4966) );
  OR2_X1 U5278 ( .A1(n9404), .A2(n4990), .ZN(n4989) );
  INV_X1 U5279 ( .A(n10027), .ZN(n5176) );
  AOI21_X1 U5280 ( .B1(n4643), .B2(n4475), .A(n4857), .ZN(n4642) );
  INV_X1 U5281 ( .A(n9665), .ZN(n5837) );
  INV_X1 U5282 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U5283 ( .A1(n5365), .A2(n5009), .ZN(n5008) );
  INV_X1 U5284 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U5285 ( .A1(n5044), .A2(n5043), .ZN(n5042) );
  NAND2_X1 U5286 ( .A1(n5046), .A2(n5045), .ZN(n5044) );
  OAI21_X1 U5287 ( .B1(n8427), .B2(n8446), .A(n5048), .ZN(n5043) );
  INV_X1 U5288 ( .A(n8427), .ZN(n5046) );
  NAND2_X1 U5289 ( .A1(n7394), .A2(n7393), .ZN(n7472) );
  NOR2_X1 U5290 ( .A1(n8417), .A2(n5032), .ZN(n5031) );
  INV_X1 U5291 ( .A(n8412), .ZN(n5032) );
  NAND2_X1 U5292 ( .A1(n8394), .A2(n8533), .ZN(n8536) );
  NAND2_X1 U5293 ( .A1(n5019), .A2(n5015), .ZN(n7148) );
  AND2_X1 U5294 ( .A1(n7112), .A2(n5018), .ZN(n5015) );
  INV_X1 U5295 ( .A(n5138), .ZN(n5018) );
  INV_X1 U5296 ( .A(n6424), .ZN(n6688) );
  OR2_X1 U5297 ( .A1(n6767), .A2(n6919), .ZN(n6027) );
  INV_X2 U5298 ( .A(n6422), .ZN(n6680) );
  INV_X1 U5299 ( .A(n7588), .ZN(n4729) );
  NAND2_X1 U5300 ( .A1(n8838), .A2(n8837), .ZN(n6070) );
  INV_X1 U5301 ( .A(n6004), .ZN(n6695) );
  NAND2_X1 U5302 ( .A1(n6642), .A2(n6641), .ZN(n6652) );
  INV_X1 U5303 ( .A(n6643), .ZN(n6642) );
  OR2_X1 U5304 ( .A1(n6604), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6613) );
  INV_X1 U5305 ( .A(n8612), .ZN(n8584) );
  INV_X1 U5306 ( .A(n9081), .ZN(n9104) );
  NAND2_X1 U5307 ( .A1(n6743), .A2(n5001), .ZN(n5000) );
  NOR2_X1 U5308 ( .A1(n8674), .A2(n5002), .ZN(n5001) );
  INV_X1 U5309 ( .A(n8676), .ZN(n5002) );
  NAND2_X2 U5310 ( .A1(n8662), .A2(n8646), .ZN(n8601) );
  OR2_X1 U5311 ( .A1(n8790), .A2(n7363), .ZN(n6445) );
  NAND2_X1 U5312 ( .A1(n6755), .A2(n7307), .ZN(n10124) );
  NAND2_X1 U5313 ( .A1(n6765), .A2(n6764), .ZN(n6771) );
  XNOR2_X1 U5314 ( .A(n8775), .B(n9169), .ZN(n8610) );
  NAND2_X1 U5315 ( .A1(n4889), .A2(n7017), .ZN(n10125) );
  NAND2_X1 U5316 ( .A1(n6750), .A2(n8713), .ZN(n9008) );
  NAND2_X1 U5317 ( .A1(n7914), .A2(n8675), .ZN(n6743) );
  NAND2_X1 U5318 ( .A1(n7826), .A2(n8618), .ZN(n7914) );
  INV_X1 U5319 ( .A(n10125), .ZN(n9090) );
  OR2_X1 U5320 ( .A1(n6697), .A2(n6754), .ZN(n7307) );
  AND2_X1 U5321 ( .A1(n6992), .A2(n6892), .ZN(n7020) );
  NAND2_X1 U5322 ( .A1(n5051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6711) );
  XNOR2_X1 U5323 ( .A(n5952), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7162) );
  OR2_X1 U5324 ( .A1(n5946), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5928) );
  INV_X1 U5325 ( .A(n4683), .ZN(n4682) );
  OAI21_X1 U5326 ( .B1(n9388), .B2(n6303), .A(n9355), .ZN(n4683) );
  NAND2_X1 U5327 ( .A1(n4652), .A2(n5727), .ZN(n9687) );
  OAI21_X1 U5328 ( .B1(n9734), .B2(n4838), .A(n4835), .ZN(n4652) );
  AOI21_X1 U5329 ( .B1(n4837), .B2(n4841), .A(n4836), .ZN(n4835) );
  NOR2_X1 U5330 ( .A1(n5597), .A2(n4649), .ZN(n4648) );
  INV_X1 U5331 ( .A(n5576), .ZN(n4649) );
  OR2_X1 U5332 ( .A1(n8297), .A2(n8300), .ZN(n7317) );
  AND2_X1 U5333 ( .A1(n5154), .A2(n5798), .ZN(n5111) );
  NAND2_X1 U5334 ( .A1(n6345), .A2(n8260), .ZN(n9885) );
  NAND2_X1 U5335 ( .A1(n4461), .A2(n6873), .ZN(n5336) );
  AND2_X1 U5336 ( .A1(n5866), .A2(n7999), .ZN(n5867) );
  INV_X1 U5337 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U5338 ( .A1(n5564), .A2(n5563), .ZN(n5587) );
  INV_X1 U5339 ( .A(n9082), .ZN(n8466) );
  OR2_X1 U5340 ( .A1(n10172), .A2(n8762), .ZN(n10122) );
  AND2_X1 U5341 ( .A1(n9435), .A2(n6325), .ZN(n9265) );
  AND2_X1 U5342 ( .A1(n9262), .A2(n9263), .ZN(n6325) );
  AOI211_X1 U5343 ( .C1(n8630), .C2(n8629), .A(n10119), .B(n8628), .ZN(n8636)
         );
  INV_X1 U5344 ( .A(n8130), .ZN(n4807) );
  OAI21_X1 U5345 ( .B1(n8126), .B2(n8125), .A(n8297), .ZN(n8127) );
  NAND2_X1 U5346 ( .A1(n4576), .A2(n8666), .ZN(n8668) );
  OAI21_X1 U5347 ( .B1(n4514), .B2(n4578), .A(n4577), .ZN(n4576) );
  OAI21_X1 U5348 ( .B1(n8670), .B2(n4517), .A(n4896), .ZN(n4895) );
  AOI21_X1 U5349 ( .B1(n8673), .B2(n6697), .A(n8672), .ZN(n4896) );
  OAI21_X1 U5350 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n4713) );
  INV_X1 U5351 ( .A(n4580), .ZN(n4579) );
  OAI21_X1 U5352 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n4580) );
  AND2_X1 U5353 ( .A1(n8716), .A2(n4574), .ZN(n4870) );
  NOR2_X1 U5354 ( .A1(n4723), .A2(n4575), .ZN(n4574) );
  OR2_X1 U5355 ( .A1(n5144), .A2(n8705), .ZN(n4866) );
  NOR3_X1 U5356 ( .A1(n8703), .A2(n8712), .A3(n4523), .ZN(n4867) );
  NOR2_X1 U5357 ( .A1(n8708), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U5358 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U5359 ( .A1(n4879), .A2(n4524), .ZN(n4874) );
  NOR2_X1 U5360 ( .A1(n4872), .A2(n4871), .ZN(n4879) );
  INV_X1 U5361 ( .A(n8730), .ZN(n4872) );
  NAND2_X1 U5362 ( .A1(n8245), .A2(n4629), .ZN(n4628) );
  AND2_X1 U5363 ( .A1(n8242), .A2(n8243), .ZN(n4629) );
  OR3_X1 U5364 ( .A1(n8238), .A2(n8237), .A3(n8236), .ZN(n8241) );
  OR2_X1 U5365 ( .A1(n9196), .A2(n9000), .ZN(n8617) );
  NOR2_X1 U5366 ( .A1(n8601), .A2(n4995), .ZN(n4994) );
  INV_X1 U5367 ( .A(n8645), .ZN(n4995) );
  NOR2_X1 U5368 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5887) );
  INV_X1 U5369 ( .A(n8211), .ZN(n8216) );
  INV_X1 U5370 ( .A(n8285), .ZN(n4815) );
  NOR2_X1 U5371 ( .A1(n9338), .A2(n7821), .ZN(n5136) );
  NAND2_X1 U5372 ( .A1(n9325), .A2(n5372), .ZN(n8122) );
  NAND2_X1 U5373 ( .A1(n4787), .A2(n4791), .ZN(n7615) );
  AOI21_X1 U5374 ( .B1(n4793), .B2(n8305), .A(n4792), .ZN(n4791) );
  INV_X1 U5375 ( .A(n5797), .ZN(n4793) );
  INV_X1 U5376 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10466) );
  INV_X1 U5377 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5559) );
  OAI21_X1 U5378 ( .B1(n5748), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4635), .ZN(
        n5362) );
  NAND2_X1 U5379 ( .A1(n5748), .A2(n6889), .ZN(n4635) );
  INV_X1 U5380 ( .A(n8963), .ZN(n4823) );
  INV_X1 U5381 ( .A(n8755), .ZN(n4821) );
  NOR3_X1 U5382 ( .A1(n8609), .A2(n4880), .A3(n8990), .ZN(n4822) );
  AND2_X1 U5383 ( .A1(n8580), .A2(n8579), .ZN(n8737) );
  AND2_X1 U5384 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  OR2_X1 U5385 ( .A1(n6412), .A2(n6402), .ZN(n6403) );
  NOR2_X1 U5386 ( .A1(n7186), .A2(n5148), .ZN(n5940) );
  NOR2_X1 U5387 ( .A1(n8857), .A2(n6535), .ZN(n4779) );
  OR2_X1 U5388 ( .A1(n8857), .A2(n10381), .ZN(n4777) );
  NAND2_X1 U5389 ( .A1(n6664), .A2(n6663), .ZN(n6675) );
  INV_X1 U5390 ( .A(n6665), .ZN(n6664) );
  INV_X1 U5391 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U5392 ( .A1(n8793), .A2(n7016), .ZN(n8625) );
  NAND2_X1 U5393 ( .A1(n8625), .A2(n10116), .ZN(n10118) );
  OR2_X1 U5394 ( .A1(n6714), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U5395 ( .A1(n5098), .A2(n8589), .ZN(n5097) );
  NAND2_X1 U5396 ( .A1(n6611), .A2(n9029), .ZN(n5098) );
  INV_X1 U5397 ( .A(n9054), .ZN(n8401) );
  OR2_X1 U5398 ( .A1(n9219), .A2(n8466), .ZN(n8695) );
  INV_X1 U5399 ( .A(n6201), .ZN(n4969) );
  INV_X1 U5400 ( .A(n7457), .ZN(n6121) );
  OR2_X1 U5401 ( .A1(n6163), .A2(n7683), .ZN(n6168) );
  NOR2_X1 U5402 ( .A1(n4476), .A2(n4509), .ZN(n4978) );
  NOR2_X1 U5403 ( .A1(n5447), .A2(n7133), .ZN(n4625) );
  NAND2_X1 U5404 ( .A1(n6289), .A2(n6290), .ZN(n4705) );
  AND2_X1 U5405 ( .A1(n8254), .A2(n4630), .ZN(n8256) );
  NOR2_X1 U5406 ( .A1(n9749), .A2(n4631), .ZN(n4630) );
  OR3_X1 U5407 ( .A1(n9855), .A2(n8252), .A3(n9838), .ZN(n8253) );
  AND2_X1 U5408 ( .A1(n8212), .A2(n8115), .ZN(n8343) );
  NOR2_X1 U5409 ( .A1(n9689), .A2(n6359), .ZN(n5835) );
  NAND2_X1 U5410 ( .A1(n4958), .A2(n4956), .ZN(n8281) );
  NOR2_X1 U5411 ( .A1(n5775), .A2(n4957), .ZN(n4956) );
  INV_X1 U5412 ( .A(n5765), .ZN(n4957) );
  NOR2_X1 U5413 ( .A1(n4843), .A2(n5707), .ZN(n4842) );
  INV_X1 U5414 ( .A(n5687), .ZN(n4843) );
  INV_X1 U5415 ( .A(n9475), .ZN(n6305) );
  INV_X1 U5416 ( .A(n8168), .ZN(n5105) );
  INV_X1 U5417 ( .A(n5107), .ZN(n5106) );
  INV_X1 U5418 ( .A(n8335), .ZN(n4759) );
  AND2_X1 U5419 ( .A1(n4639), .A2(n4555), .ZN(n4643) );
  OR2_X1 U5420 ( .A1(n4645), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U5421 ( .A1(n4641), .A2(n4644), .ZN(n4640) );
  NOR2_X1 U5422 ( .A1(n9842), .A2(n9867), .ZN(n5125) );
  OR2_X1 U5423 ( .A1(n5501), .A2(n7481), .ZN(n5525) );
  NOR2_X1 U5424 ( .A1(n4848), .A2(n8245), .ZN(n4650) );
  INV_X1 U5425 ( .A(n5430), .ZN(n4848) );
  NAND2_X1 U5426 ( .A1(n5430), .A2(n4847), .ZN(n4846) );
  INV_X1 U5427 ( .A(n5406), .ZN(n4847) );
  INV_X1 U5428 ( .A(n7722), .ZN(n4801) );
  OAI21_X1 U5429 ( .B1(n7720), .B2(n4801), .A(n8122), .ZN(n4800) );
  AND2_X1 U5430 ( .A1(n7516), .A2(n4466), .ZN(n5117) );
  NAND2_X1 U5431 ( .A1(n5232), .A2(n7692), .ZN(n5798) );
  NAND2_X1 U5432 ( .A1(n9494), .A2(n7516), .ZN(n7616) );
  NAND2_X1 U5433 ( .A1(n8305), .A2(n5797), .ZN(n7367) );
  NAND2_X1 U5434 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5265) );
  NAND2_X1 U5435 ( .A1(n7615), .A2(n7616), .ZN(n7721) );
  INV_X1 U5436 ( .A(SI_15_), .ZN(n10453) );
  AOI21_X1 U5437 ( .B1(n4947), .B2(n4949), .A(n4945), .ZN(n4944) );
  INV_X1 U5438 ( .A(n5710), .ZN(n4945) );
  AND2_X1 U5439 ( .A1(n5743), .A2(n5714), .ZN(n5728) );
  AND2_X1 U5440 ( .A1(n5710), .A2(n5694), .ZN(n5708) );
  AND2_X1 U5441 ( .A1(n5690), .A2(n5678), .ZN(n5688) );
  INV_X1 U5442 ( .A(n5649), .ZN(n4964) );
  AND2_X1 U5443 ( .A1(n5674), .A2(n5657), .ZN(n5672) );
  NAND2_X1 U5444 ( .A1(n4940), .A2(n4938), .ZN(n5583) );
  NAND2_X1 U5445 ( .A1(n4474), .A2(n4530), .ZN(n4938) );
  OR2_X1 U5446 ( .A1(n5473), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5474) );
  OR2_X1 U5447 ( .A1(n5397), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U5448 ( .A1(n5275), .A2(n5216), .ZN(n4935) );
  NOR2_X1 U5449 ( .A1(n5911), .A2(n5055), .ZN(n5912) );
  INV_X1 U5450 ( .A(n7097), .ZN(n5017) );
  INV_X1 U5451 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U5452 ( .A1(n4492), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5453 ( .A1(n5013), .A2(n4501), .ZN(n4665) );
  OR2_X1 U5454 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  AOI211_X1 U5455 ( .C1(n7868), .C2(n8783), .A(n7867), .B(n8590), .ZN(n7873)
         );
  NAND2_X1 U5456 ( .A1(n4518), .A2(n7558), .ZN(n4666) );
  NAND2_X1 U5457 ( .A1(n8524), .A2(n8412), .ZN(n8454) );
  XOR2_X1 U5458 ( .A(n7016), .B(n7111), .Z(n7090) );
  OR2_X1 U5459 ( .A1(n8760), .A2(n6754), .ZN(n4885) );
  AND2_X1 U5460 ( .A1(n8759), .A2(n8762), .ZN(n4881) );
  XNOR2_X1 U5461 ( .A(n7185), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U5462 ( .A1(n4619), .A2(n4618), .ZN(n7191) );
  NAND2_X1 U5463 ( .A1(n7185), .A2(n6413), .ZN(n4618) );
  OR2_X1 U5464 ( .A1(n7185), .A2(n6413), .ZN(n4619) );
  OR2_X1 U5465 ( .A1(n5940), .A2(n6038), .ZN(n5941) );
  NAND2_X1 U5466 ( .A1(n4901), .A2(n5941), .ZN(n8801) );
  AND2_X1 U5467 ( .A1(n4902), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5468 ( .A1(n7068), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6012) );
  AND2_X1 U5469 ( .A1(n7063), .A2(n6040), .ZN(n8796) );
  NAND2_X1 U5470 ( .A1(n8796), .A2(n8795), .ZN(n8794) );
  NAND2_X1 U5471 ( .A1(n7203), .A2(n4908), .ZN(n4906) );
  NOR2_X1 U5472 ( .A1(n10083), .A2(n10303), .ZN(n4908) );
  INV_X1 U5473 ( .A(n10083), .ZN(n4904) );
  AND2_X1 U5474 ( .A1(n4907), .A2(n4909), .ZN(n10082) );
  NAND2_X1 U5475 ( .A1(n7203), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U5476 ( .A1(n10097), .A2(n6048), .ZN(n7159) );
  NAND2_X1 U5477 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  OR2_X1 U5478 ( .A1(n5959), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5964) );
  INV_X1 U5479 ( .A(n4728), .ZN(n4727) );
  OAI21_X1 U5480 ( .B1(n4729), .B2(n6058), .A(n6062), .ZN(n4728) );
  OAI21_X1 U5481 ( .B1(n7520), .B2(n4769), .A(n4765), .ZN(n4772) );
  NAND2_X1 U5482 ( .A1(n7587), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4769) );
  INV_X1 U5483 ( .A(n4766), .ZN(n4765) );
  OAI21_X1 U5484 ( .B1(n6021), .B2(n4767), .A(n4773), .ZN(n4766) );
  INV_X1 U5485 ( .A(n4562), .ZN(n4920) );
  AOI21_X1 U5486 ( .B1(n8917), .B2(n4917), .A(n4916), .ZN(n4915) );
  INV_X1 U5487 ( .A(n8918), .ZN(n4916) );
  AOI21_X1 U5488 ( .B1(n4985), .B2(n4982), .A(n8586), .ZN(n4980) );
  INV_X1 U5489 ( .A(n4982), .ZN(n4981) );
  NOR2_X1 U5490 ( .A1(n8727), .A2(n8724), .ZN(n4982) );
  OR2_X1 U5491 ( .A1(n6652), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6665) );
  INV_X1 U5492 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n4824) );
  INV_X1 U5493 ( .A(n4826), .ZN(n4825) );
  INV_X1 U5494 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5495 ( .A1(n6376), .A2(n4831), .ZN(n6602) );
  OR2_X1 U5496 ( .A1(n6497), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6517) );
  INV_X1 U5497 ( .A(n8661), .ZN(n4997) );
  OR3_X1 U5498 ( .A1(n6787), .A2(n6993), .A3(n6727), .ZN(n6760) );
  NAND2_X1 U5499 ( .A1(n6804), .A2(n6803), .ZN(n8733) );
  INV_X1 U5500 ( .A(n8776), .ZN(n8966) );
  OR2_X1 U5501 ( .A1(n8727), .A2(n8586), .ZN(n8963) );
  OR2_X1 U5502 ( .A1(n8510), .A2(n8779), .ZN(n5058) );
  CLKBUF_X1 U5503 ( .A(n8997), .Z(n4614) );
  OAI21_X1 U5504 ( .B1(n9074), .B2(n8688), .A(n4596), .ZN(n4595) );
  AND2_X1 U5505 ( .A1(n6746), .A2(n8691), .ZN(n4596) );
  AND2_X1 U5506 ( .A1(n9089), .A2(n5067), .ZN(n5066) );
  NAND2_X1 U5507 ( .A1(n7580), .A2(n5004), .ZN(n7826) );
  AND2_X1 U5508 ( .A1(n6742), .A2(n8620), .ZN(n5004) );
  INV_X1 U5509 ( .A(n5079), .ZN(n5078) );
  NAND2_X1 U5510 ( .A1(n7581), .A2(n7870), .ZN(n7580) );
  NAND2_X1 U5511 ( .A1(n4608), .A2(n7869), .ZN(n4607) );
  INV_X1 U5512 ( .A(n6816), .ZN(n6599) );
  CLKBUF_X1 U5513 ( .A(n7423), .Z(n7424) );
  NAND2_X1 U5514 ( .A1(n7810), .A2(n7797), .ZN(n10172) );
  INV_X1 U5515 ( .A(n8029), .ZN(n5891) );
  XNOR2_X1 U5516 ( .A(n5905), .B(n5056), .ZN(n7844) );
  NAND2_X1 U5517 ( .A1(n5901), .A2(n5885), .ZN(n5904) );
  CLKBUF_X1 U5518 ( .A(n6002), .Z(n6003) );
  INV_X1 U5519 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U5520 ( .A1(n5054), .A2(n5052), .ZN(n5883) );
  INV_X1 U5521 ( .A(n5053), .ZN(n5052) );
  OR2_X1 U5522 ( .A1(n5901), .A2(n5055), .ZN(n5054) );
  OAI21_X1 U5523 ( .B1(n4504), .B2(n5055), .A(n6703), .ZN(n5053) );
  XNOR2_X1 U5524 ( .A(n5972), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6525) );
  INV_X1 U5525 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5929) );
  INV_X1 U5526 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5943) );
  INV_X1 U5527 ( .A(n4698), .ZN(n4697) );
  OAI21_X1 U5528 ( .B1(n9329), .B2(n4700), .A(n4699), .ZN(n4698) );
  INV_X1 U5529 ( .A(n9414), .ZN(n4699) );
  INV_X1 U5530 ( .A(n4502), .ZN(n4700) );
  OR2_X1 U5531 ( .A1(n4701), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5532 ( .A1(n4701), .A2(n4703), .ZN(n4694) );
  AND2_X1 U5533 ( .A1(n6122), .A2(n6121), .ZN(n6329) );
  INV_X1 U5534 ( .A(n6224), .ZN(n4690) );
  NAND2_X1 U5535 ( .A1(n4689), .A2(n6224), .ZN(n4688) );
  INV_X1 U5536 ( .A(n9340), .ZN(n4689) );
  NAND2_X1 U5537 ( .A1(n4500), .A2(n4990), .ZN(n4988) );
  OAI21_X1 U5538 ( .B1(n6129), .B2(n6326), .A(n6131), .ZN(n7240) );
  INV_X1 U5539 ( .A(n4625), .ZN(n5483) );
  INV_X1 U5540 ( .A(n4705), .ZN(n4703) );
  INV_X1 U5541 ( .A(n4702), .ZN(n4701) );
  OAI21_X1 U5542 ( .B1(n9329), .B2(n4703), .A(n6293), .ZN(n4702) );
  NAND2_X1 U5543 ( .A1(n7356), .A2(n6156), .ZN(n7492) );
  OR2_X1 U5544 ( .A1(n6352), .A2(n8357), .ZN(n6350) );
  NAND2_X1 U5545 ( .A1(n8205), .A2(n4585), .ZN(n4810) );
  AND2_X1 U5546 ( .A1(n4812), .A2(n8220), .ZN(n4811) );
  AOI21_X1 U5547 ( .B1(n8200), .B2(n5151), .A(n8199), .ZN(n8205) );
  AND2_X1 U5548 ( .A1(n5726), .A2(n5725), .ZN(n9359) );
  NAND2_X1 U5549 ( .A1(n5325), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5312) );
  AOI22_X1 U5550 ( .A1(n7480), .A2(n7479), .B1(n7484), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n7665) );
  INV_X1 U5551 ( .A(n9972), .ZN(n9654) );
  OR2_X1 U5552 ( .A1(n5753), .A2(n5752), .ZN(n5766) );
  INV_X1 U5553 ( .A(n9661), .ZN(n4859) );
  INV_X1 U5554 ( .A(n9734), .ZN(n5686) );
  AND2_X1 U5555 ( .A1(n9698), .A2(n8273), .ZN(n9717) );
  INV_X1 U5556 ( .A(n8227), .ZN(n5814) );
  NAND2_X1 U5557 ( .A1(n9770), .A2(n8335), .ZN(n8278) );
  NAND2_X1 U5558 ( .A1(n5107), .A2(n8278), .ZN(n9743) );
  OAI21_X1 U5559 ( .B1(n9818), .B2(n4475), .A(n4643), .ZN(n9775) );
  AOI21_X1 U5560 ( .B1(n5577), .B2(n4648), .A(n4506), .ZN(n4647) );
  OR2_X1 U5561 ( .A1(n9808), .A2(n10006), .ZN(n4473) );
  AND2_X1 U5562 ( .A1(n8321), .A2(n8326), .ZN(n9863) );
  AOI21_X1 U5563 ( .B1(n4851), .B2(n4853), .A(n4526), .ZN(n4850) );
  NAND2_X1 U5564 ( .A1(n7718), .A2(n5392), .ZN(n7698) );
  NAND2_X1 U5565 ( .A1(n7698), .A2(n7697), .ZN(n7696) );
  NOR2_X1 U5566 ( .A1(n7508), .A2(n7692), .ZN(n7507) );
  NAND2_X1 U5567 ( .A1(n7372), .A2(n5797), .ZN(n4790) );
  INV_X1 U5568 ( .A(n10067), .ZN(n7548) );
  AND2_X1 U5569 ( .A1(n6338), .A2(n6337), .ZN(n7449) );
  OAI21_X1 U5570 ( .B1(n9668), .B2(n9885), .A(n5840), .ZN(n5841) );
  NOR2_X1 U5571 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U5572 ( .A1(n7751), .A2(n6847), .ZN(n5615) );
  AND2_X1 U5573 ( .A1(n5865), .A2(n5864), .ZN(n6101) );
  OR2_X1 U5574 ( .A1(n7317), .A2(n8223), .ZN(n5865) );
  XNOR2_X1 U5575 ( .A(n4928), .B(n6846), .ZN(n9244) );
  OAI21_X1 U5576 ( .B1(n6844), .B2(n6843), .A(n6842), .ZN(n4928) );
  XNOR2_X1 U5577 ( .A(n6844), .B(n6843), .ZN(n8575) );
  XNOR2_X1 U5578 ( .A(n5846), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5873) );
  XNOR2_X1 U5579 ( .A(n5872), .B(n5871), .ZN(n7852) );
  NAND2_X1 U5580 ( .A1(n4959), .A2(n4960), .ZN(n5650) );
  NOR2_X1 U5581 ( .A1(n5008), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5007) );
  NOR2_X1 U5582 ( .A1(n5260), .A2(n5008), .ZN(n5519) );
  XNOR2_X1 U5583 ( .A(n4601), .B(n4600), .ZN(n6888) );
  INV_X1 U5584 ( .A(n5374), .ZN(n4600) );
  AND2_X1 U5585 ( .A1(n5244), .A2(n5229), .ZN(n6948) );
  XNOR2_X1 U5586 ( .A(n5217), .B(n5240), .ZN(n6870) );
  AND2_X1 U5587 ( .A1(n4935), .A2(n4452), .ZN(n5217) );
  INV_X1 U5588 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5187) );
  NOR2_X1 U5589 ( .A1(n8460), .A2(n5021), .ZN(n5020) );
  INV_X1 U5590 ( .A(n8396), .ZN(n5021) );
  AOI21_X1 U5591 ( .B1(n5042), .B2(n4480), .A(n8555), .ZN(n5038) );
  NAND2_X1 U5592 ( .A1(n5042), .A2(n5047), .ZN(n5041) );
  NAND2_X1 U5593 ( .A1(n8427), .A2(n8446), .ZN(n5047) );
  AOI21_X1 U5594 ( .B1(n5031), .B2(n8522), .A(n5029), .ZN(n5028) );
  INV_X1 U5595 ( .A(n5031), .ZN(n5030) );
  INV_X1 U5596 ( .A(n8416), .ZN(n5029) );
  AOI21_X1 U5597 ( .B1(n5023), .B2(n5025), .A(n4511), .ZN(n5022) );
  NAND2_X1 U5598 ( .A1(n8560), .A2(n5023), .ZN(n4677) );
  AND2_X1 U5599 ( .A1(n6636), .A2(n6635), .ZN(n8984) );
  XNOR2_X1 U5600 ( .A(n4818), .B(n8612), .ZN(n8614) );
  OAI211_X1 U5601 ( .C1(n6680), .C2(n9224), .A(n6579), .B(n6578), .ZN(n9092)
         );
  OR2_X1 U5602 ( .A1(n7928), .A2(n6436), .ZN(n6441) );
  OR2_X1 U5603 ( .A1(n6680), .A2(n6438), .ZN(n6439) );
  NAND2_X1 U5604 ( .A1(n6059), .A2(n6058), .ZN(n7589) );
  AND2_X1 U5605 ( .A1(n4911), .A2(n4910), .ZN(n7595) );
  XNOR2_X1 U5606 ( .A(n4772), .B(n4771), .ZN(n8812) );
  NAND2_X1 U5607 ( .A1(n8843), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4783) );
  OAI21_X1 U5608 ( .B1(n6070), .B2(n4737), .A(n4735), .ZN(n8859) );
  INV_X1 U5609 ( .A(n10088), .ZN(n8922) );
  INV_X1 U5610 ( .A(n6094), .ZN(n4776) );
  XNOR2_X1 U5611 ( .A(n4745), .B(n4744), .ZN(n4743) );
  INV_X1 U5612 ( .A(n6096), .ZN(n4744) );
  AOI21_X1 U5613 ( .B1(n8925), .B2(n8932), .A(n8927), .ZN(n4745) );
  NAND2_X1 U5614 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  INV_X1 U5615 ( .A(n6097), .ZN(n4742) );
  NAND2_X1 U5616 ( .A1(n10099), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4741) );
  OAI21_X1 U5617 ( .B1(n8948), .B2(n10124), .A(n4529), .ZN(n8950) );
  NAND2_X1 U5618 ( .A1(n6783), .A2(n6782), .ZN(n8954) );
  NOR2_X1 U5619 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  INV_X1 U5620 ( .A(n10115), .ZN(n8992) );
  INV_X1 U5621 ( .A(n10141), .ZN(n10144) );
  NAND2_X1 U5622 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U5623 ( .A1(n8776), .A2(n9090), .ZN(n6699) );
  INV_X1 U5624 ( .A(n8733), .ZN(n8953) );
  OR2_X1 U5625 ( .A1(n7005), .A2(n6791), .ZN(n6797) );
  AND2_X1 U5626 ( .A1(n7307), .A2(n6991), .ZN(n6791) );
  NAND2_X1 U5627 ( .A1(n6713), .A2(n6712), .ZN(n6884) );
  NAND2_X1 U5628 ( .A1(n4974), .A2(n4972), .ZN(n9327) );
  AOI21_X1 U5629 ( .B1(n4471), .B2(n4483), .A(n4973), .ZN(n4972) );
  INV_X1 U5630 ( .A(n9395), .ZN(n4973) );
  NAND2_X1 U5631 ( .A1(n9327), .A2(n9329), .ZN(n9328) );
  AND2_X1 U5632 ( .A1(n5701), .A2(n5719), .ZN(n9722) );
  NAND2_X1 U5633 ( .A1(n7258), .A2(n7259), .ZN(n5003) );
  NAND2_X1 U5634 ( .A1(n4681), .A2(n6316), .ZN(n4680) );
  NOR2_X2 U5635 ( .A1(n6350), .A2(n6339), .ZN(n9434) );
  OR2_X1 U5636 ( .A1(n9964), .A2(n8292), .ZN(n6339) );
  INV_X1 U5637 ( .A(n7798), .ZN(n8358) );
  OR2_X1 U5638 ( .A1(n9298), .A2(n5721), .ZN(n5669) );
  AND3_X1 U5639 ( .A1(n5237), .A2(n5239), .A3(n5236), .ZN(n4761) );
  INV_X1 U5640 ( .A(n7510), .ZN(n9495) );
  NAND2_X1 U5641 ( .A1(n5349), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5297) );
  OAI21_X1 U5642 ( .B1(n9551), .B2(n9560), .A(n6931), .ZN(n9584) );
  NAND2_X1 U5643 ( .A1(n4604), .A2(n5830), .ZN(n9659) );
  AND2_X1 U5644 ( .A1(n9662), .A2(n6106), .ZN(n9673) );
  NAND2_X1 U5645 ( .A1(n4861), .A2(n5741), .ZN(n6105) );
  NAND2_X1 U5646 ( .A1(n9901), .A2(n10071), .ZN(n4657) );
  INV_X1 U5647 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4808) );
  XNOR2_X1 U5648 ( .A(n5869), .B(n5868), .ZN(n7798) );
  INV_X1 U5649 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U5650 ( .A1(n5587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U5651 ( .A1(n8659), .A2(n8658), .ZN(n4578) );
  INV_X1 U5652 ( .A(n8667), .ZN(n4577) );
  NAND2_X1 U5653 ( .A1(n8659), .A2(n8656), .ZN(n4886) );
  AND2_X1 U5654 ( .A1(n8127), .A2(n4803), .ZN(n4589) );
  AND2_X1 U5655 ( .A1(n8131), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5656 ( .A1(n8125), .A2(n8130), .ZN(n4806) );
  AOI21_X1 U5657 ( .B1(n4897), .B2(n4894), .A(n8683), .ZN(n4893) );
  INV_X1 U5658 ( .A(n4895), .ZN(n4894) );
  NAND2_X1 U5659 ( .A1(n5068), .A2(n8682), .ZN(n4892) );
  NOR2_X1 U5660 ( .A1(n8591), .A2(n8590), .ZN(n8670) );
  NAND2_X1 U5661 ( .A1(n8715), .A2(n6697), .ZN(n4575) );
  AND2_X1 U5662 ( .A1(n4713), .A2(n4889), .ZN(n4712) );
  INV_X1 U5663 ( .A(n4869), .ZN(n4868) );
  INV_X1 U5664 ( .A(n8709), .ZN(n4722) );
  INV_X1 U5665 ( .A(n8725), .ZN(n4877) );
  NAND2_X1 U5666 ( .A1(n4531), .A2(n8726), .ZN(n4878) );
  AOI21_X1 U5667 ( .B1(n8162), .B2(n4495), .A(n9838), .ZN(n8174) );
  NOR2_X1 U5668 ( .A1(n4794), .A2(n4789), .ZN(n4788) );
  INV_X1 U5669 ( .A(n8304), .ZN(n4789) );
  INV_X1 U5670 ( .A(n8305), .ZN(n4794) );
  INV_X1 U5671 ( .A(n5798), .ZN(n4792) );
  INV_X1 U5672 ( .A(n8423), .ZN(n5050) );
  INV_X1 U5673 ( .A(n7864), .ZN(n5014) );
  NAND2_X1 U5674 ( .A1(n4876), .A2(n4874), .ZN(n4873) );
  NAND2_X1 U5675 ( .A1(n8739), .A2(n8736), .ZN(n4718) );
  INV_X1 U5676 ( .A(n7013), .ZN(n6793) );
  AND2_X1 U5677 ( .A1(n8244), .A2(n4627), .ZN(n8248) );
  NOR2_X1 U5678 ( .A1(n4628), .A2(n8246), .ZN(n4627) );
  NAND2_X1 U5679 ( .A1(n5814), .A2(n4510), .ZN(n4631) );
  INV_X1 U5680 ( .A(n9776), .ZN(n4632) );
  NAND2_X1 U5681 ( .A1(n8275), .A2(n8297), .ZN(n4587) );
  INV_X1 U5682 ( .A(n4648), .ZN(n4644) );
  INV_X1 U5683 ( .A(n5609), .ZN(n4641) );
  INV_X1 U5684 ( .A(n4647), .ZN(n4645) );
  NOR2_X1 U5685 ( .A1(n6835), .A2(n4927), .ZN(n4926) );
  INV_X1 U5686 ( .A(n4948), .ZN(n4947) );
  OAI21_X1 U5687 ( .B1(n5688), .B2(n4949), .A(n5708), .ZN(n4948) );
  INV_X1 U5688 ( .A(n5690), .ZN(n4949) );
  INV_X1 U5689 ( .A(n5512), .ZN(n4939) );
  AND2_X1 U5690 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  INV_X1 U5691 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5534) );
  INV_X1 U5692 ( .A(n5532), .ZN(n5533) );
  INV_X1 U5693 ( .A(n4710), .ZN(n4709) );
  OAI21_X1 U5694 ( .B1(n4952), .B2(n4953), .A(n4711), .ZN(n4710) );
  NAND2_X1 U5695 ( .A1(n5881), .A2(n4609), .ZN(n5913) );
  AND2_X1 U5696 ( .A1(n5100), .A2(n5955), .ZN(n4609) );
  NAND2_X1 U5697 ( .A1(n7092), .A2(n10126), .ZN(n7088) );
  OR2_X1 U5698 ( .A1(n7561), .A2(n5014), .ZN(n5013) );
  INV_X1 U5699 ( .A(n7111), .ZN(n7868) );
  INV_X1 U5700 ( .A(n5035), .ZN(n5034) );
  OAI21_X1 U5701 ( .B1(n8400), .B2(n5036), .A(n8471), .ZN(n5035) );
  OR2_X1 U5702 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U5703 ( .A1(n9161), .A2(n8577), .ZN(n4610) );
  OR2_X1 U5704 ( .A1(n6412), .A2(n10472), .ZN(n6395) );
  NAND2_X1 U5705 ( .A1(n4726), .A2(n8819), .ZN(n4725) );
  NAND2_X1 U5706 ( .A1(n4727), .A2(n4729), .ZN(n4726) );
  NAND2_X1 U5707 ( .A1(n7587), .A2(n4768), .ZN(n4767) );
  AOI21_X1 U5708 ( .B1(n4735), .B2(n4737), .A(n4734), .ZN(n4733) );
  INV_X1 U5709 ( .A(n8858), .ZN(n4734) );
  NAND2_X1 U5710 ( .A1(n4565), .A2(n6574), .ZN(n4564) );
  INV_X1 U5711 ( .A(n5993), .ZN(n4565) );
  AOI21_X1 U5712 ( .B1(n5094), .B2(n8731), .A(n4538), .ZN(n5093) );
  OR2_X1 U5713 ( .A1(n6675), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U5714 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  INV_X1 U5715 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n4828) );
  INV_X1 U5716 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n4827) );
  AND2_X1 U5717 ( .A1(n6375), .A2(n4832), .ZN(n4831) );
  INV_X1 U5718 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4832) );
  INV_X1 U5719 ( .A(n4496), .ZN(n6376) );
  NOR2_X1 U5720 ( .A1(n6548), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4829) );
  NOR2_X1 U5721 ( .A1(n6517), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4833) );
  INV_X1 U5722 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10263) );
  INV_X1 U5723 ( .A(n7383), .ZN(n4568) );
  OR2_X1 U5724 ( .A1(n6714), .A2(n6726), .ZN(n6792) );
  NOR2_X1 U5725 ( .A1(n9169), .A2(n8742), .ZN(n4591) );
  OR2_X1 U5726 ( .A1(n8451), .A2(n8966), .ZN(n8734) );
  AND2_X1 U5727 ( .A1(n8717), .A2(n8988), .ZN(n8996) );
  OR2_X1 U5728 ( .A1(n9060), .A2(n8542), .ZN(n9021) );
  NAND2_X1 U5729 ( .A1(n5068), .A2(n6565), .ZN(n5067) );
  NOR2_X1 U5730 ( .A1(n5069), .A2(n5064), .ZN(n5063) );
  INV_X1 U5731 ( .A(n6554), .ZN(n5064) );
  INV_X1 U5732 ( .A(n6565), .ZN(n5069) );
  NOR2_X1 U5733 ( .A1(n8684), .A2(n4999), .ZN(n4998) );
  INV_X1 U5734 ( .A(n8681), .ZN(n4999) );
  INV_X1 U5735 ( .A(n8662), .ZN(n4992) );
  INV_X1 U5736 ( .A(n4597), .ZN(n5141) );
  OR2_X1 U5737 ( .A1(n5967), .A2(n5920), .ZN(n5975) );
  NAND2_X1 U5738 ( .A1(n5937), .A2(n4865), .ZN(n4674) );
  INV_X1 U5739 ( .A(n6232), .ZN(n4990) );
  NOR2_X1 U5740 ( .A1(n5542), .A2(n5541), .ZN(n4623) );
  NAND2_X1 U5741 ( .A1(n6118), .A2(n6122), .ZN(n5012) );
  NAND2_X1 U5742 ( .A1(n8202), .A2(n9698), .ZN(n8200) );
  INV_X1 U5743 ( .A(n8198), .ZN(n8199) );
  AOI21_X1 U5744 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8198) );
  NAND2_X1 U5745 ( .A1(n4813), .A2(n8210), .ZN(n4812) );
  INV_X1 U5746 ( .A(n4814), .ZN(n4813) );
  AOI21_X1 U5747 ( .B1(n4503), .B2(n9663), .A(n4484), .ZN(n4814) );
  OR2_X1 U5748 ( .A1(n6359), .A2(n9266), .ZN(n8280) );
  NAND2_X1 U5749 ( .A1(n4842), .A2(n4840), .ZN(n4839) );
  INV_X1 U5750 ( .A(n5150), .ZN(n4840) );
  OR2_X1 U5751 ( .A1(n9706), .A2(n9359), .ZN(n8261) );
  NAND2_X1 U5752 ( .A1(n5130), .A2(n9979), .ZN(n5128) );
  NOR2_X1 U5753 ( .A1(n9357), .A2(n9736), .ZN(n5130) );
  OR2_X1 U5754 ( .A1(n9736), .A2(n9358), .ZN(n8263) );
  NAND2_X1 U5755 ( .A1(n9752), .A2(n5815), .ZN(n8168) );
  OR2_X1 U5756 ( .A1(n9781), .A2(n5122), .ZN(n5121) );
  NAND2_X1 U5757 ( .A1(n9995), .A2(n10003), .ZN(n5122) );
  NAND2_X1 U5758 ( .A1(n4624), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5663) );
  INV_X1 U5759 ( .A(n4624), .ZN(n5642) );
  NAND2_X1 U5760 ( .A1(n5523), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5542) );
  INV_X1 U5761 ( .A(n5525), .ZN(n5523) );
  INV_X1 U5762 ( .A(n4852), .ZN(n4851) );
  OAI21_X1 U5763 ( .B1(n5466), .B2(n4853), .A(n5489), .ZN(n4852) );
  INV_X1 U5764 ( .A(n5467), .ZN(n4853) );
  AND2_X1 U5765 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .ZN(n5480) );
  INV_X1 U5766 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5382) );
  XNOR2_X1 U5767 ( .A(n9493), .B(n4466), .ZN(n7610) );
  NAND2_X1 U5768 ( .A1(n9496), .A2(n10067), .ZN(n8304) );
  NAND2_X1 U5769 ( .A1(n5833), .A2(n5126), .ZN(n9865) );
  NAND2_X1 U5770 ( .A1(n7706), .A2(n5136), .ZN(n8081) );
  AND2_X1 U5771 ( .A1(n8121), .A2(n8122), .ZN(n7740) );
  INV_X1 U5772 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5988) );
  INV_X1 U5773 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10464) );
  INV_X1 U5774 ( .A(SI_17_), .ZN(n10421) );
  INV_X1 U5775 ( .A(SI_11_), .ZN(n10356) );
  AOI21_X1 U5776 ( .B1(n4962), .B2(n5599), .A(n4961), .ZN(n4960) );
  INV_X1 U5777 ( .A(n5634), .ZN(n4961) );
  INV_X1 U5778 ( .A(SI_20_), .ZN(n10268) );
  NAND2_X1 U5779 ( .A1(n5584), .A2(n10487), .ZN(n5598) );
  INV_X1 U5780 ( .A(n5578), .ZN(n5582) );
  NAND2_X1 U5781 ( .A1(n4937), .A2(n5512), .ZN(n5551) );
  NAND2_X1 U5782 ( .A1(n5413), .A2(n10356), .ZN(n5432) );
  AND2_X1 U5783 ( .A1(n4936), .A2(n5373), .ZN(n4930) );
  NAND2_X1 U5784 ( .A1(n5358), .A2(n5357), .ZN(n4936) );
  NAND2_X1 U5785 ( .A1(n4934), .A2(n5359), .ZN(n4931) );
  OR2_X1 U5786 ( .A1(n4464), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5190) );
  INV_X1 U5787 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5186) );
  XNOR2_X1 U5788 ( .A(n7084), .B(n7111), .ZN(n7108) );
  INV_X1 U5789 ( .A(n5048), .ZN(n5045) );
  NAND2_X1 U5790 ( .A1(n6369), .A2(n6368), .ZN(n6491) );
  AND2_X1 U5791 ( .A1(n8486), .A2(n5024), .ZN(n5023) );
  OR2_X1 U5792 ( .A1(n8559), .A2(n5025), .ZN(n5024) );
  INV_X1 U5793 ( .A(n8387), .ZN(n5025) );
  INV_X1 U5794 ( .A(n8413), .ZN(n8502) );
  NAND2_X1 U5795 ( .A1(n5037), .A2(n8400), .ZN(n8513) );
  INV_X1 U5796 ( .A(n8515), .ZN(n5037) );
  NOR2_X1 U5797 ( .A1(n8059), .A2(n5027), .ZN(n5026) );
  INV_X1 U5798 ( .A(n8055), .ZN(n5027) );
  INV_X1 U5799 ( .A(n4833), .ZN(n6528) );
  INV_X1 U5800 ( .A(n8790), .ZN(n7146) );
  AND2_X1 U5801 ( .A1(n8381), .A2(n9103), .ZN(n8382) );
  AND2_X1 U5802 ( .A1(n4819), .A2(n4636), .ZN(n4818) );
  NOR2_X1 U5803 ( .A1(n8611), .A2(n4637), .ZN(n4636) );
  NOR2_X1 U5804 ( .A1(n4820), .A2(n8754), .ZN(n4819) );
  AND2_X1 U5805 ( .A1(n7933), .A2(n7932), .ZN(n8941) );
  OR2_X1 U5806 ( .A1(n6424), .A2(n7311), .ZN(n6406) );
  NAND2_X1 U5807 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n6411), .ZN(n4603) );
  NAND2_X1 U5808 ( .A1(n4570), .A2(n4569), .ZN(n6032) );
  NAND2_X1 U5809 ( .A1(n6695), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5810 ( .A1(n7190), .A2(n7191), .ZN(n7189) );
  NAND2_X1 U5811 ( .A1(n4739), .A2(n4738), .ZN(n7063) );
  INV_X1 U5812 ( .A(n7066), .ZN(n4738) );
  NAND2_X1 U5813 ( .A1(n8804), .A2(n6013), .ZN(n6014) );
  NAND2_X1 U5814 ( .A1(n4731), .A2(n4730), .ZN(n10097) );
  INV_X1 U5815 ( .A(n10093), .ZN(n4730) );
  NAND2_X1 U5816 ( .A1(n4912), .A2(n5963), .ZN(n7523) );
  AND2_X1 U5817 ( .A1(n5979), .A2(n8862), .ZN(n8844) );
  NAND2_X1 U5818 ( .A1(n8844), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8863) );
  INV_X1 U5819 ( .A(n8846), .ZN(n4737) );
  NAND2_X1 U5820 ( .A1(n5982), .A2(n8876), .ZN(n5983) );
  NAND2_X1 U5821 ( .A1(n4785), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5822 ( .A1(n4778), .A2(n4777), .ZN(n4781) );
  NAND2_X1 U5823 ( .A1(n8879), .A2(n5983), .ZN(n8889) );
  NOR2_X1 U5824 ( .A1(n8927), .A2(n8926), .ZN(n8931) );
  NOR2_X1 U5825 ( .A1(n8742), .A2(n10127), .ZN(n6781) );
  NAND2_X1 U5826 ( .A1(n6376), .A2(n6375), .ZN(n6584) );
  NAND2_X1 U5827 ( .A1(n4829), .A2(n6374), .ZN(n6568) );
  INV_X1 U5828 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6374) );
  INV_X1 U5829 ( .A(n4829), .ZN(n6558) );
  NAND2_X1 U5830 ( .A1(n4833), .A2(n6371), .ZN(n6538) );
  INV_X1 U5831 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U5832 ( .A1(n6373), .A2(n6372), .ZN(n6548) );
  INV_X1 U5833 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6372) );
  INV_X1 U5834 ( .A(n6538), .ZN(n6373) );
  AND2_X1 U5835 ( .A1(n4512), .A2(n6370), .ZN(n4834) );
  INV_X1 U5836 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6370) );
  INV_X1 U5837 ( .A(n6469), .ZN(n6369) );
  AOI21_X1 U5838 ( .B1(n5089), .B2(n5087), .A(n4508), .ZN(n5086) );
  NAND2_X1 U5839 ( .A1(n6367), .A2(n6366), .ZN(n6457) );
  INV_X1 U5840 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6366) );
  INV_X1 U5841 ( .A(n6446), .ZN(n6367) );
  OR2_X1 U5842 ( .A1(n6457), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U5843 ( .A1(n10225), .A2(n10263), .ZN(n6446) );
  INV_X1 U5844 ( .A(n8792), .ZN(n7406) );
  INV_X1 U5845 ( .A(n8610), .ZN(n4616) );
  AND2_X1 U5846 ( .A1(n6697), .A2(n6729), .ZN(n6762) );
  NOR2_X1 U5847 ( .A1(n8941), .A2(n8940), .ZN(n9159) );
  INV_X1 U5848 ( .A(n6698), .ZN(n10127) );
  INV_X1 U5849 ( .A(n6751), .ZN(n9012) );
  AND2_X1 U5850 ( .A1(n5096), .A2(n5097), .ZN(n9010) );
  CLKBUF_X1 U5851 ( .A(n9020), .Z(n9050) );
  CLKBUF_X1 U5852 ( .A(n9026), .Z(n9066) );
  NAND2_X1 U5853 ( .A1(n8695), .A2(n8694), .ZN(n9065) );
  INV_X1 U5854 ( .A(n5075), .ZN(n5074) );
  INV_X1 U5855 ( .A(n10151), .ZN(n10174) );
  INV_X1 U5856 ( .A(n10172), .ZN(n10161) );
  OR2_X1 U5857 ( .A1(n6790), .A2(n6789), .ZN(n6991) );
  INV_X1 U5858 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6381) );
  INV_X1 U5859 ( .A(n5916), .ZN(n5959) );
  OR2_X1 U5860 ( .A1(n5925), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U5861 ( .A1(n7568), .A2(n7569), .ZN(n7943) );
  AOI21_X1 U5862 ( .B1(n4971), .B2(n6191), .A(n4969), .ZN(n4968) );
  INV_X2 U5863 ( .A(n6317), .ZN(n6331) );
  NAND2_X1 U5864 ( .A1(n4566), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5346) );
  INV_X1 U5865 ( .A(n5234), .ZN(n4566) );
  INV_X1 U5866 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5345) );
  OR2_X1 U5867 ( .A1(n5346), .A2(n5345), .ZN(n5383) );
  NAND2_X1 U5868 ( .A1(n6223), .A2(n9340), .ZN(n9343) );
  INV_X1 U5869 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7133) );
  INV_X1 U5870 ( .A(n9476), .ZN(n9358) );
  NAND2_X1 U5871 ( .A1(n5661), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5700) );
  INV_X1 U5872 ( .A(n5663), .ZN(n5661) );
  OR2_X1 U5873 ( .A1(n5604), .A2(n9397), .ZN(n5616) );
  NAND2_X1 U5874 ( .A1(n5592), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5604) );
  INV_X1 U5875 ( .A(n5593), .ZN(n5592) );
  INV_X1 U5876 ( .A(n4978), .ZN(n4977) );
  AND2_X1 U5877 ( .A1(n6280), .A2(n9306), .ZN(n6281) );
  NAND2_X1 U5878 ( .A1(n4978), .A2(n4976), .ZN(n4975) );
  OR2_X1 U5879 ( .A1(n6275), .A2(n6274), .ZN(n6280) );
  NAND2_X1 U5880 ( .A1(n9343), .A2(n6224), .ZN(n9403) );
  NAND2_X1 U5881 ( .A1(n9403), .A2(n9404), .ZN(n9402) );
  AND2_X1 U5882 ( .A1(n5824), .A2(n8292), .ZN(n9426) );
  NAND2_X1 U5883 ( .A1(n5424), .A2(n5423), .ZN(n5447) );
  AND2_X1 U5884 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5423) );
  INV_X1 U5885 ( .A(n5422), .ZN(n5424) );
  OR2_X1 U5886 ( .A1(n5383), .A2(n5382), .ZN(n5422) );
  INV_X1 U5887 ( .A(n4623), .ZN(n5571) );
  NAND2_X1 U5888 ( .A1(n4623), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5593) );
  INV_X1 U5889 ( .A(n9493), .ZN(n7511) );
  NAND2_X1 U5890 ( .A1(n4682), .A2(n6303), .ZN(n4681) );
  NOR2_X1 U5891 ( .A1(n4633), .A2(n8257), .ZN(n5147) );
  INV_X1 U5892 ( .A(n9457), .ZN(n9369) );
  AOI21_X1 U5893 ( .B1(n9691), .B2(n5767), .A(n5740), .ZN(n9438) );
  AND4_X1 U5894 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n8013)
         );
  AND4_X1 U5895 ( .A1(n5405), .A2(n5404), .A3(n5403), .A4(n5402), .ZN(n7728)
         );
  AND4_X1 U5896 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), .ZN(n7741)
         );
  AND2_X1 U5897 ( .A1(n5351), .A2(n4540), .ZN(n5372) );
  AND4_X1 U5898 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n5232)
         );
  AND4_X1 U5899 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n7510)
         );
  AND4_X1 U5900 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n7260)
         );
  AND4_X1 U5901 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n7250)
         );
  NAND2_X1 U5902 ( .A1(n6924), .A2(n6923), .ZN(n9523) );
  AOI22_X1 U5903 ( .A1(n6977), .A2(n6976), .B1(n6975), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n6978) );
  OR2_X1 U5904 ( .A1(n7042), .A2(n7043), .ZN(n7040) );
  OR2_X1 U5905 ( .A1(n7126), .A2(n7127), .ZN(n7224) );
  AOI22_X1 U5906 ( .A1(n7130), .A2(n7129), .B1(n7128), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7131) );
  OR2_X1 U5907 ( .A1(n7227), .A2(n7226), .ZN(n7343) );
  AND2_X1 U5908 ( .A1(n9514), .A2(n8292), .ZN(n9457) );
  AND2_X1 U5909 ( .A1(n5754), .A2(n5766), .ZN(n9675) );
  NOR2_X1 U5910 ( .A1(n8259), .A2(n5109), .ZN(n5108) );
  INV_X1 U5911 ( .A(n8272), .ZN(n5109) );
  INV_X1 U5912 ( .A(n4842), .ZN(n4841) );
  NOR2_X1 U5913 ( .A1(n9735), .A2(n5129), .ZN(n9720) );
  INV_X1 U5914 ( .A(n5130), .ZN(n5129) );
  NAND2_X1 U5915 ( .A1(n4758), .A2(n4757), .ZN(n4753) );
  NOR2_X1 U5916 ( .A1(n9735), .A2(n9736), .ZN(n9719) );
  AOI21_X1 U5917 ( .B1(n4478), .B2(n4856), .A(n4528), .ZN(n4855) );
  NOR3_X1 U5918 ( .A1(n4473), .A2(n9781), .A3(n9791), .ZN(n9778) );
  NOR2_X1 U5919 ( .A1(n4473), .A2(n9791), .ZN(n9777) );
  NOR2_X1 U5920 ( .A1(n9943), .A2(n5124), .ZN(n5123) );
  INV_X1 U5921 ( .A(n5125), .ZN(n5124) );
  NAND2_X1 U5922 ( .A1(n9860), .A2(n5531), .ZN(n9837) );
  NOR2_X1 U5923 ( .A1(n5134), .A2(n9963), .ZN(n5132) );
  AND2_X1 U5924 ( .A1(n7706), .A2(n5133), .ZN(n8080) );
  AND2_X1 U5925 ( .A1(n8249), .A2(n8145), .ZN(n5102) );
  NAND2_X1 U5926 ( .A1(n8079), .A2(n5466), .ZN(n8078) );
  NAND2_X1 U5927 ( .A1(n7699), .A2(n8314), .ZN(n4764) );
  AND2_X1 U5928 ( .A1(n4846), .A2(n5431), .ZN(n4845) );
  NAND2_X1 U5929 ( .A1(n4477), .A2(n7958), .ZN(n5114) );
  AOI21_X1 U5930 ( .B1(n4799), .B2(n4801), .A(n4797), .ZN(n4796) );
  INV_X1 U5931 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U5932 ( .A1(n8304), .A2(n5795), .ZN(n8229) );
  OR2_X1 U5933 ( .A1(n7444), .A2(n5787), .ZN(n7817) );
  NAND2_X1 U5934 ( .A1(n6124), .A2(n4588), .ZN(n7246) );
  INV_X1 U5935 ( .A(n9878), .ZN(n9858) );
  AND2_X1 U5936 ( .A1(n8260), .A2(n8223), .ZN(n7457) );
  AND2_X1 U5937 ( .A1(n8290), .A2(n6856), .ZN(n9895) );
  AND2_X1 U5938 ( .A1(n8356), .A2(n6345), .ZN(n9964) );
  AND2_X1 U5939 ( .A1(n7852), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6864) );
  XNOR2_X1 U5940 ( .A(n5735), .B(n5734), .ZN(n8445) );
  NAND4_X1 U5941 ( .A1(n5112), .A2(n5113), .A3(n5166), .A4(n4453), .ZN(n5221)
         );
  INV_X1 U5942 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U5943 ( .A1(n5845), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U5944 ( .A1(n4946), .A2(n5690), .ZN(n5709) );
  NAND2_X1 U5945 ( .A1(n5562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5564) );
  INV_X1 U5946 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5563) );
  XNOR2_X1 U5947 ( .A(n4714), .B(n5554), .ZN(n7292) );
  OAI21_X1 U5948 ( .B1(n5551), .B2(n5553), .A(n5555), .ZN(n4714) );
  NAND2_X1 U5949 ( .A1(n5519), .A2(n5784), .ZN(n5538) );
  AND2_X1 U5950 ( .A1(n5497), .A2(n5477), .ZN(n7484) );
  NAND2_X1 U5951 ( .A1(n4950), .A2(n4951), .ZN(n5469) );
  NAND2_X1 U5952 ( .A1(n5434), .A2(n4953), .ZN(n4950) );
  OR2_X1 U5953 ( .A1(n5438), .A2(n5437), .ZN(n5440) );
  NAND2_X1 U5954 ( .A1(n4935), .A2(n4933), .ZN(n5360) );
  INV_X1 U5955 ( .A(n4934), .ZN(n4933) );
  INV_X1 U5956 ( .A(n5258), .ZN(n5226) );
  XNOR2_X1 U5957 ( .A(n5205), .B(SI_3_), .ZN(n5335) );
  OAI21_X1 U5958 ( .B1(n4464), .B2(n4622), .A(n4621), .ZN(n5288) );
  NAND2_X1 U5959 ( .A1(n5748), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4621) );
  XNOR2_X1 U5960 ( .A(n8454), .B(n8502), .ZN(n8503) );
  INV_X1 U5961 ( .A(n5019), .ZN(n7110) );
  NAND2_X1 U5962 ( .A1(n8536), .A2(n8396), .ZN(n8461) );
  OR2_X1 U5963 ( .A1(n6816), .A2(n6393), .ZN(n5059) );
  NAND2_X1 U5964 ( .A1(n8513), .A2(n8403), .ZN(n8470) );
  NAND2_X1 U5965 ( .A1(n4659), .A2(n7874), .ZN(n7877) );
  AND2_X1 U5966 ( .A1(n6389), .A2(n6388), .ZN(n9001) );
  NAND2_X1 U5967 ( .A1(n8558), .A2(n8387), .ZN(n8487) );
  OAI21_X1 U5968 ( .B1(n4599), .B2(n5025), .A(n5023), .ZN(n8485) );
  NAND2_X1 U5969 ( .A1(n7148), .A2(n7147), .ZN(n4670) );
  NAND2_X1 U5970 ( .A1(n6392), .A2(n6391), .ZN(n8510) );
  NAND2_X1 U5971 ( .A1(n7558), .A2(n7557), .ZN(n4667) );
  NAND2_X1 U5972 ( .A1(n7560), .A2(n7561), .ZN(n7865) );
  AOI21_X1 U5973 ( .B1(n9035), .B2(n6688), .A(n6617), .ZN(n8527) );
  INV_X1 U5974 ( .A(n8561), .ZN(n8541) );
  NAND2_X1 U5975 ( .A1(n8056), .A2(n8055), .ZN(n8058) );
  INV_X1 U5976 ( .A(n8409), .ZN(n8523) );
  INV_X1 U5977 ( .A(n8553), .ZN(n8568) );
  NAND2_X1 U5978 ( .A1(n4599), .A2(n8559), .ZN(n8558) );
  NAND2_X1 U5979 ( .A1(n7000), .A2(n6999), .ZN(n8565) );
  OR2_X1 U5980 ( .A1(n8761), .A2(n4885), .ZN(n4883) );
  NAND2_X1 U5981 ( .A1(n6671), .A2(n6670), .ZN(n8776) );
  INV_X1 U5982 ( .A(n9001), .ZN(n8779) );
  INV_X1 U5983 ( .A(n8984), .ZN(n9014) );
  NAND2_X1 U5984 ( .A1(n6626), .A2(n6625), .ZN(n9032) );
  NAND2_X1 U5985 ( .A1(n6598), .A2(n6597), .ZN(n9054) );
  NAND2_X1 U5986 ( .A1(n6609), .A2(n6608), .ZN(n9067) );
  NAND2_X1 U5987 ( .A1(n6590), .A2(n6589), .ZN(n9082) );
  OAI211_X1 U5988 ( .C1(n7928), .C2(n9144), .A(n6571), .B(n6570), .ZN(n9081)
         );
  OR2_X1 U5989 ( .A1(n6424), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6428) );
  XNOR2_X1 U5990 ( .A(n6032), .B(n6393), .ZN(n7180) );
  AND2_X1 U5991 ( .A1(n5941), .A2(n4902), .ZN(n7067) );
  NAND2_X1 U5992 ( .A1(n8794), .A2(n6043), .ZN(n7213) );
  XNOR2_X1 U5993 ( .A(n6014), .B(n7205), .ZN(n7202) );
  NAND2_X1 U5994 ( .A1(n4906), .A2(n4903), .ZN(n10081) );
  NAND2_X1 U5995 ( .A1(n7157), .A2(n6051), .ZN(n7276) );
  OAI21_X1 U5996 ( .B1(n6059), .B2(n4729), .A(n4727), .ZN(n8820) );
  OAI21_X1 U5997 ( .B1(n8812), .B2(n10316), .A(n4770), .ZN(n8825) );
  NAND2_X1 U5998 ( .A1(n6070), .A2(n6069), .ZN(n8845) );
  AND2_X1 U5999 ( .A1(n6031), .A2(n6030), .ZN(n8928) );
  NAND2_X1 U6000 ( .A1(n6665), .A2(n6653), .ZN(n8969) );
  NAND2_X1 U6001 ( .A1(n5000), .A2(n8681), .ZN(n9099) );
  NAND2_X1 U6002 ( .A1(n4996), .A2(n8645), .ZN(n7800) );
  OR2_X1 U6003 ( .A1(n7424), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U6004 ( .A1(n5090), .A2(n6445), .ZN(n7413) );
  INV_X1 U6005 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10225) );
  INV_X1 U6006 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10472) );
  INV_X1 U6007 ( .A(n10111), .ZN(n9109) );
  NAND2_X1 U6008 ( .A1(n10141), .A2(n6770), .ZN(n10115) );
  NAND2_X1 U6009 ( .A1(n8571), .A2(n8570), .ZN(n9112) );
  AOI21_X1 U6010 ( .B1(n8575), .B2(n6486), .A(n8574), .ZN(n9164) );
  AND2_X1 U6011 ( .A1(n8959), .A2(n10162), .ZN(n4571) );
  INV_X1 U6012 ( .A(n8970), .ZN(n6657) );
  NAND2_X1 U6013 ( .A1(n4983), .A2(n8722), .ZN(n8962) );
  NAND2_X1 U6014 ( .A1(n4979), .A2(n4984), .ZN(n4983) );
  NAND2_X1 U6015 ( .A1(n4979), .A2(n4479), .ZN(n8978) );
  NAND2_X1 U6016 ( .A1(n4614), .A2(n8717), .ZN(n8989) );
  NAND2_X1 U6017 ( .A1(n6630), .A2(n6629), .ZN(n9190) );
  NAND2_X1 U6018 ( .A1(n6619), .A2(n6618), .ZN(n9196) );
  NAND2_X1 U6019 ( .A1(n6583), .A2(n6582), .ZN(n9219) );
  NAND2_X1 U6020 ( .A1(n9100), .A2(n9101), .ZN(n5065) );
  NAND2_X1 U6021 ( .A1(n6743), .A2(n8676), .ZN(n8006) );
  NAND2_X1 U6022 ( .A1(n7580), .A2(n8620), .ZN(n7828) );
  NAND2_X1 U6023 ( .A1(n5077), .A2(n5081), .ZN(n7829) );
  NAND2_X1 U6024 ( .A1(n6513), .A2(n5078), .ZN(n5077) );
  AND2_X1 U6025 ( .A1(n6767), .A2(n6766), .ZN(n6892) );
  INV_X1 U6026 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8028) );
  XNOR2_X1 U6027 ( .A(n5882), .B(n5886), .ZN(n8029) );
  INV_X1 U6028 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7997) );
  OR2_X1 U6029 ( .A1(n6711), .A2(n6703), .ZN(n5884) );
  INV_X1 U6030 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10302) );
  INV_X1 U6031 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10313) );
  INV_X1 U6032 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5899) );
  INV_X1 U6033 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8364) );
  INV_X1 U6034 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10312) );
  INV_X1 U6035 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7352) );
  INV_X1 U6036 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7351) );
  INV_X1 U6037 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7257) );
  INV_X1 U6038 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6967) );
  INV_X1 U6039 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U6040 ( .A1(n5931), .A2(n5951), .ZN(n6871) );
  NAND2_X1 U6041 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4900) );
  NAND2_X1 U6042 ( .A1(n5937), .A2(n5936), .ZN(n4898) );
  NAND2_X1 U6043 ( .A1(n5937), .A2(n5055), .ZN(n4899) );
  NAND2_X1 U6044 ( .A1(n4695), .A2(n4692), .ZN(n9296) );
  NAND2_X1 U6045 ( .A1(n4697), .A2(n4700), .ZN(n4693) );
  AND2_X1 U6046 ( .A1(n7239), .A2(n6133), .ZN(n8437) );
  NAND2_X1 U6047 ( .A1(n9386), .A2(n6304), .ZN(n9354) );
  AND2_X1 U6048 ( .A1(n4552), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U6049 ( .A1(n4505), .A2(n4690), .ZN(n4687) );
  NAND2_X1 U6050 ( .A1(n9387), .A2(n9388), .ZN(n9386) );
  NAND2_X1 U6051 ( .A1(n7568), .A2(n4970), .ZN(n4967) );
  NAND2_X1 U6052 ( .A1(n4691), .A2(n4701), .ZN(n9413) );
  OR2_X1 U6053 ( .A1(n9327), .A2(n4703), .ZN(n4691) );
  OAI21_X1 U6054 ( .B1(n9387), .B2(n6303), .A(n4682), .ZN(n9353) );
  NAND2_X1 U6055 ( .A1(n6355), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9462) );
  NAND2_X1 U6056 ( .A1(n5706), .A2(n5705), .ZN(n9475) );
  NAND2_X1 U6057 ( .A1(n9722), .A2(n5767), .ZN(n5706) );
  INV_X1 U6058 ( .A(n5372), .ZN(n9492) );
  INV_X1 U6059 ( .A(n5232), .ZN(n9494) );
  NAND2_X1 U6060 ( .A1(n9533), .A2(n9534), .ZN(n9554) );
  OAI21_X1 U6061 ( .B1(n9604), .B2(n9599), .A(n6934), .ZN(n9602) );
  OR2_X1 U6062 ( .A1(n6973), .A2(n6974), .ZN(n7031) );
  NOR2_X1 U6063 ( .A1(n7668), .A2(n7667), .ZN(n7893) );
  OR2_X1 U6064 ( .A1(n7888), .A2(n7889), .ZN(n9616) );
  OR2_X1 U6065 ( .A1(n9619), .A2(n9618), .ZN(n9629) );
  AOI21_X1 U6066 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9627), .A(n9625), .ZN(
        n9626) );
  AOI211_X1 U6067 ( .C1(n9651), .C2(n9654), .A(n9885), .B(n9653), .ZN(n9896)
         );
  AOI21_X1 U6068 ( .B1(n4493), .B2(n9686), .A(n4859), .ZN(n4858) );
  NAND2_X1 U6069 ( .A1(n9684), .A2(n9878), .ZN(n4750) );
  NAND2_X1 U6070 ( .A1(n4844), .A2(n5687), .ZN(n9718) );
  NAND2_X1 U6071 ( .A1(n5686), .A2(n5150), .ZN(n4844) );
  OAI21_X1 U6072 ( .B1(n9775), .B2(n4478), .A(n5622), .ZN(n9759) );
  AND2_X1 U6073 ( .A1(n8278), .A2(n8268), .ZN(n9760) );
  NAND2_X1 U6074 ( .A1(n4646), .A2(n4647), .ZN(n9790) );
  NAND2_X1 U6075 ( .A1(n9818), .A2(n4648), .ZN(n4646) );
  NAND2_X1 U6076 ( .A1(n5509), .A2(n5508), .ZN(n9862) );
  NAND2_X1 U6077 ( .A1(n7696), .A2(n5406), .ZN(n7813) );
  AND2_X1 U6078 ( .A1(n5110), .A2(n8310), .ZN(n7700) );
  OR2_X1 U6079 ( .A1(n10063), .A2(n5780), .ZN(n9814) );
  NAND2_X1 U6080 ( .A1(n10053), .A2(n7459), .ZN(n10049) );
  OR2_X1 U6081 ( .A1(n10063), .A2(n7817), .ZN(n7459) );
  NAND2_X1 U6082 ( .A1(n7450), .A2(n9829), .ZN(n9850) );
  INV_X1 U6083 ( .A(n9829), .ZN(n10052) );
  INV_X1 U6084 ( .A(n7650), .ZN(n7653) );
  NAND2_X1 U6085 ( .A1(n6870), .A2(n6847), .ZN(n4862) );
  NOR2_X1 U6086 ( .A1(n9896), .A2(n9895), .ZN(n9969) );
  INV_X1 U6087 ( .A(n5841), .ZN(n5842) );
  INV_X1 U6088 ( .A(n9706), .ZN(n9979) );
  INV_X1 U6089 ( .A(n9418), .ZN(n9995) );
  INV_X1 U6090 ( .A(n9781), .ZN(n9999) );
  AOI21_X1 U6091 ( .B1(n5589), .B2(P2_DATAO_REG_8__SCAN_IN), .A(n4763), .ZN(
        n4762) );
  AND2_X1 U6092 ( .A1(n4459), .A2(n6975), .ZN(n4763) );
  AND2_X1 U6093 ( .A1(n6904), .A2(n6864), .ZN(n10020) );
  NAND2_X1 U6094 ( .A1(n5218), .A2(n5219), .ZN(n5174) );
  INV_X1 U6095 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10285) );
  CLKBUF_X1 U6096 ( .A(n5825), .Z(n10031) );
  INV_X1 U6097 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8101) );
  INV_X1 U6098 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8088) );
  INV_X1 U6099 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8000) );
  OAI21_X1 U6100 ( .B1(n5776), .B2(n5169), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5850) );
  INV_X1 U6101 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10288) );
  INV_X1 U6102 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7752) );
  INV_X1 U6103 ( .A(n8223), .ZN(n8303) );
  INV_X1 U6104 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7535) );
  INV_X1 U6105 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7430) );
  INV_X1 U6106 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6968) );
  INV_X1 U6107 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10266) );
  INV_X1 U6108 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10265) );
  AND2_X1 U6109 ( .A1(n5307), .A2(n5331), .ZN(n9520) );
  NOR2_X4 U6110 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7778) );
  NAND2_X1 U6111 ( .A1(n5041), .A2(n8557), .ZN(n5040) );
  OAI22_X1 U6112 ( .A1(n7520), .A2(n7808), .B1(n6021), .B2(n6478), .ZN(n7586)
         );
  AND2_X1 U6113 ( .A1(n4783), .A2(n4786), .ZN(n8856) );
  NAND2_X1 U6114 ( .A1(n4481), .A2(n10092), .ZN(n4582) );
  AOI21_X1 U6115 ( .B1(n4743), .B2(n8883), .A(n4740), .ZN(n6098) );
  INV_X1 U6116 ( .A(n5083), .ZN(n5082) );
  OAI21_X1 U6117 ( .B1(n8950), .B2(n8949), .A(n10141), .ZN(n5084) );
  OAI21_X1 U6118 ( .B1(n8953), .B2(n10111), .A(n8952), .ZN(n5083) );
  OR2_X1 U6119 ( .A1(n8953), .A2(n9135), .ZN(n5146) );
  INV_X1 U6120 ( .A(n6757), .ZN(n6758) );
  OAI21_X1 U6121 ( .B1(n9172), .B2(n9147), .A(n6756), .ZN(n6757) );
  OAI22_X1 U6122 ( .A1(n8953), .A2(n9211), .B1(n10178), .B2(n6822), .ZN(n6823)
         );
  OR2_X1 U6123 ( .A1(n9172), .A2(n9234), .ZN(n4605) );
  AND2_X1 U6124 ( .A1(n6344), .A2(n9434), .ZN(n6363) );
  NAND2_X1 U6125 ( .A1(n5003), .A2(n6151), .ZN(n7358) );
  OR2_X1 U6126 ( .A1(n8360), .A2(n8359), .ZN(n4563) );
  NAND2_X1 U6127 ( .A1(n8212), .A2(n9940), .ZN(n6857) );
  NOR2_X1 U6128 ( .A1(n6114), .A2(n6116), .ZN(n6117) );
  NOR2_X1 U6129 ( .A1(n10077), .A2(n6115), .ZN(n6116) );
  OAI21_X1 U6130 ( .B1(n9973), .B2(n4655), .A(n4653), .ZN(P1_U3549) );
  INV_X1 U6131 ( .A(n10077), .ZN(n4655) );
  AOI21_X1 U6132 ( .B1(n9690), .B2(n9940), .A(n4654), .ZN(n4653) );
  NOR2_X1 U6133 ( .A1(n10077), .A2(n10394), .ZN(n4654) );
  INV_X1 U6134 ( .A(n6828), .ZN(n6829) );
  OAI22_X1 U6135 ( .A1(n9677), .A2(n10017), .B1(n10074), .B2(n6827), .ZN(n6828) );
  OR2_X1 U6136 ( .A1(n10074), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U6137 ( .A1(n9973), .A2(n10074), .ZN(n4749) );
  AND2_X1 U6138 ( .A1(n8281), .A2(n8285), .ZN(n9663) );
  OAI211_X1 U6139 ( .C1(n5316), .C2(n9561), .A(n5279), .B(n5278), .ZN(n7496)
         );
  AND2_X1 U6140 ( .A1(n4975), .A2(n6281), .ZN(n4471) );
  AND3_X1 U6141 ( .A1(n9663), .A2(n8286), .A3(n4836), .ZN(n4472) );
  INV_X1 U6142 ( .A(n8784), .ZN(n7869) );
  INV_X1 U6143 ( .A(n7428), .ZN(n5780) );
  OR2_X1 U6144 ( .A1(n5558), .A2(n5557), .ZN(n4474) );
  OR2_X1 U6145 ( .A1(n4645), .A2(n5609), .ZN(n4475) );
  OR2_X1 U6146 ( .A1(n6275), .A2(n6273), .ZN(n4476) );
  AND2_X1 U6147 ( .A1(n5117), .A2(n5115), .ZN(n4477) );
  NOR2_X1 U6148 ( .A1(n9781), .A2(n9479), .ZN(n4478) );
  NAND2_X1 U6149 ( .A1(n8975), .A2(n8970), .ZN(n8729) );
  XNOR2_X1 U6150 ( .A(n5470), .B(SI_13_), .ZN(n5468) );
  OR2_X1 U6151 ( .A1(n8718), .A2(n8720), .ZN(n4479) );
  OR2_X1 U6152 ( .A1(n8427), .A2(n5045), .ZN(n4480) );
  XNOR2_X1 U6153 ( .A(n8915), .B(n8914), .ZN(n4481) );
  NAND2_X1 U6154 ( .A1(n4862), .A2(n4522), .ZN(n7692) );
  INV_X1 U6155 ( .A(n7692), .ZN(n7516) );
  AND2_X1 U6156 ( .A1(n4977), .A2(n4557), .ZN(n4483) );
  INV_X1 U6157 ( .A(n5145), .ZN(n5094) );
  AND2_X1 U6158 ( .A1(n4815), .A2(n8123), .ZN(n4484) );
  OR2_X1 U6159 ( .A1(n9180), .A2(n8778), .ZN(n4485) );
  OR2_X1 U6160 ( .A1(n8759), .A2(n6754), .ZN(n4486) );
  OR2_X1 U6161 ( .A1(n4867), .A2(n4866), .ZN(n4487) );
  NAND2_X1 U6162 ( .A1(n8280), .A2(n8192), .ZN(n8258) );
  INV_X1 U6163 ( .A(n8258), .ZN(n4634) );
  AND2_X1 U6164 ( .A1(n4471), .A2(n4557), .ZN(n4488) );
  AND2_X1 U6165 ( .A1(n8587), .A2(n8722), .ZN(n8726) );
  INV_X1 U6166 ( .A(n8726), .ZN(n4880) );
  NAND2_X1 U6167 ( .A1(n5116), .A2(n5117), .ZN(n7622) );
  NAND2_X1 U6168 ( .A1(n5116), .A2(n4477), .ZN(n5118) );
  AND3_X1 U6169 ( .A1(n4912), .A2(n5963), .A3(P2_REG2_REG_9__SCAN_IN), .ZN(
        n4489) );
  AND2_X1 U6170 ( .A1(n7592), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4490) );
  AND2_X1 U6171 ( .A1(n5980), .A2(n5924), .ZN(n7106) );
  INV_X1 U6172 ( .A(n7106), .ZN(n4785) );
  AND3_X1 U6173 ( .A1(n4825), .A2(n6377), .A3(n4824), .ZN(n4491) );
  INV_X1 U6174 ( .A(n7810), .ZN(n7011) );
  NAND2_X1 U6175 ( .A1(n5013), .A2(n5014), .ZN(n4492) );
  AND2_X1 U6176 ( .A1(n8258), .A2(n5741), .ZN(n4493) );
  NAND2_X1 U6177 ( .A1(n9402), .A2(n6232), .ZN(n9275) );
  OR2_X1 U6178 ( .A1(n5260), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n4494) );
  AND2_X1 U6179 ( .A1(n4581), .A2(n4579), .ZN(n4495) );
  OR2_X1 U6180 ( .A1(n6568), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4496) );
  OR2_X1 U6181 ( .A1(n6620), .A2(n4826), .ZN(n4497) );
  OR2_X1 U6182 ( .A1(n5553), .A2(n5558), .ZN(n4498) );
  OAI211_X1 U6183 ( .C1(n6816), .C2(n7185), .A(n6419), .B(n6418), .ZN(n10150)
         );
  OAI21_X1 U6184 ( .B1(n7492), .B2(n6168), .A(n6167), .ZN(n7568) );
  AND2_X1 U6185 ( .A1(n7390), .A2(n8788), .ZN(n4499) );
  AND2_X1 U6186 ( .A1(n6243), .A2(n4989), .ZN(n4500) );
  NAND4_X2 U6187 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n9498)
         );
  NAND2_X1 U6188 ( .A1(n7556), .A2(n7805), .ZN(n4501) );
  OAI21_X1 U6189 ( .B1(n9380), .B2(n4977), .A(n4471), .ZN(n9394) );
  AND2_X1 U6190 ( .A1(n4705), .A2(n4704), .ZN(n4502) );
  AOI21_X1 U6191 ( .B1(n8478), .B2(n8479), .A(n8420), .ZN(n8547) );
  OAI21_X1 U6192 ( .B1(n9818), .B2(n5577), .A(n5576), .ZN(n9801) );
  NAND2_X1 U6193 ( .A1(n5065), .A2(n6565), .ZN(n9088) );
  AND2_X1 U6194 ( .A1(n8204), .A2(n8297), .ZN(n4503) );
  AND2_X1 U6195 ( .A1(n5885), .A2(n5056), .ZN(n4504) );
  NAND2_X1 U6196 ( .A1(n5419), .A2(n5418), .ZN(n7821) );
  AND2_X1 U6197 ( .A1(n4500), .A2(n4688), .ZN(n4505) );
  AND2_X1 U6198 ( .A1(n10006), .A2(n9481), .ZN(n4506) );
  INV_X1 U6199 ( .A(n7909), .ZN(n4608) );
  INV_X1 U6200 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5368) );
  XOR2_X1 U6201 ( .A(n10150), .B(n7111), .Z(n4507) );
  AND2_X1 U6202 ( .A1(n8789), .A2(n6739), .ZN(n4508) );
  AND2_X1 U6203 ( .A1(n9378), .A2(n9377), .ZN(n4509) );
  AND3_X1 U6204 ( .A1(n9789), .A2(n9804), .A3(n4632), .ZN(n4510) );
  NAND2_X1 U6205 ( .A1(n8409), .A2(n8408), .ZN(n8524) );
  AND2_X1 U6206 ( .A1(n8389), .A2(n9081), .ZN(n4511) );
  AND2_X1 U6207 ( .A1(n6490), .A2(n6368), .ZN(n4512) );
  INV_X1 U6208 ( .A(n5127), .ZN(n9689) );
  NOR3_X1 U6209 ( .A1(n9735), .A2(n9690), .A3(n5128), .ZN(n5127) );
  AND3_X1 U6210 ( .A1(n5844), .A2(n5843), .A3(n5842), .ZN(n4513) );
  AND2_X1 U6211 ( .A1(n8153), .A2(n8156), .ZN(n8249) );
  AND3_X1 U6212 ( .A1(n8657), .A2(n8656), .A3(n8655), .ZN(n4514) );
  OR2_X1 U6213 ( .A1(n9190), .A2(n8984), .ZN(n8717) );
  INV_X1 U6214 ( .A(n9357), .ZN(n9983) );
  NAND2_X1 U6215 ( .A1(n6674), .A2(n6673), .ZN(n9169) );
  AND2_X1 U6216 ( .A1(n8737), .A2(n4610), .ZN(n4515) );
  NAND2_X1 U6217 ( .A1(n5567), .A2(n5566), .ZN(n9943) );
  INV_X1 U6218 ( .A(n5131), .ZN(n9688) );
  INV_X1 U6219 ( .A(n5575), .ZN(n6852) );
  OR2_X1 U6220 ( .A1(n8701), .A2(n4889), .ZN(n4516) );
  OR2_X1 U6221 ( .A1(n8673), .A2(n6697), .ZN(n4517) );
  AND2_X1 U6222 ( .A1(n8588), .A2(n8988), .ZN(n8720) );
  INV_X1 U6223 ( .A(n8720), .ZN(n4723) );
  AND2_X1 U6224 ( .A1(n4492), .A2(n7557), .ZN(n4518) );
  AOI22_X1 U6225 ( .A1(n9472), .A2(n9457), .B1(n6856), .B2(n9470), .ZN(n5830)
         );
  OR2_X1 U6226 ( .A1(n9983), .A2(n6305), .ZN(n4519) );
  NAND2_X1 U6227 ( .A1(n5226), .A2(n5225), .ZN(n5260) );
  NAND2_X1 U6228 ( .A1(n9418), .A2(n9478), .ZN(n4520) );
  NAND2_X1 U6229 ( .A1(n6186), .A2(n9320), .ZN(n4521) );
  AND2_X1 U6230 ( .A1(n9180), .A2(n8985), .ZN(n8723) );
  NOR2_X1 U6231 ( .A1(n5513), .A2(n4942), .ZN(n4941) );
  AND2_X1 U6232 ( .A1(n5231), .A2(n5230), .ZN(n4522) );
  OR2_X1 U6233 ( .A1(n5372), .A2(n9325), .ZN(n8121) );
  INV_X1 U6234 ( .A(n8121), .ZN(n4797) );
  OR2_X1 U6235 ( .A1(n9023), .A2(n8702), .ZN(n4523) );
  AND2_X1 U6236 ( .A1(n4878), .A2(n4877), .ZN(n4524) );
  OR2_X1 U6237 ( .A1(n6620), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n4525) );
  INV_X1 U6238 ( .A(n6293), .ZN(n4704) );
  NOR2_X1 U6239 ( .A1(n9963), .A2(n9486), .ZN(n4526) );
  AND2_X1 U6240 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4527) );
  NOR2_X1 U6241 ( .A1(n9418), .A2(n9478), .ZN(n4528) );
  INV_X1 U6242 ( .A(n4954), .ZN(n4953) );
  AND2_X1 U6243 ( .A1(n6820), .A2(n6819), .ZN(n4529) );
  OR2_X1 U6244 ( .A1(n4498), .A2(n4939), .ZN(n4530) );
  INV_X1 U6245 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10022) );
  INV_X1 U6246 ( .A(n5134), .ZN(n5133) );
  NAND2_X1 U6247 ( .A1(n5136), .A2(n5135), .ZN(n5134) );
  NOR2_X1 U6248 ( .A1(n8721), .A2(n6697), .ZN(n4531) );
  NOR2_X1 U6249 ( .A1(n9169), .A2(n8775), .ZN(n4532) );
  NAND2_X1 U6250 ( .A1(n6369), .A2(n4512), .ZN(n4533) );
  NAND2_X1 U6251 ( .A1(n9328), .A2(n4502), .ZN(n4534) );
  OR2_X1 U6252 ( .A1(n9972), .A2(n8123), .ZN(n4535) );
  OR2_X1 U6253 ( .A1(n4473), .A2(n5121), .ZN(n4536) );
  INV_X1 U6254 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U6255 ( .A1(n4839), .A2(n4519), .ZN(n4838) );
  NAND2_X1 U6256 ( .A1(n6191), .A2(n4966), .ZN(n4537) );
  NOR2_X1 U6257 ( .A1(n6806), .A2(n8742), .ZN(n4538) );
  INV_X1 U6258 ( .A(n4971), .ZN(n4970) );
  NAND2_X1 U6259 ( .A1(n7569), .A2(n4521), .ZN(n4971) );
  INV_X1 U6260 ( .A(n4985), .ZN(n4984) );
  NAND2_X1 U6261 ( .A1(n4479), .A2(n8587), .ZN(n4985) );
  INV_X1 U6262 ( .A(n4857), .ZN(n4856) );
  NAND2_X1 U6263 ( .A1(n5622), .A2(n4520), .ZN(n4857) );
  INV_X1 U6264 ( .A(n8731), .ZN(n4871) );
  NAND2_X1 U6265 ( .A1(n8261), .A2(n8272), .ZN(n9704) );
  INV_X1 U6266 ( .A(n9704), .ZN(n4836) );
  OR2_X1 U6267 ( .A1(n9180), .A2(n8985), .ZN(n8722) );
  XNOR2_X1 U6268 ( .A(n5355), .B(SI_7_), .ZN(n5358) );
  AND2_X1 U6269 ( .A1(n7875), .A2(n8782), .ZN(n4539) );
  AND3_X1 U6270 ( .A1(n5354), .A2(n5352), .A3(n5353), .ZN(n4540) );
  INV_X1 U6271 ( .A(n8330), .ZN(n4757) );
  AND2_X1 U6272 ( .A1(n4960), .A2(n4964), .ZN(n4541) );
  AND2_X1 U6273 ( .A1(n5093), .A2(n6659), .ZN(n4542) );
  AND2_X1 U6274 ( .A1(n9039), .A2(n9065), .ZN(n4543) );
  AND2_X1 U6275 ( .A1(n9180), .A2(n8778), .ZN(n4544) );
  OAI21_X1 U6276 ( .B1(n4955), .B2(n4954), .A(n5457), .ZN(n4952) );
  OR2_X1 U6277 ( .A1(n9185), .A2(n9001), .ZN(n4545) );
  AND2_X1 U6278 ( .A1(n9855), .A2(n5508), .ZN(n4546) );
  AND2_X1 U6279 ( .A1(n4876), .A2(n4720), .ZN(n4547) );
  AND2_X1 U6280 ( .A1(n8262), .A2(n8191), .ZN(n9686) );
  NAND2_X1 U6281 ( .A1(n8426), .A2(n8776), .ZN(n4548) );
  OR2_X1 U6282 ( .A1(n4470), .A2(n6897), .ZN(n4549) );
  INV_X1 U6283 ( .A(n8403), .ZN(n5036) );
  AND2_X1 U6284 ( .A1(n4474), .A2(n4941), .ZN(n4550) );
  NOR2_X1 U6285 ( .A1(n5624), .A2(n4963), .ZN(n4962) );
  AND2_X1 U6286 ( .A1(n6153), .A2(n6151), .ZN(n4551) );
  AND2_X1 U6287 ( .A1(n6251), .A2(n4988), .ZN(n4552) );
  INV_X1 U6288 ( .A(n5433), .ZN(n4955) );
  NAND2_X1 U6289 ( .A1(n6871), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4553) );
  AND2_X1 U6290 ( .A1(n5219), .A2(n4808), .ZN(n4554) );
  NAND2_X1 U6291 ( .A1(n10003), .A2(n5812), .ZN(n4555) );
  INV_X1 U6292 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5911) );
  INV_X1 U6293 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5167) );
  INV_X1 U6294 ( .A(n7265), .ZN(n7266) );
  NAND2_X1 U6295 ( .A1(n7264), .A2(n10108), .ZN(n7265) );
  INV_X1 U6296 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10304) );
  OR2_X1 U6297 ( .A1(n10063), .A2(n7451), .ZN(n9891) );
  INV_X1 U6298 ( .A(n6514), .ZN(n4771) );
  NAND2_X1 U6299 ( .A1(n7865), .A2(n7864), .ZN(n7902) );
  AND2_X1 U6300 ( .A1(n7705), .A2(n7709), .ZN(n7706) );
  NAND2_X1 U6301 ( .A1(n7706), .A2(n8052), .ZN(n7818) );
  AND2_X1 U6302 ( .A1(n5916), .A2(n5881), .ZN(n5901) );
  AND2_X1 U6303 ( .A1(n5833), .A2(n5125), .ZN(n4556) );
  AND2_X1 U6304 ( .A1(n6715), .A2(n6920), .ZN(n7013) );
  NAND2_X1 U6305 ( .A1(n7971), .A2(n8145), .ZN(n8076) );
  NAND2_X1 U6306 ( .A1(n4447), .A2(n6554), .ZN(n9100) );
  NAND2_X1 U6307 ( .A1(n4651), .A2(n4845), .ZN(n7982) );
  NAND2_X1 U6308 ( .A1(n8078), .A2(n5467), .ZN(n8022) );
  INV_X1 U6309 ( .A(n9377), .ZN(n4976) );
  OR2_X1 U6310 ( .A1(n6288), .A2(n6287), .ZN(n4557) );
  INV_X1 U6311 ( .A(n8975), .ZN(n8777) );
  AOI21_X1 U6312 ( .B1(n8969), .B2(n6688), .A(n6656), .ZN(n8975) );
  INV_X1 U6313 ( .A(n6478), .ZN(n4768) );
  AND2_X1 U6314 ( .A1(n5961), .A2(n5964), .ZN(n6478) );
  AND2_X1 U6315 ( .A1(n4667), .A2(n4501), .ZN(n7560) );
  NAND2_X1 U6316 ( .A1(n6683), .A2(n6682), .ZN(n8775) );
  INV_X1 U6317 ( .A(n8778), .ZN(n8985) );
  NAND2_X1 U6318 ( .A1(n6649), .A2(n6648), .ZN(n8778) );
  NOR2_X1 U6319 ( .A1(n4470), .A2(n8377), .ZN(n4558) );
  NAND2_X1 U6320 ( .A1(n7706), .A2(n5132), .ZN(n8017) );
  AND2_X1 U6321 ( .A1(n4664), .A2(n5137), .ZN(n4559) );
  INV_X1 U6322 ( .A(n4736), .ZN(n4735) );
  OAI21_X1 U6323 ( .B1(n4737), .B2(n6069), .A(n6073), .ZN(n4736) );
  AND2_X1 U6324 ( .A1(n4831), .A2(n4830), .ZN(n4560) );
  INV_X1 U6325 ( .A(n8555), .ZN(n8557) );
  INV_X1 U6326 ( .A(n8082), .ZN(n5135) );
  NAND2_X1 U6327 ( .A1(n5522), .A2(n5521), .ZN(n9867) );
  OAI21_X1 U6328 ( .B1(n7111), .B2(n4678), .A(n10117), .ZN(n7092) );
  NOR2_X1 U6329 ( .A1(n7320), .A2(n7460), .ZN(n7248) );
  AND2_X1 U6330 ( .A1(n7248), .A2(n10046), .ZN(n4561) );
  XNOR2_X1 U6331 ( .A(n5949), .B(n6868), .ZN(n7203) );
  INV_X1 U6332 ( .A(n7508), .ZN(n5116) );
  NAND2_X1 U6333 ( .A1(n5796), .A2(n8304), .ZN(n7372) );
  XOR2_X1 U6334 ( .A(n7106), .B(P2_REG2_REG_14__SCAN_IN), .Z(n4562) );
  INV_X1 U6335 ( .A(n9325), .ZN(n5115) );
  XNOR2_X1 U6336 ( .A(n5011), .B(n5010), .ZN(n7428) );
  INV_X1 U6337 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6684) );
  INV_X1 U6338 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4863) );
  AND2_X1 U6339 ( .A1(n8365), .A2(n8612), .ZN(n8763) );
  AND2_X1 U6340 ( .A1(n8365), .A2(n8584), .ZN(n8762) );
  INV_X1 U6341 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n4923) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4622) );
  INV_X1 U6343 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n4917) );
  AOI21_X2 U6344 ( .B1(n9080), .B2(n9077), .A(n6580), .ZN(n9026) );
  INV_X2 U6345 ( .A(n6738), .ZN(n5087) );
  XNOR2_X2 U6346 ( .A(n8638), .B(n8790), .ZN(n6738) );
  NAND2_X1 U6347 ( .A1(n6545), .A2(n6544), .ZN(n8003) );
  NAND2_X1 U6348 ( .A1(n5208), .A2(n5207), .ZN(n5257) );
  NAND2_X1 U6349 ( .A1(n4592), .A2(n4871), .ZN(n5095) );
  NAND2_X1 U6350 ( .A1(n6477), .A2(n6476), .ZN(n7420) );
  NAND2_X1 U6351 ( .A1(n4913), .A2(n6478), .ZN(n4912) );
  NOR2_X2 U6352 ( .A1(n5953), .A2(n7162), .ZN(n7283) );
  NAND2_X1 U6353 ( .A1(n6393), .A2(n4603), .ZN(n5933) );
  NAND2_X1 U6354 ( .A1(n5973), .A2(n8829), .ZN(n8834) );
  NAND2_X1 U6355 ( .A1(n4914), .A2(n4915), .ZN(n8921) );
  NOR2_X1 U6356 ( .A1(n7174), .A2(n10472), .ZN(n7173) );
  NAND2_X1 U6357 ( .A1(n7286), .A2(n5142), .ZN(n5962) );
  OAI211_X1 U6358 ( .C1(n6099), .C2(n10088), .A(n4774), .B(n6098), .ZN(
        P2_U3201) );
  OAI21_X1 U6359 ( .B1(n8362), .B2(n8361), .A(n4563), .ZN(P1_U3242) );
  NOR3_X1 U6360 ( .A1(n8920), .A2(n8919), .A3(n8918), .ZN(n8924) );
  NAND2_X1 U6361 ( .A1(n8865), .A2(n4602), .ZN(n5982) );
  NAND2_X1 U6362 ( .A1(n4625), .A2(n5480), .ZN(n5501) );
  NAND2_X1 U6363 ( .A1(n8902), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U6364 ( .A1(n5978), .A2(n6535), .ZN(n5979) );
  XNOR2_X1 U6365 ( .A(n4617), .B(n4616), .ZN(n6702) );
  OR2_X1 U6366 ( .A1(n6695), .A2(n6394), .ZN(n4570) );
  INV_X1 U6367 ( .A(n10094), .ZN(n4731) );
  INV_X1 U6368 ( .A(n7065), .ZN(n4739) );
  AND3_X2 U6369 ( .A1(n4590), .A2(n4626), .A3(n4482), .ZN(n5955) );
  AOI21_X1 U6370 ( .B1(n6059), .B2(n4727), .A(n4725), .ZN(n4724) );
  NAND2_X1 U6371 ( .A1(n7181), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U6372 ( .A1(n5095), .A2(n5094), .ZN(n4617) );
  OR2_X1 U6373 ( .A1(n6401), .A2(n6394), .ZN(n6396) );
  NAND2_X1 U6374 ( .A1(n6420), .A2(n10119), .ZN(n10134) );
  NAND3_X1 U6375 ( .A1(n9026), .A2(n8589), .A3(n5099), .ZN(n5096) );
  AOI21_X2 U6376 ( .B1(n9008), .B2(n9012), .A(n8704), .ZN(n8997) );
  AND2_X2 U6377 ( .A1(n4572), .A2(n4929), .ZN(n5394) );
  NAND3_X1 U6378 ( .A1(n4932), .A2(n4931), .A3(n4930), .ZN(n4572) );
  OAI21_X4 U6379 ( .B1(n5412), .B2(n5411), .A(n5410), .ZN(n5434) );
  NAND2_X1 U6380 ( .A1(n4677), .A2(n5022), .ZN(n8495) );
  INV_X1 U6381 ( .A(n6445), .ZN(n5085) );
  INV_X1 U6382 ( .A(n7085), .ZN(n8793) );
  AND2_X1 U6383 ( .A1(n4676), .A2(n4675), .ZN(n4590) );
  AOI21_X1 U6384 ( .B1(n4994), .B2(n4997), .A(n4992), .ZN(n4991) );
  XNOR2_X2 U6385 ( .A(n5287), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U6386 ( .A1(n8671), .A2(n8670), .ZN(n4897) );
  OAI21_X1 U6387 ( .B1(n4893), .B2(n4892), .A(n8690), .ZN(n4891) );
  NAND2_X1 U6388 ( .A1(n7409), .A2(n7085), .ZN(n10116) );
  NOR2_X1 U6389 ( .A1(n8741), .A2(n8740), .ZN(n8758) );
  AOI21_X1 U6390 ( .B1(n8699), .B2(n6697), .A(n8702), .ZN(n4869) );
  NOR2_X1 U6391 ( .A1(n8744), .A2(n8743), .ZN(n8761) );
  OAI21_X1 U6392 ( .B1(n8158), .B2(n8317), .A(n8157), .ZN(n4581) );
  NAND2_X1 U6393 ( .A1(n8147), .A2(n8297), .ZN(n4584) );
  NOR2_X1 U6394 ( .A1(n8203), .A2(n4586), .ZN(n4585) );
  AOI21_X1 U6395 ( .B1(n8190), .B2(n8189), .A(n8188), .ZN(n8202) );
  NAND3_X1 U6396 ( .A1(n8938), .A2(n8937), .A3(n4582), .ZN(P2_U3200) );
  NAND2_X1 U6397 ( .A1(n4905), .A2(n4904), .ZN(n4903) );
  NAND2_X1 U6398 ( .A1(n4921), .A2(n4920), .ZN(n8865) );
  NOR2_X1 U6399 ( .A1(n5954), .A2(n7283), .ZN(n7160) );
  NAND2_X1 U6400 ( .A1(n8834), .A2(n5974), .ZN(n5977) );
  NAND2_X1 U6401 ( .A1(n7593), .A2(n7592), .ZN(n4911) );
  INV_X1 U6402 ( .A(n4909), .ZN(n4905) );
  NAND2_X1 U6403 ( .A1(n4922), .A2(n8862), .ZN(n4921) );
  XNOR2_X2 U6404 ( .A(n5220), .B(n5219), .ZN(n5824) );
  NAND2_X1 U6405 ( .A1(n4584), .A2(n4583), .ZN(n8158) );
  NAND2_X1 U6406 ( .A1(n8139), .A2(n8123), .ZN(n4583) );
  AND2_X2 U6407 ( .A1(n5303), .A2(n5162), .ZN(n5165) );
  NAND3_X1 U6408 ( .A1(n8210), .A2(n9663), .A3(n4587), .ZN(n4586) );
  NAND2_X1 U6409 ( .A1(n4798), .A2(n7722), .ZN(n7739) );
  NAND2_X1 U6410 ( .A1(n7249), .A2(n8234), .ZN(n5101) );
  NAND2_X1 U6411 ( .A1(n8128), .A2(n4589), .ZN(n4802) );
  AOI21_X2 U6412 ( .B1(n6802), .B2(n8610), .A(n4591), .ZN(n8576) );
  AND2_X1 U6413 ( .A1(n8637), .A2(n8651), .ZN(n7379) );
  NAND2_X1 U6414 ( .A1(n5495), .A2(n4550), .ZN(n4940) );
  INV_X1 U6415 ( .A(n4606), .ZN(n8964) );
  OAI21_X2 U6416 ( .B1(n5583), .B2(n5582), .A(n5581), .ZN(n5600) );
  NAND2_X1 U6417 ( .A1(n8003), .A2(n8674), .ZN(n6555) );
  AOI21_X1 U6418 ( .B1(n5075), .B2(n5079), .A(n4539), .ZN(n5073) );
  AOI21_X1 U6419 ( .B1(n6702), .B2(n9094), .A(n6701), .ZN(n9165) );
  NAND2_X1 U6420 ( .A1(n5073), .A2(n5074), .ZN(n5071) );
  AND2_X1 U6421 ( .A1(n5071), .A2(n8672), .ZN(n5070) );
  OAI21_X1 U6422 ( .B1(n6779), .B2(n6778), .A(n9094), .ZN(n6783) );
  NAND2_X1 U6423 ( .A1(n5199), .A2(n5200), .ZN(n4924) );
  NAND2_X1 U6424 ( .A1(n6516), .A2(n6515), .ZN(n7993) );
  INV_X1 U6425 ( .A(n5081), .ZN(n5076) );
  INV_X1 U6426 ( .A(n6777), .ZN(n4592) );
  NAND2_X1 U6427 ( .A1(n8964), .A2(n6658), .ZN(n6660) );
  OAI21_X1 U6428 ( .B1(n8973), .B2(n4544), .A(n4485), .ZN(n4606) );
  NAND3_X1 U6429 ( .A1(n4594), .A2(n4593), .A3(n8631), .ZN(n7380) );
  NAND2_X1 U6430 ( .A1(n8626), .A2(n8632), .ZN(n4593) );
  NAND3_X1 U6431 ( .A1(n8632), .A2(n8623), .A3(n8625), .ZN(n4594) );
  NAND2_X1 U6432 ( .A1(n7412), .A2(n8596), .ZN(n10103) );
  NAND2_X1 U6433 ( .A1(n4993), .A2(n4991), .ZN(n7635) );
  NAND4_X1 U6434 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5056), .ZN(n4597)
         );
  NAND2_X1 U6435 ( .A1(n4598), .A2(n8637), .ZN(n7234) );
  NAND2_X1 U6436 ( .A1(n7379), .A2(n7380), .ZN(n4598) );
  INV_X1 U6437 ( .A(n4674), .ZN(n4626) );
  AND2_X2 U6438 ( .A1(n8407), .A2(n8406), .ZN(n8409) );
  AOI21_X2 U6439 ( .B1(n9854), .B2(n9863), .A(n5807), .ZN(n9839) );
  NAND2_X2 U6440 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  INV_X1 U6441 ( .A(n9659), .ZN(n9658) );
  NAND2_X1 U6442 ( .A1(n8515), .A2(n8403), .ZN(n5033) );
  OAI21_X1 U6443 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5458) );
  NAND3_X1 U6444 ( .A1(n4931), .A2(n4932), .A3(n4936), .ZN(n4601) );
  XNOR2_X2 U6445 ( .A(n5932), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U6446 ( .A1(n5057), .A2(n4545), .ZN(n8973) );
  NAND2_X1 U6447 ( .A1(n5831), .A2(n9878), .ZN(n4604) );
  NAND3_X1 U6448 ( .A1(n9171), .A2(n9170), .A3(n4605), .ZN(P2_U3455) );
  NAND2_X1 U6449 ( .A1(n8576), .A2(n8752), .ZN(n4611) );
  NAND2_X1 U6450 ( .A1(n7234), .A2(n5087), .ZN(n7233) );
  NAND2_X1 U6451 ( .A1(n8997), .A2(n4987), .ZN(n4986) );
  INV_X1 U6452 ( .A(n8433), .ZN(n6384) );
  NAND3_X1 U6453 ( .A1(n4613), .A2(n4708), .A3(n5471), .ZN(n5492) );
  NAND2_X1 U6454 ( .A1(n5434), .A2(n4709), .ZN(n4613) );
  NAND2_X1 U6455 ( .A1(n5257), .A2(n5256), .ZN(n5275) );
  NAND2_X1 U6456 ( .A1(n6380), .A2(n6381), .ZN(n9245) );
  INV_X1 U6457 ( .A(n9101), .ZN(n5068) );
  INV_X1 U6458 ( .A(n5095), .ZN(n6779) );
  NAND2_X1 U6459 ( .A1(n8982), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U6460 ( .A1(n9168), .A2(n9167), .ZN(n9171) );
  NAND2_X1 U6461 ( .A1(n4749), .A2(n4748), .ZN(n9974) );
  OR2_X2 U6462 ( .A1(n9781), .A2(n8255), .ZN(n8118) );
  CLKBUF_X1 U6463 ( .A(n10118), .Z(n4620) );
  OAI21_X1 U6464 ( .B1(n4782), .B2(n8843), .A(n4781), .ZN(n4780) );
  NAND2_X1 U6465 ( .A1(n4780), .A2(n4784), .ZN(n6024) );
  INV_X1 U6466 ( .A(n6881), .ZN(n5061) );
  NOR2_X4 U6467 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5936) );
  XNOR2_X1 U6468 ( .A(n6026), .B(n4776), .ZN(n4775) );
  NAND2_X1 U6469 ( .A1(n4775), .A2(n10092), .ZN(n4774) );
  INV_X1 U6470 ( .A(n4758), .ZN(n4755) );
  AND3_X1 U6471 ( .A1(n6395), .A2(n6397), .A3(n6396), .ZN(n6399) );
  OAI21_X1 U6472 ( .B1(n9063), .B2(n9065), .A(n8695), .ZN(n9020) );
  OAI21_X1 U6473 ( .B1(n8765), .B2(n4817), .A(n8764), .ZN(n4816) );
  OAI21_X2 U6474 ( .B1(n7420), .B2(n7637), .A(n6511), .ZN(n6513) );
  NAND2_X1 U6475 ( .A1(n9165), .A2(n10178), .ZN(n9168) );
  NAND2_X1 U6476 ( .A1(n5280), .A2(n9495), .ZN(n8305) );
  NAND4_X1 U6477 ( .A1(n4634), .A2(n8340), .A3(n9686), .A4(n4472), .ZN(n4633)
         );
  NAND3_X1 U6478 ( .A1(n8752), .A2(n8610), .A3(n8731), .ZN(n4637) );
  INV_X2 U6479 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6480 ( .A1(n9818), .A2(n4643), .ZN(n4638) );
  NAND2_X1 U6481 ( .A1(n4642), .A2(n4638), .ZN(n4854) );
  NAND2_X1 U6482 ( .A1(n7698), .A2(n4650), .ZN(n4651) );
  INV_X1 U6483 ( .A(n7982), .ZN(n5453) );
  OAI21_X1 U6484 ( .B1(n8236), .B2(n5248), .A(n7610), .ZN(n5249) );
  OAI211_X2 U6485 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_29__SCAN_IN), 
        .A(n4809), .B(n4658), .ZN(n10027) );
  NAND2_X1 U6486 ( .A1(n4666), .A2(n4559), .ZN(n4659) );
  AND2_X2 U6487 ( .A1(n4662), .A2(n4660), .ZN(n8056) );
  OR2_X1 U6488 ( .A1(n7874), .A2(n4661), .ZN(n4660) );
  INV_X1 U6489 ( .A(n7876), .ZN(n4661) );
  NAND2_X1 U6490 ( .A1(n4666), .A2(n4663), .ZN(n4662) );
  AND3_X1 U6491 ( .A1(n4664), .A2(n7876), .A3(n5137), .ZN(n4663) );
  NAND2_X1 U6492 ( .A1(n4669), .A2(n4668), .ZN(n7269) );
  OR2_X1 U6493 ( .A1(n7267), .A2(n7266), .ZN(n4668) );
  NAND3_X1 U6494 ( .A1(n7265), .A2(n7148), .A3(n7147), .ZN(n4669) );
  XNOR2_X1 U6495 ( .A(n4671), .B(n4670), .ZN(n7155) );
  INV_X1 U6496 ( .A(n7267), .ZN(n4671) );
  NAND4_X1 U6497 ( .A1(n4482), .A2(n4673), .A3(n4676), .A4(n4675), .ZN(n4672)
         );
  NAND3_X1 U6498 ( .A1(n6411), .A2(n4865), .A3(n5937), .ZN(n5925) );
  INV_X1 U6499 ( .A(n8495), .ZN(n8391) );
  INV_X1 U6500 ( .A(n7312), .ZN(n4678) );
  INV_X1 U6501 ( .A(n4679), .ZN(n9435) );
  NAND3_X1 U6502 ( .A1(n4537), .A2(n4684), .A3(n4968), .ZN(n6198) );
  NAND3_X1 U6503 ( .A1(n7492), .A2(n6167), .A3(n6191), .ZN(n4684) );
  NAND2_X1 U6504 ( .A1(n6223), .A2(n4505), .ZN(n4685) );
  NAND2_X1 U6505 ( .A1(n4685), .A2(n4686), .ZN(n9364) );
  NAND2_X1 U6506 ( .A1(n9327), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U6507 ( .A1(n7778), .A2(n5186), .ZN(n4707) );
  NAND2_X1 U6508 ( .A1(n4952), .A2(n4709), .ZN(n4708) );
  INV_X1 U6509 ( .A(n4952), .ZN(n4951) );
  INV_X1 U6510 ( .A(n5468), .ZN(n4711) );
  OAI21_X1 U6511 ( .B1(n4868), .B2(n4712), .A(n4516), .ZN(n8712) );
  NAND2_X1 U6512 ( .A1(n7119), .A2(n6486), .ZN(n4717) );
  INV_X1 U6513 ( .A(n9073), .ZN(n8685) );
  NAND3_X1 U6514 ( .A1(n4875), .A2(n4547), .A3(n4487), .ZN(n4719) );
  NAND2_X1 U6515 ( .A1(n5454), .A2(n5432), .ZN(n4954) );
  MUX2_X1 U6516 ( .A(n10457), .B(n6960), .S(n6390), .Z(n5413) );
  INV_X1 U6517 ( .A(n4724), .ZN(n6066) );
  INV_X1 U6518 ( .A(n6070), .ZN(n4732) );
  OAI21_X1 U6519 ( .B1(n4732), .B2(n4736), .A(n4733), .ZN(n6077) );
  INV_X2 U6520 ( .A(n6695), .ZN(n6089) );
  NOR2_X2 U6521 ( .A1(n4747), .A2(n4746), .ZN(n5888) );
  NAND3_X1 U6522 ( .A1(n5878), .A2(n5895), .A3(n5880), .ZN(n4746) );
  NAND4_X1 U6523 ( .A1(n5984), .A2(n5893), .A3(n4965), .A4(n5879), .ZN(n4747)
         );
  AND2_X2 U6524 ( .A1(n5119), .A2(n5168), .ZN(n5218) );
  AND3_X2 U6525 ( .A1(n4751), .A2(n5781), .A3(n5166), .ZN(n5168) );
  AND2_X2 U6526 ( .A1(n5517), .A2(n5518), .ZN(n5166) );
  OAI21_X1 U6527 ( .B1(n9802), .B2(n4755), .A(n4752), .ZN(n9728) );
  AND2_X1 U6528 ( .A1(n5103), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U6529 ( .A1(n4756), .A2(n4754), .ZN(n5818) );
  NAND2_X1 U6530 ( .A1(n4755), .A2(n5103), .ZN(n4754) );
  NAND3_X1 U6531 ( .A1(n9802), .A2(n5103), .A3(n8330), .ZN(n4756) );
  NOR2_X2 U6532 ( .A1(n5104), .A2(n4759), .ZN(n4758) );
  AND2_X1 U6533 ( .A1(n4760), .A2(n8122), .ZN(n8243) );
  XNOR2_X1 U6534 ( .A(n6038), .B(n6010), .ZN(n7068) );
  NAND2_X1 U6535 ( .A1(n7202), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U6536 ( .A1(n8805), .A2(n8806), .ZN(n8804) );
  NAND2_X1 U6537 ( .A1(n4772), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U6538 ( .A1(n7591), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4773) );
  NAND2_X1 U6539 ( .A1(n6023), .A2(n8848), .ZN(n4786) );
  INV_X1 U6540 ( .A(n4786), .ZN(n4782) );
  NAND2_X1 U6541 ( .A1(n6023), .A2(n4779), .ZN(n4778) );
  XNOR2_X1 U6542 ( .A(n6024), .B(n6556), .ZN(n8871) );
  XNOR2_X1 U6543 ( .A(n6022), .B(n8848), .ZN(n8843) );
  NAND2_X1 U6544 ( .A1(n5796), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U6545 ( .A1(n7721), .A2(n4799), .ZN(n4795) );
  NAND2_X1 U6546 ( .A1(n4795), .A2(n4796), .ZN(n8126) );
  NAND2_X1 U6547 ( .A1(n7721), .A2(n7720), .ZN(n4798) );
  NAND2_X1 U6548 ( .A1(n4802), .A2(n4805), .ZN(n8137) );
  NOR2_X1 U6549 ( .A1(n4807), .A2(n4804), .ZN(n4803) );
  INV_X1 U6550 ( .A(n8140), .ZN(n4804) );
  NAND2_X1 U6551 ( .A1(n8127), .A2(n8128), .ZN(n8141) );
  NAND2_X1 U6552 ( .A1(n4810), .A2(n4811), .ZN(n8221) );
  NAND2_X1 U6553 ( .A1(n4816), .A2(n8772), .ZN(P2_U3296) );
  NAND3_X1 U6554 ( .A1(n4884), .A2(n4486), .A3(n4883), .ZN(n4817) );
  NAND3_X1 U6555 ( .A1(n4823), .A2(n4822), .A3(n4821), .ZN(n4820) );
  NAND2_X1 U6556 ( .A1(n6378), .A2(n4491), .ZN(n6643) );
  NAND2_X1 U6557 ( .A1(n6378), .A2(n6377), .ZN(n6620) );
  NAND2_X1 U6558 ( .A1(n6376), .A2(n4560), .ZN(n6604) );
  NAND2_X1 U6559 ( .A1(n6369), .A2(n4834), .ZN(n6497) );
  OAI21_X1 U6560 ( .B1(n5686), .B2(n4841), .A(n4837), .ZN(n9703) );
  NAND2_X1 U6561 ( .A1(n8079), .A2(n4851), .ZN(n4849) );
  NAND2_X1 U6562 ( .A1(n4849), .A2(n4850), .ZN(n9883) );
  NAND2_X1 U6563 ( .A1(n4854), .A2(n4855), .ZN(n9750) );
  NAND2_X1 U6564 ( .A1(n5509), .A2(n4546), .ZN(n9860) );
  OR2_X1 U6565 ( .A1(n9687), .A2(n9686), .ZN(n4861) );
  NAND2_X1 U6566 ( .A1(n4860), .A2(n4858), .ZN(n9664) );
  NAND2_X1 U6567 ( .A1(n9687), .A2(n4493), .ZN(n4860) );
  XNOR2_X2 U6568 ( .A(n4864), .B(n4863), .ZN(n8433) );
  NOR2_X1 U6569 ( .A1(n4880), .A2(n4870), .ZN(n4875) );
  NAND3_X1 U6570 ( .A1(n8730), .A2(n8963), .A3(n8731), .ZN(n4876) );
  OR2_X1 U6571 ( .A1(n8761), .A2(n8760), .ZN(n4882) );
  NAND2_X1 U6572 ( .A1(n4882), .A2(n4881), .ZN(n4884) );
  AOI21_X1 U6573 ( .B1(n8643), .B2(n8642), .A(n4886), .ZN(n8650) );
  NAND2_X1 U6574 ( .A1(n5940), .A2(n6038), .ZN(n4902) );
  NAND3_X1 U6575 ( .A1(n4911), .A2(n4910), .A3(n5966), .ZN(n5968) );
  NAND3_X1 U6576 ( .A1(n4912), .A2(n5963), .A3(n4490), .ZN(n4910) );
  INV_X1 U6577 ( .A(n5962), .ZN(n4913) );
  INV_X1 U6578 ( .A(n5994), .ZN(n8902) );
  NAND2_X1 U6579 ( .A1(n5994), .A2(n8917), .ZN(n4914) );
  NAND3_X1 U6580 ( .A1(n4918), .A2(P2_REG2_REG_15__SCAN_IN), .A3(n5983), .ZN(
        n8879) );
  NAND2_X1 U6581 ( .A1(n4918), .A2(n5983), .ZN(n8877) );
  INV_X1 U6582 ( .A(n5982), .ZN(n4919) );
  NAND2_X1 U6583 ( .A1(n5979), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6584 ( .A1(n5798), .A2(n7616), .ZN(n8236) );
  NAND2_X1 U6585 ( .A1(n5201), .A2(n4924), .ZN(n5204) );
  XNOR2_X1 U6586 ( .A(n4924), .B(n5299), .ZN(n5302) );
  NAND2_X1 U6587 ( .A1(n5763), .A2(n5762), .ZN(n6836) );
  NAND2_X1 U6588 ( .A1(n4925), .A2(n6834), .ZN(n6844) );
  NAND2_X1 U6589 ( .A1(n5763), .A2(n4926), .ZN(n4925) );
  INV_X1 U6590 ( .A(n5762), .ZN(n4927) );
  NAND2_X1 U6591 ( .A1(n5374), .A2(n5373), .ZN(n4929) );
  NAND2_X1 U6592 ( .A1(n4452), .A2(n5241), .ZN(n4934) );
  NAND3_X1 U6593 ( .A1(n5216), .A2(n5359), .A3(n5275), .ZN(n4932) );
  NAND3_X1 U6594 ( .A1(n4535), .A2(n8207), .A3(n8208), .ZN(n8211) );
  NAND2_X1 U6595 ( .A1(n5495), .A2(n4941), .ZN(n4937) );
  NAND2_X1 U6596 ( .A1(n5495), .A2(n5494), .ZN(n5514) );
  NAND2_X1 U6597 ( .A1(n5689), .A2(n4947), .ZN(n4943) );
  NAND2_X1 U6598 ( .A1(n4943), .A2(n4944), .ZN(n5729) );
  NAND2_X1 U6599 ( .A1(n5689), .A2(n5688), .ZN(n4946) );
  NAND2_X1 U6600 ( .A1(n5600), .A2(n4962), .ZN(n4959) );
  NAND2_X1 U6601 ( .A1(n4959), .A2(n4541), .ZN(n5652) );
  NAND2_X1 U6602 ( .A1(n9380), .A2(n4488), .ZN(n4974) );
  OAI21_X1 U6603 ( .B1(n9380), .B2(n9378), .A(n9377), .ZN(n9303) );
  CLKBUF_X1 U6604 ( .A(n4986), .Z(n4979) );
  OAI21_X2 U6605 ( .B1(n4986), .B2(n4981), .A(n4980), .ZN(n6776) );
  NAND2_X1 U6606 ( .A1(n7423), .A2(n4994), .ZN(n4993) );
  NAND2_X1 U6607 ( .A1(n5003), .A2(n4551), .ZN(n7356) );
  AND4_X2 U6608 ( .A1(n5888), .A2(n5100), .A3(n5955), .A4(n5909), .ZN(n6380)
         );
  INV_X1 U6609 ( .A(n5260), .ZN(n5006) );
  NAND2_X1 U6610 ( .A1(n5005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND3_X1 U6611 ( .A1(n5784), .A2(n5006), .A3(n5007), .ZN(n5005) );
  NAND2_X2 U6612 ( .A1(n5012), .A2(n6904), .ZN(n6326) );
  NAND2_X2 U6613 ( .A1(n7472), .A2(n7471), .ZN(n7558) );
  NAND2_X1 U6614 ( .A1(n5016), .A2(n5017), .ZN(n5019) );
  INV_X1 U6615 ( .A(n7096), .ZN(n5016) );
  NOR2_X1 U6616 ( .A1(n7110), .A2(n5138), .ZN(n7113) );
  NAND2_X1 U6617 ( .A1(n8056), .A2(n5026), .ZN(n8106) );
  NAND2_X1 U6618 ( .A1(n5033), .A2(n5034), .ZN(n8407) );
  NAND2_X1 U6619 ( .A1(n8424), .A2(n5038), .ZN(n5039) );
  OAI211_X1 U6620 ( .C1(n8424), .C2(n5040), .A(n8432), .B(n5039), .ZN(P2_U3160) );
  NAND2_X1 U6621 ( .A1(n8424), .A2(n8423), .ZN(n8447) );
  NAND3_X1 U6622 ( .A1(n5881), .A2(n5916), .A3(n4504), .ZN(n5051) );
  OR2_X1 U6623 ( .A1(n6430), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6624 ( .A1(n5062), .A2(n5066), .ZN(n6573) );
  NAND2_X1 U6625 ( .A1(n6555), .A2(n5063), .ZN(n5062) );
  OAI21_X1 U6626 ( .B1(n6513), .B2(n5074), .A(n5073), .ZN(n7912) );
  NAND2_X1 U6627 ( .A1(n5072), .A2(n5070), .ZN(n6545) );
  NAND2_X1 U6628 ( .A1(n6513), .A2(n5073), .ZN(n5072) );
  NAND2_X1 U6629 ( .A1(n6513), .A2(n6512), .ZN(n7578) );
  OR2_X1 U6630 ( .A1(n6524), .A2(n5080), .ZN(n5079) );
  INV_X1 U6631 ( .A(n6512), .ZN(n5080) );
  OR2_X1 U6632 ( .A1(n7993), .A2(n8783), .ZN(n5081) );
  NAND2_X1 U6633 ( .A1(n5084), .A2(n5082), .ZN(P2_U3204) );
  NOR2_X1 U6634 ( .A1(n6456), .A2(n5085), .ZN(n5089) );
  NAND2_X1 U6635 ( .A1(n7235), .A2(n6738), .ZN(n5090) );
  INV_X1 U6636 ( .A(n5089), .ZN(n5088) );
  NAND2_X1 U6637 ( .A1(n10105), .A2(n8595), .ZN(n6466) );
  NAND2_X1 U6638 ( .A1(n6660), .A2(n4542), .ZN(n5091) );
  NAND2_X1 U6639 ( .A1(n6660), .A2(n6659), .ZN(n6777) );
  NAND2_X1 U6640 ( .A1(n5091), .A2(n5092), .ZN(n6808) );
  NAND3_X1 U6641 ( .A1(n5096), .A2(n9011), .A3(n5097), .ZN(n6627) );
  NAND3_X1 U6642 ( .A1(n5888), .A2(n5955), .A3(n5141), .ZN(n5908) );
  XNOR2_X2 U6643 ( .A(n8376), .B(n5320), .ZN(n8234) );
  INV_X1 U6644 ( .A(n5816), .ZN(n5104) );
  NAND2_X1 U6645 ( .A1(n5820), .A2(n5108), .ZN(n6108) );
  NAND2_X1 U6646 ( .A1(n5820), .A2(n8272), .ZN(n9683) );
  NAND2_X1 U6647 ( .A1(n6108), .A2(n8262), .ZN(n5821) );
  NAND3_X1 U6648 ( .A1(n5112), .A2(n5166), .A3(n5113), .ZN(n5776) );
  INV_X1 U6649 ( .A(n5168), .ZN(n5777) );
  INV_X1 U6650 ( .A(n5118), .ZN(n7726) );
  INV_X1 U6651 ( .A(n5169), .ZN(n5120) );
  NAND2_X1 U6652 ( .A1(n5833), .A2(n5123), .ZN(n9808) );
  INV_X1 U6653 ( .A(n5833), .ZN(n9864) );
  INV_X1 U6654 ( .A(n9867), .ZN(n5126) );
  NOR2_X1 U6655 ( .A1(n9735), .A2(n5128), .ZN(n5131) );
  OAI21_X1 U6656 ( .B1(n4464), .B2(n6866), .A(n5300), .ZN(n5301) );
  AND3_X1 U6657 ( .A1(n8208), .A2(n5147), .A3(n8291), .ZN(n8295) );
  AND2_X1 U6658 ( .A1(n5953), .A2(n7162), .ZN(n5954) );
  XNOR2_X1 U6659 ( .A(n5729), .B(n5728), .ZN(n8099) );
  XNOR2_X1 U6660 ( .A(n5759), .B(n5758), .ZN(n8379) );
  AND2_X2 U6661 ( .A1(n8433), .A2(n8369), .ZN(n6422) );
  OAI211_X1 U6662 ( .C1(n6711), .C2(n6710), .A(n6709), .B(n6708), .ZN(n6714)
         );
  INV_X1 U6663 ( .A(n6709), .ZN(n8100) );
  CLKBUF_X1 U6664 ( .A(n7431), .Z(n7434) );
  OR2_X1 U6665 ( .A1(n6453), .A2(n6898), .ZN(n6419) );
  AND2_X1 U6666 ( .A1(n6816), .A2(n6696), .ZN(n7017) );
  CLKBUF_X1 U6667 ( .A(n7402), .Z(n10131) );
  OAI21_X1 U6668 ( .B1(n5748), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n5211), .ZN(
        n5214) );
  NAND2_X1 U6669 ( .A1(n5748), .A2(n6875), .ZN(n5211) );
  NAND2_X1 U6670 ( .A1(n5748), .A2(n6878), .ZN(n5189) );
  AND2_X1 U6671 ( .A1(n7420), .A2(n7419), .ZN(n7638) );
  AND2_X1 U6672 ( .A1(n6777), .A2(n8731), .ZN(n6778) );
  NAND2_X1 U6673 ( .A1(n6102), .A2(n10077), .ZN(n5876) );
  AND2_X2 U6674 ( .A1(n5181), .A2(n5176), .ZN(n5349) );
  NAND2_X1 U6675 ( .A1(n4561), .A2(n10067), .ZN(n7371) );
  INV_X1 U6676 ( .A(n5835), .ZN(n6111) );
  NAND2_X1 U6677 ( .A1(n5835), .A2(n5837), .ZN(n9651) );
  INV_X1 U6678 ( .A(n7371), .ZN(n5832) );
  NAND2_X1 U6679 ( .A1(n5832), .A2(n5280), .ZN(n7508) );
  XNOR2_X1 U6680 ( .A(n6125), .B(n6329), .ZN(n6134) );
  NAND2_X1 U6681 ( .A1(n9244), .A2(n6847), .ZN(n6851) );
  INV_X1 U6682 ( .A(n10017), .ZN(n6861) );
  AND2_X2 U6683 ( .A1(n6101), .A2(n6100), .ZN(n10074) );
  INV_X1 U6684 ( .A(n9961), .ZN(n9940) );
  AND2_X2 U6685 ( .A1(n6101), .A2(n5874), .ZN(n10077) );
  AND2_X1 U6686 ( .A1(n7988), .A2(n7866), .ZN(n5137) );
  AND2_X1 U6687 ( .A1(n7109), .A2(n8791), .ZN(n5138) );
  AND2_X1 U6688 ( .A1(n5146), .A2(n6825), .ZN(n5139) );
  NAND2_X1 U6689 ( .A1(n5780), .A2(n7798), .ZN(n8297) );
  OR2_X1 U6690 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5140) );
  NAND2_X2 U6691 ( .A1(n6771), .A2(n10123), .ZN(n10141) );
  INV_X1 U6692 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5188) );
  INV_X1 U6693 ( .A(n7255), .ZN(n5989) );
  INV_X1 U6694 ( .A(n8378), .ZN(n10024) );
  OR2_X1 U6695 ( .A1(n6487), .A2(n7537), .ZN(n5142) );
  AND4_X1 U6696 ( .A1(n5995), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n5143)
         );
  OR2_X1 U6697 ( .A1(n8704), .A2(n6697), .ZN(n5144) );
  AND2_X1 U6698 ( .A1(n8957), .A2(n8966), .ZN(n5145) );
  AND2_X1 U6699 ( .A1(n7185), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U6700 ( .A1(n9677), .A2(n9961), .ZN(n6114) );
  INV_X1 U6701 ( .A(n9211), .ZN(n6799) );
  AND2_X1 U6702 ( .A1(n8711), .A2(n6749), .ZN(n5149) );
  NAND2_X1 U6703 ( .A1(n9736), .A2(n9476), .ZN(n5150) );
  INV_X1 U6704 ( .A(n9729), .ZN(n5817) );
  NOR2_X1 U6705 ( .A1(n8275), .A2(n8193), .ZN(n5151) );
  AND2_X1 U6706 ( .A1(n9338), .A2(n9488), .ZN(n5152) );
  OR2_X1 U6707 ( .A1(n9338), .A2(n9488), .ZN(n5153) );
  INV_X1 U6708 ( .A(n8208), .ZN(n8225) );
  INV_X1 U6709 ( .A(n9094), .ZN(n10132) );
  NAND2_X1 U6710 ( .A1(n6687), .A2(n6789), .ZN(n9094) );
  AND2_X1 U6711 ( .A1(n8140), .A2(n8243), .ZN(n5154) );
  OR2_X1 U6712 ( .A1(n6760), .A2(n6734), .ZN(n10187) );
  INV_X1 U6713 ( .A(n9838), .ZN(n5808) );
  INV_X1 U6714 ( .A(n8451), .ZN(n8957) );
  INV_X1 U6715 ( .A(n8249), .ZN(n5466) );
  INV_X1 U6716 ( .A(n8297), .ZN(n8123) );
  NOR2_X1 U6717 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  AND2_X1 U6718 ( .A1(n9021), .A2(n8695), .ZN(n8696) );
  INV_X1 U6719 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5880) );
  NOR2_X1 U6720 ( .A1(n5837), .A2(n10066), .ZN(n5838) );
  OR2_X1 U6721 ( .A1(n7985), .A2(n8784), .ZN(n7866) );
  OR2_X1 U6722 ( .A1(n6504), .A2(n7756), .ZN(n5966) );
  NOR2_X1 U6723 ( .A1(n9305), .A2(n9304), .ZN(n6273) );
  AOI22_X1 U6724 ( .A1(n8214), .A2(n8213), .B1(n8287), .B2(n8212), .ZN(n8215)
         );
  INV_X1 U6725 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5170) );
  AND2_X1 U6726 ( .A1(n8798), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U6727 ( .A1(n10118), .A2(n7403), .ZN(n7402) );
  INV_X1 U6728 ( .A(n8598), .ZN(n6476) );
  OAI22_X1 U6729 ( .A1(n6124), .A2(n4455), .B1(n4588), .B2(n6317), .ZN(n6125)
         );
  OR2_X1 U6730 ( .A1(n6245), .A2(n9451), .ZN(n6250) );
  INV_X1 U6731 ( .A(n8217), .ZN(n8218) );
  INV_X1 U6732 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5233) );
  INV_X1 U6733 ( .A(n8326), .ZN(n5807) );
  AND2_X1 U6734 ( .A1(n7714), .A2(n7715), .ZN(n5371) );
  NAND2_X1 U6735 ( .A1(n5317), .A2(n10055), .ZN(n5319) );
  INV_X1 U6736 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5172) );
  INV_X1 U6737 ( .A(SI_24_), .ZN(n10292) );
  INV_X1 U6738 ( .A(SI_19_), .ZN(n10487) );
  NOR2_X1 U6739 ( .A1(n5533), .A2(SI_16_), .ZN(n5553) );
  INV_X1 U6740 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5225) );
  INV_X1 U6741 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5909) );
  NOR2_X1 U6742 ( .A1(n8975), .A2(n10125), .ZN(n6780) );
  AND2_X1 U6743 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  NOR2_X1 U6744 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  INV_X1 U6745 ( .A(n9789), .ZN(n9786) );
  INV_X1 U6746 ( .A(n9663), .ZN(n8206) );
  INV_X1 U6747 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5658) );
  AND2_X1 U6748 ( .A1(n5389), .A2(n7723), .ZN(n5390) );
  INV_X1 U6749 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U6750 ( .A1(n8104), .A2(n8111), .ZN(n8105) );
  INV_X1 U6751 ( .A(n9032), .ZN(n9000) );
  NAND2_X1 U6752 ( .A1(n7145), .A2(n7146), .ZN(n7147) );
  INV_X1 U6753 ( .A(n4507), .ZN(n7086) );
  INV_X1 U6754 ( .A(n8780), .ZN(n9103) );
  AND2_X1 U6755 ( .A1(n10102), .A2(n8655), .ZN(n8596) );
  NOR2_X1 U6756 ( .A1(n6884), .A2(n6793), .ZN(n6787) );
  CLKBUF_X1 U6757 ( .A(n9245), .Z(n9249) );
  AOI21_X1 U6758 ( .B1(n5916), .B2(n5143), .A(n5055), .ZN(n5896) );
  AND2_X1 U6759 ( .A1(n9436), .A2(n9437), .ZN(n6316) );
  INV_X1 U6760 ( .A(n8343), .ZN(n8291) );
  OR2_X1 U6761 ( .A1(n9441), .A2(n5721), .ZN(n5726) );
  INV_X1 U6762 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7481) );
  AND2_X1 U6763 ( .A1(n8228), .A2(n9771), .ZN(n9789) );
  INV_X1 U6764 ( .A(n9426), .ZN(n9455) );
  AND2_X1 U6765 ( .A1(n7798), .A2(n8303), .ZN(n6345) );
  INV_X1 U6766 ( .A(n9885), .ZN(n9843) );
  NAND2_X1 U6767 ( .A1(n5849), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U6768 ( .A(n5579), .B(SI_18_), .ZN(n5578) );
  INV_X1 U6769 ( .A(n8563), .ZN(n8539) );
  AND2_X1 U6770 ( .A1(n7020), .A2(n7007), .ZN(n8561) );
  NAND2_X1 U6771 ( .A1(n7006), .A2(n10123), .ZN(n8553) );
  AND4_X1 U6772 ( .A1(n6543), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(n8111)
         );
  INV_X1 U6773 ( .A(n10095), .ZN(n8883) );
  INV_X1 U6774 ( .A(n7207), .ZN(n10099) );
  AND2_X1 U6775 ( .A1(n7141), .A2(n8766), .ZN(n10092) );
  OAI21_X1 U6776 ( .B1(n9172), .B2(n10115), .A(n6772), .ZN(n6773) );
  INV_X1 U6777 ( .A(n10123), .ZN(n9096) );
  INV_X1 U6778 ( .A(n9135), .ZN(n9154) );
  INV_X1 U6779 ( .A(n8996), .ZN(n8998) );
  AND2_X1 U6780 ( .A1(n8762), .A2(n7797), .ZN(n10151) );
  NAND2_X1 U6781 ( .A1(n10124), .A2(n10174), .ZN(n10162) );
  NAND2_X1 U6782 ( .A1(n5891), .A2(n5890), .ZN(n6767) );
  XNOR2_X1 U6783 ( .A(n5903), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U6784 ( .A(n5965), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U6785 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  INV_X1 U6786 ( .A(n9460), .ZN(n9444) );
  OR2_X1 U6787 ( .A1(n7317), .A2(n6348), .ZN(n9829) );
  INV_X1 U6788 ( .A(n9462), .ZN(n9442) );
  INV_X1 U6789 ( .A(n9412), .ZN(n9465) );
  AOI21_X1 U6790 ( .B1(n9675), .B2(n5767), .A(n5757), .ZN(n9266) );
  INV_X1 U6791 ( .A(n5767), .ZN(n5721) );
  AND4_X1 U6792 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n9456)
         );
  INV_X1 U6793 ( .A(n9636), .ZN(n9592) );
  INV_X1 U6794 ( .A(n9633), .ZN(n9632) );
  AND2_X1 U6795 ( .A1(n8178), .A2(n8330), .ZN(n9804) );
  NAND2_X1 U6796 ( .A1(n5823), .A2(n8296), .ZN(n9878) );
  INV_X1 U6797 ( .A(n9891), .ZN(n10054) );
  INV_X1 U6798 ( .A(n8444), .ZN(n10055) );
  NAND2_X1 U6799 ( .A1(n5873), .A2(n5852), .ZN(n6914) );
  XNOR2_X1 U6800 ( .A(n5850), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7999) );
  AND2_X1 U6801 ( .A1(n5416), .A2(n5399), .ZN(n7032) );
  INV_X1 U6802 ( .A(n8565), .ZN(n8063) );
  AND2_X1 U6803 ( .A1(n7004), .A2(n7003), .ZN(n8555) );
  INV_X1 U6804 ( .A(n8527), .ZN(n9043) );
  OR2_X1 U6805 ( .A1(n6027), .A2(P2_U3151), .ZN(n8929) );
  OR2_X1 U6806 ( .A1(P2_U3150), .A2(n6028), .ZN(n7207) );
  INV_X1 U6807 ( .A(n10092), .ZN(n8939) );
  INV_X1 U6808 ( .A(n6773), .ZN(n6774) );
  OR2_X1 U6809 ( .A1(n6997), .A2(n6768), .ZN(n10123) );
  OR2_X1 U6810 ( .A1(n6771), .A2(n10122), .ZN(n10111) );
  NAND2_X1 U6811 ( .A1(n10189), .A2(n10162), .ZN(n9147) );
  NAND2_X1 U6812 ( .A1(n10189), .A2(n10161), .ZN(n9135) );
  INV_X2 U6813 ( .A(n10187), .ZN(n10189) );
  INV_X1 U6814 ( .A(n6823), .ZN(n6824) );
  NAND2_X1 U6815 ( .A1(n10178), .A2(n10162), .ZN(n9234) );
  NAND2_X1 U6816 ( .A1(n10178), .A2(n10161), .ZN(n9211) );
  AND2_X1 U6817 ( .A1(n6797), .A2(n6796), .ZN(n10180) );
  INV_X2 U6818 ( .A(n10180), .ZN(n10178) );
  AND2_X1 U6819 ( .A1(n6892), .A2(n6714), .ZN(n6918) );
  INV_X1 U6820 ( .A(n6918), .ZN(n6913) );
  INV_X1 U6821 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10429) );
  INV_X1 U6822 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6960) );
  INV_X1 U6823 ( .A(n9643), .ZN(n10038) );
  AOI21_X1 U6824 ( .B1(n9265), .B2(n6363), .A(n6362), .ZN(n6364) );
  AND2_X1 U6825 ( .A1(n6349), .A2(n9829), .ZN(n9412) );
  INV_X1 U6826 ( .A(n9434), .ZN(n9467) );
  INV_X1 U6827 ( .A(n9359), .ZN(n9474) );
  OR2_X1 U6828 ( .A1(n6936), .A2(n6935), .ZN(n10041) );
  OR2_X1 U6829 ( .A1(n6936), .A2(n6907), .ZN(n9643) );
  OR2_X1 U6830 ( .A1(n10063), .A2(n7458), .ZN(n10053) );
  INV_X1 U6831 ( .A(n10049), .ZN(n9852) );
  NAND2_X1 U6832 ( .A1(n4655), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5875) );
  INV_X1 U6833 ( .A(n9690), .ZN(n9975) );
  INV_X1 U6834 ( .A(n7821), .ZN(n8052) );
  INV_X1 U6835 ( .A(n10074), .ZN(n10072) );
  NAND2_X1 U6836 ( .A1(n10020), .A2(n6914), .ZN(n10223) );
  INV_X1 U6837 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10440) );
  INV_X1 U6838 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10457) );
  INV_X2 U6839 ( .A(n8929), .ZN(P2_U3893) );
  INV_X1 U6840 ( .A(n9469), .ZN(P1_U3973) );
  OAI21_X1 U6841 ( .B1(n6830), .B2(n4655), .A(n6117), .ZN(P1_U3550) );
  NOR2_X1 U6842 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5161) );
  NOR2_X1 U6843 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5160) );
  NOR2_X1 U6844 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5159) );
  NOR2_X1 U6845 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5162) );
  NOR2_X1 U6846 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5163) );
  NOR2_X2 U6847 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5224) );
  NOR3_X1 U6848 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6849 ( .A1(n4458), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6850 ( .A1(n4456), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5184) );
  INV_X1 U6851 ( .A(n5175), .ZN(n5181) );
  INV_X1 U6852 ( .A(n5265), .ZN(n5177) );
  NAND2_X1 U6853 ( .A1(n5177), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5267) );
  INV_X1 U6854 ( .A(n5267), .ZN(n5178) );
  NAND2_X1 U6855 ( .A1(n5178), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5234) );
  INV_X1 U6856 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6857 ( .A1(n5267), .A2(n5179), .ZN(n5180) );
  AND2_X1 U6858 ( .A1(n5234), .A2(n5180), .ZN(n7691) );
  NAND2_X1 U6859 ( .A1(n5349), .A2(n7691), .ZN(n5183) );
  NAND2_X1 U6860 ( .A1(n5325), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5182) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U6862 ( .A1(n5190), .A2(n5189), .ZN(n5205) );
  NAND2_X1 U6863 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5191) );
  INV_X1 U6864 ( .A(SI_1_), .ZN(n5194) );
  INV_X1 U6865 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6882) );
  AOI21_X1 U6866 ( .B1(n5191), .B2(n5194), .A(n6882), .ZN(n5193) );
  NOR2_X1 U6867 ( .A1(n5191), .A2(n5194), .ZN(n5192) );
  OAI21_X1 U6868 ( .B1(n5193), .B2(n5192), .A(n5748), .ZN(n5200) );
  NAND2_X1 U6869 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6870 ( .A1(n5195), .A2(n5194), .ZN(n5197) );
  INV_X1 U6871 ( .A(n5195), .ZN(n5196) );
  AOI22_X1 U6872 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n5197), .B1(n5196), .B2(
        SI_1_), .ZN(n5198) );
  OR2_X1 U6873 ( .A1(n5748), .A2(n5198), .ZN(n5199) );
  INV_X1 U6874 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U6875 ( .A1(n5748), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5300) );
  INV_X1 U6876 ( .A(SI_2_), .ZN(n5299) );
  OAI211_X1 U6877 ( .C1(n5748), .C2(n6866), .A(n5300), .B(n5299), .ZN(n5201)
         );
  INV_X1 U6878 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U6879 ( .A1(n5748), .A2(n6897), .ZN(n5202) );
  OAI211_X1 U6880 ( .C1(n5748), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5202), .B(
        SI_2_), .ZN(n5203) );
  NAND2_X1 U6881 ( .A1(n5204), .A2(n5203), .ZN(n5334) );
  NAND2_X1 U6882 ( .A1(n5335), .A2(n5334), .ZN(n5208) );
  INV_X1 U6883 ( .A(n5205), .ZN(n5206) );
  NAND2_X1 U6884 ( .A1(n5206), .A2(SI_3_), .ZN(n5207) );
  INV_X1 U6885 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6867) );
  INV_X1 U6886 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6880) );
  MUX2_X1 U6887 ( .A(n6867), .B(n6880), .S(n5748), .Z(n5209) );
  XNOR2_X1 U6888 ( .A(n5209), .B(SI_4_), .ZN(n5256) );
  INV_X1 U6889 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6890 ( .A1(n5210), .A2(SI_4_), .ZN(n5274) );
  INV_X1 U6891 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6869) );
  INV_X1 U6892 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6875) );
  INV_X1 U6893 ( .A(n5214), .ZN(n5212) );
  NAND2_X1 U6894 ( .A1(n5212), .A2(SI_5_), .ZN(n5213) );
  AND2_X1 U6895 ( .A1(n5213), .A2(n5274), .ZN(n5216) );
  INV_X1 U6896 ( .A(n5213), .ZN(n5215) );
  XNOR2_X1 U6897 ( .A(n5214), .B(SI_5_), .ZN(n5276) );
  MUX2_X1 U6898 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5748), .Z(n5242) );
  OAI21_X1 U6899 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6900 ( .A1(n5845), .A2(n5222), .ZN(n5223) );
  INV_X2 U6901 ( .A(n5336), .ZN(n6847) );
  INV_X1 U6902 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10264) );
  OR2_X1 U6903 ( .A1(n4469), .A2(n10264), .ZN(n5231) );
  NAND2_X1 U6904 ( .A1(n5303), .A2(n5224), .ZN(n5258) );
  NAND2_X1 U6905 ( .A1(n4494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5228) );
  INV_X1 U6906 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6907 ( .A1(n5228), .A2(n5227), .ZN(n5244) );
  OR2_X1 U6908 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND2_X1 U6909 ( .A1(n4465), .A2(n6948), .ZN(n5230) );
  NAND2_X1 U6910 ( .A1(n5232), .A2(n7516), .ZN(n7611) );
  INV_X1 U6911 ( .A(n7611), .ZN(n5248) );
  NAND2_X1 U6912 ( .A1(n4458), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6913 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  AND2_X1 U6914 ( .A1(n5346), .A2(n5235), .ZN(n7570) );
  NAND2_X1 U6915 ( .A1(n5767), .A2(n7570), .ZN(n5238) );
  NAND2_X1 U6916 ( .A1(n4457), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6917 ( .A1(n5325), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5236) );
  INV_X1 U6918 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6919 ( .A1(n5242), .A2(SI_6_), .ZN(n5356) );
  NAND2_X1 U6920 ( .A1(n5360), .A2(n5356), .ZN(n5243) );
  MUX2_X1 U6921 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4464), .Z(n5355) );
  XNOR2_X1 U6922 ( .A(n5243), .B(n5358), .ZN(n6893) );
  NAND2_X1 U6923 ( .A1(n6893), .A2(n6847), .ZN(n5247) );
  NAND2_X1 U6924 ( .A1(n5244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5245) );
  XNOR2_X1 U6925 ( .A(n5245), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9598) );
  AOI22_X1 U6926 ( .A1(n5589), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4465), .B2(
        n9598), .ZN(n5246) );
  INV_X1 U6927 ( .A(n5249), .ZN(n5344) );
  NAND2_X1 U6928 ( .A1(n4457), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5255) );
  INV_X1 U6929 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10043) );
  INV_X1 U6930 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6931 ( .A1(n10043), .A2(n5250), .ZN(n5251) );
  AND2_X1 U6932 ( .A1(n5251), .A2(n5265), .ZN(n7547) );
  NAND2_X1 U6933 ( .A1(n5349), .A2(n7547), .ZN(n5254) );
  NAND2_X1 U6934 ( .A1(n5325), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6935 ( .A1(n4458), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5252) );
  INV_X1 U6936 ( .A(n7260), .ZN(n9496) );
  XNOR2_X1 U6937 ( .A(n5257), .B(n5256), .ZN(n6879) );
  OR2_X1 U6938 ( .A1(n5336), .A2(n6879), .ZN(n5264) );
  OR2_X1 U6939 ( .A1(n4470), .A2(n6880), .ZN(n5263) );
  NAND2_X1 U6940 ( .A1(n5258), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5259) );
  MUX2_X1 U6941 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5259), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5261) );
  AND2_X1 U6942 ( .A1(n5261), .A2(n5260), .ZN(n9547) );
  NAND2_X1 U6943 ( .A1(n4459), .A2(n9547), .ZN(n5262) );
  NAND2_X1 U6944 ( .A1(n7260), .A2(n7548), .ZN(n5795) );
  NAND2_X1 U6945 ( .A1(n7260), .A2(n10067), .ZN(n7368) );
  INV_X1 U6946 ( .A(n7368), .ZN(n5281) );
  NAND2_X1 U6947 ( .A1(n4458), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6948 ( .A1(n4456), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5270) );
  INV_X1 U6949 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U6950 ( .A1(n5265), .A2(n10267), .ZN(n5266) );
  AND2_X1 U6951 ( .A1(n5267), .A2(n5266), .ZN(n7603) );
  NAND2_X1 U6952 ( .A1(n5349), .A2(n7603), .ZN(n5269) );
  NAND2_X1 U6953 ( .A1(n5325), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6954 ( .A1(n5260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5272) );
  MUX2_X1 U6955 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5272), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5273) );
  NAND2_X1 U6956 ( .A1(n5273), .A2(n4494), .ZN(n9561) );
  OR2_X1 U6957 ( .A1(n4469), .A2(n6875), .ZN(n5279) );
  NAND2_X1 U6958 ( .A1(n5275), .A2(n5274), .ZN(n5277) );
  XNOR2_X1 U6959 ( .A(n5277), .B(n5276), .ZN(n6874) );
  OR2_X1 U6960 ( .A1(n5336), .A2(n6874), .ZN(n5278) );
  NAND2_X1 U6961 ( .A1(n7510), .A2(n7496), .ZN(n5797) );
  OAI21_X1 U6962 ( .B1(n8229), .B2(n5281), .A(n7367), .ZN(n5282) );
  INV_X1 U6963 ( .A(n5282), .ZN(n5341) );
  NAND2_X1 U6964 ( .A1(n5326), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6965 ( .A1(n5349), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6966 ( .A1(n5325), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6967 ( .A1(n5350), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5283) );
  AND4_X4 U6968 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n6124)
         );
  OR2_X1 U6969 ( .A1(n4468), .A2(n6882), .ZN(n5294) );
  NAND2_X1 U6970 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5287) );
  NAND2_X1 U6971 ( .A1(n5588), .A2(n9502), .ZN(n5293) );
  XNOR2_X1 U6972 ( .A(n5288), .B(SI_1_), .ZN(n5291) );
  MUX2_X1 U6973 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5748), .Z(n5289) );
  NAND2_X1 U6974 ( .A1(n5289), .A2(SI_0_), .ZN(n5290) );
  XNOR2_X1 U6975 ( .A(n5291), .B(n5290), .ZN(n6881) );
  OR2_X1 U6976 ( .A1(n5336), .A2(n6881), .ZN(n5292) );
  NAND2_X1 U6977 ( .A1(n5325), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6978 ( .A1(n5350), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6979 ( .A1(n5326), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6980 ( .A1(n7246), .A2(n9498), .ZN(n5310) );
  XNOR2_X1 U6981 ( .A(n5302), .B(n5301), .ZN(n6898) );
  OR2_X1 U6982 ( .A1(n5336), .A2(n6898), .ZN(n5309) );
  INV_X1 U6983 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6984 ( .A1(n5304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5306) );
  INV_X1 U6985 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6986 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  NAND2_X1 U6987 ( .A1(n5306), .A2(n5305), .ZN(n5331) );
  NAND2_X1 U6988 ( .A1(n5588), .A2(n9520), .ZN(n5308) );
  NAND2_X1 U6989 ( .A1(n5310), .A2(n8376), .ZN(n5324) );
  NAND2_X1 U6990 ( .A1(n5349), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6991 ( .A1(n5326), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6992 ( .A1(n5350), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5311) );
  NAND4_X2 U6993 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n7323)
         );
  NAND2_X1 U6994 ( .A1(n6873), .A2(SI_0_), .ZN(n5315) );
  XNOR2_X1 U6995 ( .A(n5315), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U6996 ( .A1(n7323), .A2(n7452), .ZN(n7319) );
  INV_X1 U6997 ( .A(n6124), .ZN(n5317) );
  NAND2_X1 U6998 ( .A1(n9498), .A2(n7460), .ZN(n5318) );
  NAND3_X1 U6999 ( .A1(n7319), .A2(n5319), .A3(n5318), .ZN(n5323) );
  INV_X1 U7000 ( .A(n7246), .ZN(n5321) );
  NAND2_X1 U7001 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  NAND3_X1 U7002 ( .A1(n5324), .A2(n5323), .A3(n5322), .ZN(n7295) );
  NAND2_X1 U7003 ( .A1(n5349), .A2(n10043), .ZN(n5330) );
  NAND2_X1 U7004 ( .A1(n4456), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U7005 ( .A1(n5325), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U7006 ( .A1(n4458), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U7007 ( .A1(n5331), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5333) );
  INV_X1 U7008 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U7009 ( .A(n5333), .B(n5332), .ZN(n9535) );
  OR2_X1 U7010 ( .A1(n4470), .A2(n6878), .ZN(n5338) );
  XNOR2_X1 U7011 ( .A(n5335), .B(n5334), .ZN(n6877) );
  OR2_X1 U7012 ( .A1(n5336), .A2(n6877), .ZN(n5337) );
  OAI211_X1 U7013 ( .C1(n5316), .C2(n9535), .A(n5338), .B(n5337), .ZN(n7301)
         );
  NAND2_X1 U7014 ( .A1(n7250), .A2(n7301), .ZN(n5792) );
  INV_X1 U7015 ( .A(n7250), .ZN(n9497) );
  NAND2_X1 U7016 ( .A1(n9497), .A2(n10046), .ZN(n5793) );
  NAND2_X1 U7017 ( .A1(n5792), .A2(n5793), .ZN(n8230) );
  NAND2_X1 U7018 ( .A1(n7295), .A2(n8230), .ZN(n7294) );
  NAND2_X1 U7019 ( .A1(n7250), .A2(n10046), .ZN(n7366) );
  AND2_X1 U7020 ( .A1(n7368), .A2(n7366), .ZN(n5339) );
  NAND2_X1 U7021 ( .A1(n7294), .A2(n5339), .ZN(n5340) );
  NAND2_X1 U7022 ( .A1(n5341), .A2(n5340), .ZN(n7369) );
  NAND2_X1 U7023 ( .A1(n7510), .A2(n5280), .ZN(n7505) );
  AND2_X1 U7024 ( .A1(n7611), .A2(n7505), .ZN(n5342) );
  NAND2_X1 U7025 ( .A1(n7369), .A2(n5342), .ZN(n5343) );
  NAND2_X1 U7026 ( .A1(n5344), .A2(n5343), .ZN(n7613) );
  NAND2_X1 U7027 ( .A1(n7511), .A2(n4466), .ZN(n7714) );
  NAND2_X1 U7028 ( .A1(n4458), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U7029 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  NAND2_X1 U7030 ( .A1(n5383), .A2(n5347), .ZN(n9318) );
  INV_X1 U7031 ( .A(n9318), .ZN(n5348) );
  NAND2_X1 U7032 ( .A1(n5349), .A2(n5348), .ZN(n5353) );
  NAND2_X1 U7033 ( .A1(n4457), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U7034 ( .A1(n5325), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U7035 ( .A1(n5355), .A2(SI_7_), .ZN(n5357) );
  AND2_X1 U7036 ( .A1(n5356), .A2(n5357), .ZN(n5359) );
  INV_X1 U7037 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6891) );
  INV_X1 U7038 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6889) );
  INV_X1 U7039 ( .A(SI_8_), .ZN(n5361) );
  NAND2_X1 U7040 ( .A1(n5362), .A2(n5361), .ZN(n5373) );
  INV_X1 U7041 ( .A(n5362), .ZN(n5363) );
  NAND2_X1 U7042 ( .A1(n5363), .A2(SI_8_), .ZN(n5364) );
  NAND2_X1 U7043 ( .A1(n5373), .A2(n5364), .ZN(n5374) );
  NAND2_X1 U7044 ( .A1(n6888), .A2(n6847), .ZN(n5370) );
  NOR2_X1 U7045 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5365) );
  INV_X1 U7046 ( .A(n5519), .ZN(n5366) );
  NAND2_X1 U7047 ( .A1(n5366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5367) );
  MUX2_X1 U7048 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5367), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5369) );
  NAND2_X1 U7049 ( .A1(n5519), .A2(n5368), .ZN(n5397) );
  NAND2_X1 U7050 ( .A1(n5369), .A2(n5397), .ZN(n6940) );
  INV_X1 U7051 ( .A(n6940), .ZN(n6975) );
  OR2_X1 U7052 ( .A1(n9492), .A2(n9325), .ZN(n7715) );
  NAND2_X1 U7053 ( .A1(n7613), .A2(n5371), .ZN(n5391) );
  NAND2_X1 U7054 ( .A1(n7740), .A2(n7715), .ZN(n5389) );
  INV_X1 U7055 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6896) );
  MUX2_X1 U7056 ( .A(n6896), .B(n10265), .S(n6873), .Z(n5376) );
  INV_X1 U7057 ( .A(SI_9_), .ZN(n5375) );
  NAND2_X1 U7058 ( .A1(n5376), .A2(n5375), .ZN(n5395) );
  INV_X1 U7059 ( .A(n5376), .ZN(n5377) );
  NAND2_X1 U7060 ( .A1(n5377), .A2(SI_9_), .ZN(n5378) );
  AND2_X2 U7061 ( .A1(n5395), .A2(n5378), .ZN(n5393) );
  XNOR2_X1 U7062 ( .A(n5394), .B(n5393), .ZN(n6895) );
  NAND2_X1 U7063 ( .A1(n6895), .A2(n6847), .ZN(n5381) );
  NAND2_X1 U7064 ( .A1(n5397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5379) );
  XNOR2_X1 U7065 ( .A(n5379), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7029) );
  AOI22_X1 U7066 ( .A1(n5589), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4465), .B2(
        n7029), .ZN(n5380) );
  NAND2_X1 U7067 ( .A1(n5381), .A2(n5380), .ZN(n7727) );
  NAND2_X1 U7068 ( .A1(n4457), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U7069 ( .A1(n4458), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U7070 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  AND2_X1 U7071 ( .A1(n5422), .A2(n5384), .ZN(n7949) );
  NAND2_X1 U7072 ( .A1(n5767), .A2(n7949), .ZN(n5386) );
  NAND2_X1 U7073 ( .A1(n5325), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5385) );
  OR2_X1 U7074 ( .A1(n7727), .A2(n7741), .ZN(n8129) );
  NAND2_X1 U7075 ( .A1(n7727), .A2(n7741), .ZN(n8140) );
  NAND2_X1 U7076 ( .A1(n8129), .A2(n8140), .ZN(n7723) );
  NAND2_X1 U7077 ( .A1(n5391), .A2(n5390), .ZN(n7718) );
  INV_X1 U7078 ( .A(n7741), .ZN(n9491) );
  OR2_X1 U7079 ( .A1(n7727), .A2(n9491), .ZN(n5392) );
  MUX2_X1 U7080 ( .A(n6910), .B(n10266), .S(n6873), .Z(n5408) );
  XNOR2_X1 U7081 ( .A(n5408), .B(SI_10_), .ZN(n5407) );
  XNOR2_X1 U7082 ( .A(n5412), .B(n5407), .ZN(n6909) );
  NAND2_X1 U7083 ( .A1(n6909), .A2(n6847), .ZN(n5401) );
  NAND2_X1 U7084 ( .A1(n5438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5398) );
  INV_X1 U7085 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7086 ( .A1(n5398), .A2(n5436), .ZN(n5416) );
  OR2_X1 U7087 ( .A1(n5398), .A2(n5436), .ZN(n5399) );
  AOI22_X1 U7088 ( .A1(n5589), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4465), .B2(
        n7032), .ZN(n5400) );
  NAND2_X1 U7089 ( .A1(n4458), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U7090 ( .A1(n4456), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5404) );
  XNOR2_X1 U7091 ( .A(n5422), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U7092 ( .A1(n5767), .A2(n7708), .ZN(n5403) );
  NAND2_X1 U7093 ( .A1(n5325), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5402) );
  OR2_X1 U7094 ( .A1(n7968), .A2(n7728), .ZN(n8311) );
  NAND2_X1 U7095 ( .A1(n7968), .A2(n7728), .ZN(n8130) );
  NAND2_X1 U7096 ( .A1(n8311), .A2(n8130), .ZN(n7697) );
  INV_X1 U7097 ( .A(n7728), .ZN(n9490) );
  OR2_X1 U7098 ( .A1(n7968), .A2(n9490), .ZN(n5406) );
  INV_X1 U7099 ( .A(n5407), .ZN(n5411) );
  INV_X1 U7100 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U7101 ( .A1(n5409), .A2(SI_10_), .ZN(n5410) );
  INV_X1 U7102 ( .A(n5413), .ZN(n5414) );
  NAND2_X1 U7103 ( .A1(n5414), .A2(SI_11_), .ZN(n5415) );
  NAND2_X1 U7104 ( .A1(n5432), .A2(n5415), .ZN(n5433) );
  XNOR2_X1 U7105 ( .A(n5434), .B(n5433), .ZN(n6959) );
  NAND2_X1 U7106 ( .A1(n6959), .A2(n6847), .ZN(n5419) );
  NAND2_X1 U7107 ( .A1(n5416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5417) );
  XNOR2_X1 U7108 ( .A(n5417), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7128) );
  AOI22_X1 U7109 ( .A1(n5589), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4465), .B2(
        n7128), .ZN(n5418) );
  NAND2_X1 U7110 ( .A1(n4458), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5429) );
  INV_X1 U7111 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5421) );
  INV_X1 U7112 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U7113 ( .B1(n5422), .B2(n5421), .A(n5420), .ZN(n5425) );
  AND2_X1 U7114 ( .A1(n5425), .A2(n5447), .ZN(n8046) );
  NAND2_X1 U7115 ( .A1(n5767), .A2(n8046), .ZN(n5428) );
  NAND2_X1 U7116 ( .A1(n4457), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U7117 ( .A1(n5325), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5426) );
  NAND4_X1 U7118 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9489)
         );
  NAND2_X1 U7119 ( .A1(n7821), .A2(n9489), .ZN(n5430) );
  OR2_X1 U7120 ( .A1(n7821), .A2(n9489), .ZN(n5431) );
  MUX2_X1 U7121 ( .A(n6967), .B(n6968), .S(n5748), .Z(n5455) );
  XNOR2_X1 U7122 ( .A(n5455), .B(SI_12_), .ZN(n5454) );
  XNOR2_X1 U7123 ( .A(n5458), .B(n5454), .ZN(n6966) );
  NAND2_X1 U7124 ( .A1(n6966), .A2(n6847), .ZN(n5446) );
  INV_X1 U7125 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U7126 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NAND2_X1 U7127 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5439) );
  MUX2_X1 U7128 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5439), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5443) );
  INV_X1 U7129 ( .A(n5440), .ZN(n5442) );
  INV_X1 U7130 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7131 ( .A1(n5442), .A2(n5441), .ZN(n5473) );
  NAND2_X1 U7132 ( .A1(n5443), .A2(n5473), .ZN(n7222) );
  OAI22_X1 U7133 ( .A1(n4469), .A2(n6968), .B1(n5316), .B2(n7222), .ZN(n5444)
         );
  INV_X1 U7134 ( .A(n5444), .ZN(n5445) );
  NAND2_X1 U7135 ( .A1(n4458), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7136 ( .A1(n5447), .A2(n7133), .ZN(n5448) );
  AND2_X1 U7137 ( .A1(n5483), .A2(n5448), .ZN(n7977) );
  NAND2_X1 U7138 ( .A1(n5767), .A2(n7977), .ZN(n5451) );
  NAND2_X1 U7139 ( .A1(n4457), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5450) );
  INV_X1 U7140 ( .A(n5325), .ZN(n5575) );
  NAND2_X1 U7141 ( .A1(n6852), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5449) );
  NAND4_X1 U7142 ( .A1(n5452), .A2(n5451), .A3(n5450), .A4(n5449), .ZN(n9488)
         );
  INV_X1 U7143 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U7144 ( .A1(n5456), .A2(SI_12_), .ZN(n5457) );
  MUX2_X1 U7145 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6873), .Z(n5470) );
  XNOR2_X1 U7146 ( .A(n5469), .B(n5468), .ZN(n6985) );
  NAND2_X1 U7147 ( .A1(n6985), .A2(n6847), .ZN(n5461) );
  NAND2_X1 U7148 ( .A1(n5473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5459) );
  XNOR2_X1 U7149 ( .A(n5459), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7341) );
  AOI22_X1 U7150 ( .A1(n5589), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7341), .B2(
        n4465), .ZN(n5460) );
  NAND2_X1 U7151 ( .A1(n4458), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7152 ( .A1(n4457), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5464) );
  XNOR2_X1 U7153 ( .A(n5483), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n9409) );
  NAND2_X1 U7154 ( .A1(n5767), .A2(n9409), .ZN(n5463) );
  NAND2_X1 U7155 ( .A1(n6852), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5462) );
  OR2_X1 U7156 ( .A1(n8082), .A2(n8013), .ZN(n8153) );
  NAND2_X1 U7157 ( .A1(n8082), .A2(n8013), .ZN(n8156) );
  INV_X1 U7158 ( .A(n8013), .ZN(n9487) );
  OR2_X1 U7159 ( .A1(n8082), .A2(n9487), .ZN(n5467) );
  NAND2_X1 U7160 ( .A1(n5470), .A2(SI_13_), .ZN(n5471) );
  BUF_X1 U7161 ( .A(n5492), .Z(n5472) );
  MUX2_X1 U7162 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6873), .Z(n5493) );
  XNOR2_X1 U7163 ( .A(n5493), .B(SI_14_), .ZN(n5490) );
  XNOR2_X1 U7164 ( .A(n5472), .B(n5490), .ZN(n7105) );
  NAND2_X1 U7165 ( .A1(n7105), .A2(n6847), .ZN(n5479) );
  NAND2_X1 U7166 ( .A1(n5474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5476) );
  INV_X1 U7167 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7168 ( .A1(n5476), .A2(n5475), .ZN(n5497) );
  OR2_X1 U7169 ( .A1(n5476), .A2(n5475), .ZN(n5477) );
  AOI22_X1 U7170 ( .A1(n7484), .A2(n4459), .B1(n5589), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5478) );
  NAND2_X2 U7171 ( .A1(n5479), .A2(n5478), .ZN(n9963) );
  NAND2_X1 U7172 ( .A1(n4458), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5488) );
  INV_X1 U7173 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5482) );
  INV_X1 U7174 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5481) );
  OAI21_X1 U7175 ( .B1(n5483), .B2(n5482), .A(n5481), .ZN(n5484) );
  AND2_X1 U7176 ( .A1(n5501), .A2(n5484), .ZN(n9283) );
  NAND2_X1 U7177 ( .A1(n5767), .A2(n9283), .ZN(n5487) );
  NAND2_X1 U7178 ( .A1(n4456), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7179 ( .A1(n6852), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5485) );
  NAND4_X1 U7180 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n9486)
         );
  NAND2_X1 U7181 ( .A1(n9963), .A2(n9486), .ZN(n5489) );
  INV_X1 U7182 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U7183 ( .A1(n5492), .A2(n5491), .ZN(n5495) );
  NAND2_X1 U7184 ( .A1(n5493), .A2(SI_14_), .ZN(n5494) );
  MUX2_X1 U7185 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6873), .Z(n5510) );
  XNOR2_X1 U7186 ( .A(n5510), .B(SI_15_), .ZN(n5496) );
  XNOR2_X1 U7187 ( .A(n5514), .B(n5496), .ZN(n7119) );
  NAND2_X1 U7188 ( .A1(n7119), .A2(n6847), .ZN(n5500) );
  NAND2_X1 U7189 ( .A1(n5497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U7190 ( .A(n5498), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7672) );
  AOI22_X1 U7191 ( .A1(n7672), .A2(n4459), .B1(n5589), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7192 ( .A1(n5501), .A2(n7481), .ZN(n5502) );
  AND2_X1 U7193 ( .A1(n5525), .A2(n5502), .ZN(n9888) );
  NAND2_X1 U7194 ( .A1(n5767), .A2(n9888), .ZN(n5506) );
  NAND2_X1 U7195 ( .A1(n4458), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7196 ( .A1(n4456), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7197 ( .A1(n6852), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5503) );
  NAND4_X1 U7198 ( .A1(n5506), .A2(n5505), .A3(n5504), .A4(n5503), .ZN(n9485)
         );
  NAND2_X1 U7199 ( .A1(n9886), .A2(n9485), .ZN(n5507) );
  NAND2_X1 U7200 ( .A1(n9883), .A2(n5507), .ZN(n5509) );
  OR2_X1 U7201 ( .A1(n9886), .A2(n9485), .ZN(n5508) );
  AND2_X1 U7202 ( .A1(n5510), .A2(SI_15_), .ZN(n5513) );
  INV_X1 U7203 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U7204 ( .A1(n5511), .A2(n10453), .ZN(n5512) );
  MUX2_X1 U7205 ( .A(n7257), .B(n10440), .S(n6873), .Z(n5532) );
  XNOR2_X1 U7206 ( .A(n5532), .B(SI_16_), .ZN(n5515) );
  XNOR2_X1 U7207 ( .A(n5551), .B(n5515), .ZN(n7254) );
  NAND2_X1 U7208 ( .A1(n7254), .A2(n6847), .ZN(n5522) );
  INV_X1 U7209 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5516) );
  AND3_X1 U7210 ( .A1(n5518), .A2(n5517), .A3(n5516), .ZN(n5784) );
  NAND2_X1 U7211 ( .A1(n5538), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5520) );
  XNOR2_X1 U7212 ( .A(n5520), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7884) );
  AOI22_X1 U7213 ( .A1(n5589), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4465), .B2(
        n7884), .ZN(n5521) );
  NAND2_X1 U7214 ( .A1(n4458), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7215 ( .A1(n4456), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5529) );
  INV_X1 U7216 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7217 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  AND2_X1 U7218 ( .A1(n5542), .A2(n5526), .ZN(n9868) );
  NAND2_X1 U7219 ( .A1(n5767), .A2(n9868), .ZN(n5528) );
  NAND2_X1 U7220 ( .A1(n6852), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5527) );
  OR2_X1 U7221 ( .A1(n9867), .A2(n9456), .ZN(n8321) );
  NAND2_X1 U7222 ( .A1(n9867), .A2(n9456), .ZN(n8326) );
  INV_X1 U7223 ( .A(n9456), .ZN(n9484) );
  NAND2_X1 U7224 ( .A1(n9867), .A2(n9484), .ZN(n5531) );
  NAND2_X1 U7225 ( .A1(n5533), .A2(SI_16_), .ZN(n5555) );
  MUX2_X1 U7226 ( .A(n7351), .B(n5534), .S(n6873), .Z(n5535) );
  NAND2_X1 U7227 ( .A1(n5535), .A2(n10421), .ZN(n5552) );
  INV_X1 U7228 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U7229 ( .A1(n5536), .A2(SI_17_), .ZN(n5537) );
  NAND2_X1 U7230 ( .A1(n5552), .A2(n5537), .ZN(n5554) );
  NAND2_X1 U7231 ( .A1(n7292), .A2(n6847), .ZN(n5540) );
  XNOR2_X1 U7232 ( .A(n5561), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9614) );
  AOI22_X1 U7233 ( .A1(n5589), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4459), .B2(
        n9614), .ZN(n5539) );
  INV_X1 U7234 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7235 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  AND2_X1 U7236 ( .A1(n5571), .A2(n5543), .ZN(n9846) );
  NAND2_X1 U7237 ( .A1(n5767), .A2(n9846), .ZN(n5547) );
  NAND2_X1 U7238 ( .A1(n4458), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7239 ( .A1(n4456), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7240 ( .A1(n6852), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5544) );
  NAND4_X1 U7241 ( .A1(n5547), .A2(n5546), .A3(n5545), .A4(n5544), .ZN(n9483)
         );
  OR2_X1 U7242 ( .A1(n9842), .A2(n9483), .ZN(n5548) );
  NAND2_X1 U7243 ( .A1(n9837), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7244 ( .A1(n9842), .A2(n9483), .ZN(n5549) );
  NAND2_X1 U7245 ( .A1(n5550), .A2(n5549), .ZN(n9818) );
  INV_X1 U7246 ( .A(n5552), .ZN(n5558) );
  INV_X1 U7247 ( .A(n5554), .ZN(n5556) );
  MUX2_X1 U7248 ( .A(n7352), .B(n5559), .S(n6873), .Z(n5579) );
  XNOR2_X1 U7249 ( .A(n5583), .B(n5578), .ZN(n7315) );
  NAND2_X1 U7250 ( .A1(n7315), .A2(n6847), .ZN(n5567) );
  INV_X1 U7251 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7252 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  OR2_X1 U7253 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  AND2_X1 U7254 ( .A1(n5587), .A2(n5565), .ZN(n9627) );
  AOI22_X1 U7255 ( .A1(n5589), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4459), .B2(
        n9627), .ZN(n5566) );
  INV_X1 U7256 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U7257 ( .A1(n4458), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7258 ( .A1(n4456), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5568) );
  AND2_X1 U7259 ( .A1(n5569), .A2(n5568), .ZN(n5574) );
  INV_X1 U7260 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7261 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  NAND2_X1 U7262 ( .A1(n5593), .A2(n5572), .ZN(n9828) );
  OR2_X1 U7263 ( .A1(n9828), .A2(n5721), .ZN(n5573) );
  OAI211_X1 U7264 ( .C1(n5575), .C2(n9617), .A(n5574), .B(n5573), .ZN(n9482)
         );
  AND2_X1 U7265 ( .A1(n9943), .A2(n9482), .ZN(n5577) );
  OR2_X1 U7266 ( .A1(n9943), .A2(n9482), .ZN(n5576) );
  INV_X1 U7267 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7268 ( .A1(n5580), .A2(SI_18_), .ZN(n5581) );
  MUX2_X1 U7269 ( .A(n10312), .B(n7430), .S(n6873), .Z(n5584) );
  INV_X1 U7270 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7271 ( .A1(n5585), .A2(SI_19_), .ZN(n5586) );
  NAND2_X1 U7272 ( .A1(n5598), .A2(n5586), .ZN(n5599) );
  XNOR2_X1 U7273 ( .A(n5600), .B(n5599), .ZN(n7427) );
  NAND2_X1 U7274 ( .A1(n7427), .A2(n6847), .ZN(n5591) );
  AOI22_X1 U7275 ( .A1(n5589), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5780), .B2(
        n4465), .ZN(n5590) );
  INV_X1 U7276 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10368) );
  INV_X1 U7277 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U7278 ( .A1(n5593), .A2(n10257), .ZN(n5594) );
  NAND2_X1 U7279 ( .A1(n5604), .A2(n5594), .ZN(n9811) );
  OR2_X1 U7280 ( .A1(n9811), .A2(n5721), .ZN(n5596) );
  AOI22_X1 U7281 ( .A1(n4456), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n6852), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7282 ( .C1(n5771), .C2(n10368), .A(n5596), .B(n5595), .ZN(n9481)
         );
  NOR2_X1 U7283 ( .A1(n10006), .A2(n9481), .ZN(n5597) );
  MUX2_X1 U7284 ( .A(n8364), .B(n7535), .S(n6873), .Z(n5626) );
  XNOR2_X1 U7285 ( .A(n5626), .B(SI_20_), .ZN(n5601) );
  NAND2_X1 U7286 ( .A1(n8363), .A2(n6847), .ZN(n5603) );
  OR2_X1 U7287 ( .A1(n4470), .A2(n7535), .ZN(n5602) );
  INV_X1 U7288 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5608) );
  INV_X1 U7289 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U7290 ( .A1(n5604), .A2(n9397), .ZN(n5605) );
  NAND2_X1 U7291 ( .A1(n5616), .A2(n5605), .ZN(n9794) );
  OR2_X1 U7292 ( .A1(n9794), .A2(n5721), .ZN(n5607) );
  AOI22_X1 U7293 ( .A1(n4458), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4457), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U7294 ( .C1(n5575), .C2(n5608), .A(n5607), .B(n5606), .ZN(n9480)
         );
  AND2_X1 U7295 ( .A1(n9791), .A2(n9480), .ZN(n5609) );
  OAI21_X1 U7296 ( .B1(n5625), .B2(n10268), .A(n5626), .ZN(n5611) );
  NAND2_X1 U7297 ( .A1(n5625), .A2(n10268), .ZN(n5610) );
  NAND2_X1 U7298 ( .A1(n5611), .A2(n5610), .ZN(n5613) );
  MUX2_X1 U7299 ( .A(n10313), .B(n7752), .S(n6873), .Z(n5629) );
  XNOR2_X1 U7300 ( .A(n5629), .B(SI_21_), .ZN(n5612) );
  OR2_X1 U7302 ( .A1(n4469), .A2(n7752), .ZN(n5614) );
  NAND2_X2 U7303 ( .A1(n5615), .A2(n5614), .ZN(n9781) );
  INV_X1 U7304 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U7305 ( .A1(n5616), .A2(n9333), .ZN(n5617) );
  NAND2_X1 U7306 ( .A1(n5642), .A2(n5617), .ZN(n9330) );
  INV_X1 U7307 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U7308 ( .A1(n6852), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7309 ( .A1(n4457), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7310 ( .C1(n5771), .C2(n9930), .A(n5619), .B(n5618), .ZN(n5620)
         );
  INV_X1 U7311 ( .A(n5620), .ZN(n5621) );
  OAI21_X1 U7312 ( .B1(n9330), .B2(n5721), .A(n5621), .ZN(n9479) );
  NAND2_X1 U7313 ( .A1(n9781), .A2(n9479), .ZN(n5622) );
  INV_X1 U7314 ( .A(SI_21_), .ZN(n5627) );
  AOI22_X1 U7315 ( .A1(n10268), .A2(n5626), .B1(n5629), .B2(n5627), .ZN(n5623)
         );
  INV_X1 U7316 ( .A(n5623), .ZN(n5624) );
  INV_X1 U7317 ( .A(n5626), .ZN(n5631) );
  NAND2_X1 U7318 ( .A1(n5631), .A2(SI_20_), .ZN(n5628) );
  NAND2_X1 U7319 ( .A1(n5628), .A2(n5627), .ZN(n5633) );
  INV_X1 U7320 ( .A(n5629), .ZN(n5632) );
  AND2_X1 U7321 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5630) );
  AOI22_X1 U7322 ( .A1(n5633), .A2(n5632), .B1(n5631), .B2(n5630), .ZN(n5634)
         );
  MUX2_X1 U7323 ( .A(n10302), .B(n10288), .S(n6873), .Z(n5636) );
  INV_X1 U7324 ( .A(SI_22_), .ZN(n5635) );
  NAND2_X1 U7325 ( .A1(n5636), .A2(n5635), .ZN(n5651) );
  INV_X1 U7326 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U7327 ( .A1(n5637), .A2(SI_22_), .ZN(n5638) );
  NAND2_X1 U7328 ( .A1(n5651), .A2(n5638), .ZN(n5649) );
  XNOR2_X1 U7329 ( .A(n5650), .B(n5649), .ZN(n7796) );
  NAND2_X1 U7330 ( .A1(n7796), .A2(n6847), .ZN(n5640) );
  OR2_X1 U7331 ( .A1(n4470), .A2(n10288), .ZN(n5639) );
  INV_X1 U7332 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7333 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  AND2_X1 U7334 ( .A1(n5663), .A2(n5643), .ZN(n9764) );
  NAND2_X1 U7335 ( .A1(n9764), .A2(n5767), .ZN(n5648) );
  INV_X1 U7336 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U7337 ( .A1(n4457), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7338 ( .A1(n6852), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5644) );
  OAI211_X1 U7339 ( .C1(n9924), .C2(n5771), .A(n5645), .B(n5644), .ZN(n5646)
         );
  INV_X1 U7340 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7341 ( .A1(n5648), .A2(n5647), .ZN(n9478) );
  NAND2_X1 U7342 ( .A1(n5652), .A2(n5651), .ZN(n5673) );
  INV_X1 U7343 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5653) );
  MUX2_X1 U7344 ( .A(n5653), .B(n5658), .S(n6873), .Z(n5655) );
  INV_X1 U7345 ( .A(SI_23_), .ZN(n5654) );
  NAND2_X1 U7346 ( .A1(n5655), .A2(n5654), .ZN(n5674) );
  INV_X1 U7347 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7348 ( .A1(n5656), .A2(SI_23_), .ZN(n5657) );
  NAND2_X1 U7349 ( .A1(n7843), .A2(n6847), .ZN(n5660) );
  OR2_X1 U7350 ( .A1(n4470), .A2(n5658), .ZN(n5659) );
  INV_X1 U7351 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7352 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  NAND2_X1 U7353 ( .A1(n5700), .A2(n5664), .ZN(n9298) );
  INV_X1 U7354 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U7355 ( .A1(n6852), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7356 ( .A1(n4457), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U7357 ( .C1(n5771), .C2(n9919), .A(n5666), .B(n5665), .ZN(n5667)
         );
  INV_X1 U7358 ( .A(n5667), .ZN(n5668) );
  NAND2_X2 U7359 ( .A1(n5669), .A2(n5668), .ZN(n9477) );
  NOR2_X1 U7360 ( .A1(n9752), .A2(n9477), .ZN(n5671) );
  NAND2_X1 U7361 ( .A1(n9752), .A2(n9477), .ZN(n5670) );
  NAND2_X1 U7362 ( .A1(n5673), .A2(n5672), .ZN(n5675) );
  NAND2_X1 U7363 ( .A1(n5675), .A2(n5674), .ZN(n5689) );
  MUX2_X1 U7364 ( .A(n7997), .B(n8000), .S(n6873), .Z(n5676) );
  NAND2_X1 U7365 ( .A1(n5676), .A2(n10292), .ZN(n5690) );
  INV_X1 U7366 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7367 ( .A1(n5677), .A2(SI_24_), .ZN(n5678) );
  XNOR2_X1 U7368 ( .A(n5689), .B(n5688), .ZN(n7996) );
  NAND2_X1 U7369 ( .A1(n7996), .A2(n6847), .ZN(n5680) );
  OR2_X1 U7370 ( .A1(n4470), .A2(n8000), .ZN(n5679) );
  XNOR2_X1 U7371 ( .A(n5700), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U7372 ( .A1(n9737), .A2(n5767), .ZN(n5685) );
  INV_X1 U7373 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U7374 ( .A1(n6852), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7375 ( .A1(n4456), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5681) );
  OAI211_X1 U7376 ( .C1(n5771), .C2(n10341), .A(n5682), .B(n5681), .ZN(n5683)
         );
  INV_X1 U7377 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7378 ( .A1(n5685), .A2(n5684), .ZN(n9476) );
  OR2_X1 U7379 ( .A1(n9736), .A2(n9476), .ZN(n5687) );
  MUX2_X1 U7380 ( .A(n8028), .B(n8088), .S(n6873), .Z(n5692) );
  INV_X1 U7381 ( .A(SI_25_), .ZN(n5691) );
  NAND2_X1 U7382 ( .A1(n5692), .A2(n5691), .ZN(n5710) );
  INV_X1 U7383 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7384 ( .A1(n5693), .A2(SI_25_), .ZN(n5694) );
  XNOR2_X1 U7385 ( .A(n5709), .B(n5708), .ZN(n8027) );
  NAND2_X1 U7386 ( .A1(n8027), .A2(n6847), .ZN(n5696) );
  OR2_X1 U7387 ( .A1(n4469), .A2(n8088), .ZN(n5695) );
  INV_X1 U7388 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5698) );
  INV_X1 U7389 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5697) );
  OAI21_X1 U7390 ( .B1(n5700), .B2(n5698), .A(n5697), .ZN(n5701) );
  NAND2_X1 U7391 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5699) );
  INV_X1 U7392 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U7393 ( .A1(n6852), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7394 ( .A1(n4457), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U7395 ( .C1(n5771), .C2(n9909), .A(n5703), .B(n5702), .ZN(n5704)
         );
  INV_X1 U7396 ( .A(n5704), .ZN(n5705) );
  NOR2_X1 U7397 ( .A1(n9357), .A2(n9475), .ZN(n5707) );
  MUX2_X1 U7398 ( .A(n10429), .B(n8101), .S(n6873), .Z(n5712) );
  INV_X1 U7399 ( .A(SI_26_), .ZN(n5711) );
  NAND2_X1 U7400 ( .A1(n5712), .A2(n5711), .ZN(n5743) );
  INV_X1 U7401 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7402 ( .A1(n5713), .A2(SI_26_), .ZN(n5714) );
  NAND2_X1 U7403 ( .A1(n8099), .A2(n6847), .ZN(n5716) );
  OR2_X1 U7404 ( .A1(n4470), .A2(n8101), .ZN(n5715) );
  INV_X1 U7405 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7406 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NAND2_X1 U7407 ( .A1(n5753), .A2(n5720), .ZN(n9441) );
  INV_X1 U7408 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U7409 ( .A1(n6852), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7410 ( .A1(n4457), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5722) );
  OAI211_X1 U7411 ( .C1(n5771), .C2(n10437), .A(n5723), .B(n5722), .ZN(n5724)
         );
  INV_X1 U7412 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U7413 ( .A1(n9706), .A2(n9359), .ZN(n8272) );
  NAND2_X1 U7414 ( .A1(n9706), .A2(n9474), .ZN(n5727) );
  NAND2_X1 U7415 ( .A1(n5729), .A2(n5728), .ZN(n5747) );
  NAND2_X1 U7416 ( .A1(n5747), .A2(n5743), .ZN(n5735) );
  INV_X1 U7417 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5730) );
  MUX2_X1 U7418 ( .A(n5730), .B(n10285), .S(n6873), .Z(n5732) );
  INV_X1 U7419 ( .A(SI_27_), .ZN(n5731) );
  NAND2_X1 U7420 ( .A1(n5732), .A2(n5731), .ZN(n5742) );
  INV_X1 U7421 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7422 ( .A1(n5733), .A2(SI_27_), .ZN(n5744) );
  AND2_X1 U7423 ( .A1(n5742), .A2(n5744), .ZN(n5734) );
  NAND2_X1 U7424 ( .A1(n8445), .A2(n6847), .ZN(n5737) );
  OR2_X1 U7425 ( .A1(n4469), .A2(n10285), .ZN(n5736) );
  XNOR2_X1 U7426 ( .A(n5753), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9691) );
  INV_X1 U7427 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U7428 ( .A1(n4457), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7429 ( .A1(n6852), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5738) );
  OAI211_X1 U7430 ( .C1(n5771), .C2(n10394), .A(n5739), .B(n5738), .ZN(n5740)
         );
  NAND2_X1 U7431 ( .A1(n9690), .A2(n9438), .ZN(n8191) );
  INV_X1 U7432 ( .A(n9438), .ZN(n9473) );
  OR2_X1 U7433 ( .A1(n9690), .A2(n9473), .ZN(n5741) );
  AND2_X1 U7434 ( .A1(n5743), .A2(n5742), .ZN(n5746) );
  INV_X1 U7435 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5749) );
  INV_X1 U7436 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8380) );
  MUX2_X1 U7437 ( .A(n5749), .B(n8380), .S(n6873), .Z(n5761) );
  XNOR2_X1 U7438 ( .A(n5761), .B(SI_28_), .ZN(n5758) );
  NAND2_X1 U7439 ( .A1(n8379), .A2(n6847), .ZN(n5751) );
  OR2_X1 U7440 ( .A1(n4470), .A2(n8380), .ZN(n5750) );
  INV_X1 U7441 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9269) );
  INV_X1 U7442 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10328) );
  OAI21_X1 U7443 ( .B1(n5753), .B2(n9269), .A(n10328), .ZN(n5754) );
  NAND2_X1 U7444 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n5752) );
  INV_X1 U7445 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7446 ( .A1(n6852), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7447 ( .A1(n4456), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5755) );
  OAI211_X1 U7448 ( .C1(n5771), .C2(n6115), .A(n5756), .B(n5755), .ZN(n5757)
         );
  NAND2_X1 U7449 ( .A1(n6359), .A2(n9266), .ZN(n8192) );
  INV_X1 U7450 ( .A(n9662), .ZN(n5788) );
  NAND2_X1 U7451 ( .A1(n5759), .A2(n5758), .ZN(n5763) );
  INV_X1 U7452 ( .A(SI_28_), .ZN(n5760) );
  NAND2_X1 U7453 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  INV_X1 U7454 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8368) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10287) );
  MUX2_X1 U7456 ( .A(n8368), .B(n10287), .S(n6873), .Z(n6832) );
  XNOR2_X1 U7457 ( .A(n6832), .B(SI_29_), .ZN(n5764) );
  OR2_X1 U7458 ( .A1(n4469), .A2(n10287), .ZN(n5765) );
  INV_X1 U7459 ( .A(n5766), .ZN(n9660) );
  NAND2_X1 U7460 ( .A1(n9660), .A2(n5767), .ZN(n5774) );
  INV_X1 U7461 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7462 ( .A1(n5325), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7463 ( .A1(n4456), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5768) );
  OAI211_X1 U7464 ( .C1(n5771), .C2(n5770), .A(n5769), .B(n5768), .ZN(n5772)
         );
  INV_X1 U7465 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U7466 ( .A1(n5774), .A2(n5773), .ZN(n9471) );
  INV_X1 U7467 ( .A(n9471), .ZN(n5775) );
  NAND2_X1 U7468 ( .A1(n9665), .A2(n5775), .ZN(n8285) );
  NAND2_X1 U7469 ( .A1(n5776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7470 ( .A1(n5777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5778) );
  INV_X1 U7471 ( .A(n8292), .ZN(n5779) );
  INV_X1 U7472 ( .A(n6345), .ZN(n7059) );
  NAND2_X1 U7473 ( .A1(n5779), .A2(n7059), .ZN(n7444) );
  INV_X1 U7474 ( .A(n5781), .ZN(n5782) );
  NOR2_X1 U7475 ( .A1(n5782), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5783) );
  NAND3_X1 U7476 ( .A1(n5006), .A2(n5784), .A3(n5783), .ZN(n5785) );
  NAND2_X1 U7477 ( .A1(n5785), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7478 ( .A1(n7428), .A2(n8358), .ZN(n6122) );
  AND2_X1 U7479 ( .A1(n8356), .A2(n6122), .ZN(n5787) );
  NAND3_X1 U7480 ( .A1(n5788), .A2(n9663), .A3(n10071), .ZN(n5844) );
  NAND2_X1 U7481 ( .A1(n8235), .A2(n7326), .ZN(n5790) );
  NAND2_X1 U7482 ( .A1(n6124), .A2(n10055), .ZN(n5789) );
  NAND2_X1 U7483 ( .A1(n5790), .A2(n5789), .ZN(n7249) );
  NAND2_X1 U7484 ( .A1(n5320), .A2(n7460), .ZN(n5791) );
  INV_X1 U7485 ( .A(n5792), .ZN(n5794) );
  NAND2_X1 U7486 ( .A1(n7550), .A2(n5795), .ZN(n5796) );
  INV_X1 U7487 ( .A(n8243), .ZN(n5799) );
  NAND3_X1 U7488 ( .A1(n8129), .A2(n8121), .A3(n5799), .ZN(n5800) );
  NAND2_X1 U7489 ( .A1(n5800), .A2(n8140), .ZN(n8307) );
  NAND2_X1 U7490 ( .A1(n9493), .A2(n4466), .ZN(n7722) );
  AND2_X1 U7491 ( .A1(n8121), .A2(n7722), .ZN(n8239) );
  AND3_X1 U7492 ( .A1(n8239), .A2(n8129), .A3(n7616), .ZN(n5801) );
  OR2_X1 U7493 ( .A1(n8307), .A2(n5801), .ZN(n8310) );
  INV_X1 U7494 ( .A(n7697), .ZN(n8245) );
  INV_X1 U7495 ( .A(n9489), .ZN(n5802) );
  NAND2_X1 U7496 ( .A1(n7821), .A2(n5802), .ZN(n8133) );
  AND2_X1 U7497 ( .A1(n8133), .A2(n8130), .ZN(n8314) );
  OR2_X1 U7498 ( .A1(n7821), .A2(n5802), .ZN(n8144) );
  XNOR2_X1 U7499 ( .A(n9338), .B(n9488), .ZN(n8247) );
  INV_X1 U7500 ( .A(n9488), .ZN(n8132) );
  OR2_X1 U7501 ( .A1(n9338), .A2(n8132), .ZN(n8145) );
  INV_X1 U7502 ( .A(n9486), .ZN(n5803) );
  NAND2_X1 U7503 ( .A1(n9963), .A2(n5803), .ZN(n8155) );
  NAND2_X1 U7504 ( .A1(n9874), .A2(n8155), .ZN(n8251) );
  INV_X1 U7505 ( .A(n8156), .ZN(n5804) );
  NOR2_X1 U7506 ( .A1(n8251), .A2(n5804), .ZN(n8149) );
  INV_X1 U7507 ( .A(n9485), .ZN(n9370) );
  OR2_X1 U7508 ( .A1(n9886), .A2(n9370), .ZN(n8320) );
  NAND2_X1 U7509 ( .A1(n9886), .A2(n9370), .ZN(n8154) );
  NAND2_X1 U7510 ( .A1(n8320), .A2(n8154), .ZN(n9884) );
  INV_X1 U7511 ( .A(n9874), .ZN(n5805) );
  NOR2_X1 U7512 ( .A1(n9884), .A2(n5805), .ZN(n5806) );
  INV_X1 U7513 ( .A(n9483), .ZN(n9371) );
  OR2_X1 U7514 ( .A1(n9842), .A2(n9371), .ZN(n8163) );
  NAND2_X1 U7515 ( .A1(n9842), .A2(n9371), .ZN(n8175) );
  NAND2_X1 U7516 ( .A1(n8163), .A2(n8175), .ZN(n9838) );
  NAND2_X1 U7517 ( .A1(n9839), .A2(n5808), .ZN(n9819) );
  INV_X1 U7518 ( .A(n9482), .ZN(n5809) );
  OR2_X1 U7519 ( .A1(n9943), .A2(n5809), .ZN(n8177) );
  NAND2_X1 U7520 ( .A1(n9943), .A2(n5809), .ZN(n8176) );
  NAND2_X1 U7521 ( .A1(n8177), .A2(n8176), .ZN(n9820) );
  INV_X1 U7522 ( .A(n8163), .ZN(n9821) );
  NOR2_X1 U7523 ( .A1(n9820), .A2(n9821), .ZN(n5810) );
  NAND2_X1 U7524 ( .A1(n9819), .A2(n5810), .ZN(n9823) );
  NAND2_X1 U7525 ( .A1(n9823), .A2(n8176), .ZN(n9803) );
  INV_X1 U7526 ( .A(n9481), .ZN(n5811) );
  OR2_X1 U7527 ( .A1(n10006), .A2(n5811), .ZN(n8178) );
  NAND2_X1 U7528 ( .A1(n10006), .A2(n5811), .ZN(n8330) );
  INV_X1 U7529 ( .A(n9479), .ZN(n8255) );
  NAND2_X1 U7530 ( .A1(n10003), .A2(n9480), .ZN(n9771) );
  AND2_X1 U7531 ( .A1(n8118), .A2(n9771), .ZN(n8335) );
  INV_X1 U7532 ( .A(n9480), .ZN(n5812) );
  AND2_X1 U7533 ( .A1(n9791), .A2(n5812), .ZN(n8165) );
  NAND2_X1 U7534 ( .A1(n8118), .A2(n8165), .ZN(n5813) );
  NAND2_X1 U7535 ( .A1(n9781), .A2(n8255), .ZN(n8183) );
  AND2_X1 U7536 ( .A1(n5813), .A2(n8183), .ZN(n8268) );
  INV_X1 U7537 ( .A(n9478), .ZN(n6291) );
  OR2_X1 U7538 ( .A1(n9418), .A2(n6291), .ZN(n9744) );
  NAND2_X1 U7539 ( .A1(n9418), .A2(n6291), .ZN(n8167) );
  NAND2_X1 U7540 ( .A1(n9744), .A2(n8167), .ZN(n8227) );
  INV_X1 U7541 ( .A(n9477), .ZN(n5815) );
  OR2_X1 U7542 ( .A1(n9752), .A2(n5815), .ZN(n8169) );
  INV_X1 U7543 ( .A(n9744), .ZN(n8116) );
  NAND2_X1 U7544 ( .A1(n9736), .A2(n9358), .ZN(n8270) );
  NAND2_X1 U7545 ( .A1(n8263), .A2(n8270), .ZN(n9729) );
  NAND2_X1 U7546 ( .A1(n5818), .A2(n5817), .ZN(n9731) );
  NAND2_X1 U7547 ( .A1(n9731), .A2(n8263), .ZN(n9713) );
  NAND2_X1 U7548 ( .A1(n9357), .A2(n6305), .ZN(n8273) );
  INV_X1 U7549 ( .A(n9698), .ZN(n8265) );
  NOR2_X1 U7550 ( .A1(n9704), .A2(n8265), .ZN(n5819) );
  NAND2_X1 U7551 ( .A1(n5821), .A2(n4634), .ZN(n6107) );
  NAND2_X1 U7552 ( .A1(n6107), .A2(n8280), .ZN(n5822) );
  XNOR2_X1 U7553 ( .A(n5822), .B(n8206), .ZN(n5831) );
  NAND2_X1 U7554 ( .A1(n5780), .A2(n8358), .ZN(n5823) );
  NAND2_X1 U7555 ( .A1(n8300), .A2(n8223), .ZN(n8296) );
  INV_X1 U7556 ( .A(n9266), .ZN(n9472) );
  INV_X1 U7557 ( .A(n5824), .ZN(n9514) );
  INV_X1 U7558 ( .A(P1_B_REG_SCAN_IN), .ZN(n10459) );
  OR2_X1 U7559 ( .A1(n10031), .A2(n10459), .ZN(n5826) );
  AND2_X1 U7560 ( .A1(n9426), .A2(n5826), .ZN(n6856) );
  NAND2_X1 U7561 ( .A1(n4458), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7562 ( .A1(n5325), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7563 ( .A1(n4456), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5827) );
  NAND3_X1 U7564 ( .A1(n5829), .A2(n5828), .A3(n5827), .ZN(n9470) );
  NAND2_X1 U7565 ( .A1(n4588), .A2(n7321), .ZN(n7320) );
  INV_X1 U7566 ( .A(n7968), .ZN(n7709) );
  INV_X1 U7567 ( .A(n9963), .ZN(n8021) );
  INV_X1 U7568 ( .A(n9943), .ZN(n9831) );
  INV_X1 U7569 ( .A(n5834), .ZN(n9735) );
  NAND2_X1 U7570 ( .A1(n9665), .A2(n6111), .ZN(n5836) );
  NAND2_X1 U7571 ( .A1(n9651), .A2(n5836), .ZN(n9668) );
  INV_X1 U7572 ( .A(n10071), .ZN(n9968) );
  NAND2_X1 U7573 ( .A1(n6359), .A2(n9472), .ZN(n9661) );
  NOR3_X1 U7574 ( .A1(n8206), .A2(n9968), .A3(n9661), .ZN(n5839) );
  INV_X1 U7575 ( .A(n9964), .ZN(n10066) );
  NAND4_X1 U7576 ( .A1(n9662), .A2(n8206), .A3(n10071), .A4(n9661), .ZN(n5843)
         );
  OR2_X1 U7577 ( .A1(n5845), .A2(n5847), .ZN(n5848) );
  NAND2_X1 U7578 ( .A1(n8090), .A2(P1_B_REG_SCAN_IN), .ZN(n5851) );
  MUX2_X1 U7579 ( .A(n5851), .B(P1_B_REG_SCAN_IN), .S(n7999), .Z(n5852) );
  INV_X1 U7580 ( .A(n5873), .ZN(n8103) );
  NAND2_X1 U7581 ( .A1(n8103), .A2(n8090), .ZN(n6915) );
  OAI21_X1 U7582 ( .B1(n6914), .B2(P1_D_REG_1__SCAN_IN), .A(n6915), .ZN(n6336)
         );
  INV_X1 U7583 ( .A(n6914), .ZN(n5863) );
  NOR2_X1 U7584 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n10228) );
  NOR4_X1 U7585 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5855) );
  NOR4_X1 U7586 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5854) );
  NOR4_X1 U7587 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5853) );
  AND4_X1 U7588 ( .A1(n10228), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n5861)
         );
  NOR4_X1 U7589 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5859) );
  NOR4_X1 U7590 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5858) );
  NOR4_X1 U7591 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5857) );
  NOR4_X1 U7592 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5856) );
  AND4_X1 U7593 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n5860)
         );
  NAND2_X1 U7594 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7595 ( .A1(n5863), .A2(n5862), .ZN(n6337) );
  AND2_X1 U7596 ( .A1(n6336), .A2(n6337), .ZN(n5864) );
  NAND2_X1 U7597 ( .A1(n8356), .A2(n8292), .ZN(n6353) );
  INV_X1 U7598 ( .A(n8090), .ZN(n5866) );
  NAND2_X1 U7599 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U7600 ( .A1(n5870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7601 ( .A1(n6353), .A2(n10020), .ZN(n7242) );
  OAI22_X1 U7602 ( .A1(n6914), .A2(P1_D_REG_0__SCAN_IN), .B1(n5873), .B2(n7999), .ZN(n7447) );
  NOR2_X1 U7603 ( .A1(n7242), .A2(n7447), .ZN(n5874) );
  NAND2_X1 U7604 ( .A1(n5876), .A2(n5875), .ZN(P1_U3551) );
  NOR2_X1 U7605 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5879) );
  NOR2_X1 U7606 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5878) );
  NAND2_X1 U7607 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7608 ( .A1(n5884), .A2(n5883), .ZN(n7998) );
  NAND2_X1 U7609 ( .A1(n5908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7610 ( .A(n5889), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6709) );
  NOR2_X1 U7611 ( .A1(n7998), .A2(n8100), .ZN(n5890) );
  NOR2_X1 U7612 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5892) );
  AND2_X1 U7613 ( .A1(n5984), .A2(n5892), .ZN(n5995) );
  NOR2_X1 U7614 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5894) );
  INV_X1 U7615 ( .A(n5896), .ZN(n6685) );
  AND2_X1 U7616 ( .A1(n6684), .A2(n10304), .ZN(n5897) );
  NAND2_X1 U7617 ( .A1(n6685), .A2(n5897), .ZN(n5898) );
  NAND2_X1 U7618 ( .A1(n5898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  INV_X1 U7619 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7620 ( .A1(n5902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7621 ( .A1(n6767), .A2(n6697), .ZN(n5906) );
  NAND2_X1 U7622 ( .A1(n5904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7623 ( .A1(n5906), .A2(n7844), .ZN(n6029) );
  NAND2_X1 U7624 ( .A1(n10466), .A2(n5911), .ZN(n5907) );
  NAND2_X1 U7625 ( .A1(n6029), .A2(n6816), .ZN(n5915) );
  NAND2_X1 U7626 ( .A1(n5915), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7627 ( .A(n7844), .ZN(n6919) );
  INV_X1 U7628 ( .A(n5964), .ZN(n5918) );
  INV_X1 U7629 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7630 ( .A1(n5918), .A2(n5917), .ZN(n5967) );
  INV_X1 U7631 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5969) );
  INV_X1 U7632 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7633 ( .A1(n5969), .A2(n5919), .ZN(n5920) );
  INV_X1 U7634 ( .A(n5975), .ZN(n5922) );
  INV_X1 U7635 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7636 ( .A1(n5922), .A2(n5921), .ZN(n5997) );
  NAND2_X1 U7637 ( .A1(n5997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  INV_X1 U7638 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7639 ( .A1(n5987), .A2(n5923), .ZN(n5980) );
  OR2_X1 U7640 ( .A1(n5987), .A2(n5923), .ZN(n5924) );
  INV_X1 U7641 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10412) );
  INV_X1 U7642 ( .A(n5942), .ZN(n5926) );
  NAND2_X1 U7643 ( .A1(n5926), .A2(n5943), .ZN(n5946) );
  NAND2_X1 U7644 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  MUX2_X1 U7645 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5927), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5931) );
  INV_X1 U7646 ( .A(n5928), .ZN(n5930) );
  NAND2_X1 U7647 ( .A1(n5930), .A2(n5929), .ZN(n5951) );
  INV_X1 U7648 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U7649 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5932) );
  NAND2_X1 U7650 ( .A1(n5936), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7651 ( .A1(n5933), .A2(n5934), .ZN(n7174) );
  INV_X1 U7652 ( .A(n5934), .ZN(n5935) );
  NAND2_X1 U7653 ( .A1(n5925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5938) );
  MUX2_X1 U7654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5938), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5939) );
  NAND2_X1 U7655 ( .A1(n5939), .A2(n5942), .ZN(n7071) );
  NAND2_X1 U7656 ( .A1(n5942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5944) );
  XNOR2_X1 U7657 ( .A(n8798), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U7658 ( .A1(n5946), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5948) );
  INV_X1 U7659 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7660 ( .A(n5948), .B(n5947), .ZN(n6868) );
  INV_X1 U7661 ( .A(n5949), .ZN(n5950) );
  XNOR2_X1 U7662 ( .A(n6871), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U7663 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  INV_X1 U7664 ( .A(n5955), .ZN(n5956) );
  NAND2_X1 U7665 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  MUX2_X1 U7666 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5957), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5958) );
  NAND2_X1 U7667 ( .A1(n5958), .A2(n5959), .ZN(n7281) );
  INV_X1 U7668 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7537) );
  XNOR2_X1 U7669 ( .A(n7281), .B(n7537), .ZN(n7282) );
  OAI21_X1 U7670 ( .B1(n7284), .B2(n7283), .A(n7282), .ZN(n7286) );
  INV_X1 U7671 ( .A(n7281), .ZN(n6487) );
  NAND2_X1 U7672 ( .A1(n5959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5960) );
  MUX2_X1 U7673 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5960), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5961) );
  INV_X1 U7674 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7524) );
  INV_X1 U7675 ( .A(n5963), .ZN(n7593) );
  NAND2_X1 U7676 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7677 ( .A(n6504), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7592) );
  INV_X1 U7678 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U7679 ( .A1(n5967), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5970) );
  XNOR2_X1 U7680 ( .A(n5970), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6514) );
  OAI21_X1 U7681 ( .B1(n5968), .B2(n4771), .A(n8830), .ZN(n8815) );
  INV_X1 U7682 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U7683 ( .A1(n8832), .A2(n8830), .ZN(n5973) );
  NAND2_X1 U7684 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  NAND2_X1 U7685 ( .A1(n5971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7686 ( .A(n6525), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8829) );
  INV_X1 U7687 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7831) );
  OR2_X1 U7688 ( .A1(n6525), .A2(n7831), .ZN(n5974) );
  NAND2_X1 U7689 ( .A1(n5975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5976) );
  XNOR2_X1 U7690 ( .A(n5976), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6535) );
  INV_X1 U7691 ( .A(n6535), .ZN(n8848) );
  NAND2_X1 U7692 ( .A1(n5977), .A2(n8848), .ZN(n8862) );
  INV_X1 U7693 ( .A(n5977), .ZN(n5978) );
  NAND2_X1 U7694 ( .A1(n5980), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U7695 ( .A(n5981), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6556) );
  INV_X1 U7696 ( .A(n6556), .ZN(n8876) );
  INV_X1 U7697 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9107) );
  INV_X1 U7698 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7699 ( .A1(n5985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7700 ( .A1(n5987), .A2(n5986), .ZN(n5991) );
  XNOR2_X1 U7701 ( .A(n5991), .B(n5988), .ZN(n7255) );
  XNOR2_X1 U7702 ( .A(n7255), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8890) );
  INV_X1 U7703 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U7704 ( .A1(n5989), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5990) );
  OAI21_X1 U7705 ( .B1(n5991), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7706 ( .A(n5992), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6574) );
  INV_X1 U7707 ( .A(n6574), .ZN(n8906) );
  INV_X1 U7708 ( .A(n5995), .ZN(n5996) );
  OAI21_X1 U7709 ( .B1(n5997), .B2(n5996), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5998) );
  XNOR2_X1 U7710 ( .A(n5998), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6581) );
  INV_X1 U7711 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9069) );
  OR2_X1 U7712 ( .A1(n6581), .A2(n9069), .ZN(n6000) );
  NAND2_X1 U7713 ( .A1(n6581), .A2(n9069), .ZN(n5999) );
  AND2_X1 U7714 ( .A1(n6000), .A2(n5999), .ZN(n8918) );
  NAND2_X1 U7715 ( .A1(n8921), .A2(n6000), .ZN(n6001) );
  XNOR2_X1 U7716 ( .A(n8612), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7717 ( .A(n6001), .B(n6095), .ZN(n6099) );
  NOR2_X1 U7718 ( .A1(n6003), .A2(P2_U3151), .ZN(n9252) );
  AND2_X1 U7719 ( .A1(n6029), .A2(n9252), .ZN(n7141) );
  NAND2_X1 U7720 ( .A1(n7141), .A2(n6695), .ZN(n10088) );
  XNOR2_X1 U7721 ( .A(n8612), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6094) );
  INV_X1 U7722 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6413) );
  AND2_X1 U7723 ( .A1(n5936), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6006) );
  INV_X1 U7724 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U7725 ( .A1(n6411), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6005) );
  OAI22_X1 U7726 ( .A1(n6006), .A2(n6393), .B1(n5936), .B2(n6005), .ZN(n7172)
         );
  NAND2_X1 U7727 ( .A1(n7172), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6008) );
  INV_X1 U7728 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7729 ( .A1(n6008), .A2(n6007), .ZN(n7190) );
  NAND2_X1 U7730 ( .A1(n7185), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7731 ( .A1(n6010), .A2(n7071), .ZN(n6011) );
  NAND2_X1 U7732 ( .A1(n6012), .A2(n6011), .ZN(n8805) );
  INV_X1 U7733 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6436) );
  MUX2_X1 U7734 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6436), .S(n8798), .Z(n8806)
         );
  NAND2_X1 U7735 ( .A1(n8798), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6013) );
  INV_X1 U7736 ( .A(n6868), .ZN(n7205) );
  NAND2_X1 U7737 ( .A1(n6014), .A2(n6868), .ZN(n6015) );
  NAND2_X1 U7738 ( .A1(n6016), .A2(n6015), .ZN(n10079) );
  MUX2_X1 U7739 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10185), .S(n6871), .Z(n10080) );
  NAND2_X1 U7740 ( .A1(n10079), .A2(n10080), .ZN(n10078) );
  NAND2_X1 U7741 ( .A1(n6871), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7742 ( .A1(n10078), .A2(n6017), .ZN(n6018) );
  XNOR2_X1 U7743 ( .A(n6018), .B(n7162), .ZN(n7156) );
  NAND2_X1 U7744 ( .A1(n7156), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6020) );
  INV_X1 U7745 ( .A(n7162), .ZN(n6900) );
  NAND2_X1 U7746 ( .A1(n6018), .A2(n6900), .ZN(n6019) );
  INV_X1 U7747 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7502) );
  XNOR2_X1 U7748 ( .A(n7281), .B(n7502), .ZN(n7278) );
  INV_X1 U7749 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U7750 ( .A(n6504), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7587) );
  INV_X1 U7751 ( .A(n6504), .ZN(n7591) );
  INV_X1 U7752 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10316) );
  XNOR2_X1 U7753 ( .A(n6525), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8826) );
  INV_X1 U7754 ( .A(n6525), .ZN(n8828) );
  AOI22_X1 U7755 ( .A1(n8825), .A2(n8826), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n8828), .ZN(n6022) );
  INV_X1 U7756 ( .A(n6022), .ZN(n6023) );
  XOR2_X1 U7757 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7106), .Z(n8857) );
  INV_X1 U7758 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9153) );
  AOI22_X1 U7759 ( .A1(n8871), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n8876), .B2(
        n6024), .ZN(n8886) );
  XOR2_X1 U7760 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n7255), .Z(n8887) );
  INV_X1 U7761 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9144) );
  OAI22_X1 U7762 ( .A1(n8886), .A2(n8887), .B1(n9144), .B2(n7255), .ZN(n6025)
         );
  XNOR2_X1 U7763 ( .A(n6025), .B(n6574), .ZN(n8901) );
  AOI22_X1 U7764 ( .A1(n8901), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8906), .B2(
        n6025), .ZN(n8914) );
  XOR2_X1 U7765 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n6581), .Z(n8915) );
  INV_X1 U7766 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9138) );
  OAI22_X1 U7767 ( .A1(n8914), .A2(n8915), .B1(n6581), .B2(n9138), .ZN(n6026)
         );
  INV_X1 U7768 ( .A(n6027), .ZN(n6028) );
  NAND2_X1 U7769 ( .A1(n6028), .A2(n9252), .ZN(n6031) );
  NOR2_X1 U7770 ( .A1(n6089), .A2(P2_U3151), .ZN(n9255) );
  NAND3_X1 U7771 ( .A1(n6029), .A2(n9255), .A3(n6003), .ZN(n6030) );
  NAND2_X1 U7772 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8464) );
  OAI21_X1 U7773 ( .B1(n8928), .B2(n8612), .A(n8464), .ZN(n6097) );
  INV_X1 U7774 ( .A(n6581), .ZN(n8932) );
  INV_X1 U7775 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6400) );
  MUX2_X1 U7776 ( .A(n6402), .B(n6400), .S(n8766), .Z(n7139) );
  NAND2_X1 U7777 ( .A1(n7139), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7181) );
  INV_X1 U7778 ( .A(n6393), .ZN(n7171) );
  NAND2_X1 U7779 ( .A1(n6032), .A2(n7171), .ZN(n6033) );
  NAND2_X1 U7780 ( .A1(n7179), .A2(n6033), .ZN(n7199) );
  MUX2_X1 U7781 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6089), .Z(n6035) );
  INV_X1 U7782 ( .A(n7185), .ZN(n6034) );
  XNOR2_X1 U7783 ( .A(n6035), .B(n6034), .ZN(n7198) );
  NAND2_X1 U7784 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U7785 ( .A1(n6035), .A2(n7185), .ZN(n6036) );
  NAND2_X1 U7786 ( .A1(n7197), .A2(n6036), .ZN(n7065) );
  MUX2_X1 U7787 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6089), .Z(n6037) );
  XNOR2_X1 U7788 ( .A(n6037), .B(n7071), .ZN(n7066) );
  INV_X1 U7789 ( .A(n6037), .ZN(n6039) );
  NAND2_X1 U7790 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  MUX2_X1 U7791 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6089), .Z(n6042) );
  INV_X1 U7792 ( .A(n8798), .ZN(n6041) );
  XNOR2_X1 U7793 ( .A(n6042), .B(n6041), .ZN(n8795) );
  NAND2_X1 U7794 ( .A1(n6042), .A2(n8798), .ZN(n6043) );
  MUX2_X1 U7795 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6089), .Z(n6044) );
  XNOR2_X1 U7796 ( .A(n6044), .B(n7205), .ZN(n7212) );
  NAND2_X1 U7797 ( .A1(n7213), .A2(n7212), .ZN(n7211) );
  NAND2_X1 U7798 ( .A1(n6044), .A2(n6868), .ZN(n6045) );
  NAND2_X1 U7799 ( .A1(n7211), .A2(n6045), .ZN(n10094) );
  MUX2_X1 U7800 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6089), .Z(n6046) );
  XNOR2_X1 U7801 ( .A(n6046), .B(n6871), .ZN(n10093) );
  INV_X1 U7802 ( .A(n6046), .ZN(n6047) );
  INV_X1 U7803 ( .A(n6871), .ZN(n10084) );
  NAND2_X1 U7804 ( .A1(n6047), .A2(n10084), .ZN(n6048) );
  MUX2_X1 U7805 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6089), .Z(n6049) );
  XNOR2_X1 U7806 ( .A(n6049), .B(n7162), .ZN(n7158) );
  INV_X1 U7807 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7808 ( .A1(n6050), .A2(n7162), .ZN(n6051) );
  MUX2_X1 U7809 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8766), .Z(n6052) );
  XNOR2_X1 U7810 ( .A(n6052), .B(n6487), .ZN(n7277) );
  NAND2_X1 U7811 ( .A1(n7276), .A2(n7277), .ZN(n6055) );
  INV_X1 U7812 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7813 ( .A1(n6053), .A2(n6487), .ZN(n6054) );
  NAND2_X1 U7814 ( .A1(n6055), .A2(n6054), .ZN(n7522) );
  MUX2_X1 U7815 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6089), .Z(n6056) );
  XNOR2_X1 U7816 ( .A(n6056), .B(n6478), .ZN(n7521) );
  NAND2_X1 U7817 ( .A1(n7522), .A2(n7521), .ZN(n6059) );
  INV_X1 U7818 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7819 ( .A1(n6057), .A2(n6478), .ZN(n6058) );
  MUX2_X1 U7820 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6089), .Z(n6060) );
  XNOR2_X1 U7821 ( .A(n6060), .B(n6504), .ZN(n7588) );
  INV_X1 U7822 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7823 ( .A1(n6061), .A2(n6504), .ZN(n6062) );
  MUX2_X1 U7824 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8766), .Z(n6063) );
  XNOR2_X1 U7825 ( .A(n6063), .B(n6514), .ZN(n8819) );
  INV_X1 U7826 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7827 ( .A1(n6064), .A2(n6514), .ZN(n6065) );
  NAND2_X1 U7828 ( .A1(n6066), .A2(n6065), .ZN(n8838) );
  MUX2_X1 U7829 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6089), .Z(n6067) );
  XNOR2_X1 U7830 ( .A(n6067), .B(n6525), .ZN(n8837) );
  INV_X1 U7831 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7832 ( .A1(n6068), .A2(n6525), .ZN(n6069) );
  MUX2_X1 U7833 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6089), .Z(n6071) );
  XNOR2_X1 U7834 ( .A(n6071), .B(n6535), .ZN(n8846) );
  INV_X1 U7835 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7836 ( .A1(n6072), .A2(n6535), .ZN(n6073) );
  MUX2_X1 U7837 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6089), .Z(n6074) );
  XNOR2_X1 U7838 ( .A(n7106), .B(n6074), .ZN(n8858) );
  INV_X1 U7839 ( .A(n6074), .ZN(n6075) );
  NAND2_X1 U7840 ( .A1(n7106), .A2(n6075), .ZN(n6076) );
  NAND2_X1 U7841 ( .A1(n6077), .A2(n6076), .ZN(n8873) );
  MUX2_X1 U7842 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6089), .Z(n6078) );
  XNOR2_X1 U7843 ( .A(n6556), .B(n6078), .ZN(n8872) );
  NAND2_X1 U7844 ( .A1(n8873), .A2(n8872), .ZN(n6081) );
  INV_X1 U7845 ( .A(n6078), .ZN(n6079) );
  NAND2_X1 U7846 ( .A1(n6556), .A2(n6079), .ZN(n6080) );
  NAND2_X1 U7847 ( .A1(n6081), .A2(n6080), .ZN(n8891) );
  MUX2_X1 U7848 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6089), .Z(n6082) );
  XNOR2_X1 U7849 ( .A(n7255), .B(n6082), .ZN(n8892) );
  NAND2_X1 U7850 ( .A1(n8891), .A2(n8892), .ZN(n6085) );
  INV_X1 U7851 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7852 ( .A1(n7255), .A2(n6083), .ZN(n6084) );
  NAND2_X1 U7853 ( .A1(n6085), .A2(n6084), .ZN(n8903) );
  MUX2_X1 U7854 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8766), .Z(n6086) );
  XNOR2_X1 U7855 ( .A(n6574), .B(n6086), .ZN(n8904) );
  INV_X1 U7856 ( .A(n6086), .ZN(n6087) );
  AND2_X1 U7857 ( .A1(n6574), .A2(n6087), .ZN(n6088) );
  INV_X1 U7858 ( .A(n6093), .ZN(n6091) );
  MUX2_X1 U7859 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6089), .Z(n6092) );
  INV_X1 U7860 ( .A(n6092), .ZN(n6090) );
  NAND2_X1 U7861 ( .A1(n6091), .A2(n6090), .ZN(n8925) );
  AND2_X1 U7862 ( .A1(n6093), .A2(n6092), .ZN(n8927) );
  MUX2_X1 U7863 ( .A(n6095), .B(n6094), .S(n8766), .Z(n6096) );
  NAND2_X1 U7864 ( .A1(P2_U3893), .A2(n6003), .ZN(n10095) );
  INV_X1 U7865 ( .A(n7447), .ZN(n10021) );
  NOR2_X1 U7866 ( .A1(n10021), .A2(n7242), .ZN(n6100) );
  NAND2_X1 U7867 ( .A1(n6102), .A2(n10074), .ZN(n6104) );
  NAND2_X1 U7868 ( .A1(n10072), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7869 ( .A1(n6104), .A2(n6103), .ZN(P1_U3519) );
  NAND2_X1 U7870 ( .A1(n6105), .A2(n4634), .ZN(n6106) );
  NAND3_X1 U7871 ( .A1(n6108), .A2(n8262), .A3(n8258), .ZN(n6109) );
  NAND3_X1 U7872 ( .A1(n6107), .A2(n9878), .A3(n6109), .ZN(n6110) );
  AOI22_X1 U7873 ( .A1(n9473), .A2(n9457), .B1(n9471), .B2(n9426), .ZN(n6357)
         );
  AOI21_X1 U7874 ( .B1(n6359), .B2(n9689), .A(n9885), .ZN(n6112) );
  NAND2_X1 U7875 ( .A1(n6112), .A2(n6111), .ZN(n9674) );
  NAND2_X1 U7876 ( .A1(n9682), .A2(n9674), .ZN(n6113) );
  INV_X1 U7877 ( .A(n6359), .ZN(n9677) );
  NAND2_X1 U7878 ( .A1(n10077), .A2(n9964), .ZN(n9961) );
  NAND2_X1 U7879 ( .A1(n8356), .A2(n6121), .ZN(n6118) );
  OAI22_X1 U7880 ( .A1(n9999), .A2(n4455), .B1(n8255), .B2(n6326), .ZN(n6290)
         );
  NAND2_X1 U7881 ( .A1(n9781), .A2(n6331), .ZN(n6120) );
  NAND2_X1 U7882 ( .A1(n9479), .A2(n6141), .ZN(n6119) );
  NAND2_X1 U7883 ( .A1(n6120), .A2(n6119), .ZN(n6123) );
  XNOR2_X1 U7884 ( .A(n6123), .B(n6318), .ZN(n6289) );
  OAI22_X1 U7885 ( .A1(n6124), .A2(n6326), .B1(n4588), .B2(n4455), .ZN(n6135)
         );
  XNOR2_X1 U7886 ( .A(n6134), .B(n6135), .ZN(n8438) );
  AND2_X1 U7887 ( .A1(n7452), .A2(n6331), .ZN(n6126) );
  AOI21_X1 U7888 ( .B1(n7323), .B2(n6141), .A(n6126), .ZN(n6132) );
  INV_X1 U7889 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6127) );
  OR2_X1 U7890 ( .A1(n6904), .A2(n6127), .ZN(n6128) );
  NAND2_X1 U7891 ( .A1(n6132), .A2(n6128), .ZN(n7241) );
  INV_X1 U7892 ( .A(n7323), .ZN(n6129) );
  INV_X1 U7893 ( .A(n6904), .ZN(n6130) );
  AOI22_X1 U7894 ( .A1(n7452), .A2(n6141), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6130), .ZN(n6131) );
  NAND2_X1 U7895 ( .A1(n7241), .A2(n7240), .ZN(n7239) );
  NAND2_X1 U7896 ( .A1(n6132), .A2(n6329), .ZN(n6133) );
  NAND2_X1 U7897 ( .A1(n8438), .A2(n8437), .ZN(n8436) );
  INV_X1 U7898 ( .A(n6134), .ZN(n6136) );
  OR2_X1 U7899 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  NAND2_X1 U7900 ( .A1(n8436), .A2(n6137), .ZN(n8371) );
  NAND2_X1 U7901 ( .A1(n9498), .A2(n6141), .ZN(n6139) );
  NAND2_X1 U7902 ( .A1(n7460), .A2(n6331), .ZN(n6138) );
  NAND2_X1 U7903 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  XNOR2_X1 U7904 ( .A(n6140), .B(n6318), .ZN(n6142) );
  AOI22_X1 U7905 ( .A1(n9498), .A2(n6307), .B1(n6141), .B2(n7460), .ZN(n6143)
         );
  XNOR2_X1 U7906 ( .A(n6142), .B(n6143), .ZN(n8370) );
  NAND2_X1 U7907 ( .A1(n8371), .A2(n8370), .ZN(n6146) );
  INV_X1 U7908 ( .A(n6142), .ZN(n6144) );
  NAND2_X1 U7909 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  NAND2_X1 U7910 ( .A1(n6146), .A2(n6145), .ZN(n7258) );
  OAI22_X1 U7911 ( .A1(n7250), .A2(n4455), .B1(n10046), .B2(n6317), .ZN(n6147)
         );
  XNOR2_X1 U7912 ( .A(n6147), .B(n6329), .ZN(n6148) );
  OAI22_X1 U7913 ( .A1(n7250), .A2(n6326), .B1(n10046), .B2(n4455), .ZN(n6149)
         );
  XNOR2_X1 U7914 ( .A(n6148), .B(n6149), .ZN(n7259) );
  INV_X1 U7915 ( .A(n6148), .ZN(n6150) );
  OR2_X1 U7916 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  OAI22_X1 U7917 ( .A1(n7260), .A2(n4455), .B1(n10067), .B2(n6317), .ZN(n6152)
         );
  XNOR2_X1 U7918 ( .A(n6152), .B(n6318), .ZN(n6155) );
  OAI22_X1 U7919 ( .A1(n7260), .A2(n6326), .B1(n10067), .B2(n4455), .ZN(n6154)
         );
  XNOR2_X1 U7920 ( .A(n6155), .B(n6154), .ZN(n7359) );
  INV_X1 U7921 ( .A(n7359), .ZN(n6153) );
  NAND2_X1 U7922 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  OAI22_X1 U7923 ( .A1(n7510), .A2(n4455), .B1(n5280), .B2(n6317), .ZN(n6157)
         );
  XNOR2_X1 U7924 ( .A(n6157), .B(n6318), .ZN(n7687) );
  OR2_X1 U7925 ( .A1(n7510), .A2(n6326), .ZN(n6159) );
  NAND2_X1 U7926 ( .A1(n7496), .A2(n6141), .ZN(n6158) );
  NAND2_X1 U7927 ( .A1(n6159), .A2(n6158), .ZN(n7491) );
  AND2_X1 U7928 ( .A1(n7687), .A2(n7491), .ZN(n6163) );
  OAI22_X1 U7929 ( .A1(n5232), .A2(n4455), .B1(n7516), .B2(n6317), .ZN(n6160)
         );
  XNOR2_X1 U7930 ( .A(n6160), .B(n6318), .ZN(n6164) );
  OR2_X1 U7931 ( .A1(n5232), .A2(n6326), .ZN(n6162) );
  NAND2_X1 U7932 ( .A1(n7692), .A2(n6141), .ZN(n6161) );
  NAND2_X1 U7933 ( .A1(n6162), .A2(n6161), .ZN(n7682) );
  AND2_X1 U7934 ( .A1(n6164), .A2(n7682), .ZN(n7683) );
  OAI21_X1 U7935 ( .B1(n7687), .B2(n7491), .A(n7682), .ZN(n6166) );
  INV_X1 U7936 ( .A(n6164), .ZN(n7685) );
  INV_X1 U7937 ( .A(n7687), .ZN(n7493) );
  NOR2_X1 U7938 ( .A1(n7491), .A2(n7682), .ZN(n6165) );
  AOI22_X1 U7939 ( .A1(n6166), .A2(n7685), .B1(n7493), .B2(n6165), .ZN(n6167)
         );
  NAND2_X1 U7940 ( .A1(n9493), .A2(n6141), .ZN(n6169) );
  OAI21_X1 U7941 ( .B1(n4466), .B2(n6317), .A(n6169), .ZN(n6170) );
  XNOR2_X1 U7942 ( .A(n6170), .B(n6329), .ZN(n6173) );
  OR2_X1 U7943 ( .A1(n4466), .A2(n4455), .ZN(n6172) );
  NAND2_X1 U7944 ( .A1(n9493), .A2(n6307), .ZN(n6171) );
  AND2_X1 U7945 ( .A1(n6172), .A2(n6171), .ZN(n6174) );
  NAND2_X1 U7946 ( .A1(n6173), .A2(n6174), .ZN(n7942) );
  INV_X1 U7947 ( .A(n6173), .ZN(n6176) );
  INV_X1 U7948 ( .A(n6174), .ZN(n6175) );
  NAND2_X1 U7949 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  AND2_X1 U7950 ( .A1(n7942), .A2(n6177), .ZN(n7569) );
  NAND2_X1 U7951 ( .A1(n9325), .A2(n6331), .ZN(n6179) );
  NAND2_X1 U7952 ( .A1(n9492), .A2(n6141), .ZN(n6178) );
  NAND2_X1 U7953 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  XNOR2_X1 U7954 ( .A(n6180), .B(n6318), .ZN(n6186) );
  NAND2_X1 U7955 ( .A1(n9325), .A2(n6141), .ZN(n6182) );
  NAND2_X1 U7956 ( .A1(n9492), .A2(n6307), .ZN(n6181) );
  NAND2_X1 U7957 ( .A1(n6182), .A2(n6181), .ZN(n9320) );
  NAND2_X1 U7958 ( .A1(n7727), .A2(n6331), .ZN(n6184) );
  OR2_X1 U7959 ( .A1(n7741), .A2(n4455), .ZN(n6183) );
  NAND2_X1 U7960 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  XNOR2_X1 U7961 ( .A(n6185), .B(n6318), .ZN(n6192) );
  AOI22_X1 U7962 ( .A1(n7727), .A2(n6141), .B1(n6307), .B2(n9491), .ZN(n6193)
         );
  XNOR2_X1 U7963 ( .A(n6192), .B(n6193), .ZN(n7947) );
  INV_X1 U7964 ( .A(n6186), .ZN(n7945) );
  NAND2_X1 U7965 ( .A1(n7942), .A2(n9320), .ZN(n6189) );
  INV_X1 U7966 ( .A(n7942), .ZN(n6188) );
  INV_X1 U7967 ( .A(n9320), .ZN(n6187) );
  AOI22_X1 U7968 ( .A1(n7945), .A2(n6189), .B1(n6188), .B2(n6187), .ZN(n6190)
         );
  AND2_X1 U7969 ( .A1(n7947), .A2(n6190), .ZN(n6191) );
  INV_X1 U7970 ( .A(n6192), .ZN(n6194) );
  OR2_X1 U7971 ( .A1(n6194), .A2(n6193), .ZN(n6201) );
  NAND2_X1 U7972 ( .A1(n7968), .A2(n6331), .ZN(n6196) );
  OR2_X1 U7973 ( .A1(n7728), .A2(n4455), .ZN(n6195) );
  NAND2_X1 U7974 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  XNOR2_X1 U7975 ( .A(n6197), .B(n6318), .ZN(n6200) );
  NAND2_X1 U7976 ( .A1(n6198), .A2(n6200), .ZN(n7961) );
  NOR2_X1 U7977 ( .A1(n7728), .A2(n6326), .ZN(n6199) );
  AOI21_X1 U7978 ( .B1(n7968), .B2(n6141), .A(n6199), .ZN(n7960) );
  NAND2_X1 U7979 ( .A1(n7961), .A2(n7960), .ZN(n7959) );
  INV_X1 U7980 ( .A(n6200), .ZN(n6202) );
  AND2_X1 U7981 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  NAND2_X1 U7982 ( .A1(n7946), .A2(n6203), .ZN(n8037) );
  NAND2_X1 U7983 ( .A1(n7959), .A2(n8037), .ZN(n6213) );
  NAND2_X1 U7984 ( .A1(n7821), .A2(n6331), .ZN(n6205) );
  NAND2_X1 U7985 ( .A1(n9489), .A2(n6141), .ZN(n6204) );
  NAND2_X1 U7986 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  XNOR2_X1 U7987 ( .A(n6206), .B(n6329), .ZN(n6208) );
  AND2_X1 U7988 ( .A1(n9489), .A2(n6307), .ZN(n6207) );
  AOI21_X1 U7989 ( .B1(n7821), .B2(n6141), .A(n6207), .ZN(n6209) );
  NAND2_X1 U7990 ( .A1(n6208), .A2(n6209), .ZN(n9339) );
  INV_X1 U7991 ( .A(n6208), .ZN(n6211) );
  INV_X1 U7992 ( .A(n6209), .ZN(n6210) );
  NAND2_X1 U7993 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  AND2_X1 U7994 ( .A1(n9339), .A2(n6212), .ZN(n8038) );
  NAND2_X1 U7995 ( .A1(n6213), .A2(n8038), .ZN(n8041) );
  NAND2_X1 U7996 ( .A1(n8041), .A2(n9339), .ZN(n6223) );
  NAND2_X1 U7997 ( .A1(n9338), .A2(n6331), .ZN(n6215) );
  NAND2_X1 U7998 ( .A1(n9488), .A2(n6141), .ZN(n6214) );
  NAND2_X1 U7999 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  XNOR2_X1 U8000 ( .A(n6216), .B(n6329), .ZN(n6218) );
  AND2_X1 U8001 ( .A1(n9488), .A2(n6307), .ZN(n6217) );
  AOI21_X1 U8002 ( .B1(n9338), .B2(n6141), .A(n6217), .ZN(n6219) );
  NAND2_X1 U8003 ( .A1(n6218), .A2(n6219), .ZN(n6224) );
  INV_X1 U8004 ( .A(n6218), .ZN(n6221) );
  INV_X1 U8005 ( .A(n6219), .ZN(n6220) );
  NAND2_X1 U8006 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  AND2_X1 U8007 ( .A1(n6224), .A2(n6222), .ZN(n9340) );
  NAND2_X1 U8008 ( .A1(n8082), .A2(n6331), .ZN(n6226) );
  OR2_X1 U8009 ( .A1(n8013), .A2(n4455), .ZN(n6225) );
  NAND2_X1 U8010 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  XNOR2_X1 U8011 ( .A(n6227), .B(n6318), .ZN(n6229) );
  NOR2_X1 U8012 ( .A1(n8013), .A2(n6326), .ZN(n6228) );
  AOI21_X1 U8013 ( .B1(n8082), .B2(n6141), .A(n6228), .ZN(n6230) );
  XNOR2_X1 U8014 ( .A(n6229), .B(n6230), .ZN(n9404) );
  INV_X1 U8015 ( .A(n6229), .ZN(n6231) );
  NAND2_X1 U8016 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  NAND2_X1 U8017 ( .A1(n9886), .A2(n6331), .ZN(n6234) );
  NAND2_X1 U8018 ( .A1(n9485), .A2(n6141), .ZN(n6233) );
  NAND2_X1 U8019 ( .A1(n6234), .A2(n6233), .ZN(n6235) );
  XNOR2_X1 U8020 ( .A(n6235), .B(n6318), .ZN(n9452) );
  NAND2_X1 U8021 ( .A1(n9886), .A2(n6141), .ZN(n6237) );
  NAND2_X1 U8022 ( .A1(n9485), .A2(n6307), .ZN(n6236) );
  NAND2_X1 U8023 ( .A1(n6237), .A2(n6236), .ZN(n9451) );
  NAND2_X1 U8024 ( .A1(n9963), .A2(n6141), .ZN(n6239) );
  NAND2_X1 U8025 ( .A1(n9486), .A2(n6307), .ZN(n6238) );
  NAND2_X1 U8026 ( .A1(n6239), .A2(n6238), .ZN(n6244) );
  NAND2_X1 U8027 ( .A1(n9963), .A2(n6331), .ZN(n6241) );
  NAND2_X1 U8028 ( .A1(n9486), .A2(n6141), .ZN(n6240) );
  NAND2_X1 U8029 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  XNOR2_X1 U8030 ( .A(n6242), .B(n6318), .ZN(n9276) );
  AOI22_X1 U8031 ( .A1(n9452), .A2(n9451), .B1(n6244), .B2(n9276), .ZN(n6243)
         );
  INV_X1 U8032 ( .A(n9276), .ZN(n9278) );
  INV_X1 U8033 ( .A(n6244), .ZN(n9279) );
  AND2_X1 U8034 ( .A1(n9278), .A2(n9279), .ZN(n6248) );
  INV_X1 U8035 ( .A(n6248), .ZN(n6245) );
  INV_X1 U8036 ( .A(n9451), .ZN(n6247) );
  INV_X1 U8037 ( .A(n9452), .ZN(n6246) );
  OAI21_X1 U8038 ( .B1(n6248), .B2(n6247), .A(n6246), .ZN(n6249) );
  NOR2_X1 U8039 ( .A1(n9456), .A2(n4455), .ZN(n6252) );
  AOI21_X1 U8040 ( .B1(n9867), .B2(n6331), .A(n6252), .ZN(n6253) );
  XNOR2_X1 U8041 ( .A(n6253), .B(n6318), .ZN(n6256) );
  NOR2_X1 U8042 ( .A1(n9456), .A2(n6326), .ZN(n6254) );
  AOI21_X1 U8043 ( .B1(n9867), .B2(n6141), .A(n6254), .ZN(n6255) );
  OR2_X1 U8044 ( .A1(n6256), .A2(n6255), .ZN(n9366) );
  AND2_X1 U8045 ( .A1(n6256), .A2(n6255), .ZN(n9365) );
  NAND2_X1 U8046 ( .A1(n9842), .A2(n6331), .ZN(n6258) );
  NAND2_X1 U8047 ( .A1(n9483), .A2(n6141), .ZN(n6257) );
  NAND2_X1 U8048 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  XNOR2_X1 U8049 ( .A(n6259), .B(n6329), .ZN(n6262) );
  AND2_X1 U8050 ( .A1(n9483), .A2(n6307), .ZN(n6260) );
  AOI21_X1 U8051 ( .B1(n9842), .B2(n6141), .A(n6260), .ZN(n6261) );
  NOR2_X1 U8052 ( .A1(n6262), .A2(n6261), .ZN(n9378) );
  NAND2_X1 U8053 ( .A1(n6262), .A2(n6261), .ZN(n9377) );
  NAND2_X1 U8054 ( .A1(n10006), .A2(n6331), .ZN(n6264) );
  NAND2_X1 U8055 ( .A1(n9481), .A2(n6141), .ZN(n6263) );
  NAND2_X1 U8056 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  XNOR2_X1 U8057 ( .A(n6265), .B(n6318), .ZN(n6276) );
  NAND2_X1 U8058 ( .A1(n10006), .A2(n6141), .ZN(n6267) );
  NAND2_X1 U8059 ( .A1(n9481), .A2(n6307), .ZN(n6266) );
  NAND2_X1 U8060 ( .A1(n6267), .A2(n6266), .ZN(n6277) );
  NAND2_X1 U8061 ( .A1(n6276), .A2(n6277), .ZN(n9307) );
  NAND2_X1 U8062 ( .A1(n9943), .A2(n6331), .ZN(n6269) );
  NAND2_X1 U8063 ( .A1(n9482), .A2(n6141), .ZN(n6268) );
  NAND2_X1 U8064 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  XNOR2_X1 U8065 ( .A(n6270), .B(n6329), .ZN(n9305) );
  NAND2_X1 U8066 ( .A1(n9943), .A2(n6141), .ZN(n6272) );
  NAND2_X1 U8067 ( .A1(n9482), .A2(n6307), .ZN(n6271) );
  AND2_X1 U8068 ( .A1(n6272), .A2(n6271), .ZN(n9304) );
  INV_X1 U8069 ( .A(n9307), .ZN(n6275) );
  NAND2_X1 U8070 ( .A1(n9305), .A2(n9304), .ZN(n6274) );
  INV_X1 U8071 ( .A(n6276), .ZN(n6279) );
  INV_X1 U8072 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U8073 ( .A1(n6279), .A2(n6278), .ZN(n9306) );
  NAND2_X1 U8074 ( .A1(n9791), .A2(n6331), .ZN(n6283) );
  NAND2_X1 U8075 ( .A1(n9480), .A2(n6141), .ZN(n6282) );
  NAND2_X1 U8076 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  XNOR2_X1 U8077 ( .A(n6284), .B(n6318), .ZN(n6288) );
  NAND2_X1 U8078 ( .A1(n9791), .A2(n6141), .ZN(n6286) );
  NAND2_X1 U8079 ( .A1(n9480), .A2(n6307), .ZN(n6285) );
  NAND2_X1 U8080 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  NAND2_X1 U8081 ( .A1(n6288), .A2(n6287), .ZN(n9395) );
  XOR2_X1 U8082 ( .A(n6290), .B(n6289), .Z(n9329) );
  OAI22_X1 U8083 ( .A1(n9995), .A2(n6317), .B1(n6291), .B2(n4455), .ZN(n6292)
         );
  XNOR2_X1 U8084 ( .A(n6292), .B(n6318), .ZN(n6293) );
  AOI22_X1 U8085 ( .A1(n9418), .A2(n6141), .B1(n6307), .B2(n9478), .ZN(n9414)
         );
  NAND2_X1 U8086 ( .A1(n9752), .A2(n6331), .ZN(n6295) );
  NAND2_X1 U8087 ( .A1(n9477), .A2(n6141), .ZN(n6294) );
  NAND2_X1 U8088 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U8089 ( .A(n6296), .B(n6329), .ZN(n6299) );
  AND2_X1 U8090 ( .A1(n9477), .A2(n6307), .ZN(n6297) );
  AOI21_X1 U8091 ( .B1(n9752), .B2(n6141), .A(n6297), .ZN(n6298) );
  NOR2_X1 U8092 ( .A1(n6299), .A2(n6298), .ZN(n9294) );
  NAND2_X1 U8093 ( .A1(n6299), .A2(n6298), .ZN(n9292) );
  AOI22_X1 U8094 ( .A1(n9736), .A2(n6331), .B1(n6141), .B2(n9476), .ZN(n6300)
         );
  XOR2_X1 U8095 ( .A(n6318), .B(n6300), .Z(n6302) );
  INV_X1 U8096 ( .A(n9736), .ZN(n9987) );
  OAI22_X1 U8097 ( .A1(n9987), .A2(n4455), .B1(n9358), .B2(n6326), .ZN(n6301)
         );
  NOR2_X1 U8098 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  AOI21_X1 U8099 ( .B1(n6302), .B2(n6301), .A(n6303), .ZN(n9388) );
  INV_X1 U8100 ( .A(n6303), .ZN(n6304) );
  OAI22_X1 U8101 ( .A1(n9983), .A2(n6317), .B1(n6305), .B2(n4455), .ZN(n6306)
         );
  XNOR2_X1 U8102 ( .A(n6306), .B(n6318), .ZN(n6313) );
  AND2_X1 U8103 ( .A1(n9475), .A2(n6307), .ZN(n6308) );
  AOI21_X1 U8104 ( .B1(n9357), .B2(n6141), .A(n6308), .ZN(n6314) );
  XNOR2_X1 U8105 ( .A(n6313), .B(n6314), .ZN(n9355) );
  NAND2_X1 U8106 ( .A1(n9706), .A2(n6331), .ZN(n6310) );
  NAND2_X1 U8107 ( .A1(n9474), .A2(n6141), .ZN(n6309) );
  NAND2_X1 U8108 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  XNOR2_X1 U8109 ( .A(n6311), .B(n6318), .ZN(n6324) );
  NOR2_X1 U8110 ( .A1(n9359), .A2(n6326), .ZN(n6312) );
  AOI21_X1 U8111 ( .B1(n9706), .B2(n6141), .A(n6312), .ZN(n6322) );
  XNOR2_X1 U8112 ( .A(n6324), .B(n6322), .ZN(n9436) );
  INV_X1 U8113 ( .A(n6313), .ZN(n6315) );
  NAND2_X1 U8114 ( .A1(n6315), .A2(n6314), .ZN(n9437) );
  OAI22_X1 U8115 ( .A1(n9975), .A2(n6317), .B1(n9438), .B2(n4455), .ZN(n6319)
         );
  XNOR2_X1 U8116 ( .A(n6319), .B(n6318), .ZN(n6321) );
  OAI22_X1 U8117 ( .A1(n9975), .A2(n4455), .B1(n9438), .B2(n6326), .ZN(n6320)
         );
  NOR2_X1 U8118 ( .A1(n6321), .A2(n6320), .ZN(n6343) );
  AOI21_X1 U8119 ( .B1(n6321), .B2(n6320), .A(n6343), .ZN(n9262) );
  INV_X1 U8120 ( .A(n6322), .ZN(n6323) );
  NAND2_X1 U8121 ( .A1(n6324), .A2(n6323), .ZN(n9263) );
  INV_X1 U8122 ( .A(n9265), .ZN(n6342) );
  INV_X1 U8123 ( .A(n6343), .ZN(n6341) );
  NAND2_X1 U8124 ( .A1(n6359), .A2(n6141), .ZN(n6328) );
  OR2_X1 U8125 ( .A1(n9266), .A2(n6326), .ZN(n6327) );
  NAND2_X1 U8126 ( .A1(n6328), .A2(n6327), .ZN(n6330) );
  XNOR2_X1 U8127 ( .A(n6330), .B(n6329), .ZN(n6335) );
  NAND2_X1 U8128 ( .A1(n6359), .A2(n6331), .ZN(n6332) );
  OAI21_X1 U8129 ( .B1(n9266), .B2(n4455), .A(n6332), .ZN(n6334) );
  XNOR2_X1 U8130 ( .A(n6335), .B(n6334), .ZN(n6344) );
  INV_X1 U8131 ( .A(n6344), .ZN(n6340) );
  INV_X1 U8132 ( .A(n6336), .ZN(n6338) );
  NAND2_X1 U8133 ( .A1(n7449), .A2(n10021), .ZN(n6352) );
  INV_X1 U8134 ( .A(n10020), .ZN(n8357) );
  NAND4_X1 U8135 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n9434), .ZN(n6365)
         );
  NAND3_X1 U8136 ( .A1(n6344), .A2(n6343), .A3(n9434), .ZN(n6361) );
  INV_X1 U8137 ( .A(n6350), .ZN(n6347) );
  NAND2_X1 U8138 ( .A1(n6345), .A2(n8300), .ZN(n7451) );
  INV_X1 U8139 ( .A(n7451), .ZN(n6346) );
  NAND2_X1 U8140 ( .A1(n6347), .A2(n6346), .ZN(n6349) );
  NAND2_X1 U8141 ( .A1(n10020), .A2(n8303), .ZN(n6348) );
  NOR2_X2 U8142 ( .A1(n6350), .A2(n8356), .ZN(n9460) );
  NAND2_X1 U8143 ( .A1(n8300), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7533) );
  NAND2_X1 U8144 ( .A1(n9964), .A2(n7533), .ZN(n6351) );
  NAND2_X1 U8145 ( .A1(n6352), .A2(n6351), .ZN(n7243) );
  AND3_X1 U8146 ( .A1(n6353), .A2(n6904), .A3(n7852), .ZN(n6354) );
  NAND2_X1 U8147 ( .A1(n7243), .A2(n6354), .ZN(n6355) );
  AOI22_X1 U8148 ( .A1(n9675), .A2(n9442), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6356) );
  OAI21_X1 U8149 ( .B1(n6357), .B2(n9444), .A(n6356), .ZN(n6358) );
  AOI21_X1 U8150 ( .B1(n6359), .B2(n9465), .A(n6358), .ZN(n6360) );
  NAND2_X1 U8151 ( .A1(n6365), .A2(n6364), .ZN(P1_U3220) );
  INV_X1 U8152 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6735) );
  INV_X1 U8153 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6375) );
  INV_X1 U8154 ( .A(n6613), .ZN(n6378) );
  INV_X1 U8155 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U8156 ( .A1(n4497), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8157 ( .A1(n6643), .A2(n6379), .ZN(n8987) );
  NAND2_X2 U8158 ( .A1(n6384), .A2(n6383), .ZN(n6424) );
  NAND2_X1 U8159 ( .A1(n8987), .A2(n6688), .ZN(n6389) );
  INV_X1 U8160 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U8161 ( .A1(n7927), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8162 ( .A1(n4467), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6385) );
  OAI211_X1 U8163 ( .C1(n7928), .C2(n10284), .A(n6386), .B(n6385), .ZN(n6387)
         );
  INV_X1 U8164 ( .A(n6387), .ZN(n6388) );
  INV_X2 U8165 ( .A(n6453), .ZN(n6486) );
  NAND2_X1 U8166 ( .A1(n7996), .A2(n6486), .ZN(n6392) );
  NAND2_X1 U8167 ( .A1(n6672), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6391) );
  INV_X1 U8168 ( .A(n8510), .ZN(n9185) );
  INV_X1 U8169 ( .A(n7016), .ZN(n7409) );
  NAND2_X1 U8170 ( .A1(n6422), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6397) );
  INV_X1 U8171 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6394) );
  INV_X1 U8172 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7170) );
  OR2_X1 U8173 ( .A1(n6424), .A2(n7170), .ZN(n6398) );
  NAND2_X1 U8174 ( .A1(n6422), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6405) );
  OR2_X1 U8175 ( .A1(n6401), .A2(n6400), .ZN(n6404) );
  INV_X1 U8176 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U8177 ( .A1(n6407), .A2(n6406), .ZN(n6736) );
  INV_X1 U8178 ( .A(SI_0_), .ZN(n6408) );
  OR2_X1 U8179 ( .A1(n4464), .A2(n6408), .ZN(n6410) );
  INV_X1 U8180 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6409) );
  XNOR2_X1 U8181 ( .A(n6410), .B(n6409), .ZN(n9260) );
  MUX2_X1 U8182 ( .A(n6411), .B(n9260), .S(n6816), .Z(n7312) );
  NAND2_X1 U8183 ( .A1(n7404), .A2(n4678), .ZN(n7403) );
  NAND2_X1 U8184 ( .A1(n10126), .A2(n7016), .ZN(n10129) );
  NAND2_X1 U8185 ( .A1(n7402), .A2(n10129), .ZN(n6420) );
  NAND2_X1 U8186 ( .A1(n6422), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6417) );
  OR2_X1 U8187 ( .A1(n6424), .A2(n7184), .ZN(n6416) );
  INV_X1 U8188 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10143) );
  OR2_X1 U8189 ( .A1(n6412), .A2(n10143), .ZN(n6415) );
  OR2_X1 U8190 ( .A1(n6401), .A2(n6413), .ZN(n6414) );
  OR2_X1 U8191 ( .A1(n6430), .A2(n6866), .ZN(n6418) );
  NAND2_X1 U8192 ( .A1(n7383), .A2(n10150), .ZN(n8631) );
  NAND2_X1 U8193 ( .A1(n8632), .A2(n8631), .ZN(n10119) );
  NAND2_X1 U8194 ( .A1(n7406), .A2(n4567), .ZN(n6421) );
  NAND2_X1 U8195 ( .A1(n10134), .A2(n6421), .ZN(n7381) );
  INV_X1 U8196 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6423) );
  OR2_X1 U8197 ( .A1(n6680), .A2(n6423), .ZN(n6429) );
  INV_X1 U8198 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6425) );
  OR2_X1 U8199 ( .A1(n6401), .A2(n6425), .ZN(n6426) );
  OR2_X1 U8200 ( .A1(n6453), .A2(n6877), .ZN(n6432) );
  OR2_X1 U8201 ( .A1(n6430), .A2(n5188), .ZN(n6431) );
  OAI211_X1 U8202 ( .C1(n6816), .C2(n7071), .A(n6432), .B(n6431), .ZN(n7084)
         );
  NAND2_X1 U8203 ( .A1(n8791), .A2(n7084), .ZN(n6433) );
  NAND2_X1 U8204 ( .A1(n7381), .A2(n6433), .ZN(n6435) );
  OR2_X1 U8205 ( .A1(n8791), .A2(n7084), .ZN(n6434) );
  NAND2_X1 U8206 ( .A1(n4467), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8207 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6437) );
  AND2_X1 U8208 ( .A1(n6446), .A2(n6437), .ZN(n7629) );
  OR2_X1 U8209 ( .A1(n6424), .A2(n7629), .ZN(n6440) );
  INV_X1 U8210 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6438) );
  NAND4_X4 U8211 ( .A1(n6442), .A2(n6441), .A3(n6440), .A4(n6439), .ZN(n8790)
         );
  OR2_X1 U8212 ( .A1(n6453), .A2(n6879), .ZN(n6444) );
  OR2_X1 U8213 ( .A1(n6430), .A2(n6867), .ZN(n6443) );
  NAND2_X1 U8214 ( .A1(n7927), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6452) );
  INV_X1 U8215 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10303) );
  OR2_X1 U8216 ( .A1(n4451), .A2(n10303), .ZN(n6451) );
  NAND2_X1 U8217 ( .A1(n6446), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6447) );
  AND2_X1 U8218 ( .A1(n6457), .A2(n6447), .ZN(n7149) );
  OR2_X1 U8219 ( .A1(n6424), .A2(n7149), .ZN(n6450) );
  INV_X1 U8220 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8221 ( .A1(n7928), .A2(n6448), .ZN(n6449) );
  NAND4_X1 U8222 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n8789)
         );
  OR2_X1 U8223 ( .A1(n6874), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8224 ( .A1(n4463), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U8225 ( .A1(n8789), .A2(n6739), .ZN(n6456) );
  NAND2_X1 U8226 ( .A1(n4467), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8227 ( .A1(n6457), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6458) );
  AND2_X1 U8228 ( .A1(n6469), .A2(n6458), .ZN(n10110) );
  OR2_X1 U8229 ( .A1(n6424), .A2(n10110), .ZN(n6462) );
  INV_X1 U8230 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6459) );
  OR2_X1 U8231 ( .A1(n6680), .A2(n6459), .ZN(n6461) );
  OR2_X1 U8232 ( .A1(n7928), .A2(n10185), .ZN(n6460) );
  NAND4_X1 U8233 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n8788)
         );
  NAND2_X1 U8234 ( .A1(n6870), .A2(n6486), .ZN(n6465) );
  AOI22_X1 U8235 ( .A1(n6672), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10084), .B2(
        n6599), .ZN(n6464) );
  NAND2_X1 U8236 ( .A1(n6465), .A2(n6464), .ZN(n7268) );
  OR2_X1 U8237 ( .A1(n8788), .A2(n7268), .ZN(n8595) );
  NAND2_X1 U8238 ( .A1(n8788), .A2(n7268), .ZN(n8594) );
  NAND2_X1 U8239 ( .A1(n6466), .A2(n8594), .ZN(n7435) );
  INV_X1 U8240 ( .A(n7435), .ZN(n6477) );
  NAND2_X1 U8241 ( .A1(n6893), .A2(n6486), .ZN(n6468) );
  AOI22_X1 U8242 ( .A1(n6672), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7162), .B2(
        n6599), .ZN(n6467) );
  NAND2_X1 U8243 ( .A1(n6468), .A2(n6467), .ZN(n7392) );
  NAND2_X1 U8244 ( .A1(n4467), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6475) );
  OR2_X1 U8245 ( .A1(n6680), .A2(n10179), .ZN(n6474) );
  NAND2_X1 U8246 ( .A1(n6469), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6470) );
  AND2_X1 U8247 ( .A1(n6491), .A2(n6470), .ZN(n7439) );
  OR2_X1 U8248 ( .A1(n6424), .A2(n7439), .ZN(n6473) );
  INV_X1 U8249 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6471) );
  OR2_X1 U8250 ( .A1(n7928), .A2(n6471), .ZN(n6472) );
  NAND4_X1 U8251 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n8787)
         );
  INV_X1 U8252 ( .A(n8787), .ZN(n10109) );
  OR2_X1 U8253 ( .A1(n7392), .A2(n10109), .ZN(n8660) );
  NAND2_X1 U8254 ( .A1(n7392), .A2(n10109), .ZN(n8644) );
  NAND2_X1 U8255 ( .A1(n6895), .A2(n6486), .ZN(n6480) );
  AOI22_X1 U8256 ( .A1(n6672), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6478), .B2(
        n6599), .ZN(n6479) );
  NAND2_X1 U8257 ( .A1(n6480), .A2(n6479), .ZN(n7559) );
  NAND2_X1 U8258 ( .A1(n6677), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6485) );
  OR2_X1 U8259 ( .A1(n4612), .A2(n7524), .ZN(n6484) );
  NAND2_X1 U8260 ( .A1(n4533), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6481) );
  AND2_X1 U8261 ( .A1(n6497), .A2(n6481), .ZN(n7920) );
  OR2_X1 U8262 ( .A1(n6424), .A2(n7920), .ZN(n6483) );
  INV_X1 U8263 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10370) );
  OR2_X1 U8264 ( .A1(n6680), .A2(n10370), .ZN(n6482) );
  NAND2_X1 U8265 ( .A1(n7559), .A2(n7862), .ZN(n8646) );
  NAND2_X1 U8266 ( .A1(n6888), .A2(n6486), .ZN(n6489) );
  AOI22_X1 U8267 ( .A1(n6672), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6487), .B2(
        n6599), .ZN(n6488) );
  NAND2_X1 U8268 ( .A1(n4467), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6496) );
  OR2_X1 U8269 ( .A1(n7928), .A2(n7502), .ZN(n6495) );
  XNOR2_X1 U8270 ( .A(n6491), .B(n6490), .ZN(n7539) );
  OR2_X1 U8271 ( .A1(n6424), .A2(n7539), .ZN(n6494) );
  INV_X1 U8272 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6492) );
  OR2_X1 U8273 ( .A1(n6680), .A2(n6492), .ZN(n6493) );
  NAND4_X1 U8274 ( .A1(n6496), .A2(n6495), .A3(n6494), .A4(n6493), .ZN(n8786)
         );
  AND2_X1 U8275 ( .A1(n7541), .A2(n8786), .ZN(n6507) );
  INV_X1 U8276 ( .A(n6507), .ZN(n7801) );
  NAND2_X1 U8277 ( .A1(n8601), .A2(n7801), .ZN(n7637) );
  NAND2_X1 U8278 ( .A1(n6677), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6503) );
  OR2_X1 U8279 ( .A1(n4612), .A2(n7756), .ZN(n6502) );
  NAND2_X1 U8280 ( .A1(n6497), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6498) );
  AND2_X1 U8281 ( .A1(n6517), .A2(n6498), .ZN(n7907) );
  OR2_X1 U8282 ( .A1(n6424), .A2(n7907), .ZN(n6501) );
  INV_X1 U8283 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6499) );
  OR2_X1 U8284 ( .A1(n6680), .A2(n6499), .ZN(n6500) );
  NAND4_X1 U8285 ( .A1(n6503), .A2(n6502), .A3(n6501), .A4(n6500), .ZN(n8784)
         );
  NAND2_X1 U8286 ( .A1(n6909), .A2(n6486), .ZN(n6506) );
  AOI22_X1 U8287 ( .A1(n6672), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6504), .B2(
        n6599), .ZN(n6505) );
  OR2_X1 U8288 ( .A1(n7541), .A2(n7805), .ZN(n8661) );
  NAND2_X1 U8289 ( .A1(n7541), .A2(n7805), .ZN(n8645) );
  NOR2_X1 U8290 ( .A1(n8599), .A2(n6507), .ZN(n6509) );
  NOR2_X1 U8291 ( .A1(n7559), .A2(n8785), .ZN(n6508) );
  AOI21_X1 U8292 ( .B1(n8601), .B2(n6509), .A(n6508), .ZN(n7636) );
  OR2_X1 U8293 ( .A1(n7392), .A2(n8787), .ZN(n7419) );
  OR2_X1 U8294 ( .A1(n7637), .A2(n7419), .ZN(n6510) );
  NAND2_X1 U8295 ( .A1(n7909), .A2(n8784), .ZN(n6512) );
  NAND2_X1 U8296 ( .A1(n6959), .A2(n6486), .ZN(n6516) );
  AOI22_X1 U8297 ( .A1(n6672), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6514), .B2(
        n6599), .ZN(n6515) );
  NAND2_X1 U8298 ( .A1(n4467), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6523) );
  OR2_X1 U8299 ( .A1(n7928), .A2(n10316), .ZN(n6522) );
  NAND2_X1 U8300 ( .A1(n6517), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6518) );
  AND2_X1 U8301 ( .A1(n6528), .A2(n6518), .ZN(n7991) );
  OR2_X1 U8302 ( .A1(n6424), .A2(n7991), .ZN(n6521) );
  INV_X1 U8303 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6519) );
  OR2_X1 U8304 ( .A1(n6680), .A2(n6519), .ZN(n6520) );
  NAND4_X1 U8305 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n8783)
         );
  AND2_X1 U8306 ( .A1(n7993), .A2(n8783), .ZN(n6524) );
  NAND2_X1 U8307 ( .A1(n6966), .A2(n6486), .ZN(n6527) );
  AOI22_X1 U8308 ( .A1(n6672), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6525), .B2(
        n6599), .ZN(n6526) );
  NAND2_X1 U8309 ( .A1(n4467), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6533) );
  INV_X1 U8310 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10478) );
  OR2_X1 U8311 ( .A1(n7928), .A2(n10478), .ZN(n6532) );
  NAND2_X1 U8312 ( .A1(n6528), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6529) );
  AND2_X1 U8313 ( .A1(n6538), .A2(n6529), .ZN(n7878) );
  OR2_X1 U8314 ( .A1(n6424), .A2(n7878), .ZN(n6531) );
  INV_X1 U8315 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10400) );
  OR2_X1 U8316 ( .A1(n6680), .A2(n10400), .ZN(n6530) );
  NAND4_X1 U8317 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n8782)
         );
  NOR2_X1 U8318 ( .A1(n7875), .A2(n8782), .ZN(n6534) );
  NAND2_X1 U8319 ( .A1(n6985), .A2(n6486), .ZN(n6537) );
  AOI22_X1 U8320 ( .A1(n6672), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6535), .B2(
        n6599), .ZN(n6536) );
  NAND2_X1 U8321 ( .A1(n4467), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6543) );
  INV_X1 U8322 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10381) );
  OR2_X1 U8323 ( .A1(n7928), .A2(n10381), .ZN(n6542) );
  NAND2_X1 U8324 ( .A1(n6538), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6539) );
  AND2_X1 U8325 ( .A1(n6548), .A2(n6539), .ZN(n8062) );
  OR2_X1 U8326 ( .A1(n6424), .A2(n8062), .ZN(n6541) );
  INV_X1 U8327 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7917) );
  OR2_X1 U8328 ( .A1(n6680), .A2(n7917), .ZN(n6540) );
  OR2_X1 U8329 ( .A1(n8065), .A2(n8111), .ZN(n8676) );
  NAND2_X1 U8330 ( .A1(n8065), .A2(n8111), .ZN(n8675) );
  NAND2_X1 U8331 ( .A1(n8676), .A2(n8675), .ZN(n8672) );
  INV_X1 U8332 ( .A(n8111), .ZN(n8781) );
  NAND2_X1 U8333 ( .A1(n8065), .A2(n8781), .ZN(n6544) );
  NAND2_X1 U8334 ( .A1(n7105), .A2(n6486), .ZN(n6547) );
  AOI22_X1 U8335 ( .A1(n7106), .A2(n6599), .B1(n6672), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8336 ( .A1(n6548), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8337 ( .A1(n6558), .A2(n6549), .ZN(n8108) );
  NAND2_X1 U8338 ( .A1(n6688), .A2(n8108), .ZN(n6553) );
  OR2_X1 U8339 ( .A1(n4612), .A2(n10412), .ZN(n6552) );
  OR2_X1 U8340 ( .A1(n7928), .A2(n9153), .ZN(n6551) );
  INV_X1 U8341 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9238) );
  OR2_X1 U8342 ( .A1(n6680), .A2(n9238), .ZN(n6550) );
  NAND4_X1 U8343 ( .A1(n6553), .A2(n6552), .A3(n6551), .A4(n6550), .ZN(n8780)
         );
  XNOR2_X1 U8344 ( .A(n9239), .B(n9103), .ZN(n8674) );
  NAND2_X1 U8345 ( .A1(n9239), .A2(n8780), .ZN(n6554) );
  AOI22_X1 U8346 ( .A1(n6556), .A2(n6599), .B1(n6672), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6557) );
  INV_X1 U8347 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U8348 ( .A1(n6558), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8349 ( .A1(n6568), .A2(n6559), .ZN(n9105) );
  NAND2_X1 U8350 ( .A1(n9105), .A2(n6688), .ZN(n6563) );
  NAND2_X1 U8351 ( .A1(n6677), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8352 ( .A1(n4467), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6560) );
  AND2_X1 U8353 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  OAI211_X1 U8354 ( .C1(n6680), .C2(n6564), .A(n6563), .B(n6562), .ZN(n9091)
         );
  INV_X1 U8355 ( .A(n9091), .ZN(n8489) );
  NAND2_X1 U8356 ( .A1(n9149), .A2(n8489), .ZN(n6744) );
  NAND2_X1 U8357 ( .A1(n9073), .A2(n6744), .ZN(n9101) );
  NAND2_X1 U8358 ( .A1(n9149), .A2(n9091), .ZN(n6565) );
  NAND2_X1 U8359 ( .A1(n7254), .A2(n6486), .ZN(n6567) );
  AOI22_X1 U8360 ( .A1(n7255), .A2(n6599), .B1(P1_DATAO_REG_16__SCAN_IN), .B2(
        n6672), .ZN(n6566) );
  NAND2_X1 U8361 ( .A1(n6568), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8362 ( .A1(n4496), .A2(n6569), .ZN(n9095) );
  NAND2_X1 U8363 ( .A1(n9095), .A2(n6688), .ZN(n6571) );
  AOI22_X1 U8364 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n4467), .B1(n7927), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6570) );
  OR2_X1 U8365 ( .A1(n9231), .A2(n9104), .ZN(n8687) );
  NAND2_X1 U8366 ( .A1(n9231), .A2(n9104), .ZN(n9076) );
  NAND2_X1 U8367 ( .A1(n8687), .A2(n9076), .ZN(n9089) );
  NAND2_X1 U8368 ( .A1(n9231), .A2(n9081), .ZN(n6572) );
  NAND2_X1 U8369 ( .A1(n7292), .A2(n6486), .ZN(n6576) );
  AOI22_X1 U8370 ( .A1(n6574), .A2(n6599), .B1(n6672), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6575) );
  INV_X1 U8371 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U8372 ( .A1(n4496), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U8373 ( .A1(n6584), .A2(n6577), .ZN(n9084) );
  NAND2_X1 U8374 ( .A1(n9084), .A2(n6688), .ZN(n6579) );
  AOI22_X1 U8375 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n6677), .B1(n4467), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6578) );
  INV_X1 U8376 ( .A(n9092), .ZN(n8392) );
  OR2_X1 U8377 ( .A1(n9225), .A2(n8392), .ZN(n8691) );
  NAND2_X1 U8378 ( .A1(n9225), .A2(n8392), .ZN(n8693) );
  NAND2_X1 U8379 ( .A1(n8691), .A2(n8693), .ZN(n9077) );
  AND2_X1 U8380 ( .A1(n9225), .A2(n9092), .ZN(n6580) );
  NAND2_X1 U8381 ( .A1(n7315), .A2(n6486), .ZN(n6583) );
  AOI22_X1 U8382 ( .A1(n6581), .A2(n6599), .B1(n6672), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U8383 ( .A1(n6584), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U8384 ( .A1(n6602), .A2(n6585), .ZN(n9070) );
  NAND2_X1 U8385 ( .A1(n9070), .A2(n6688), .ZN(n6590) );
  NAND2_X1 U8386 ( .A1(n7927), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U8387 ( .A1(n4467), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6586) );
  OAI211_X1 U8388 ( .C1(n7928), .C2(n9138), .A(n6587), .B(n6586), .ZN(n6588)
         );
  INV_X1 U8389 ( .A(n6588), .ZN(n6589) );
  NAND2_X1 U8390 ( .A1(n9219), .A2(n8466), .ZN(n8694) );
  NAND2_X1 U8391 ( .A1(n8363), .A2(n6486), .ZN(n6592) );
  NAND2_X1 U8392 ( .A1(n6672), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6591) );
  NAND2_X2 U8393 ( .A1(n6592), .A2(n6591), .ZN(n6610) );
  NAND2_X1 U8394 ( .A1(n6604), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8395 ( .A1(n6613), .A2(n6593), .ZN(n9046) );
  NAND2_X1 U8396 ( .A1(n9046), .A2(n6688), .ZN(n6598) );
  INV_X1 U8397 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U8398 ( .A1(n6677), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8399 ( .A1(n7927), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6594) );
  OAI211_X1 U8400 ( .C1(n4612), .C2(n9045), .A(n6595), .B(n6594), .ZN(n6596)
         );
  INV_X1 U8401 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U8402 ( .A1(n6610), .A2(n8401), .ZN(n8710) );
  NAND2_X1 U8403 ( .A1(n7427), .A2(n6486), .ZN(n6601) );
  AOI22_X1 U8404 ( .A1(n6672), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8584), .B2(
        n6599), .ZN(n6600) );
  NAND2_X1 U8405 ( .A1(n6602), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8406 ( .A1(n6604), .A2(n6603), .ZN(n9059) );
  NAND2_X1 U8407 ( .A1(n9059), .A2(n6688), .ZN(n6609) );
  INV_X1 U8408 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U8409 ( .A1(n6677), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8410 ( .A1(n7927), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6605) );
  OAI211_X1 U8411 ( .C1(n4612), .C2(n10366), .A(n6606), .B(n6605), .ZN(n6607)
         );
  INV_X1 U8412 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8413 ( .A1(n9060), .A2(n9067), .ZN(n9039) );
  INV_X1 U8414 ( .A(n9067), .ZN(n8542) );
  NAND2_X1 U8415 ( .A1(n9060), .A2(n8542), .ZN(n6747) );
  NAND2_X1 U8416 ( .A1(n9021), .A2(n6747), .ZN(n9052) );
  OR2_X1 U8417 ( .A1(n9219), .A2(n9082), .ZN(n9053) );
  NAND2_X1 U8418 ( .A1(n9052), .A2(n9053), .ZN(n9027) );
  NAND3_X1 U8419 ( .A1(n9041), .A2(n9039), .A3(n9027), .ZN(n6611) );
  OR2_X1 U8420 ( .A1(n6610), .A2(n9054), .ZN(n9029) );
  NOR2_X1 U8421 ( .A1(n6430), .A2(n10313), .ZN(n6612) );
  NAND2_X1 U8422 ( .A1(n6613), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U8423 ( .A1(n6620), .A2(n6614), .ZN(n9035) );
  INV_X1 U8424 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9201) );
  NAND2_X1 U8425 ( .A1(n4467), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8426 ( .A1(n6677), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6615) );
  OAI211_X1 U8427 ( .C1(n9201), .C2(n6680), .A(n6616), .B(n6615), .ZN(n6617)
         );
  OR2_X1 U8428 ( .A1(n8472), .A2(n9043), .ZN(n8711) );
  NAND2_X1 U8429 ( .A1(n8472), .A2(n9043), .ZN(n8713) );
  NAND2_X1 U8430 ( .A1(n8711), .A2(n8713), .ZN(n8589) );
  NAND2_X1 U8431 ( .A1(n8472), .A2(n8527), .ZN(n9011) );
  NAND2_X1 U8432 ( .A1(n7796), .A2(n6486), .ZN(n6619) );
  OR2_X1 U8433 ( .A1(n6430), .A2(n10302), .ZN(n6618) );
  NAND2_X1 U8434 ( .A1(n6620), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U8435 ( .A1(n4525), .A2(n6621), .ZN(n9017) );
  NAND2_X1 U8436 ( .A1(n9017), .A2(n6688), .ZN(n6626) );
  INV_X1 U8437 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U8438 ( .A1(n6677), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8439 ( .A1(n4467), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6622) );
  OAI211_X1 U8440 ( .C1(n9195), .C2(n6680), .A(n6623), .B(n6622), .ZN(n6624)
         );
  INV_X1 U8441 ( .A(n6624), .ZN(n6625) );
  NAND2_X1 U8442 ( .A1(n9196), .A2(n9000), .ZN(n8715) );
  NAND2_X1 U8443 ( .A1(n8617), .A2(n8715), .ZN(n6751) );
  NAND2_X1 U8444 ( .A1(n6627), .A2(n6751), .ZN(n9009) );
  OR2_X1 U8445 ( .A1(n9196), .A2(n9032), .ZN(n6628) );
  NAND2_X1 U8446 ( .A1(n7843), .A2(n6486), .ZN(n6630) );
  NAND2_X1 U8447 ( .A1(n6672), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U8448 ( .A1(n4525), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8449 ( .A1(n4497), .A2(n6631), .ZN(n9005) );
  NAND2_X1 U8450 ( .A1(n9005), .A2(n6688), .ZN(n6636) );
  INV_X1 U8451 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U8452 ( .A1(n4467), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8453 ( .A1(n6677), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6632) );
  OAI211_X1 U8454 ( .C1(n6680), .C2(n10497), .A(n6633), .B(n6632), .ZN(n6634)
         );
  INV_X1 U8455 ( .A(n6634), .ZN(n6635) );
  NAND2_X1 U8456 ( .A1(n9190), .A2(n9014), .ZN(n6638) );
  NOR2_X1 U8457 ( .A1(n9190), .A2(n9014), .ZN(n6637) );
  NAND2_X1 U8458 ( .A1(n8027), .A2(n6486), .ZN(n6640) );
  NAND2_X1 U8459 ( .A1(n4463), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6639) );
  INV_X1 U8460 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8461 ( .A1(n6643), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8462 ( .A1(n6652), .A2(n6644), .ZN(n8977) );
  NAND2_X1 U8463 ( .A1(n8977), .A2(n6688), .ZN(n6649) );
  INV_X1 U8464 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U8465 ( .A1(n4467), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8466 ( .A1(n6677), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6645) );
  OAI211_X1 U8467 ( .C1(n6680), .C2(n9179), .A(n6646), .B(n6645), .ZN(n6647)
         );
  INV_X1 U8468 ( .A(n6647), .ZN(n6648) );
  INV_X1 U8469 ( .A(n9180), .ZN(n9118) );
  NAND2_X1 U8470 ( .A1(n8099), .A2(n6486), .ZN(n6651) );
  OR2_X1 U8471 ( .A1(n6430), .A2(n10429), .ZN(n6650) );
  NAND2_X1 U8472 ( .A1(n6652), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6653) );
  INV_X1 U8473 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U8474 ( .A1(n6677), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8475 ( .A1(n7927), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6654) );
  OAI211_X1 U8476 ( .C1(n4612), .C2(n8968), .A(n6655), .B(n6654), .ZN(n6656)
         );
  NAND2_X1 U8477 ( .A1(n6657), .A2(n8975), .ZN(n6658) );
  NAND2_X1 U8478 ( .A1(n8970), .A2(n8777), .ZN(n6659) );
  NAND2_X1 U8479 ( .A1(n8445), .A2(n6486), .ZN(n6662) );
  NAND2_X1 U8480 ( .A1(n6672), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6661) );
  INV_X1 U8481 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8482 ( .A1(n6665), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8483 ( .A1(n6675), .A2(n6666), .ZN(n8955) );
  NAND2_X1 U8484 ( .A1(n8955), .A2(n6688), .ZN(n6671) );
  INV_X1 U8485 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U8486 ( .A1(n6677), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U8487 ( .A1(n4467), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6667) );
  OAI211_X1 U8488 ( .C1(n10371), .C2(n6680), .A(n6668), .B(n6667), .ZN(n6669)
         );
  INV_X1 U8489 ( .A(n6669), .ZN(n6670) );
  NAND2_X1 U8490 ( .A1(n8451), .A2(n8966), .ZN(n8735) );
  NAND2_X1 U8491 ( .A1(n8379), .A2(n6486), .ZN(n6674) );
  NAND2_X1 U8492 ( .A1(n6672), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8493 ( .A1(n6675), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8494 ( .A1(n8942), .A2(n6676), .ZN(n8428) );
  NAND2_X1 U8495 ( .A1(n8428), .A2(n6688), .ZN(n6683) );
  INV_X1 U8496 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U8497 ( .A1(n4467), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8498 ( .A1(n6677), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6678) );
  OAI211_X1 U8499 ( .C1(n9166), .C2(n6680), .A(n6679), .B(n6678), .ZN(n6681)
         );
  INV_X1 U8500 ( .A(n6681), .ZN(n6682) );
  NAND2_X1 U8501 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  OR2_X1 U8502 ( .A1(n7810), .A2(n8365), .ZN(n6687) );
  NAND2_X1 U8503 ( .A1(n8771), .A2(n8584), .ZN(n6789) );
  INV_X1 U8504 ( .A(n8942), .ZN(n6689) );
  NAND2_X1 U8505 ( .A1(n6689), .A2(n6688), .ZN(n7933) );
  INV_X1 U8506 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U8507 ( .A1(n4467), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8508 ( .A1(n7927), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6691) );
  OAI211_X1 U8509 ( .C1(n10300), .C2(n7928), .A(n6692), .B(n6691), .ZN(n6693)
         );
  INV_X1 U8510 ( .A(n6693), .ZN(n6694) );
  NAND2_X1 U8511 ( .A1(n7933), .A2(n6694), .ZN(n8774) );
  INV_X1 U8512 ( .A(n6003), .ZN(n8767) );
  NAND2_X1 U8513 ( .A1(n8767), .A2(n6695), .ZN(n6696) );
  NAND2_X1 U8514 ( .A1(n8774), .A2(n6698), .ZN(n6700) );
  NAND2_X1 U8515 ( .A1(n8029), .A2(n8100), .ZN(n6713) );
  NAND2_X1 U8516 ( .A1(n6703), .A2(P2_B_REG_SCAN_IN), .ZN(n6706) );
  INV_X1 U8517 ( .A(P2_B_REG_SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8518 ( .A1(n6704), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6705) );
  NAND3_X1 U8519 ( .A1(n6706), .A2(n6705), .A3(P2_IR_REG_25__SCAN_IN), .ZN(
        n6710) );
  OAI21_X1 U8520 ( .B1(n6706), .B2(P2_IR_REG_25__SCAN_IN), .A(n6705), .ZN(
        n6707) );
  NAND2_X1 U8521 ( .A1(n6711), .A2(n6707), .ZN(n6708) );
  OR2_X1 U8522 ( .A1(n6714), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U8523 ( .A1(n7998), .A2(n8100), .ZN(n6920) );
  OAI211_X1 U8524 ( .C1(n8763), .C2(n6697), .A(n6767), .B(n7844), .ZN(n6993)
         );
  NOR2_X1 U8525 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n6719) );
  NOR4_X1 U8526 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6718) );
  NOR4_X1 U8527 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6717) );
  NOR4_X1 U8528 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6716) );
  NAND4_X1 U8529 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6725)
         );
  NOR4_X1 U8530 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6723) );
  NOR4_X1 U8531 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6722) );
  NOR4_X1 U8532 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6721) );
  NOR4_X1 U8533 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6720) );
  NAND4_X1 U8534 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6724)
         );
  NOR2_X1 U8535 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  NAND2_X1 U8536 ( .A1(n6792), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6727) );
  INV_X1 U8537 ( .A(n8771), .ZN(n7797) );
  NAND2_X1 U8538 ( .A1(n10151), .A2(n7810), .ZN(n6768) );
  NAND2_X1 U8539 ( .A1(n6768), .A2(n7013), .ZN(n6730) );
  XNOR2_X1 U8540 ( .A(n6728), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8613) );
  AND2_X1 U8541 ( .A1(n8771), .A2(n8612), .ZN(n6752) );
  NAND2_X1 U8542 ( .A1(n8613), .A2(n6752), .ZN(n6729) );
  NAND2_X1 U8543 ( .A1(n6730), .A2(n6762), .ZN(n6733) );
  INV_X1 U8544 ( .A(n6762), .ZN(n6731) );
  NAND2_X1 U8545 ( .A1(n6884), .A2(n6731), .ZN(n6732) );
  NAND2_X1 U8546 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  MUX2_X1 U8547 ( .A(n6735), .B(n9165), .S(n10189), .Z(n6759) );
  INV_X1 U8548 ( .A(n6736), .ZN(n6737) );
  INV_X1 U8549 ( .A(n10116), .ZN(n8626) );
  NAND2_X1 U8550 ( .A1(n8791), .A2(n10157), .ZN(n8651) );
  OR2_X1 U8551 ( .A1(n8790), .A2(n8638), .ZN(n8652) );
  NAND2_X1 U8552 ( .A1(n7233), .A2(n8652), .ZN(n7412) );
  INV_X1 U8553 ( .A(n6739), .ZN(n6740) );
  OR2_X1 U8554 ( .A1(n8789), .A2(n6740), .ZN(n10102) );
  NAND2_X1 U8555 ( .A1(n8789), .A2(n6740), .ZN(n8655) );
  INV_X1 U8556 ( .A(n7268), .ZN(n10167) );
  OR2_X1 U8557 ( .A1(n10167), .A2(n8788), .ZN(n8658) );
  AND2_X1 U8558 ( .A1(n8658), .A2(n10102), .ZN(n8642) );
  NAND2_X1 U8559 ( .A1(n10103), .A2(n8642), .ZN(n6741) );
  NAND2_X1 U8560 ( .A1(n10167), .A2(n8788), .ZN(n8656) );
  NAND2_X1 U8561 ( .A1(n6741), .A2(n8656), .ZN(n7432) );
  NAND2_X1 U8562 ( .A1(n7432), .A2(n8598), .ZN(n7431) );
  NAND2_X1 U8563 ( .A1(n7431), .A2(n8660), .ZN(n7423) );
  OR2_X1 U8564 ( .A1(n7909), .A2(n7869), .ZN(n8663) );
  NAND2_X1 U8565 ( .A1(n7909), .A2(n7869), .ZN(n8666) );
  NAND2_X1 U8566 ( .A1(n8663), .A2(n8666), .ZN(n7639) );
  INV_X1 U8567 ( .A(n8783), .ZN(n7904) );
  NAND2_X1 U8568 ( .A1(n4615), .A2(n7904), .ZN(n8620) );
  INV_X1 U8569 ( .A(n8782), .ZN(n8053) );
  OR2_X1 U8570 ( .A1(n7875), .A2(n8053), .ZN(n8618) );
  NAND2_X1 U8571 ( .A1(n7875), .A2(n8053), .ZN(n8621) );
  NAND2_X1 U8572 ( .A1(n8618), .A2(n8621), .ZN(n8591) );
  INV_X1 U8573 ( .A(n8591), .ZN(n6742) );
  NAND2_X1 U8574 ( .A1(n9239), .A2(n9103), .ZN(n8681) );
  INV_X1 U8575 ( .A(n6744), .ZN(n8684) );
  INV_X1 U8576 ( .A(n9076), .ZN(n8688) );
  INV_X1 U8577 ( .A(n9231), .ZN(n8493) );
  NAND2_X1 U8578 ( .A1(n9073), .A2(n9104), .ZN(n6745) );
  AOI22_X1 U8579 ( .A1(n8493), .A2(n6745), .B1(n8685), .B2(n9081), .ZN(n6746)
         );
  NAND2_X1 U8580 ( .A1(n9024), .A2(n9021), .ZN(n8700) );
  NAND2_X1 U8581 ( .A1(n6747), .A2(n9054), .ZN(n6748) );
  INV_X1 U8582 ( .A(n6747), .ZN(n8702) );
  AOI22_X1 U8583 ( .A1(n6610), .A2(n6748), .B1(n8702), .B2(n8401), .ZN(n6749)
         );
  INV_X1 U8584 ( .A(n8617), .ZN(n8704) );
  NAND2_X1 U8585 ( .A1(n8510), .A2(n9001), .ZN(n8588) );
  NAND2_X1 U8586 ( .A1(n9190), .A2(n8984), .ZN(n8988) );
  NOR2_X1 U8587 ( .A1(n8510), .A2(n9001), .ZN(n8718) );
  NOR2_X1 U8588 ( .A1(n8970), .A2(n8975), .ZN(n8727) );
  XNOR2_X1 U8589 ( .A(n6802), .B(n8610), .ZN(n9172) );
  OR2_X1 U8590 ( .A1(n8763), .A2(n6752), .ZN(n6753) );
  AND2_X1 U8591 ( .A1(n6753), .A2(n10172), .ZN(n6755) );
  INV_X1 U8592 ( .A(n8763), .ZN(n6754) );
  NAND2_X1 U8593 ( .A1(n9169), .A2(n9154), .ZN(n6756) );
  NAND2_X1 U8594 ( .A1(n6759), .A2(n6758), .ZN(P2_U3487) );
  INV_X1 U8595 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6769) );
  INV_X1 U8596 ( .A(n6760), .ZN(n6765) );
  NAND2_X1 U8597 ( .A1(n6884), .A2(n6762), .ZN(n6761) );
  OAI21_X1 U8598 ( .B1(n7013), .B2(n6762), .A(n6761), .ZN(n6763) );
  INV_X1 U8599 ( .A(n6763), .ZN(n6764) );
  AND2_X1 U8600 ( .A1(n7844), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6766) );
  INV_X1 U8601 ( .A(n6892), .ZN(n6997) );
  MUX2_X1 U8602 ( .A(n6769), .B(n9165), .S(n10141), .Z(n6775) );
  NAND2_X1 U8603 ( .A1(n7011), .A2(n8762), .ZN(n8947) );
  NAND2_X1 U8604 ( .A1(n10124), .A2(n8947), .ZN(n6770) );
  AOI22_X1 U8605 ( .A1(n9169), .A2(n9109), .B1(n9096), .B2(n8428), .ZN(n6772)
         );
  NAND2_X1 U8606 ( .A1(n6775), .A2(n6774), .ZN(P2_U3205) );
  INV_X1 U8607 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6784) );
  XNOR2_X1 U8608 ( .A(n6776), .B(n8731), .ZN(n8959) );
  INV_X1 U8609 ( .A(n8775), .ZN(n8742) );
  MUX2_X1 U8610 ( .A(n6784), .B(n6798), .S(n10189), .Z(n6786) );
  NAND2_X1 U8611 ( .A1(n8451), .A2(n9154), .ZN(n6785) );
  NAND2_X1 U8612 ( .A1(n6786), .A2(n6785), .ZN(P2_U3486) );
  NAND2_X1 U8613 ( .A1(n6787), .A2(n6792), .ZN(n6990) );
  INV_X1 U8614 ( .A(n6990), .ZN(n6788) );
  NAND2_X1 U8615 ( .A1(n6788), .A2(n6892), .ZN(n7005) );
  AND2_X1 U8616 ( .A1(n7810), .A2(n8613), .ZN(n7012) );
  INV_X1 U8617 ( .A(n7012), .ZN(n6790) );
  AND2_X1 U8618 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  AND2_X1 U8619 ( .A1(n6697), .A2(n10172), .ZN(n6795) );
  NAND2_X1 U8620 ( .A1(n6795), .A2(n6991), .ZN(n7001) );
  NAND2_X1 U8621 ( .A1(n7001), .A2(n10122), .ZN(n6989) );
  NAND2_X1 U8622 ( .A1(n7020), .A2(n6989), .ZN(n6796) );
  MUX2_X1 U8623 ( .A(n10371), .B(n6798), .S(n10178), .Z(n6801) );
  NAND2_X1 U8624 ( .A1(n8451), .A2(n6799), .ZN(n6800) );
  NAND2_X1 U8625 ( .A1(n6801), .A2(n6800), .ZN(P2_U3454) );
  INV_X1 U8626 ( .A(n9169), .ZN(n6806) );
  NAND2_X1 U8627 ( .A1(n8367), .A2(n6486), .ZN(n6804) );
  OR2_X1 U8628 ( .A1(n6430), .A2(n8368), .ZN(n6803) );
  INV_X1 U8629 ( .A(n8774), .ZN(n6805) );
  NAND2_X1 U8630 ( .A1(n8733), .A2(n6805), .ZN(n8578) );
  NAND2_X1 U8631 ( .A1(n8752), .A2(n8578), .ZN(n6807) );
  XNOR2_X1 U8632 ( .A(n6808), .B(n6807), .ZN(n6809) );
  NAND2_X1 U8633 ( .A1(n6809), .A2(n9094), .ZN(n6820) );
  INV_X1 U8634 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8635 ( .A1(n7927), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6812) );
  INV_X1 U8636 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6810) );
  OR2_X1 U8637 ( .A1(n7928), .A2(n6810), .ZN(n6811) );
  OAI211_X1 U8638 ( .C1(n4612), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  INV_X1 U8639 ( .A(n6814), .ZN(n6815) );
  AND2_X1 U8640 ( .A1(n7933), .A2(n6815), .ZN(n8581) );
  NAND2_X1 U8641 ( .A1(n6816), .A2(P2_B_REG_SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8642 ( .A1(n6698), .A2(n6817), .ZN(n8940) );
  OAI22_X1 U8643 ( .A1(n8742), .A2(n10125), .B1(n8581), .B2(n8940), .ZN(n6818)
         );
  INV_X1 U8644 ( .A(n6818), .ZN(n6819) );
  NOR2_X1 U8645 ( .A1(n8948), .A2(n10174), .ZN(n6821) );
  INV_X1 U8646 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6822) );
  OAI21_X1 U8647 ( .B1(n6826), .B2(n10180), .A(n6824), .ZN(P2_U3456) );
  OR2_X1 U8648 ( .A1(n10189), .A2(n10300), .ZN(n6825) );
  OAI21_X1 U8649 ( .B1(n6826), .B2(n10187), .A(n5139), .ZN(P2_U3488) );
  NAND2_X1 U8650 ( .A1(n10074), .A2(n9964), .ZN(n10017) );
  INV_X1 U8651 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6827) );
  OAI21_X1 U8652 ( .B1(n6830), .B2(n10072), .A(n6829), .ZN(P1_U3518) );
  INV_X1 U8653 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10493) );
  INV_X1 U8654 ( .A(n9651), .ZN(n6841) );
  INV_X1 U8655 ( .A(SI_29_), .ZN(n6831) );
  AND2_X1 U8656 ( .A1(n6832), .A2(n6831), .ZN(n6835) );
  INV_X1 U8657 ( .A(n6832), .ZN(n6833) );
  NAND2_X1 U8658 ( .A1(n6833), .A2(SI_29_), .ZN(n6834) );
  INV_X1 U8659 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8572) );
  INV_X1 U8660 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8377) );
  MUX2_X1 U8661 ( .A(n8572), .B(n8377), .S(n6873), .Z(n6838) );
  INV_X1 U8662 ( .A(SI_30_), .ZN(n6837) );
  NAND2_X1 U8663 ( .A1(n6838), .A2(n6837), .ZN(n6842) );
  INV_X1 U8664 ( .A(n6838), .ZN(n6839) );
  NAND2_X1 U8665 ( .A1(n6839), .A2(SI_30_), .ZN(n6840) );
  NAND2_X1 U8666 ( .A1(n6842), .A2(n6840), .ZN(n6843) );
  AOI21_X2 U8667 ( .B1(n8575), .B2(n6847), .A(n4558), .ZN(n9972) );
  NAND2_X1 U8668 ( .A1(n6841), .A2(n9972), .ZN(n9652) );
  INV_X1 U8669 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9247) );
  INV_X1 U8670 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6848) );
  MUX2_X1 U8671 ( .A(n9247), .B(n6848), .S(n6873), .Z(n6845) );
  XNOR2_X1 U8672 ( .A(n6845), .B(SI_31_), .ZN(n6846) );
  OR2_X1 U8673 ( .A1(n4469), .A2(n6848), .ZN(n6850) );
  NAND2_X1 U8674 ( .A1(n4458), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8675 ( .A1(n4457), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8676 ( .A1(n6852), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6853) );
  NAND3_X1 U8677 ( .A1(n6855), .A2(n6854), .A3(n6853), .ZN(n8290) );
  AOI21_X1 U8678 ( .B1(n9646), .B2(n9843), .A(n9895), .ZN(n6859) );
  MUX2_X1 U8679 ( .A(n10493), .B(n6859), .S(n10077), .Z(n6858) );
  NAND2_X1 U8680 ( .A1(n6858), .A2(n6857), .ZN(P1_U3553) );
  INV_X1 U8681 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6860) );
  MUX2_X1 U8682 ( .A(n6860), .B(n6859), .S(n10074), .Z(n6863) );
  NAND2_X1 U8683 ( .A1(n8212), .A2(n6861), .ZN(n6862) );
  NAND2_X1 U8684 ( .A1(n6863), .A2(n6862), .ZN(P1_U3521) );
  INV_X1 U8685 ( .A(n6864), .ZN(n6865) );
  XNOR2_X1 U8686 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8687 ( .A1(n6873), .A2(P2_U3151), .ZN(n9256) );
  INV_X2 U8688 ( .A(n9256), .ZN(n9246) );
  OR2_X2 U8689 ( .A1(n6873), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9258) );
  OAI222_X1 U8690 ( .A1(n9246), .A2(n4622), .B1(P2_U3151), .B2(n7171), .C1(
        n9258), .C2(n6881), .ZN(P2_U3294) );
  OAI222_X1 U8691 ( .A1(n9246), .A2(n6866), .B1(n9258), .B2(n6898), .C1(n7185), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U8692 ( .A1(n9246), .A2(n6867), .B1(n9258), .B2(n6879), .C1(n8798), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  OAI222_X1 U8693 ( .A1(n9246), .A2(n5188), .B1(n9258), .B2(n6877), .C1(n7071), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  OAI222_X1 U8694 ( .A1(n9246), .A2(n6869), .B1(n9258), .B2(n6874), .C1(n6868), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6872) );
  INV_X1 U8696 ( .A(n6870), .ZN(n6876) );
  OAI222_X1 U8697 ( .A1(n9246), .A2(n6872), .B1(n9258), .B2(n6876), .C1(n6871), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  OR2_X2 U8698 ( .A1(n6873), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8378) );
  AND2_X1 U8699 ( .A1(n6873), .A2(P1_U3086), .ZN(n7532) );
  INV_X2 U8700 ( .A(n7532), .ZN(n10029) );
  OAI222_X1 U8701 ( .A1(n8378), .A2(n6875), .B1(n10029), .B2(n6874), .C1(
        P1_U3086), .C2(n9561), .ZN(P1_U3350) );
  INV_X1 U8702 ( .A(n6948), .ZN(n9576) );
  OAI222_X1 U8703 ( .A1(n8378), .A2(n10264), .B1(n10029), .B2(n6876), .C1(
        P1_U3086), .C2(n9576), .ZN(P1_U3349) );
  OAI222_X1 U8704 ( .A1(n8378), .A2(n6878), .B1(n10029), .B2(n6877), .C1(
        P1_U3086), .C2(n9535), .ZN(P1_U3352) );
  INV_X1 U8705 ( .A(n9547), .ZN(n6929) );
  OAI222_X1 U8706 ( .A1(n8378), .A2(n6880), .B1(n10029), .B2(n6879), .C1(
        P1_U3086), .C2(n6929), .ZN(P1_U3351) );
  INV_X1 U8707 ( .A(n9502), .ZN(n6883) );
  OAI222_X1 U8708 ( .A1(P1_U3086), .A2(n6883), .B1(n8378), .B2(n6882), .C1(
        n10029), .C2(n6881), .ZN(P1_U3354) );
  INV_X1 U8709 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6887) );
  INV_X1 U8710 ( .A(n6884), .ZN(n6885) );
  NAND2_X1 U8711 ( .A1(n6885), .A2(n6892), .ZN(n6886) );
  OAI21_X1 U8712 ( .B1(n6892), .B2(n6887), .A(n6886), .ZN(P2_U3377) );
  INV_X1 U8713 ( .A(n6888), .ZN(n6890) );
  OAI222_X1 U8714 ( .A1(n8378), .A2(n6889), .B1(n10029), .B2(n6890), .C1(
        P1_U3086), .C2(n6940), .ZN(P1_U3347) );
  OAI222_X1 U8715 ( .A1(n9246), .A2(n6891), .B1(n9258), .B2(n6890), .C1(n7281), 
        .C2(P2_U3151), .ZN(P2_U3287) );
  INV_X1 U8716 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10441) );
  NOR2_X1 U8717 ( .A1(n6918), .A2(n10441), .ZN(P2_U3249) );
  INV_X1 U8718 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10379) );
  NOR2_X1 U8719 ( .A1(n6918), .A2(n10379), .ZN(P2_U3247) );
  INV_X1 U8720 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10454) );
  NOR2_X1 U8721 ( .A1(n6918), .A2(n10454), .ZN(P2_U3253) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6894) );
  INV_X1 U8723 ( .A(n6893), .ZN(n6901) );
  INV_X1 U8724 ( .A(n9598), .ZN(n9591) );
  OAI222_X1 U8725 ( .A1(n8378), .A2(n6894), .B1(n10029), .B2(n6901), .C1(
        P1_U3086), .C2(n9591), .ZN(P1_U3348) );
  INV_X1 U8726 ( .A(n6895), .ZN(n6908) );
  OAI222_X1 U8727 ( .A1(n9258), .A2(n6908), .B1(P2_U3151), .B2(n4768), .C1(
        n6896), .C2(n9246), .ZN(P2_U3286) );
  INV_X1 U8728 ( .A(n9520), .ZN(n6899) );
  OAI222_X1 U8729 ( .A1(n6899), .A2(P1_U3086), .B1(n10029), .B2(n6898), .C1(
        n6897), .C2(n8378), .ZN(P1_U3353) );
  INV_X1 U8730 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6902) );
  OAI222_X1 U8731 ( .A1(n9246), .A2(n6902), .B1(n9258), .B2(n6901), .C1(n6900), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  INV_X1 U8732 ( .A(n7852), .ZN(n6903) );
  OR2_X1 U8733 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  NAND2_X1 U8734 ( .A1(n6905), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8735 ( .A1(n8292), .A2(n7852), .ZN(n6906) );
  NAND2_X1 U8736 ( .A1(n5316), .A2(n6906), .ZN(n6935) );
  INV_X1 U8737 ( .A(n6935), .ZN(n6907) );
  NOR2_X1 U8738 ( .A1(n10038), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8739 ( .A(n7029), .ZN(n7025) );
  OAI222_X1 U8740 ( .A1(P1_U3086), .A2(n7025), .B1(n10029), .B2(n6908), .C1(
        n10265), .C2(n8378), .ZN(P1_U3346) );
  INV_X1 U8741 ( .A(n6909), .ZN(n6911) );
  OAI222_X1 U8742 ( .A1(n9258), .A2(n6911), .B1(P2_U3151), .B2(n7591), .C1(
        n6910), .C2(n9246), .ZN(P2_U3285) );
  INV_X1 U8743 ( .A(n7032), .ZN(n7052) );
  OAI222_X1 U8744 ( .A1(P1_U3086), .A2(n7052), .B1(n10029), .B2(n6911), .C1(
        n10266), .C2(n8378), .ZN(P1_U3345) );
  NAND2_X1 U8745 ( .A1(n7323), .A2(P1_U3973), .ZN(n6912) );
  OAI21_X1 U8746 ( .B1(P1_U3973), .B2(n6409), .A(n6912), .ZN(P1_U3554) );
  AND2_X1 U8747 ( .A1(n6913), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8748 ( .A1(n6913), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8749 ( .A1(n6913), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8750 ( .A1(n6913), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8751 ( .A1(n6913), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8752 ( .A1(n6913), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8753 ( .A1(n6913), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8754 ( .A1(n6913), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8755 ( .A1(n6913), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8756 ( .A1(n6913), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8757 ( .A1(n6913), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  INV_X1 U8758 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6917) );
  INV_X1 U8759 ( .A(n10223), .ZN(n10064) );
  OAI21_X1 U8760 ( .B1(n10064), .B2(P1_D_REG_1__SCAN_IN), .A(n6915), .ZN(n6916) );
  OAI21_X1 U8761 ( .B1(n10020), .B2(n6917), .A(n6916), .ZN(P1_U3440) );
  INV_X1 U8762 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6922) );
  NOR3_X1 U8763 ( .A1(n6920), .A2(n6919), .A3(P2_U3151), .ZN(n6921) );
  AOI21_X1 U8764 ( .B1(n6913), .B2(n6922), .A(n6921), .ZN(P2_U3376) );
  AND2_X1 U8765 ( .A1(n6913), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8766 ( .A1(n6913), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8767 ( .A1(n6913), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8768 ( .A1(n6913), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8769 ( .A1(n6913), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8770 ( .A1(n6913), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8771 ( .A1(n6913), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8772 ( .A1(n6913), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8773 ( .A1(n6913), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8774 ( .A1(n6913), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8775 ( .A1(n6913), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8776 ( .A1(n6913), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8777 ( .A1(n6913), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8778 ( .A1(n6913), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8779 ( .A1(n6913), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8780 ( .A1(n6913), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  INV_X1 U8781 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9521) );
  MUX2_X1 U8782 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9521), .S(n9520), .Z(n6926)
         );
  INV_X1 U8783 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9499) );
  MUX2_X1 U8784 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9499), .S(n9502), .Z(n6924)
         );
  AND2_X1 U8785 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6923) );
  NAND2_X1 U8786 ( .A1(n9502), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U8787 ( .A1(n9523), .A2(n9522), .ZN(n6925) );
  NAND2_X1 U8788 ( .A1(n6926), .A2(n6925), .ZN(n9526) );
  NAND2_X1 U8789 ( .A1(n9520), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8790 ( .A1(n9526), .A2(n6927), .ZN(n9533) );
  INV_X1 U8791 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6928) );
  MUX2_X1 U8792 ( .A(n6928), .B(P1_REG1_REG_3__SCAN_IN), .S(n9535), .Z(n9534)
         );
  OR2_X1 U8793 ( .A1(n9535), .A2(n6928), .ZN(n9553) );
  INV_X1 U8794 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10075) );
  MUX2_X1 U8795 ( .A(n10075), .B(P1_REG1_REG_4__SCAN_IN), .S(n9547), .Z(n9552)
         );
  AOI21_X1 U8796 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9551) );
  NOR2_X1 U8797 ( .A1(n6929), .A2(n10075), .ZN(n9560) );
  INV_X1 U8798 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6930) );
  MUX2_X1 U8799 ( .A(n6930), .B(P1_REG1_REG_5__SCAN_IN), .S(n9561), .Z(n6931)
         );
  INV_X1 U8800 ( .A(n9561), .ZN(n9569) );
  NAND2_X1 U8801 ( .A1(n9569), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9583) );
  INV_X1 U8802 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6932) );
  MUX2_X1 U8803 ( .A(n6932), .B(P1_REG1_REG_6__SCAN_IN), .S(n6948), .Z(n9582)
         );
  AOI21_X1 U8804 ( .B1(n9584), .B2(n9583), .A(n9582), .ZN(n9604) );
  NOR2_X1 U8805 ( .A1(n9576), .A2(n6932), .ZN(n9599) );
  INV_X1 U8806 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6933) );
  MUX2_X1 U8807 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6933), .S(n9598), .Z(n6934)
         );
  OAI21_X1 U8808 ( .B1(n6933), .B2(n9591), .A(n9602), .ZN(n6977) );
  XNOR2_X1 U8809 ( .A(n6940), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6976) );
  XNOR2_X1 U8810 ( .A(n6977), .B(n6976), .ZN(n6958) );
  INV_X1 U8811 ( .A(n10041), .ZN(n6937) );
  NAND2_X1 U8812 ( .A1(n6937), .A2(n10031), .ZN(n9633) );
  INV_X1 U8813 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U8814 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9316) );
  OAI21_X1 U8815 ( .B1(n9643), .B2(n6938), .A(n9316), .ZN(n6939) );
  AOI21_X1 U8816 ( .B1(n9636), .B2(n6975), .A(n6939), .ZN(n6957) );
  INV_X1 U8817 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10357) );
  MUX2_X1 U8818 ( .A(n10357), .B(P1_REG2_REG_8__SCAN_IN), .S(n6940), .Z(n6955)
         );
  INV_X1 U8819 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7463) );
  MUX2_X1 U8820 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7463), .S(n9520), .Z(n9529)
         );
  INV_X1 U8821 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6941) );
  MUX2_X1 U8822 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6941), .S(n9502), .Z(n9505)
         );
  NAND2_X1 U8823 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9512) );
  INV_X1 U8824 ( .A(n9512), .ZN(n9504) );
  NAND2_X1 U8825 ( .A1(n9505), .A2(n9504), .ZN(n9503) );
  NAND2_X1 U8826 ( .A1(n9502), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8827 ( .A1(n9503), .A2(n6942), .ZN(n9528) );
  NAND2_X1 U8828 ( .A1(n9529), .A2(n9528), .ZN(n9527) );
  NAND2_X1 U8829 ( .A1(n9520), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8830 ( .A1(n9527), .A2(n6943), .ZN(n9539) );
  XNOR2_X1 U8831 ( .A(n9535), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U8832 ( .A1(n9539), .A2(n9540), .ZN(n9538) );
  INV_X1 U8833 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6944) );
  OR2_X1 U8834 ( .A1(n9535), .A2(n6944), .ZN(n6945) );
  NAND2_X1 U8835 ( .A1(n9538), .A2(n6945), .ZN(n9549) );
  INV_X1 U8836 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10293) );
  MUX2_X1 U8837 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10293), .S(n9547), .Z(n9550)
         );
  NAND2_X1 U8838 ( .A1(n9549), .A2(n9550), .ZN(n9548) );
  NAND2_X1 U8839 ( .A1(n9547), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8840 ( .A1(n9548), .A2(n6946), .ZN(n9571) );
  INV_X1 U8841 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10471) );
  MUX2_X1 U8842 ( .A(n10471), .B(P1_REG2_REG_5__SCAN_IN), .S(n9561), .Z(n9572)
         );
  NAND2_X1 U8843 ( .A1(n9571), .A2(n9572), .ZN(n9570) );
  NAND2_X1 U8844 ( .A1(n9569), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8845 ( .A1(n9570), .A2(n6947), .ZN(n9580) );
  INV_X1 U8846 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U8847 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10317), .S(n6948), .Z(n9581)
         );
  NAND2_X1 U8848 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  NAND2_X1 U8849 ( .A1(n6948), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8850 ( .A1(n9579), .A2(n6949), .ZN(n9596) );
  INV_X1 U8851 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6950) );
  MUX2_X1 U8852 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6950), .S(n9598), .Z(n9597)
         );
  NAND2_X1 U8853 ( .A1(n9596), .A2(n9597), .ZN(n9595) );
  NAND2_X1 U8854 ( .A1(n9598), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8855 ( .A1(n9595), .A2(n6951), .ZN(n6954) );
  NAND2_X1 U8856 ( .A1(n6954), .A2(n6955), .ZN(n6971) );
  INV_X1 U8857 ( .A(n10031), .ZN(n6952) );
  NAND2_X1 U8858 ( .A1(n9514), .A2(n6952), .ZN(n6953) );
  NOR2_X2 U8859 ( .A1(n10041), .A2(n6953), .ZN(n9638) );
  OAI211_X1 U8860 ( .C1(n6955), .C2(n6954), .A(n6971), .B(n9638), .ZN(n6956)
         );
  OAI211_X1 U8861 ( .C1(n6958), .C2(n9633), .A(n6957), .B(n6956), .ZN(P1_U3251) );
  INV_X1 U8862 ( .A(n6959), .ZN(n6962) );
  OAI222_X1 U8863 ( .A1(n9246), .A2(n6960), .B1(n9258), .B2(n6962), .C1(n4771), 
        .C2(P2_U3151), .ZN(P2_U3284) );
  INV_X1 U8864 ( .A(n7128), .ZN(n6961) );
  OAI222_X1 U8865 ( .A1(n8378), .A2(n10457), .B1(n10029), .B2(n6962), .C1(
        P1_U3086), .C2(n6961), .ZN(P1_U3344) );
  NAND2_X1 U8866 ( .A1(n8290), .A2(P1_U3973), .ZN(n6963) );
  OAI21_X1 U8867 ( .B1(P1_U3973), .B2(n9247), .A(n6963), .ZN(P1_U3585) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U8869 ( .A1(P2_U3893), .A2(n7404), .ZN(n6964) );
  OAI21_X1 U8870 ( .B1(P2_U3893), .B2(n6965), .A(n6964), .ZN(P2_U3491) );
  INV_X1 U8871 ( .A(n6966), .ZN(n6969) );
  OAI222_X1 U8872 ( .A1(n9258), .A2(n6969), .B1(P2_U3151), .B2(n8828), .C1(
        n6967), .C2(n9246), .ZN(P2_U3283) );
  OAI222_X1 U8873 ( .A1(P1_U3086), .A2(n7222), .B1(n10029), .B2(n6969), .C1(
        n6968), .C2(n8378), .ZN(P1_U3343) );
  XNOR2_X1 U8874 ( .A(n7029), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8875 ( .A1(n6975), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8876 ( .A1(n6971), .A2(n6970), .ZN(n6973) );
  INV_X1 U8877 ( .A(n7031), .ZN(n6972) );
  AOI21_X1 U8878 ( .B1(n6974), .B2(n6973), .A(n6972), .ZN(n6984) );
  INV_X1 U8879 ( .A(n9638), .ZN(n7900) );
  XOR2_X1 U8880 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7029), .Z(n6979) );
  NAND2_X1 U8881 ( .A1(n6978), .A2(n6979), .ZN(n7045) );
  OAI21_X1 U8882 ( .B1(n6979), .B2(n6978), .A(n7045), .ZN(n6982) );
  NAND2_X1 U8883 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U8884 ( .A1(n10038), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6980) );
  OAI211_X1 U8885 ( .C1(n9592), .C2(n7025), .A(n7952), .B(n6980), .ZN(n6981)
         );
  AOI21_X1 U8886 ( .B1(n6982), .B2(n9632), .A(n6981), .ZN(n6983) );
  OAI21_X1 U8887 ( .B1(n6984), .B2(n7900), .A(n6983), .ZN(P1_U3252) );
  INV_X1 U8888 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6986) );
  INV_X1 U8889 ( .A(n6985), .ZN(n6987) );
  INV_X1 U8890 ( .A(n7341), .ZN(n7337) );
  OAI222_X1 U8891 ( .A1(n8378), .A2(n6986), .B1(n10029), .B2(n6987), .C1(
        P1_U3086), .C2(n7337), .ZN(P1_U3342) );
  INV_X1 U8892 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6988) );
  OAI222_X1 U8893 ( .A1(n9246), .A2(n6988), .B1(n9258), .B2(n6987), .C1(n8848), 
        .C2(P2_U3151), .ZN(P2_U3282) );
  NAND2_X1 U8894 ( .A1(n6990), .A2(n6989), .ZN(n6995) );
  INV_X1 U8895 ( .A(n6991), .ZN(n7002) );
  INV_X1 U8896 ( .A(n6992), .ZN(n6998) );
  AOI21_X1 U8897 ( .B1(n7002), .B2(n6998), .A(n6993), .ZN(n6994) );
  NAND2_X1 U8898 ( .A1(n6995), .A2(n6994), .ZN(n6996) );
  NAND2_X1 U8899 ( .A1(n6996), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7000) );
  NOR2_X1 U8900 ( .A1(n6997), .A2(n7307), .ZN(n8768) );
  NAND2_X1 U8901 ( .A1(n8768), .A2(n6998), .ZN(n6999) );
  NAND2_X1 U8902 ( .A1(n8063), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7081) );
  INV_X1 U8903 ( .A(n7081), .ZN(n7010) );
  AND2_X1 U8904 ( .A1(n7404), .A2(n7312), .ZN(n8624) );
  INV_X1 U8905 ( .A(n8624), .ZN(n8622) );
  NAND2_X1 U8906 ( .A1(n10117), .A2(n8622), .ZN(n8592) );
  OR2_X1 U8907 ( .A1(n7005), .A2(n7001), .ZN(n7004) );
  NAND2_X1 U8908 ( .A1(n7020), .A2(n7002), .ZN(n7003) );
  OR2_X1 U8909 ( .A1(n7005), .A2(n10172), .ZN(n7006) );
  NOR2_X1 U8910 ( .A1(n7307), .A2(n7017), .ZN(n7007) );
  OAI22_X1 U8911 ( .A1(n8568), .A2(n7312), .B1(n10126), .B2(n8541), .ZN(n7008)
         );
  AOI21_X1 U8912 ( .B1(n8592), .B2(n8557), .A(n7008), .ZN(n7009) );
  OAI21_X1 U8913 ( .B1(n7010), .B2(n7311), .A(n7009), .ZN(P2_U3172) );
  AOI21_X1 U8914 ( .B1(n7011), .B2(n8365), .A(n8763), .ZN(n7015) );
  NAND2_X1 U8915 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  NAND2_X2 U8916 ( .A1(n7015), .A2(n7014), .ZN(n7111) );
  XOR2_X1 U8917 ( .A(n7090), .B(n10126), .Z(n7076) );
  XOR2_X1 U8918 ( .A(n7092), .B(n7076), .Z(n7024) );
  INV_X1 U8919 ( .A(n7017), .ZN(n7018) );
  NOR2_X1 U8920 ( .A1(n7307), .A2(n7018), .ZN(n7019) );
  NAND2_X1 U8921 ( .A1(n7020), .A2(n7019), .ZN(n8563) );
  AOI22_X1 U8922 ( .A1(n8539), .A2(n7404), .B1(n8561), .B2(n8792), .ZN(n7021)
         );
  OAI21_X1 U8923 ( .B1(n8568), .B2(n7016), .A(n7021), .ZN(n7022) );
  AOI21_X1 U8924 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7081), .A(n7022), .ZN(
        n7023) );
  OAI21_X1 U8925 ( .B1(n7024), .B2(n8555), .A(n7023), .ZN(P2_U3162) );
  INV_X1 U8926 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7026) );
  XOR2_X1 U8927 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7032), .Z(n7047) );
  INV_X1 U8928 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U8929 ( .A1(n7025), .A2(n10315), .ZN(n7044) );
  NAND3_X1 U8930 ( .A1(n7045), .A2(n7047), .A3(n7044), .ZN(n7046) );
  OAI21_X1 U8931 ( .B1(n7026), .B2(n7052), .A(n7046), .ZN(n7130) );
  INV_X1 U8932 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8035) );
  XNOR2_X1 U8933 ( .A(n7128), .B(n8035), .ZN(n7129) );
  XNOR2_X1 U8934 ( .A(n7130), .B(n7129), .ZN(n7039) );
  INV_X1 U8935 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8936 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8043) );
  OAI21_X1 U8937 ( .B1(n9643), .B2(n7027), .A(n8043), .ZN(n7028) );
  AOI21_X1 U8938 ( .B1(n9636), .B2(n7128), .A(n7028), .ZN(n7038) );
  OR2_X1 U8939 ( .A1(n7029), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8940 ( .A1(n7031), .A2(n7030), .ZN(n7042) );
  INV_X1 U8941 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7704) );
  MUX2_X1 U8942 ( .A(n7704), .B(P1_REG2_REG_10__SCAN_IN), .S(n7032), .Z(n7043)
         );
  NAND2_X1 U8943 ( .A1(n7032), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8944 ( .A1(n7040), .A2(n7033), .ZN(n7036) );
  INV_X1 U8945 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7034) );
  XNOR2_X1 U8946 ( .A(n7128), .B(n7034), .ZN(n7035) );
  NAND2_X1 U8947 ( .A1(n7036), .A2(n7035), .ZN(n7124) );
  OAI211_X1 U8948 ( .C1(n7036), .C2(n7035), .A(n7124), .B(n9638), .ZN(n7037)
         );
  OAI211_X1 U8949 ( .C1(n7039), .C2(n9633), .A(n7038), .B(n7037), .ZN(P1_U3254) );
  INV_X1 U8950 ( .A(n7040), .ZN(n7041) );
  AOI211_X1 U8951 ( .C1(n7043), .C2(n7042), .A(n7900), .B(n7041), .ZN(n7054)
         );
  AND2_X1 U8952 ( .A1(n7045), .A2(n7044), .ZN(n7048) );
  OAI211_X1 U8953 ( .C1(n7048), .C2(n7047), .A(n9632), .B(n7046), .ZN(n7051)
         );
  AND2_X1 U8954 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7049) );
  AOI21_X1 U8955 ( .B1(n10038), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7049), .ZN(
        n7050) );
  OAI211_X1 U8956 ( .C1(n9592), .C2(n7052), .A(n7051), .B(n7050), .ZN(n7053)
         );
  OR2_X1 U8957 ( .A1(n7054), .A2(n7053), .ZN(P1_U3253) );
  NAND2_X1 U8958 ( .A1(n7323), .A2(n7321), .ZN(n8301) );
  INV_X1 U8959 ( .A(n8301), .ZN(n7055) );
  NOR2_X1 U8960 ( .A1(n7326), .A2(n7055), .ZN(n8231) );
  INV_X1 U8961 ( .A(n8231), .ZN(n7056) );
  OAI21_X1 U8962 ( .B1(n9878), .B2(n10071), .A(n7056), .ZN(n7058) );
  NOR2_X1 U8963 ( .A1(n6124), .A2(n9455), .ZN(n7446) );
  INV_X1 U8964 ( .A(n7446), .ZN(n7057) );
  OAI211_X1 U8965 ( .C1(n7321), .C2(n7059), .A(n7058), .B(n7057), .ZN(n7061)
         );
  NAND2_X1 U8966 ( .A1(n7061), .A2(n10077), .ZN(n7060) );
  OAI21_X1 U8967 ( .B1(n10077), .B2(n6127), .A(n7060), .ZN(P1_U3522) );
  INV_X1 U8968 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U8969 ( .A1(n7061), .A2(n10074), .ZN(n7062) );
  OAI21_X1 U8970 ( .B1(n10074), .B2(n10402), .A(n7062), .ZN(P1_U3453) );
  INV_X1 U8971 ( .A(n7063), .ZN(n7064) );
  AOI21_X1 U8972 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7075) );
  OAI21_X1 U8973 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7067), .A(n8801), .ZN(
        n7070) );
  XNOR2_X1 U8974 ( .A(n7068), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7069) );
  AOI22_X1 U8975 ( .A1(n7070), .A2(n8922), .B1(n10092), .B2(n7069), .ZN(n7074)
         );
  OAI22_X1 U8976 ( .A1(n8928), .A2(n7071), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10225), .ZN(n7072) );
  AOI21_X1 U8977 ( .B1(n10099), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7072), .ZN(
        n7073) );
  OAI211_X1 U8978 ( .C1(n7075), .C2(n10095), .A(n7074), .B(n7073), .ZN(
        P2_U3185) );
  AOI22_X1 U8979 ( .A1(n7076), .A2(n7092), .B1(n10126), .B2(n7090), .ZN(n7078)
         );
  XNOR2_X1 U8980 ( .A(n8792), .B(n7086), .ZN(n7077) );
  XNOR2_X1 U8981 ( .A(n7078), .B(n7077), .ZN(n7083) );
  INV_X1 U8982 ( .A(n8791), .ZN(n10128) );
  OAI22_X1 U8983 ( .A1(n8541), .A2(n10128), .B1(n10126), .B2(n8563), .ZN(n7080) );
  NOR2_X1 U8984 ( .A1(n8568), .A2(n4567), .ZN(n7079) );
  AOI211_X1 U8985 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7081), .A(n7080), .B(
        n7079), .ZN(n7082) );
  OAI21_X1 U8986 ( .B1(n7083), .B2(n8555), .A(n7082), .ZN(P2_U3177) );
  XOR2_X1 U8987 ( .A(n8791), .B(n7108), .Z(n7097) );
  NAND2_X1 U8988 ( .A1(n7088), .A2(n8792), .ZN(n7087) );
  NAND2_X1 U8989 ( .A1(n7087), .A2(n7086), .ZN(n7095) );
  INV_X1 U8990 ( .A(n7088), .ZN(n7089) );
  NAND2_X1 U8991 ( .A1(n7089), .A2(n7406), .ZN(n7094) );
  NAND2_X1 U8992 ( .A1(n4507), .A2(n8792), .ZN(n7091) );
  OAI211_X1 U8993 ( .C1(n7092), .C2(n10126), .A(n7091), .B(n7090), .ZN(n7093)
         );
  NAND3_X1 U8994 ( .A1(n7095), .A2(n7094), .A3(n7093), .ZN(n7096) );
  AOI211_X1 U8995 ( .C1(n7097), .C2(n7096), .A(n8555), .B(n7110), .ZN(n7101)
         );
  MUX2_X1 U8996 ( .A(P2_STATE_REG_SCAN_IN), .B(n8063), .S(n10225), .Z(n7099)
         );
  AOI22_X1 U8997 ( .A1(n8539), .A2(n8792), .B1(n8561), .B2(n8790), .ZN(n7098)
         );
  OAI211_X1 U8998 ( .C1(n10157), .C2(n8568), .A(n7099), .B(n7098), .ZN(n7100)
         );
  OR2_X1 U8999 ( .A1(n7101), .A2(n7100), .ZN(P2_U3158) );
  INV_X1 U9000 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7104) );
  OAI21_X1 U9001 ( .B1(n9094), .B2(n10162), .A(n8592), .ZN(n7102) );
  OR2_X1 U9002 ( .A1(n10126), .A2(n10127), .ZN(n7308) );
  OAI211_X1 U9003 ( .C1(n10172), .C2(n7312), .A(n7102), .B(n7308), .ZN(n9158)
         );
  NAND2_X1 U9004 ( .A1(n10178), .A2(n9158), .ZN(n7103) );
  OAI21_X1 U9005 ( .B1(n10178), .B2(n7104), .A(n7103), .ZN(P2_U3390) );
  INV_X1 U9006 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10410) );
  INV_X1 U9007 ( .A(n7105), .ZN(n7107) );
  INV_X1 U9008 ( .A(n7484), .ZN(n7339) );
  OAI222_X1 U9009 ( .A1(n8378), .A2(n10410), .B1(n10029), .B2(n7107), .C1(
        P1_U3086), .C2(n7339), .ZN(P1_U3341) );
  INV_X1 U9010 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10486) );
  OAI222_X1 U9011 ( .A1(n9246), .A2(n10486), .B1(n9258), .B2(n7107), .C1(n4785), .C2(P2_U3151), .ZN(P2_U3281) );
  INV_X1 U9012 ( .A(n7108), .ZN(n7109) );
  XNOR2_X1 U9013 ( .A(n7363), .B(n4460), .ZN(n7145) );
  XNOR2_X1 U9014 ( .A(n7145), .B(n8790), .ZN(n7112) );
  OAI21_X1 U9015 ( .B1(n7113), .B2(n7112), .A(n7148), .ZN(n7114) );
  NAND2_X1 U9016 ( .A1(n7114), .A2(n8557), .ZN(n7118) );
  NAND2_X1 U9017 ( .A1(n8561), .A2(n8789), .ZN(n7115) );
  NAND2_X1 U9018 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U9019 ( .C1(n10128), .C2(n8563), .A(n7115), .B(n8797), .ZN(n7116)
         );
  AOI21_X1 U9020 ( .B1(n7363), .B2(n8553), .A(n7116), .ZN(n7117) );
  OAI211_X1 U9021 ( .C1(n7629), .C2(n8063), .A(n7118), .B(n7117), .ZN(P2_U3170) );
  INV_X1 U9022 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7120) );
  INV_X1 U9023 ( .A(n7119), .ZN(n7121) );
  OAI222_X1 U9024 ( .A1(n9246), .A2(n7120), .B1(n9258), .B2(n7121), .C1(n8876), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U9025 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7122) );
  INV_X1 U9026 ( .A(n7672), .ZN(n7664) );
  OAI222_X1 U9027 ( .A1(n8378), .A2(n7122), .B1(n10029), .B2(n7121), .C1(
        P1_U3086), .C2(n7664), .ZN(P1_U3340) );
  INV_X1 U9028 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7978) );
  XNOR2_X1 U9029 ( .A(n7222), .B(n7978), .ZN(n7127) );
  NAND2_X1 U9030 ( .A1(n7128), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7123) );
  NAND2_X1 U9031 ( .A1(n7124), .A2(n7123), .ZN(n7126) );
  INV_X1 U9032 ( .A(n7224), .ZN(n7125) );
  AOI21_X1 U9033 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n7138) );
  XNOR2_X1 U9034 ( .A(n7222), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U9035 ( .A1(n7131), .A2(n7132), .ZN(n7219) );
  OAI21_X1 U9036 ( .B1(n7132), .B2(n7131), .A(n7219), .ZN(n7136) );
  NOR2_X1 U9037 ( .A1(n7133), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9348) );
  AOI21_X1 U9038 ( .B1(n10038), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9348), .ZN(
        n7134) );
  OAI21_X1 U9039 ( .B1(n9592), .B2(n7222), .A(n7134), .ZN(n7135) );
  AOI21_X1 U9040 ( .B1(n7136), .B2(n9632), .A(n7135), .ZN(n7137) );
  OAI21_X1 U9041 ( .B1(n7138), .B2(n7900), .A(n7137), .ZN(P1_U3255) );
  INV_X1 U9042 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7144) );
  INV_X1 U9043 ( .A(n8928), .ZN(n10085) );
  AOI22_X1 U9044 ( .A1(n10085), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n7143) );
  OAI21_X1 U9045 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7139), .A(n7181), .ZN(n7140) );
  OAI21_X1 U9046 ( .B1(n8883), .B2(n7141), .A(n7140), .ZN(n7142) );
  OAI211_X1 U9047 ( .C1(n7144), .C2(n7207), .A(n7143), .B(n7142), .ZN(P2_U3182) );
  XNOR2_X1 U9048 ( .A(n6739), .B(n8107), .ZN(n7264) );
  XNOR2_X1 U9049 ( .A(n7264), .B(n8789), .ZN(n7267) );
  INV_X1 U9050 ( .A(n7149), .ZN(n7415) );
  INV_X1 U9051 ( .A(n8788), .ZN(n7152) );
  NAND2_X1 U9052 ( .A1(n8553), .A2(n6739), .ZN(n7151) );
  AND2_X1 U9053 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7204) );
  AOI21_X1 U9054 ( .B1(n8539), .B2(n8790), .A(n7204), .ZN(n7150) );
  OAI211_X1 U9055 ( .C1(n7152), .C2(n8541), .A(n7151), .B(n7150), .ZN(n7153)
         );
  AOI21_X1 U9056 ( .B1(n7415), .B2(n8565), .A(n7153), .ZN(n7154) );
  OAI21_X1 U9057 ( .B1(n7155), .B2(n8555), .A(n7154), .ZN(P2_U3167) );
  XOR2_X1 U9058 ( .A(n7156), .B(P2_REG1_REG_7__SCAN_IN), .Z(n7169) );
  OAI21_X1 U9059 ( .B1(n7159), .B2(n7158), .A(n7157), .ZN(n7167) );
  INV_X1 U9060 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7165) );
  NOR2_X1 U9061 ( .A1(n7160), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7161) );
  OAI21_X1 U9062 ( .B1(n7161), .B2(n7284), .A(n8922), .ZN(n7164) );
  AND2_X1 U9063 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7396) );
  AOI21_X1 U9064 ( .B1(n10085), .B2(n7162), .A(n7396), .ZN(n7163) );
  OAI211_X1 U9065 ( .C1(n7207), .C2(n7165), .A(n7164), .B(n7163), .ZN(n7166)
         );
  AOI21_X1 U9066 ( .B1(n8883), .B2(n7167), .A(n7166), .ZN(n7168) );
  OAI21_X1 U9067 ( .B1(n7169), .B2(n8939), .A(n7168), .ZN(P2_U3189) );
  OAI22_X1 U9068 ( .A1(n8928), .A2(n7171), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7170), .ZN(n7178) );
  XOR2_X1 U9069 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n7172), .Z(n7176) );
  AOI21_X1 U9070 ( .B1(n10472), .B2(n7174), .A(n7173), .ZN(n7175) );
  OAI22_X1 U9071 ( .A1(n8939), .A2(n7176), .B1(n7175), .B2(n10088), .ZN(n7177)
         );
  AOI211_X1 U9072 ( .C1(n10099), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7178), .B(
        n7177), .ZN(n7183) );
  OAI211_X1 U9073 ( .C1(n7181), .C2(n7180), .A(n8883), .B(n7179), .ZN(n7182)
         );
  NAND2_X1 U9074 ( .A1(n7183), .A2(n7182), .ZN(P2_U3183) );
  INV_X1 U9075 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7184) );
  OAI22_X1 U9076 ( .A1(n8928), .A2(n7185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7184), .ZN(n7196) );
  AOI21_X1 U9077 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7194) );
  OAI21_X1 U9078 ( .B1(n7191), .B2(n7190), .A(n7189), .ZN(n7192) );
  NAND2_X1 U9079 ( .A1(n10092), .A2(n7192), .ZN(n7193) );
  OAI21_X1 U9080 ( .B1(n7194), .B2(n10088), .A(n7193), .ZN(n7195) );
  AOI211_X1 U9081 ( .C1(n10099), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7196), .B(
        n7195), .ZN(n7201) );
  OAI211_X1 U9082 ( .C1(n7199), .C2(n7198), .A(n8883), .B(n7197), .ZN(n7200)
         );
  NAND2_X1 U9083 ( .A1(n7201), .A2(n7200), .ZN(P2_U3184) );
  XOR2_X1 U9084 ( .A(n7202), .B(P2_REG1_REG_5__SCAN_IN), .Z(n7216) );
  XNOR2_X1 U9085 ( .A(n7203), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7210) );
  INV_X1 U9086 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7208) );
  AOI21_X1 U9087 ( .B1(n10085), .B2(n7205), .A(n7204), .ZN(n7206) );
  OAI21_X1 U9088 ( .B1(n7208), .B2(n7207), .A(n7206), .ZN(n7209) );
  AOI21_X1 U9089 ( .B1(n7210), .B2(n8922), .A(n7209), .ZN(n7215) );
  OAI211_X1 U9090 ( .C1(n7213), .C2(n7212), .A(n7211), .B(n8883), .ZN(n7214)
         );
  OAI211_X1 U9091 ( .C1(n7216), .C2(n8939), .A(n7215), .B(n7214), .ZN(P2_U3187) );
  XOR2_X1 U9092 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7341), .Z(n7217) );
  INV_X1 U9093 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U9094 ( .A1(n7222), .A2(n10256), .ZN(n7218) );
  NAND3_X1 U9095 ( .A1(n7219), .A2(n7217), .A3(n7218), .ZN(n7336) );
  NAND2_X1 U9096 ( .A1(n7336), .A2(n9632), .ZN(n7232) );
  AOI21_X1 U9097 ( .B1(n7219), .B2(n7218), .A(n7217), .ZN(n7231) );
  INV_X1 U9098 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U9099 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9406) );
  OAI21_X1 U9100 ( .B1(n9643), .B2(n7220), .A(n9406), .ZN(n7221) );
  AOI21_X1 U9101 ( .B1(n9636), .B2(n7341), .A(n7221), .ZN(n7230) );
  NAND2_X1 U9102 ( .A1(n7222), .A2(n7978), .ZN(n7223) );
  NAND2_X1 U9103 ( .A1(n7224), .A2(n7223), .ZN(n7227) );
  INV_X1 U9104 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7225) );
  MUX2_X1 U9105 ( .A(n7225), .B(P1_REG2_REG_13__SCAN_IN), .S(n7341), .Z(n7226)
         );
  AOI21_X1 U9106 ( .B1(n7227), .B2(n7226), .A(n7900), .ZN(n7228) );
  NAND2_X1 U9107 ( .A1(n7228), .A2(n7343), .ZN(n7229) );
  OAI211_X1 U9108 ( .C1(n7232), .C2(n7231), .A(n7230), .B(n7229), .ZN(P1_U3256) );
  OAI21_X1 U9109 ( .B1(n7234), .B2(n5087), .A(n7233), .ZN(n7633) );
  INV_X1 U9110 ( .A(n8789), .ZN(n10108) );
  XNOR2_X1 U9111 ( .A(n7235), .B(n5087), .ZN(n7236) );
  OAI222_X1 U9112 ( .A1(n10127), .A2(n10108), .B1(n10125), .B2(n10128), .C1(
        n7236), .C2(n10132), .ZN(n7630) );
  AOI21_X1 U9113 ( .B1(n10162), .B2(n7633), .A(n7630), .ZN(n7365) );
  OAI22_X1 U9114 ( .A1(n9211), .A2(n8638), .B1(n6438), .B2(n10178), .ZN(n7237)
         );
  INV_X1 U9115 ( .A(n7237), .ZN(n7238) );
  OAI21_X1 U9116 ( .B1(n7365), .B2(n10180), .A(n7238), .ZN(P2_U3402) );
  OAI21_X1 U9117 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n9510) );
  NAND2_X1 U9118 ( .A1(n9465), .A2(n7452), .ZN(n7245) );
  INV_X1 U9119 ( .A(n7242), .ZN(n7448) );
  NAND2_X1 U9120 ( .A1(n7243), .A2(n7448), .ZN(n8440) );
  AOI22_X1 U9121 ( .A1(n9460), .A2(n7446), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n8440), .ZN(n7244) );
  OAI211_X1 U9122 ( .C1(n9510), .C2(n9467), .A(n7245), .B(n7244), .ZN(P1_U3232) );
  INV_X1 U9123 ( .A(n8235), .ZN(n7327) );
  NAND2_X1 U9124 ( .A1(n7327), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U9125 ( .A1(n7318), .A2(n7246), .ZN(n7247) );
  XOR2_X1 U9126 ( .A(n8234), .B(n7247), .Z(n7456) );
  AOI211_X1 U9127 ( .C1(n7460), .C2(n7320), .A(n9885), .B(n7248), .ZN(n7465)
         );
  XOR2_X1 U9128 ( .A(n8234), .B(n7249), .Z(n7252) );
  OAI22_X1 U9129 ( .A1(n7250), .A2(n9455), .B1(n6124), .B2(n9369), .ZN(n8373)
         );
  INV_X1 U9130 ( .A(n8373), .ZN(n7251) );
  OAI21_X1 U9131 ( .B1(n7252), .B2(n9858), .A(n7251), .ZN(n7466) );
  AOI211_X1 U9132 ( .C1(n7456), .C2(n10071), .A(n7465), .B(n7466), .ZN(n7355)
         );
  AOI22_X1 U9133 ( .A1(n9940), .A2(n7460), .B1(n4655), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7253) );
  OAI21_X1 U9134 ( .B1(n7355), .B2(n4655), .A(n7253), .ZN(P1_U3524) );
  INV_X1 U9135 ( .A(n7884), .ZN(n7669) );
  INV_X1 U9136 ( .A(n7254), .ZN(n7256) );
  OAI222_X1 U9137 ( .A1(P1_U3086), .A2(n7669), .B1(n10029), .B2(n7256), .C1(
        n10440), .C2(n8378), .ZN(P1_U3339) );
  OAI222_X1 U9138 ( .A1(n9246), .A2(n7257), .B1(P2_U3151), .B2(n5989), .C1(
        n9258), .C2(n7256), .ZN(P2_U3279) );
  XOR2_X1 U9139 ( .A(n7258), .B(n7259), .Z(n7263) );
  OAI22_X1 U9140 ( .A1(n5320), .A2(n9369), .B1(n7260), .B2(n9455), .ZN(n7298)
         );
  AOI22_X1 U9141 ( .A1(n9465), .A2(n7301), .B1(n9460), .B2(n7298), .ZN(n7262)
         );
  MUX2_X1 U9142 ( .A(P1_STATE_REG_SCAN_IN), .B(n9462), .S(n10043), .Z(n7261)
         );
  OAI211_X1 U9143 ( .C1(n7263), .C2(n9467), .A(n7262), .B(n7261), .ZN(P1_U3218) );
  XNOR2_X1 U9144 ( .A(n7268), .B(n8107), .ZN(n7389) );
  XNOR2_X1 U9145 ( .A(n7389), .B(n8788), .ZN(n7271) );
  INV_X1 U9146 ( .A(n7391), .ZN(n7270) );
  OAI211_X1 U9147 ( .C1(n7269), .C2(n7271), .A(n7270), .B(n8557), .ZN(n7275)
         );
  NAND2_X1 U9148 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10087) );
  OAI21_X1 U9149 ( .B1(n8563), .B2(n10108), .A(n10087), .ZN(n7273) );
  NOR2_X1 U9150 ( .A1(n8063), .A2(n10110), .ZN(n7272) );
  AOI211_X1 U9151 ( .C1(n8561), .C2(n8787), .A(n7273), .B(n7272), .ZN(n7274)
         );
  OAI211_X1 U9152 ( .C1(n10167), .C2(n8568), .A(n7275), .B(n7274), .ZN(
        P2_U3179) );
  XOR2_X1 U9153 ( .A(n7276), .B(n7277), .Z(n7291) );
  XNOR2_X1 U9154 ( .A(n7279), .B(n7278), .ZN(n7289) );
  NAND2_X1 U9155 ( .A1(n10099), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7280) );
  NAND2_X1 U9156 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n7473) );
  OAI211_X1 U9157 ( .C1(n8928), .C2(n7281), .A(n7280), .B(n7473), .ZN(n7288)
         );
  OR3_X1 U9158 ( .A1(n7284), .A2(n7283), .A3(n7282), .ZN(n7285) );
  AOI21_X1 U9159 ( .B1(n7286), .B2(n7285), .A(n10088), .ZN(n7287) );
  AOI211_X1 U9160 ( .C1(n10092), .C2(n7289), .A(n7288), .B(n7287), .ZN(n7290)
         );
  OAI21_X1 U9161 ( .B1(n7291), .B2(n10095), .A(n7290), .ZN(P2_U3190) );
  INV_X1 U9162 ( .A(n7292), .ZN(n7350) );
  AOI22_X1 U9163 ( .A1(n9614), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10024), .ZN(n7293) );
  OAI21_X1 U9164 ( .B1(n7350), .B2(n10029), .A(n7293), .ZN(P1_U3338) );
  OAI21_X1 U9165 ( .B1(n7295), .B2(n8230), .A(n7294), .ZN(n10048) );
  INV_X1 U9166 ( .A(n7248), .ZN(n7296) );
  AOI211_X1 U9167 ( .C1(n7301), .C2(n7296), .A(n9885), .B(n4561), .ZN(n10042)
         );
  XOR2_X1 U9168 ( .A(n8230), .B(n7297), .Z(n7299) );
  AOI21_X1 U9169 ( .B1(n7299), .B2(n9878), .A(n7298), .ZN(n10051) );
  INV_X1 U9170 ( .A(n10051), .ZN(n7300) );
  AOI211_X1 U9171 ( .C1(n10071), .C2(n10048), .A(n10042), .B(n7300), .ZN(n7306) );
  AOI22_X1 U9172 ( .A1(n9940), .A2(n7301), .B1(n4655), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7302) );
  OAI21_X1 U9173 ( .B1(n7306), .B2(n4655), .A(n7302), .ZN(P1_U3525) );
  INV_X1 U9174 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7303) );
  OAI22_X1 U9175 ( .A1(n10017), .A2(n10046), .B1(n10074), .B2(n7303), .ZN(
        n7304) );
  INV_X1 U9176 ( .A(n7304), .ZN(n7305) );
  OAI21_X1 U9177 ( .B1(n7306), .B2(n10072), .A(n7305), .ZN(P1_U3462) );
  NAND3_X1 U9178 ( .A1(n8592), .A2(n7307), .A3(n10172), .ZN(n7309) );
  NAND2_X1 U9179 ( .A1(n7309), .A2(n7308), .ZN(n7310) );
  MUX2_X1 U9180 ( .A(n7310), .B(P2_REG2_REG_0__SCAN_IN), .S(n10144), .Z(n7314)
         );
  OAI22_X1 U9181 ( .A1(n10111), .A2(n7312), .B1(n7311), .B2(n10123), .ZN(n7313) );
  OR2_X1 U9182 ( .A1(n7314), .A2(n7313), .ZN(P2_U3233) );
  INV_X1 U9183 ( .A(n7315), .ZN(n7353) );
  AOI22_X1 U9184 ( .A1(n9627), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10024), .ZN(n7316) );
  OAI21_X1 U9185 ( .B1(n7353), .B2(n10029), .A(n7316), .ZN(P1_U3337) );
  INV_X1 U9186 ( .A(n7317), .ZN(n8034) );
  OAI21_X1 U9187 ( .B1(n7327), .B2(n7319), .A(n7318), .ZN(n10059) );
  OAI211_X1 U9188 ( .C1(n7321), .C2(n4588), .A(n9843), .B(n7320), .ZN(n7322)
         );
  INV_X1 U9189 ( .A(n7322), .ZN(n10056) );
  INV_X1 U9190 ( .A(n7817), .ZN(n7618) );
  NAND2_X1 U9191 ( .A1(n7323), .A2(n9457), .ZN(n7325) );
  NAND2_X1 U9192 ( .A1(n9498), .A2(n9426), .ZN(n7324) );
  NAND2_X1 U9193 ( .A1(n7325), .A2(n7324), .ZN(n8441) );
  XNOR2_X1 U9194 ( .A(n7327), .B(n7326), .ZN(n7328) );
  NOR2_X1 U9195 ( .A1(n7328), .A2(n9858), .ZN(n7329) );
  AOI211_X1 U9196 ( .C1(n7618), .C2(n10059), .A(n8441), .B(n7329), .ZN(n10062)
         );
  INV_X1 U9197 ( .A(n10062), .ZN(n7330) );
  AOI211_X1 U9198 ( .C1(n8034), .C2(n10059), .A(n10056), .B(n7330), .ZN(n7335)
         );
  INV_X1 U9199 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7331) );
  OAI22_X1 U9200 ( .A1(n10017), .A2(n4588), .B1(n10074), .B2(n7331), .ZN(n7332) );
  INV_X1 U9201 ( .A(n7332), .ZN(n7333) );
  OAI21_X1 U9202 ( .B1(n7335), .B2(n10072), .A(n7333), .ZN(P1_U3456) );
  AOI22_X1 U9203 ( .A1(n9940), .A2(n10055), .B1(n4655), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7334) );
  OAI21_X1 U9204 ( .B1(n7335), .B2(n4655), .A(n7334), .ZN(P1_U3523) );
  INV_X1 U9205 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8097) );
  OAI21_X1 U9206 ( .B1(n8097), .B2(n7337), .A(n7336), .ZN(n7480) );
  INV_X1 U9207 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7338) );
  XNOR2_X1 U9208 ( .A(n7484), .B(n7338), .ZN(n7479) );
  XNOR2_X1 U9209 ( .A(n7480), .B(n7479), .ZN(n7349) );
  NOR2_X1 U9210 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5481), .ZN(n9285) );
  NOR2_X1 U9211 ( .A1(n9592), .A2(n7339), .ZN(n7340) );
  AOI211_X1 U9212 ( .C1(n10038), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9285), .B(
        n7340), .ZN(n7348) );
  NAND2_X1 U9213 ( .A1(n7341), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7342) );
  NAND2_X1 U9214 ( .A1(n7343), .A2(n7342), .ZN(n7346) );
  INV_X1 U9215 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7344) );
  MUX2_X1 U9216 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n7344), .S(n7484), .Z(n7345)
         );
  NAND2_X1 U9217 ( .A1(n7346), .A2(n7345), .ZN(n7486) );
  OAI211_X1 U9218 ( .C1(n7346), .C2(n7345), .A(n7486), .B(n9638), .ZN(n7347)
         );
  OAI211_X1 U9219 ( .C1(n7349), .C2(n9633), .A(n7348), .B(n7347), .ZN(P1_U3257) );
  OAI222_X1 U9220 ( .A1(n9246), .A2(n7351), .B1(n9258), .B2(n7350), .C1(n8906), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OAI222_X1 U9221 ( .A1(n9258), .A2(n7353), .B1(P2_U3151), .B2(n8932), .C1(
        n7352), .C2(n9246), .ZN(P2_U3277) );
  AOI22_X1 U9222 ( .A1(n6861), .A2(n7460), .B1(n10072), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n7354) );
  OAI21_X1 U9223 ( .B1(n7355), .B2(n10072), .A(n7354), .ZN(P1_U3459) );
  INV_X1 U9224 ( .A(n7356), .ZN(n7357) );
  AOI211_X1 U9225 ( .C1(n7359), .C2(n7358), .A(n9467), .B(n7357), .ZN(n7362)
         );
  AOI22_X1 U9226 ( .A1(n9426), .A2(n9495), .B1(n9497), .B2(n9457), .ZN(n7551)
         );
  AOI22_X1 U9227 ( .A1(n9465), .A2(n7548), .B1(n9442), .B2(n7547), .ZN(n7360)
         );
  NAND2_X1 U9228 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9544) );
  OAI211_X1 U9229 ( .C1(n7551), .C2(n9444), .A(n7360), .B(n9544), .ZN(n7361)
         );
  OR2_X1 U9230 ( .A1(n7362), .A2(n7361), .ZN(P1_U3230) );
  AOI22_X1 U9231 ( .A1(n9154), .A2(n7363), .B1(n10187), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n7364) );
  OAI21_X1 U9232 ( .B1(n7365), .B2(n10187), .A(n7364), .ZN(P2_U3463) );
  NAND2_X1 U9233 ( .A1(n7294), .A2(n7366), .ZN(n7546) );
  NAND2_X1 U9234 ( .A1(n7546), .A2(n8229), .ZN(n7545) );
  INV_X1 U9235 ( .A(n7367), .ZN(n8232) );
  NAND3_X1 U9236 ( .A1(n7545), .A2(n8232), .A3(n7368), .ZN(n7370) );
  NAND2_X1 U9237 ( .A1(n7370), .A2(n7369), .ZN(n7607) );
  AOI211_X1 U9238 ( .C1(n7496), .C2(n7371), .A(n9885), .B(n5116), .ZN(n7602)
         );
  XNOR2_X1 U9239 ( .A(n7372), .B(n8232), .ZN(n7373) );
  AOI22_X1 U9240 ( .A1(n9426), .A2(n9494), .B1(n9496), .B2(n9457), .ZN(n7498)
         );
  OAI21_X1 U9241 ( .B1(n7373), .B2(n9858), .A(n7498), .ZN(n7601) );
  AOI211_X1 U9242 ( .C1(n10071), .C2(n7607), .A(n7602), .B(n7601), .ZN(n7378)
         );
  INV_X1 U9243 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7374) );
  OAI22_X1 U9244 ( .A1(n10017), .A2(n5280), .B1(n10074), .B2(n7374), .ZN(n7375) );
  INV_X1 U9245 ( .A(n7375), .ZN(n7376) );
  OAI21_X1 U9246 ( .B1(n7378), .B2(n10072), .A(n7376), .ZN(P1_U3468) );
  AOI22_X1 U9247 ( .A1(n9940), .A2(n7496), .B1(n4655), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7377) );
  OAI21_X1 U9248 ( .B1(n7378), .B2(n4655), .A(n7377), .ZN(P1_U3527) );
  INV_X1 U9249 ( .A(n7379), .ZN(n8593) );
  XNOR2_X1 U9250 ( .A(n7380), .B(n8593), .ZN(n10158) );
  INV_X1 U9251 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7386) );
  XNOR2_X1 U9252 ( .A(n7381), .B(n8593), .ZN(n7385) );
  NAND2_X1 U9253 ( .A1(n8790), .A2(n6698), .ZN(n7382) );
  OAI21_X1 U9254 ( .B1(n7406), .B2(n10125), .A(n7382), .ZN(n7384) );
  AOI21_X1 U9255 ( .B1(n7385), .B2(n9094), .A(n7384), .ZN(n10156) );
  MUX2_X1 U9256 ( .A(n7386), .B(n10156), .S(n10141), .Z(n7388) );
  AOI22_X1 U9257 ( .A1(n9109), .A2(n7084), .B1(n9096), .B2(n10225), .ZN(n7387)
         );
  OAI211_X1 U9258 ( .C1(n10115), .C2(n10158), .A(n7388), .B(n7387), .ZN(
        P2_U3230) );
  INV_X1 U9259 ( .A(n7392), .ZN(n10173) );
  INV_X1 U9260 ( .A(n7389), .ZN(n7390) );
  XNOR2_X1 U9261 ( .A(n7392), .B(n8107), .ZN(n7470) );
  XNOR2_X1 U9262 ( .A(n7470), .B(n8787), .ZN(n7393) );
  OAI21_X1 U9263 ( .B1(n7394), .B2(n7393), .A(n7472), .ZN(n7395) );
  NAND2_X1 U9264 ( .A1(n7395), .A2(n8557), .ZN(n7401) );
  INV_X1 U9265 ( .A(n7439), .ZN(n7399) );
  AOI21_X1 U9266 ( .B1(n8539), .B2(n8788), .A(n7396), .ZN(n7397) );
  OAI21_X1 U9267 ( .B1(n7805), .B2(n8541), .A(n7397), .ZN(n7398) );
  AOI21_X1 U9268 ( .B1(n7399), .B2(n8565), .A(n7398), .ZN(n7400) );
  OAI211_X1 U9269 ( .C1(n10173), .C2(n8568), .A(n7401), .B(n7400), .ZN(
        P2_U3153) );
  XNOR2_X1 U9270 ( .A(n4620), .B(n8623), .ZN(n10145) );
  OAI21_X1 U9271 ( .B1(n7403), .B2(n4620), .A(n10131), .ZN(n7408) );
  NAND2_X1 U9272 ( .A1(n7404), .A2(n9090), .ZN(n7405) );
  OAI21_X1 U9273 ( .B1(n7406), .B2(n10127), .A(n7405), .ZN(n7407) );
  AOI21_X1 U9274 ( .B1(n7408), .B2(n9094), .A(n7407), .ZN(n10146) );
  MUX2_X1 U9275 ( .A(n10472), .B(n10146), .S(n10141), .Z(n7411) );
  AOI22_X1 U9276 ( .A1(n9109), .A2(n7409), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9096), .ZN(n7410) );
  OAI211_X1 U9277 ( .C1(n10145), .C2(n10115), .A(n7411), .B(n7410), .ZN(
        P2_U3232) );
  OAI21_X1 U9278 ( .B1(n7412), .B2(n8596), .A(n4450), .ZN(n10163) );
  INV_X1 U9279 ( .A(n10163), .ZN(n7418) );
  XOR2_X1 U9280 ( .A(n7413), .B(n8596), .Z(n7414) );
  AOI222_X1 U9281 ( .A1(n9094), .A2(n7414), .B1(n8788), .B2(n6698), .C1(n8790), 
        .C2(n9090), .ZN(n10165) );
  MUX2_X1 U9282 ( .A(n10303), .B(n10165), .S(n10141), .Z(n7417) );
  AOI22_X1 U9283 ( .A1(n9109), .A2(n6739), .B1(n9096), .B2(n7415), .ZN(n7416)
         );
  OAI211_X1 U9284 ( .C1(n7418), .C2(n10115), .A(n7417), .B(n7416), .ZN(
        P2_U3228) );
  NAND2_X1 U9285 ( .A1(n7638), .A2(n8599), .ZN(n7802) );
  OAI211_X1 U9286 ( .C1(n7638), .C2(n8599), .A(n7802), .B(n9094), .ZN(n7422)
         );
  AOI22_X1 U9287 ( .A1(n9090), .A2(n8787), .B1(n8785), .B2(n6698), .ZN(n7421)
         );
  AND2_X1 U9288 ( .A1(n7422), .A2(n7421), .ZN(n7538) );
  AOI22_X1 U9289 ( .A1(n6799), .A2(n7541), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10180), .ZN(n7426) );
  XNOR2_X1 U9290 ( .A(n7424), .B(n8599), .ZN(n7536) );
  INV_X1 U9291 ( .A(n9234), .ZN(n9240) );
  NAND2_X1 U9292 ( .A1(n7536), .A2(n9240), .ZN(n7425) );
  OAI211_X1 U9293 ( .C1(n7538), .C2(n10180), .A(n7426), .B(n7425), .ZN(
        P2_U3414) );
  INV_X1 U9294 ( .A(n7427), .ZN(n7429) );
  OAI222_X1 U9295 ( .A1(n9246), .A2(n10312), .B1(n9258), .B2(n7429), .C1(n8612), .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9296 ( .A1(n8378), .A2(n7430), .B1(n10029), .B2(n7429), .C1(
        P1_U3086), .C2(n7428), .ZN(P1_U3336) );
  INV_X1 U9297 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7442) );
  OR2_X1 U9298 ( .A1(n7432), .A2(n8598), .ZN(n7433) );
  NAND2_X1 U9299 ( .A1(n7434), .A2(n7433), .ZN(n10175) );
  XNOR2_X1 U9300 ( .A(n7435), .B(n8598), .ZN(n7436) );
  NAND2_X1 U9301 ( .A1(n7436), .A2(n9094), .ZN(n7438) );
  AOI22_X1 U9302 ( .A1(n9090), .A2(n8788), .B1(n8786), .B2(n6698), .ZN(n7437)
         );
  OAI211_X1 U9303 ( .C1(n10124), .C2(n10175), .A(n7438), .B(n7437), .ZN(n10177) );
  OAI22_X1 U9304 ( .A1(n10175), .A2(n8947), .B1(n7439), .B2(n10123), .ZN(n7440) );
  NOR2_X1 U9305 ( .A1(n10177), .A2(n7440), .ZN(n7441) );
  MUX2_X1 U9306 ( .A(n7442), .B(n7441), .S(n10141), .Z(n7443) );
  OAI21_X1 U9307 ( .B1(n10173), .B2(n10111), .A(n7443), .ZN(P2_U3226) );
  INV_X1 U9308 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U9309 ( .A1(n8231), .A2(n7444), .ZN(n7445) );
  AOI211_X1 U9310 ( .C1(n10052), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7446), .B(
        n7445), .ZN(n7455) );
  NAND3_X1 U9311 ( .A1(n7449), .A2(n7448), .A3(n7447), .ZN(n7450) );
  NAND2_X1 U9312 ( .A1(n10063), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U9313 ( .A1(n10057), .A2(n9843), .ZN(n9667) );
  INV_X1 U9314 ( .A(n9667), .ZN(n9645) );
  OAI21_X1 U9315 ( .B1(n9645), .B2(n10054), .A(n7452), .ZN(n7453) );
  OAI211_X1 U9316 ( .C1(n7455), .C2(n10063), .A(n7454), .B(n7453), .ZN(
        P1_U3293) );
  INV_X1 U9317 ( .A(n7456), .ZN(n7469) );
  NAND2_X1 U9318 ( .A1(n5780), .A2(n7457), .ZN(n7458) );
  NAND2_X1 U9319 ( .A1(n10054), .A2(n7460), .ZN(n7462) );
  NAND2_X1 U9320 ( .A1(n10052), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7461) );
  OAI211_X1 U9321 ( .C1(n7463), .C2(n9850), .A(n7462), .B(n7461), .ZN(n7464)
         );
  AOI21_X1 U9322 ( .B1(n10057), .B2(n7465), .A(n7464), .ZN(n7468) );
  NAND2_X1 U9323 ( .A1(n7466), .A2(n9850), .ZN(n7467) );
  OAI211_X1 U9324 ( .C1(n7469), .C2(n9852), .A(n7468), .B(n7467), .ZN(P1_U3291) );
  NAND2_X1 U9325 ( .A1(n7470), .A2(n10109), .ZN(n7471) );
  XNOR2_X1 U9326 ( .A(n7541), .B(n8107), .ZN(n7556) );
  XNOR2_X1 U9327 ( .A(n7556), .B(n8786), .ZN(n7557) );
  XOR2_X1 U9328 ( .A(n7558), .B(n7557), .Z(n7478) );
  OAI21_X1 U9329 ( .B1(n8541), .B2(n7862), .A(n7473), .ZN(n7474) );
  AOI21_X1 U9330 ( .B1(n8539), .B2(n8787), .A(n7474), .ZN(n7475) );
  OAI21_X1 U9331 ( .B1(n8063), .B2(n7539), .A(n7475), .ZN(n7476) );
  AOI21_X1 U9332 ( .B1(n7541), .B2(n8553), .A(n7476), .ZN(n7477) );
  OAI21_X1 U9333 ( .B1(n7478), .B2(n8555), .A(n7477), .ZN(P2_U3161) );
  XOR2_X1 U9334 ( .A(n7672), .B(n7665), .Z(n7666) );
  INV_X1 U9335 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10353) );
  XNOR2_X1 U9336 ( .A(n7666), .B(n10353), .ZN(n7490) );
  NOR2_X1 U9337 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7481), .ZN(n7483) );
  NOR2_X1 U9338 ( .A1(n9592), .A2(n7664), .ZN(n7482) );
  AOI211_X1 U9339 ( .C1(n10038), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7483), .B(
        n7482), .ZN(n7489) );
  NAND2_X1 U9340 ( .A1(n7484), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U9341 ( .A1(n7486), .A2(n7485), .ZN(n7673) );
  XNOR2_X1 U9342 ( .A(n7673), .B(n7664), .ZN(n7487) );
  NAND2_X1 U9343 ( .A1(n7487), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7675) );
  OAI211_X1 U9344 ( .C1(n7487), .C2(P1_REG2_REG_15__SCAN_IN), .A(n7675), .B(
        n9638), .ZN(n7488) );
  OAI211_X1 U9345 ( .C1(n7490), .C2(n9633), .A(n7489), .B(n7488), .ZN(P1_U3258) );
  INV_X1 U9346 ( .A(n7491), .ZN(n7495) );
  XNOR2_X1 U9347 ( .A(n7492), .B(n7493), .ZN(n7494) );
  NAND2_X1 U9348 ( .A1(n7494), .A2(n7495), .ZN(n7686) );
  OAI21_X1 U9349 ( .B1(n7495), .B2(n7494), .A(n7686), .ZN(n7500) );
  AOI22_X1 U9350 ( .A1(n9465), .A2(n7496), .B1(n9442), .B2(n7603), .ZN(n7497)
         );
  NAND2_X1 U9351 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9566) );
  OAI211_X1 U9352 ( .C1(n7498), .C2(n9444), .A(n7497), .B(n9566), .ZN(n7499)
         );
  AOI21_X1 U9353 ( .B1(n7500), .B2(n9434), .A(n7499), .ZN(n7501) );
  INV_X1 U9354 ( .A(n7501), .ZN(P1_U3227) );
  MUX2_X1 U9355 ( .A(n7538), .B(n7502), .S(n10187), .Z(n7504) );
  INV_X1 U9356 ( .A(n9147), .ZN(n9155) );
  AOI22_X1 U9357 ( .A1(n7536), .A2(n9155), .B1(n9154), .B2(n7541), .ZN(n7503)
         );
  NAND2_X1 U9358 ( .A1(n7504), .A2(n7503), .ZN(P2_U3467) );
  NAND2_X1 U9359 ( .A1(n7369), .A2(n7505), .ZN(n7506) );
  NAND2_X1 U9360 ( .A1(n7506), .A2(n8236), .ZN(n7612) );
  OAI21_X1 U9361 ( .B1(n7506), .B2(n8236), .A(n7612), .ZN(n7662) );
  AOI211_X1 U9362 ( .C1(n7692), .C2(n7508), .A(n9885), .B(n7507), .ZN(n7656)
         );
  XOR2_X1 U9363 ( .A(n4448), .B(n8236), .Z(n7513) );
  OAI22_X1 U9364 ( .A1(n7511), .A2(n9455), .B1(n7510), .B2(n9369), .ZN(n7690)
         );
  INV_X1 U9365 ( .A(n7690), .ZN(n7512) );
  OAI21_X1 U9366 ( .B1(n7513), .B2(n9858), .A(n7512), .ZN(n7659) );
  AOI211_X1 U9367 ( .C1(n10071), .C2(n7662), .A(n7656), .B(n7659), .ZN(n7519)
         );
  AOI22_X1 U9368 ( .A1(n9940), .A2(n7692), .B1(n4655), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7514) );
  OAI21_X1 U9369 ( .B1(n7519), .B2(n4655), .A(n7514), .ZN(P1_U3528) );
  INV_X1 U9370 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7515) );
  OAI22_X1 U9371 ( .A1(n10017), .A2(n7516), .B1(n10074), .B2(n7515), .ZN(n7517) );
  INV_X1 U9372 ( .A(n7517), .ZN(n7518) );
  OAI21_X1 U9373 ( .B1(n7519), .B2(n10072), .A(n7518), .ZN(P1_U3471) );
  XNOR2_X1 U9374 ( .A(n7520), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7531) );
  XNOR2_X1 U9375 ( .A(n7522), .B(n7521), .ZN(n7529) );
  AOI21_X1 U9376 ( .B1(n7524), .B2(n7523), .A(n4489), .ZN(n7527) );
  NAND2_X1 U9377 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7562) );
  OAI21_X1 U9378 ( .B1(n8928), .B2(n4768), .A(n7562), .ZN(n7525) );
  AOI21_X1 U9379 ( .B1(n10099), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7525), .ZN(
        n7526) );
  OAI21_X1 U9380 ( .B1(n7527), .B2(n10088), .A(n7526), .ZN(n7528) );
  AOI21_X1 U9381 ( .B1(n8883), .B2(n7529), .A(n7528), .ZN(n7530) );
  OAI21_X1 U9382 ( .B1(n7531), .B2(n8939), .A(n7530), .ZN(P2_U3191) );
  NAND2_X1 U9383 ( .A1(n8363), .A2(n7532), .ZN(n7534) );
  OAI211_X1 U9384 ( .C1(n7535), .C2(n8378), .A(n7534), .B(n7533), .ZN(P1_U3335) );
  INV_X1 U9385 ( .A(n7536), .ZN(n7544) );
  MUX2_X1 U9386 ( .A(n7538), .B(n7537), .S(n10144), .Z(n7543) );
  INV_X1 U9387 ( .A(n7539), .ZN(n7540) );
  AOI22_X1 U9388 ( .A1(n9109), .A2(n7541), .B1(n7540), .B2(n9096), .ZN(n7542)
         );
  OAI211_X1 U9389 ( .C1(n7544), .C2(n10115), .A(n7543), .B(n7542), .ZN(
        P2_U3225) );
  OAI21_X1 U9390 ( .B1(n7546), .B2(n8229), .A(n7545), .ZN(n10070) );
  OAI211_X1 U9391 ( .C1(n4561), .C2(n10067), .A(n9843), .B(n7371), .ZN(n10065)
         );
  AOI22_X1 U9392 ( .A1(n10054), .A2(n7548), .B1(n10052), .B2(n7547), .ZN(n7549) );
  OAI21_X1 U9393 ( .B1(n10065), .B2(n9814), .A(n7549), .ZN(n7554) );
  XOR2_X1 U9394 ( .A(n7550), .B(n8229), .Z(n7552) );
  OAI21_X1 U9395 ( .B1(n7552), .B2(n9858), .A(n7551), .ZN(n10068) );
  MUX2_X1 U9396 ( .A(n10068), .B(P1_REG2_REG_4__SCAN_IN), .S(n10063), .Z(n7553) );
  AOI211_X1 U9397 ( .C1(n10049), .C2(n10070), .A(n7554), .B(n7553), .ZN(n7555)
         );
  INV_X1 U9398 ( .A(n7555), .ZN(P1_U3289) );
  INV_X1 U9399 ( .A(n7559), .ZN(n7921) );
  XNOR2_X1 U9400 ( .A(n7559), .B(n8107), .ZN(n7863) );
  XNOR2_X1 U9401 ( .A(n7863), .B(n8785), .ZN(n7561) );
  OAI211_X1 U9402 ( .C1(n7560), .C2(n7561), .A(n7865), .B(n8557), .ZN(n7567)
         );
  INV_X1 U9403 ( .A(n7920), .ZN(n7565) );
  NAND2_X1 U9404 ( .A1(n8561), .A2(n8784), .ZN(n7563) );
  OAI211_X1 U9405 ( .C1(n7805), .C2(n8563), .A(n7563), .B(n7562), .ZN(n7564)
         );
  AOI21_X1 U9406 ( .B1(n7565), .B2(n8565), .A(n7564), .ZN(n7566) );
  OAI211_X1 U9407 ( .C1(n7921), .C2(n8568), .A(n7567), .B(n7566), .ZN(P2_U3171) );
  OAI21_X1 U9408 ( .B1(n7569), .B2(n7568), .A(n7943), .ZN(n7576) );
  NOR2_X1 U9409 ( .A1(n9412), .A2(n4466), .ZN(n7575) );
  INV_X1 U9410 ( .A(n7570), .ZN(n7624) );
  OR2_X1 U9411 ( .A1(n5232), .A2(n9369), .ZN(n7572) );
  NAND2_X1 U9412 ( .A1(n9492), .A2(n9426), .ZN(n7571) );
  NAND2_X1 U9413 ( .A1(n7572), .A2(n7571), .ZN(n7617) );
  NAND2_X1 U9414 ( .A1(n9460), .A2(n7617), .ZN(n7573) );
  NAND2_X1 U9415 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9590) );
  OAI211_X1 U9416 ( .C1(n9462), .C2(n7624), .A(n7573), .B(n9590), .ZN(n7574)
         );
  AOI211_X1 U9417 ( .C1(n7576), .C2(n9434), .A(n7575), .B(n7574), .ZN(n7577)
         );
  INV_X1 U9418 ( .A(n7577), .ZN(P1_U3213) );
  XNOR2_X1 U9419 ( .A(n7578), .B(n7870), .ZN(n7579) );
  AOI222_X1 U9420 ( .A1(n9094), .A2(n7579), .B1(n8782), .B2(n6698), .C1(n8784), 
        .C2(n9090), .ZN(n7785) );
  AOI22_X1 U9421 ( .A1(n4615), .A2(n9154), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n10187), .ZN(n7583) );
  OAI21_X1 U9422 ( .B1(n7581), .B2(n7870), .A(n7580), .ZN(n7784) );
  NAND2_X1 U9423 ( .A1(n7784), .A2(n9155), .ZN(n7582) );
  OAI211_X1 U9424 ( .C1(n7785), .C2(n10187), .A(n7583), .B(n7582), .ZN(
        P2_U3470) );
  AOI22_X1 U9425 ( .A1(n4615), .A2(n6799), .B1(P2_REG0_REG_11__SCAN_IN), .B2(
        n10180), .ZN(n7585) );
  NAND2_X1 U9426 ( .A1(n7784), .A2(n9240), .ZN(n7584) );
  OAI211_X1 U9427 ( .C1(n7785), .C2(n10180), .A(n7585), .B(n7584), .ZN(
        P2_U3423) );
  XOR2_X1 U9428 ( .A(n7587), .B(n7586), .Z(n7600) );
  XNOR2_X1 U9429 ( .A(n7589), .B(n7588), .ZN(n7598) );
  NAND2_X1 U9430 ( .A1(n10099), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9431 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7903) );
  OAI211_X1 U9432 ( .C1(n8928), .C2(n7591), .A(n7590), .B(n7903), .ZN(n7597)
         );
  OR3_X1 U9433 ( .A1(n4489), .A2(n7593), .A3(n7592), .ZN(n7594) );
  AOI21_X1 U9434 ( .B1(n7595), .B2(n7594), .A(n10088), .ZN(n7596) );
  AOI211_X1 U9435 ( .C1(n8883), .C2(n7598), .A(n7597), .B(n7596), .ZN(n7599)
         );
  OAI21_X1 U9436 ( .B1(n7600), .B2(n8939), .A(n7599), .ZN(P2_U3192) );
  INV_X1 U9437 ( .A(n7601), .ZN(n7609) );
  NAND2_X1 U9438 ( .A1(n7602), .A2(n10057), .ZN(n7605) );
  AOI22_X1 U9439 ( .A1(n10063), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7603), .B2(
        n10052), .ZN(n7604) );
  OAI211_X1 U9440 ( .C1(n5280), .C2(n9891), .A(n7605), .B(n7604), .ZN(n7606)
         );
  AOI21_X1 U9441 ( .B1(n10049), .B2(n7607), .A(n7606), .ZN(n7608) );
  OAI21_X1 U9442 ( .B1(n7609), .B2(n10063), .A(n7608), .ZN(P1_U3288) );
  INV_X1 U9443 ( .A(n7610), .ZN(n7720) );
  NAND3_X1 U9444 ( .A1(n7612), .A2(n7720), .A3(n7611), .ZN(n7614) );
  NAND2_X1 U9445 ( .A1(n7614), .A2(n7613), .ZN(n7648) );
  INV_X1 U9446 ( .A(n7648), .ZN(n7628) );
  XNOR2_X1 U9447 ( .A(n7721), .B(n7720), .ZN(n7620) );
  AOI21_X1 U9448 ( .B1(n7648), .B2(n7618), .A(n7617), .ZN(n7619) );
  OAI21_X1 U9449 ( .B1(n7620), .B2(n9858), .A(n7619), .ZN(n7646) );
  INV_X1 U9450 ( .A(n7646), .ZN(n7621) );
  MUX2_X1 U9451 ( .A(n6950), .B(n7621), .S(n9850), .Z(n7627) );
  OR2_X1 U9452 ( .A1(n7507), .A2(n4466), .ZN(n7623) );
  AND3_X1 U9453 ( .A1(n7622), .A2(n9843), .A3(n7623), .ZN(n7647) );
  OAI22_X1 U9454 ( .A1(n9891), .A2(n4466), .B1(n9829), .B2(n7624), .ZN(n7625)
         );
  AOI21_X1 U9455 ( .B1(n7647), .B2(n10057), .A(n7625), .ZN(n7626) );
  OAI211_X1 U9456 ( .C1(n7628), .C2(n10053), .A(n7627), .B(n7626), .ZN(
        P1_U3286) );
  OAI22_X1 U9457 ( .A1(n10111), .A2(n8638), .B1(n7629), .B2(n10123), .ZN(n7632) );
  MUX2_X1 U9458 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7630), .S(n10141), .Z(n7631)
         );
  AOI211_X1 U9459 ( .C1(n8992), .C2(n7633), .A(n7632), .B(n7631), .ZN(n7634)
         );
  INV_X1 U9460 ( .A(n7634), .ZN(P2_U3229) );
  INV_X1 U9461 ( .A(n7639), .ZN(n8603) );
  XNOR2_X1 U9462 ( .A(n7635), .B(n8603), .ZN(n7644) );
  INV_X1 U9463 ( .A(n7644), .ZN(n7754) );
  OAI21_X1 U9464 ( .B1(n7638), .B2(n7637), .A(n7636), .ZN(n7640) );
  XNOR2_X1 U9465 ( .A(n7640), .B(n7639), .ZN(n7641) );
  NAND2_X1 U9466 ( .A1(n7641), .A2(n9094), .ZN(n7643) );
  AOI22_X1 U9467 ( .A1(n9090), .A2(n8785), .B1(n8783), .B2(n6698), .ZN(n7642)
         );
  OAI211_X1 U9468 ( .C1(n7644), .C2(n10124), .A(n7643), .B(n7642), .ZN(n7753)
         );
  AOI21_X1 U9469 ( .B1(n10151), .B2(n7754), .A(n7753), .ZN(n7781) );
  AOI22_X1 U9470 ( .A1(n6799), .A2(n7909), .B1(n10180), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n7645) );
  OAI21_X1 U9471 ( .B1(n7781), .B2(n10180), .A(n7645), .ZN(P2_U3420) );
  AOI211_X1 U9472 ( .C1(n8034), .C2(n7648), .A(n7647), .B(n7646), .ZN(n7655)
         );
  INV_X1 U9473 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7649) );
  OAI22_X1 U9474 ( .A1(n10017), .A2(n4466), .B1(n10074), .B2(n7649), .ZN(n7651) );
  INV_X1 U9475 ( .A(n7651), .ZN(n7652) );
  OAI21_X1 U9476 ( .B1(n7655), .B2(n10072), .A(n7652), .ZN(P1_U3474) );
  AOI22_X1 U9477 ( .A1(n9940), .A2(n7653), .B1(n4655), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7654) );
  OAI21_X1 U9478 ( .B1(n7655), .B2(n4655), .A(n7654), .ZN(P1_U3529) );
  INV_X1 U9479 ( .A(n7656), .ZN(n7658) );
  AOI22_X1 U9480 ( .A1(n10054), .A2(n7692), .B1(n10052), .B2(n7691), .ZN(n7657) );
  OAI21_X1 U9481 ( .B1(n7658), .B2(n9814), .A(n7657), .ZN(n7661) );
  MUX2_X1 U9482 ( .A(n7659), .B(P1_REG2_REG_6__SCAN_IN), .S(n10063), .Z(n7660)
         );
  AOI211_X1 U9483 ( .C1(n10049), .C2(n7662), .A(n7661), .B(n7660), .ZN(n7663)
         );
  INV_X1 U9484 ( .A(n7663), .ZN(P1_U3287) );
  OAI22_X1 U9485 ( .A1(n7666), .A2(n10353), .B1(n7665), .B2(n7664), .ZN(n7668)
         );
  INV_X1 U9486 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U9487 ( .A1(n7669), .A2(n9954), .ZN(n7891) );
  OAI21_X1 U9488 ( .B1(n7669), .B2(n9954), .A(n7891), .ZN(n7667) );
  AOI21_X1 U9489 ( .B1(n7668), .B2(n7667), .A(n7893), .ZN(n7681) );
  NOR2_X1 U9490 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5524), .ZN(n7671) );
  NOR2_X1 U9491 ( .A1(n9592), .A2(n7669), .ZN(n7670) );
  AOI211_X1 U9492 ( .C1(n10038), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n7671), .B(
        n7670), .ZN(n7680) );
  NAND2_X1 U9493 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NAND2_X1 U9494 ( .A1(n7675), .A2(n7674), .ZN(n7678) );
  INV_X1 U9495 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7676) );
  MUX2_X1 U9496 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n7676), .S(n7884), .Z(n7677)
         );
  NAND2_X1 U9497 ( .A1(n7678), .A2(n7677), .ZN(n7886) );
  OAI211_X1 U9498 ( .C1(n7678), .C2(n7677), .A(n7886), .B(n9638), .ZN(n7679)
         );
  OAI211_X1 U9499 ( .C1(n7681), .C2(n9633), .A(n7680), .B(n7679), .ZN(P1_U3259) );
  INV_X1 U9500 ( .A(n7682), .ZN(n7684) );
  AOI21_X1 U9501 ( .B1(n7685), .B2(n7684), .A(n7683), .ZN(n7689) );
  OAI21_X1 U9502 ( .B1(n7687), .B2(n7492), .A(n7686), .ZN(n7688) );
  XOR2_X1 U9503 ( .A(n7689), .B(n7688), .Z(n7695) );
  AOI22_X1 U9504 ( .A1(n9460), .A2(n7690), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7694) );
  AOI22_X1 U9505 ( .A1(n9465), .A2(n7692), .B1(n9442), .B2(n7691), .ZN(n7693)
         );
  OAI211_X1 U9506 ( .C1(n7695), .C2(n9467), .A(n7694), .B(n7693), .ZN(P1_U3239) );
  OAI21_X1 U9507 ( .B1(n7698), .B2(n7697), .A(n7696), .ZN(n7839) );
  INV_X1 U9508 ( .A(n7839), .ZN(n7713) );
  OAI21_X1 U9509 ( .B1(n7700), .B2(n8245), .A(n7699), .ZN(n7703) );
  OR2_X1 U9510 ( .A1(n7741), .A2(n9369), .ZN(n7702) );
  NAND2_X1 U9511 ( .A1(n9489), .A2(n9426), .ZN(n7701) );
  NAND2_X1 U9512 ( .A1(n7702), .A2(n7701), .ZN(n7963) );
  AOI21_X1 U9513 ( .B1(n7703), .B2(n9878), .A(n7963), .ZN(n7836) );
  MUX2_X1 U9514 ( .A(n7836), .B(n7704), .S(n10063), .Z(n7712) );
  INV_X1 U9515 ( .A(n7705), .ZN(n7707) );
  AOI211_X1 U9516 ( .C1(n7707), .C2(n7968), .A(n9885), .B(n7706), .ZN(n7838)
         );
  INV_X1 U9517 ( .A(n7708), .ZN(n7966) );
  OAI22_X1 U9518 ( .A1(n7709), .A2(n9891), .B1(n9829), .B2(n7966), .ZN(n7710)
         );
  AOI21_X1 U9519 ( .B1(n7838), .B2(n10057), .A(n7710), .ZN(n7711) );
  OAI211_X1 U9520 ( .C1(n9852), .C2(n7713), .A(n7712), .B(n7711), .ZN(P1_U3283) );
  NAND2_X1 U9521 ( .A1(n7613), .A2(n7714), .ZN(n7738) );
  INV_X1 U9522 ( .A(n7740), .ZN(n7737) );
  NAND2_X1 U9523 ( .A1(n7738), .A2(n7737), .ZN(n7736) );
  INV_X1 U9524 ( .A(n7715), .ZN(n7716) );
  NOR2_X1 U9525 ( .A1(n7723), .A2(n7716), .ZN(n7717) );
  NAND2_X1 U9526 ( .A1(n7736), .A2(n7717), .ZN(n7719) );
  NAND2_X1 U9527 ( .A1(n7719), .A2(n7718), .ZN(n7858) );
  INV_X1 U9528 ( .A(n7858), .ZN(n7735) );
  INV_X1 U9529 ( .A(n7723), .ZN(n8242) );
  XNOR2_X1 U9530 ( .A(n8126), .B(n8242), .ZN(n7725) );
  AND2_X1 U9531 ( .A1(n9492), .A2(n9457), .ZN(n7951) );
  INV_X1 U9532 ( .A(n7951), .ZN(n7724) );
  OAI21_X1 U9533 ( .B1(n7725), .B2(n9858), .A(n7724), .ZN(n7856) );
  NAND2_X1 U9534 ( .A1(n7856), .A2(n9850), .ZN(n7734) );
  INV_X1 U9535 ( .A(n7727), .ZN(n7958) );
  XNOR2_X1 U9536 ( .A(n5118), .B(n7958), .ZN(n7729) );
  NOR2_X1 U9537 ( .A1(n7728), .A2(n9455), .ZN(n7950) );
  AOI21_X1 U9538 ( .B1(n7729), .B2(n9843), .A(n7950), .ZN(n7855) );
  INV_X1 U9539 ( .A(n7855), .ZN(n7732) );
  AOI22_X1 U9540 ( .A1(n10063), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7949), .B2(
        n10052), .ZN(n7730) );
  OAI21_X1 U9541 ( .B1(n7958), .B2(n9891), .A(n7730), .ZN(n7731) );
  AOI21_X1 U9542 ( .B1(n7732), .B2(n10057), .A(n7731), .ZN(n7733) );
  OAI211_X1 U9543 ( .C1(n9852), .C2(n7735), .A(n7734), .B(n7733), .ZN(P1_U3284) );
  OAI21_X1 U9544 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7792) );
  INV_X1 U9545 ( .A(n7792), .ZN(n7750) );
  XNOR2_X1 U9546 ( .A(n7739), .B(n7740), .ZN(n7745) );
  OR2_X1 U9547 ( .A1(n7741), .A2(n9455), .ZN(n7743) );
  NAND2_X1 U9548 ( .A1(n9493), .A2(n9457), .ZN(n7742) );
  NAND2_X1 U9549 ( .A1(n7743), .A2(n7742), .ZN(n9315) );
  INV_X1 U9550 ( .A(n9315), .ZN(n7744) );
  OAI21_X1 U9551 ( .B1(n7745), .B2(n9858), .A(n7744), .ZN(n7790) );
  INV_X1 U9552 ( .A(n7790), .ZN(n7746) );
  MUX2_X1 U9553 ( .A(n10357), .B(n7746), .S(n9850), .Z(n7749) );
  AOI211_X1 U9554 ( .C1(n9325), .C2(n7622), .A(n9885), .B(n7726), .ZN(n7791)
         );
  OAI22_X1 U9555 ( .A1(n9891), .A2(n5115), .B1(n9829), .B2(n9318), .ZN(n7747)
         );
  AOI21_X1 U9556 ( .B1(n7791), .B2(n10057), .A(n7747), .ZN(n7748) );
  OAI211_X1 U9557 ( .C1(n9852), .C2(n7750), .A(n7749), .B(n7748), .ZN(P1_U3285) );
  INV_X1 U9558 ( .A(n7751), .ZN(n7811) );
  OAI222_X1 U9559 ( .A1(n8378), .A2(n7752), .B1(n10029), .B2(n7811), .C1(n8303), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U9560 ( .A(n8947), .ZN(n10140) );
  AOI21_X1 U9561 ( .B1(n10140), .B2(n7754), .A(n7753), .ZN(n7755) );
  MUX2_X1 U9562 ( .A(n7756), .B(n7755), .S(n10141), .Z(n7758) );
  NAND2_X1 U9563 ( .A1(n7909), .A2(n9109), .ZN(n7757) );
  OAI211_X1 U9564 ( .C1(n7907), .C2(n10123), .A(n7758), .B(n7757), .ZN(
        P2_U3223) );
  INV_X1 U9565 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U9566 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7759) );
  AOI21_X1 U9567 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7759), .ZN(n10201) );
  NOR2_X1 U9568 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7760) );
  AOI21_X1 U9569 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7760), .ZN(n10204) );
  NOR2_X1 U9570 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7761) );
  AOI21_X1 U9571 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7761), .ZN(n10207) );
  NOR2_X1 U9572 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7762) );
  AOI21_X1 U9573 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7762), .ZN(n10210) );
  NOR2_X1 U9574 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7763) );
  AOI21_X1 U9575 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7763), .ZN(n10213) );
  NOR2_X1 U9576 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7764) );
  AOI21_X1 U9577 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7764), .ZN(n10216) );
  NOR2_X1 U9578 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7765) );
  AOI21_X1 U9579 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7765), .ZN(n10219) );
  NOR2_X1 U9580 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7766) );
  AOI21_X1 U9581 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7766), .ZN(n10222) );
  NOR2_X1 U9582 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7767) );
  AOI21_X1 U9583 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7767), .ZN(n10522) );
  NOR2_X1 U9584 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7768) );
  AOI21_X1 U9585 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7768), .ZN(n10528) );
  NOR2_X1 U9586 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7769) );
  AOI21_X1 U9587 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7769), .ZN(n10525) );
  NOR2_X1 U9588 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7770) );
  AOI21_X1 U9589 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n7770), .ZN(n10531) );
  NOR2_X1 U9590 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7771) );
  AOI21_X1 U9591 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7771), .ZN(n10519) );
  AND2_X1 U9592 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7772) );
  NOR2_X1 U9593 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7772), .ZN(n10191) );
  INV_X1 U9594 ( .A(n10191), .ZN(n10192) );
  INV_X1 U9595 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10194) );
  NAND3_X1 U9596 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U9597 ( .A1(n10194), .A2(n10193), .ZN(n10190) );
  NAND2_X1 U9598 ( .A1(n10192), .A2(n10190), .ZN(n10534) );
  NAND2_X1 U9599 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7773) );
  OAI21_X1 U9600 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7773), .ZN(n10533) );
  NOR2_X1 U9601 ( .A1(n10534), .A2(n10533), .ZN(n10532) );
  AOI21_X1 U9602 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10532), .ZN(n10537) );
  NAND2_X1 U9603 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7774) );
  OAI21_X1 U9604 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7774), .ZN(n10536) );
  NOR2_X1 U9605 ( .A1(n10537), .A2(n10536), .ZN(n10535) );
  AOI21_X1 U9606 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10535), .ZN(n10540) );
  NOR2_X1 U9607 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7775) );
  AOI21_X1 U9608 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7775), .ZN(n10539) );
  NAND2_X1 U9609 ( .A1(n10540), .A2(n10539), .ZN(n10538) );
  OAI21_X1 U9610 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10538), .ZN(n10518) );
  NAND2_X1 U9611 ( .A1(n10519), .A2(n10518), .ZN(n10517) );
  OAI21_X1 U9612 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10517), .ZN(n10530) );
  NAND2_X1 U9613 ( .A1(n10531), .A2(n10530), .ZN(n10529) );
  OAI21_X1 U9614 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10529), .ZN(n10524) );
  NAND2_X1 U9615 ( .A1(n10525), .A2(n10524), .ZN(n10523) );
  OAI21_X1 U9616 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10523), .ZN(n10527) );
  NAND2_X1 U9617 ( .A1(n10528), .A2(n10527), .ZN(n10526) );
  OAI21_X1 U9618 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10526), .ZN(n10521) );
  NAND2_X1 U9619 ( .A1(n10522), .A2(n10521), .ZN(n10520) );
  OAI21_X1 U9620 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10520), .ZN(n10221) );
  NAND2_X1 U9621 ( .A1(n10222), .A2(n10221), .ZN(n10220) );
  OAI21_X1 U9622 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10220), .ZN(n10218) );
  NAND2_X1 U9623 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  OAI21_X1 U9624 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10217), .ZN(n10215) );
  NAND2_X1 U9625 ( .A1(n10216), .A2(n10215), .ZN(n10214) );
  OAI21_X1 U9626 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10214), .ZN(n10212) );
  NAND2_X1 U9627 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  OAI21_X1 U9628 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10211), .ZN(n10209) );
  NAND2_X1 U9629 ( .A1(n10210), .A2(n10209), .ZN(n10208) );
  OAI21_X1 U9630 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10208), .ZN(n10206) );
  NAND2_X1 U9631 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  OAI21_X1 U9632 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10205), .ZN(n10203) );
  NAND2_X1 U9633 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  OAI21_X1 U9634 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10202), .ZN(n10200) );
  NAND2_X1 U9635 ( .A1(n10201), .A2(n10200), .ZN(n10199) );
  OAI21_X1 U9636 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10199), .ZN(n10197) );
  NOR2_X1 U9637 ( .A1(n10196), .A2(n10197), .ZN(n7776) );
  NAND2_X1 U9638 ( .A1(n10196), .A2(n10197), .ZN(n10195) );
  OAI21_X1 U9639 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7776), .A(n10195), .ZN(
        n7780) );
  NOR2_X1 U9640 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  XNOR2_X1 U9641 ( .A(n7780), .B(n7779), .ZN(ADD_1068_U4) );
  INV_X1 U9642 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7782) );
  MUX2_X1 U9643 ( .A(n7782), .B(n7781), .S(n10189), .Z(n7783) );
  OAI21_X1 U9644 ( .B1(n4608), .B2(n9135), .A(n7783), .ZN(P2_U3469) );
  INV_X1 U9645 ( .A(n7784), .ZN(n7789) );
  OAI21_X1 U9646 ( .B1(n7991), .B2(n10123), .A(n7785), .ZN(n7786) );
  NAND2_X1 U9647 ( .A1(n7786), .A2(n10141), .ZN(n7788) );
  AOI22_X1 U9648 ( .A1(n4615), .A2(n9109), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n10144), .ZN(n7787) );
  OAI211_X1 U9649 ( .C1(n7789), .C2(n10115), .A(n7788), .B(n7787), .ZN(
        P2_U3222) );
  AOI211_X1 U9650 ( .C1(n10071), .C2(n7792), .A(n7791), .B(n7790), .ZN(n7795)
         );
  AOI22_X1 U9651 ( .A1(n6861), .A2(n9325), .B1(P1_REG0_REG_8__SCAN_IN), .B2(
        n10072), .ZN(n7793) );
  OAI21_X1 U9652 ( .B1(n7795), .B2(n10072), .A(n7793), .ZN(P1_U3477) );
  AOI22_X1 U9653 ( .A1(n9940), .A2(n9325), .B1(P1_REG1_REG_8__SCAN_IN), .B2(
        n4655), .ZN(n7794) );
  OAI21_X1 U9654 ( .B1(n7795), .B2(n4655), .A(n7794), .ZN(P1_U3530) );
  INV_X1 U9655 ( .A(n7796), .ZN(n7799) );
  OAI222_X1 U9656 ( .A1(n9246), .A2(n10302), .B1(n9258), .B2(n7799), .C1(n7797), .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9657 ( .A1(n8378), .A2(n10288), .B1(n10029), .B2(n7799), .C1(
        P1_U3086), .C2(n7798), .ZN(P1_U3333) );
  XOR2_X1 U9658 ( .A(n8601), .B(n7800), .Z(n7925) );
  NAND2_X1 U9659 ( .A1(n7802), .A2(n7801), .ZN(n7803) );
  XNOR2_X1 U9660 ( .A(n7803), .B(n8601), .ZN(n7804) );
  OAI222_X1 U9661 ( .A1(n10127), .A2(n7869), .B1(n10125), .B2(n7805), .C1(
        n7804), .C2(n10132), .ZN(n7922) );
  AOI21_X1 U9662 ( .B1(n7925), .B2(n10162), .A(n7922), .ZN(n7807) );
  MUX2_X1 U9663 ( .A(n10370), .B(n7807), .S(n10178), .Z(n7806) );
  OAI21_X1 U9664 ( .B1(n7921), .B2(n9211), .A(n7806), .ZN(P2_U3417) );
  MUX2_X1 U9665 ( .A(n7808), .B(n7807), .S(n10189), .Z(n7809) );
  OAI21_X1 U9666 ( .B1(n7921), .B2(n9135), .A(n7809), .ZN(P2_U3468) );
  OAI222_X1 U9667 ( .A1(n9258), .A2(n7811), .B1(P2_U3151), .B2(n7810), .C1(
        n10313), .C2(n9246), .ZN(P2_U3274) );
  NAND2_X1 U9668 ( .A1(n8144), .A2(n8133), .ZN(n8246) );
  INV_X1 U9669 ( .A(n8246), .ZN(n7812) );
  XNOR2_X1 U9670 ( .A(n7813), .B(n7812), .ZN(n8030) );
  NAND2_X1 U9671 ( .A1(n7699), .A2(n8130), .ZN(n7814) );
  XOR2_X1 U9672 ( .A(n8246), .B(n7814), .Z(n7815) );
  NAND2_X1 U9673 ( .A1(n7815), .A2(n9878), .ZN(n7816) );
  AOI22_X1 U9674 ( .A1(n9490), .A2(n9457), .B1(n9426), .B2(n9488), .ZN(n8044)
         );
  OAI211_X1 U9675 ( .C1(n8030), .C2(n7817), .A(n7816), .B(n8044), .ZN(n8031)
         );
  NAND2_X1 U9676 ( .A1(n8031), .A2(n9850), .ZN(n7825) );
  INV_X1 U9677 ( .A(n7706), .ZN(n7820) );
  INV_X1 U9678 ( .A(n7818), .ZN(n7819) );
  AOI211_X1 U9679 ( .C1(n7821), .C2(n7820), .A(n9885), .B(n7819), .ZN(n8032)
         );
  AOI22_X1 U9680 ( .A1(n10063), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8046), .B2(
        n10052), .ZN(n7822) );
  OAI21_X1 U9681 ( .B1(n8052), .B2(n9891), .A(n7822), .ZN(n7823) );
  AOI21_X1 U9682 ( .B1(n8032), .B2(n10057), .A(n7823), .ZN(n7824) );
  OAI211_X1 U9683 ( .C1(n8030), .C2(n10053), .A(n7825), .B(n7824), .ZN(
        P1_U3282) );
  INV_X1 U9684 ( .A(n7826), .ZN(n7827) );
  AOI21_X1 U9685 ( .B1(n8591), .B2(n7828), .A(n7827), .ZN(n7849) );
  INV_X1 U9686 ( .A(n7849), .ZN(n7835) );
  XNOR2_X1 U9687 ( .A(n7829), .B(n8591), .ZN(n7830) );
  AOI222_X1 U9688 ( .A1(n9094), .A2(n7830), .B1(n8781), .B2(n6698), .C1(n8783), 
        .C2(n9090), .ZN(n7848) );
  MUX2_X1 U9689 ( .A(n7831), .B(n7848), .S(n10141), .Z(n7834) );
  INV_X1 U9690 ( .A(n7878), .ZN(n7832) );
  AOI22_X1 U9691 ( .A1(n7875), .A2(n9109), .B1(n9096), .B2(n7832), .ZN(n7833)
         );
  OAI211_X1 U9692 ( .C1(n7835), .C2(n10115), .A(n7834), .B(n7833), .ZN(
        P2_U3221) );
  INV_X1 U9693 ( .A(n7836), .ZN(n7837) );
  AOI211_X1 U9694 ( .C1(n10071), .C2(n7839), .A(n7838), .B(n7837), .ZN(n7842)
         );
  AOI22_X1 U9695 ( .A1(n7968), .A2(n6861), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n10072), .ZN(n7840) );
  OAI21_X1 U9696 ( .B1(n7842), .B2(n10072), .A(n7840), .ZN(P1_U3483) );
  AOI22_X1 U9697 ( .A1(n7968), .A2(n9940), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n4655), .ZN(n7841) );
  OAI21_X1 U9698 ( .B1(n7842), .B2(n4655), .A(n7841), .ZN(P1_U3532) );
  INV_X1 U9699 ( .A(n7843), .ZN(n7854) );
  OR2_X1 U9700 ( .A1(n7844), .A2(P2_U3151), .ZN(n8770) );
  INV_X1 U9701 ( .A(n8770), .ZN(n8764) );
  AOI21_X1 U9702 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9256), .A(n8764), .ZN(
        n7845) );
  OAI21_X1 U9703 ( .B1(n7854), .B2(n9258), .A(n7845), .ZN(P2_U3272) );
  MUX2_X1 U9704 ( .A(n10478), .B(n7848), .S(n10189), .Z(n7847) );
  AOI22_X1 U9705 ( .A1(n7849), .A2(n9155), .B1(n9154), .B2(n7875), .ZN(n7846)
         );
  NAND2_X1 U9706 ( .A1(n7847), .A2(n7846), .ZN(P2_U3471) );
  MUX2_X1 U9707 ( .A(n10400), .B(n7848), .S(n10178), .Z(n7851) );
  AOI22_X1 U9708 ( .A1(n7849), .A2(n9240), .B1(n6799), .B2(n7875), .ZN(n7850)
         );
  NAND2_X1 U9709 ( .A1(n7851), .A2(n7850), .ZN(P2_U3426) );
  OR2_X1 U9710 ( .A1(n7852), .A2(P1_U3086), .ZN(n8361) );
  NAND2_X1 U9711 ( .A1(n10024), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7853) );
  OAI211_X1 U9712 ( .C1(n7854), .C2(n10029), .A(n8361), .B(n7853), .ZN(
        P1_U3332) );
  OAI21_X1 U9713 ( .B1(n7958), .B2(n10066), .A(n7855), .ZN(n7857) );
  AOI211_X1 U9714 ( .C1(n10071), .C2(n7858), .A(n7857), .B(n7856), .ZN(n7861)
         );
  NAND2_X1 U9715 ( .A1(n10072), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7859) );
  OAI21_X1 U9716 ( .B1(n7861), .B2(n10072), .A(n7859), .ZN(P1_U3480) );
  NAND2_X1 U9717 ( .A1(n4655), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7860) );
  OAI21_X1 U9718 ( .B1(n7861), .B2(n4655), .A(n7860), .ZN(P1_U3531) );
  INV_X1 U9719 ( .A(n7875), .ZN(n7883) );
  XNOR2_X1 U9720 ( .A(n7870), .B(n8107), .ZN(n7988) );
  XOR2_X1 U9721 ( .A(n8107), .B(n7909), .Z(n7985) );
  NOR3_X1 U9722 ( .A1(n7909), .A2(n7869), .A3(n7868), .ZN(n7867) );
  INV_X1 U9723 ( .A(n7870), .ZN(n8590) );
  NOR3_X1 U9724 ( .A1(n4608), .A2(n7869), .A3(n8107), .ZN(n7871) );
  AOI211_X1 U9725 ( .C1(n8783), .C2(n8107), .A(n7871), .B(n7870), .ZN(n7872)
         );
  XNOR2_X1 U9726 ( .A(n7875), .B(n8107), .ZN(n8054) );
  XNOR2_X1 U9727 ( .A(n8054), .B(n8782), .ZN(n7876) );
  OAI211_X1 U9728 ( .C1(n7877), .C2(n7876), .A(n8056), .B(n8557), .ZN(n7882)
         );
  NAND2_X1 U9729 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8827) );
  OAI21_X1 U9730 ( .B1(n8541), .B2(n8111), .A(n8827), .ZN(n7880) );
  NOR2_X1 U9731 ( .A1(n8063), .A2(n7878), .ZN(n7879) );
  AOI211_X1 U9732 ( .C1(n8539), .C2(n8783), .A(n7880), .B(n7879), .ZN(n7881)
         );
  OAI211_X1 U9733 ( .C1(n7883), .C2(n8568), .A(n7882), .B(n7881), .ZN(P2_U3164) );
  XNOR2_X1 U9734 ( .A(n9614), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U9735 ( .A1(n7884), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9736 ( .A1(n7886), .A2(n7885), .ZN(n7888) );
  INV_X1 U9737 ( .A(n9616), .ZN(n7887) );
  AOI21_X1 U9738 ( .B1(n7889), .B2(n7888), .A(n7887), .ZN(n7901) );
  INV_X1 U9739 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U9740 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9382) );
  OAI21_X1 U9741 ( .B1(n9643), .B2(n7890), .A(n9382), .ZN(n7898) );
  INV_X1 U9742 ( .A(n7891), .ZN(n7892) );
  NOR2_X1 U9743 ( .A1(n7893), .A2(n7892), .ZN(n7895) );
  XNOR2_X1 U9744 ( .A(n9614), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7894) );
  NOR2_X1 U9745 ( .A1(n7895), .A2(n7894), .ZN(n9610) );
  AOI21_X1 U9746 ( .B1(n7895), .B2(n7894), .A(n9610), .ZN(n7896) );
  NOR2_X1 U9747 ( .A1(n7896), .A2(n9633), .ZN(n7897) );
  AOI211_X1 U9748 ( .C1(n9636), .C2(n9614), .A(n7898), .B(n7897), .ZN(n7899)
         );
  OAI21_X1 U9749 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(P1_U3260) );
  XNOR2_X1 U9750 ( .A(n7902), .B(n8784), .ZN(n7986) );
  XOR2_X1 U9751 ( .A(n7985), .B(n7986), .Z(n7911) );
  OAI21_X1 U9752 ( .B1(n8541), .B2(n7904), .A(n7903), .ZN(n7905) );
  AOI21_X1 U9753 ( .B1(n8539), .B2(n8785), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9754 ( .B1(n7907), .B2(n8063), .A(n7906), .ZN(n7908) );
  AOI21_X1 U9755 ( .B1(n7909), .B2(n8553), .A(n7908), .ZN(n7910) );
  OAI21_X1 U9756 ( .B1(n7911), .B2(n8555), .A(n7910), .ZN(P2_U3157) );
  INV_X1 U9757 ( .A(n8672), .ZN(n8604) );
  XNOR2_X1 U9758 ( .A(n7912), .B(n8604), .ZN(n7913) );
  AOI222_X1 U9759 ( .A1(n9094), .A2(n7913), .B1(n8780), .B2(n6698), .C1(n8782), 
        .C2(n9090), .ZN(n7935) );
  MUX2_X1 U9760 ( .A(n10381), .B(n7935), .S(n10189), .Z(n7916) );
  XNOR2_X1 U9761 ( .A(n7914), .B(n8672), .ZN(n7939) );
  AOI22_X1 U9762 ( .A1(n7939), .A2(n9155), .B1(n9154), .B2(n8065), .ZN(n7915)
         );
  NAND2_X1 U9763 ( .A1(n7916), .A2(n7915), .ZN(P2_U3472) );
  MUX2_X1 U9764 ( .A(n7917), .B(n7935), .S(n10178), .Z(n7919) );
  AOI22_X1 U9765 ( .A1(n7939), .A2(n9240), .B1(n6799), .B2(n8065), .ZN(n7918)
         );
  NAND2_X1 U9766 ( .A1(n7919), .A2(n7918), .ZN(P2_U3429) );
  OAI22_X1 U9767 ( .A1(n7921), .A2(n10111), .B1(n7920), .B2(n10123), .ZN(n7924) );
  MUX2_X1 U9768 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7922), .S(n10141), .Z(n7923)
         );
  AOI211_X1 U9769 ( .C1(n7925), .C2(n8992), .A(n7924), .B(n7923), .ZN(n7926)
         );
  INV_X1 U9770 ( .A(n7926), .ZN(P2_U3224) );
  INV_X1 U9771 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U9772 ( .A1(n7927), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7930) );
  INV_X1 U9773 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10498) );
  OR2_X1 U9774 ( .A1(n7928), .A2(n10498), .ZN(n7929) );
  OAI211_X1 U9775 ( .C1(n4612), .C2(n8944), .A(n7930), .B(n7929), .ZN(n7931)
         );
  INV_X1 U9776 ( .A(n7931), .ZN(n7932) );
  INV_X1 U9777 ( .A(n8941), .ZN(n8750) );
  NAND2_X1 U9778 ( .A1(n8750), .A2(P2_U3893), .ZN(n7934) );
  OAI21_X1 U9779 ( .B1(P2_U3893), .B2(n6848), .A(n7934), .ZN(P2_U3522) );
  INV_X1 U9780 ( .A(n10122), .ZN(n7937) );
  INV_X1 U9781 ( .A(n7935), .ZN(n7936) );
  AOI21_X1 U9782 ( .B1(n7937), .B2(n8065), .A(n7936), .ZN(n7941) );
  OAI22_X1 U9783 ( .A1(n10141), .A2(n4923), .B1(n8062), .B2(n10123), .ZN(n7938) );
  AOI21_X1 U9784 ( .B1(n7939), .B2(n8992), .A(n7938), .ZN(n7940) );
  OAI21_X1 U9785 ( .B1(n7941), .B2(n10144), .A(n7940), .ZN(P2_U3220) );
  NAND2_X1 U9786 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  XNOR2_X1 U9787 ( .A(n7944), .B(n7945), .ZN(n9321) );
  NOR2_X1 U9788 ( .A1(n9321), .A2(n9320), .ZN(n9319) );
  AOI21_X1 U9789 ( .B1(n7945), .B2(n7944), .A(n9319), .ZN(n7948) );
  OAI211_X1 U9790 ( .C1(n7948), .C2(n7947), .A(n9434), .B(n7946), .ZN(n7957)
         );
  INV_X1 U9791 ( .A(n7949), .ZN(n7954) );
  OAI21_X1 U9792 ( .B1(n7951), .B2(n7950), .A(n9460), .ZN(n7953) );
  OAI211_X1 U9793 ( .C1(n9462), .C2(n7954), .A(n7953), .B(n7952), .ZN(n7955)
         );
  INV_X1 U9794 ( .A(n7955), .ZN(n7956) );
  OAI211_X1 U9795 ( .C1(n7958), .C2(n9412), .A(n7957), .B(n7956), .ZN(P1_U3231) );
  INV_X1 U9796 ( .A(n7959), .ZN(n8040) );
  AOI21_X1 U9797 ( .B1(n7961), .B2(n8037), .A(n7960), .ZN(n7962) );
  AOI21_X1 U9798 ( .B1(n8040), .B2(n8037), .A(n7962), .ZN(n7970) );
  NAND2_X1 U9799 ( .A1(n9460), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U9800 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7964) );
  OAI211_X1 U9801 ( .C1(n9462), .C2(n7966), .A(n7965), .B(n7964), .ZN(n7967)
         );
  AOI21_X1 U9802 ( .B1(n7968), .B2(n9465), .A(n7967), .ZN(n7969) );
  OAI21_X1 U9803 ( .B1(n7970), .B2(n9467), .A(n7969), .ZN(P1_U3217) );
  OAI211_X1 U9804 ( .C1(n7972), .C2(n8247), .A(n7971), .B(n9878), .ZN(n7976)
         );
  OR2_X1 U9805 ( .A1(n8013), .A2(n9455), .ZN(n7974) );
  NAND2_X1 U9806 ( .A1(n9489), .A2(n9457), .ZN(n7973) );
  NAND2_X1 U9807 ( .A1(n7974), .A2(n7973), .ZN(n9349) );
  INV_X1 U9808 ( .A(n9349), .ZN(n7975) );
  AND2_X1 U9809 ( .A1(n7976), .A2(n7975), .ZN(n8069) );
  INV_X1 U9810 ( .A(n7977), .ZN(n9346) );
  OAI22_X1 U9811 ( .A1(n9850), .A2(n7978), .B1(n9346), .B2(n9829), .ZN(n7981)
         );
  AOI21_X1 U9812 ( .B1(n7818), .B2(n9338), .A(n9885), .ZN(n7979) );
  NAND2_X1 U9813 ( .A1(n7979), .A2(n8081), .ZN(n8068) );
  NOR2_X1 U9814 ( .A1(n8068), .A2(n9814), .ZN(n7980) );
  AOI211_X1 U9815 ( .C1(n10054), .C2(n9338), .A(n7981), .B(n7980), .ZN(n7984)
         );
  XNOR2_X1 U9816 ( .A(n7982), .B(n8247), .ZN(n8070) );
  OR2_X1 U9817 ( .A1(n8070), .A2(n9852), .ZN(n7983) );
  OAI211_X1 U9818 ( .C1(n8069), .C2(n10063), .A(n7984), .B(n7983), .ZN(
        P1_U3281) );
  OAI22_X1 U9819 ( .A1(n7986), .A2(n7985), .B1(n8784), .B2(n7902), .ZN(n7987)
         );
  XOR2_X1 U9820 ( .A(n7988), .B(n7987), .Z(n7995) );
  NAND2_X1 U9821 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8813) );
  OAI21_X1 U9822 ( .B1(n8541), .B2(n8053), .A(n8813), .ZN(n7989) );
  AOI21_X1 U9823 ( .B1(n8539), .B2(n8784), .A(n7989), .ZN(n7990) );
  OAI21_X1 U9824 ( .B1(n7991), .B2(n8063), .A(n7990), .ZN(n7992) );
  AOI21_X1 U9825 ( .B1(n4615), .B2(n8553), .A(n7992), .ZN(n7994) );
  OAI21_X1 U9826 ( .B1(n7995), .B2(n8555), .A(n7994), .ZN(P2_U3176) );
  INV_X1 U9827 ( .A(n7996), .ZN(n8001) );
  OAI222_X1 U9828 ( .A1(n9258), .A2(n8001), .B1(P2_U3151), .B2(n7998), .C1(
        n7997), .C2(n9246), .ZN(P2_U3271) );
  INV_X1 U9829 ( .A(n7999), .ZN(n8002) );
  OAI222_X1 U9830 ( .A1(P1_U3086), .A2(n8002), .B1(n10029), .B2(n8001), .C1(
        n8000), .C2(n8378), .ZN(P1_U3331) );
  INV_X1 U9831 ( .A(n9239), .ZN(n8679) );
  NOR2_X1 U9832 ( .A1(n8679), .A2(n10122), .ZN(n8005) );
  XNOR2_X1 U9833 ( .A(n8003), .B(n8674), .ZN(n8004) );
  OAI222_X1 U9834 ( .A1(n10127), .A2(n8489), .B1(n10125), .B2(n8111), .C1(
        n10132), .C2(n8004), .ZN(n9152) );
  AOI211_X1 U9835 ( .C1(n9096), .C2(n8108), .A(n8005), .B(n9152), .ZN(n8008)
         );
  XNOR2_X1 U9836 ( .A(n8006), .B(n8674), .ZN(n9241) );
  AOI22_X1 U9837 ( .A1(n9241), .A2(n8992), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10144), .ZN(n8007) );
  OAI21_X1 U9838 ( .B1(n8008), .B2(n10144), .A(n8007), .ZN(P2_U3219) );
  NAND2_X1 U9839 ( .A1(n8009), .A2(n8156), .ZN(n8012) );
  INV_X1 U9840 ( .A(n8010), .ZN(n8011) );
  AOI211_X1 U9841 ( .C1(n8251), .C2(n8012), .A(n9858), .B(n8011), .ZN(n8016)
         );
  OR2_X1 U9842 ( .A1(n8013), .A2(n9369), .ZN(n8015) );
  NAND2_X1 U9843 ( .A1(n9485), .A2(n9426), .ZN(n8014) );
  NAND2_X1 U9844 ( .A1(n8015), .A2(n8014), .ZN(n9284) );
  NOR2_X1 U9845 ( .A1(n8016), .A2(n9284), .ZN(n9966) );
  INV_X1 U9846 ( .A(n8080), .ZN(n8019) );
  INV_X1 U9847 ( .A(n8017), .ZN(n8018) );
  AOI211_X1 U9848 ( .C1(n9963), .C2(n8019), .A(n9885), .B(n8018), .ZN(n9962)
         );
  AOI22_X1 U9849 ( .A1(n10063), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9283), .B2(
        n10052), .ZN(n8020) );
  OAI21_X1 U9850 ( .B1(n8021), .B2(n9891), .A(n8020), .ZN(n8025) );
  INV_X1 U9851 ( .A(n8251), .ZN(n8023) );
  XNOR2_X1 U9852 ( .A(n8022), .B(n8023), .ZN(n9967) );
  NOR2_X1 U9853 ( .A1(n9967), .A2(n9852), .ZN(n8024) );
  AOI211_X1 U9854 ( .C1(n9962), .C2(n10057), .A(n8025), .B(n8024), .ZN(n8026)
         );
  OAI21_X1 U9855 ( .B1(n9966), .B2(n10063), .A(n8026), .ZN(P1_U3279) );
  INV_X1 U9856 ( .A(n8027), .ZN(n8089) );
  OAI222_X1 U9857 ( .A1(n9258), .A2(n8089), .B1(P2_U3151), .B2(n8029), .C1(
        n8028), .C2(n9246), .ZN(P2_U3270) );
  INV_X1 U9858 ( .A(n8030), .ZN(n8033) );
  AOI211_X1 U9859 ( .C1(n8034), .C2(n8033), .A(n8032), .B(n8031), .ZN(n8049)
         );
  MUX2_X1 U9860 ( .A(n8035), .B(n8049), .S(n10077), .Z(n8036) );
  OAI21_X1 U9861 ( .B1(n8052), .B2(n9961), .A(n8036), .ZN(P1_U3533) );
  INV_X1 U9862 ( .A(n8037), .ZN(n8039) );
  NOR3_X1 U9863 ( .A1(n8040), .A2(n8039), .A3(n8038), .ZN(n8042) );
  INV_X1 U9864 ( .A(n8041), .ZN(n9342) );
  OAI21_X1 U9865 ( .B1(n8042), .B2(n9342), .A(n9434), .ZN(n8048) );
  OAI21_X1 U9866 ( .B1(n9444), .B2(n8044), .A(n8043), .ZN(n8045) );
  AOI21_X1 U9867 ( .B1(n8046), .B2(n9442), .A(n8045), .ZN(n8047) );
  OAI211_X1 U9868 ( .C1(n8052), .C2(n9412), .A(n8048), .B(n8047), .ZN(P1_U3236) );
  INV_X1 U9869 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8050) );
  MUX2_X1 U9870 ( .A(n8050), .B(n8049), .S(n10074), .Z(n8051) );
  OAI21_X1 U9871 ( .B1(n8052), .B2(n10017), .A(n8051), .ZN(P1_U3486) );
  XNOR2_X1 U9872 ( .A(n8065), .B(n8107), .ZN(n8104) );
  XNOR2_X1 U9873 ( .A(n8104), .B(n8111), .ZN(n8059) );
  OR2_X1 U9874 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  INV_X1 U9875 ( .A(n8106), .ZN(n8057) );
  AOI21_X1 U9876 ( .B1(n8059), .B2(n8058), .A(n8057), .ZN(n8067) );
  AOI22_X1 U9877 ( .A1(n8561), .A2(n8780), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8061) );
  NAND2_X1 U9878 ( .A1(n8539), .A2(n8782), .ZN(n8060) );
  OAI211_X1 U9879 ( .C1(n8063), .C2(n8062), .A(n8061), .B(n8060), .ZN(n8064)
         );
  AOI21_X1 U9880 ( .B1(n8065), .B2(n8553), .A(n8064), .ZN(n8066) );
  OAI21_X1 U9881 ( .B1(n8067), .B2(n8555), .A(n8066), .ZN(P2_U3174) );
  OAI211_X1 U9882 ( .C1(n9968), .C2(n8070), .A(n8069), .B(n8068), .ZN(n8073)
         );
  MUX2_X1 U9883 ( .A(n8073), .B(P1_REG1_REG_12__SCAN_IN), .S(n4655), .Z(n8071)
         );
  AOI21_X1 U9884 ( .B1(n9940), .B2(n9338), .A(n8071), .ZN(n8072) );
  INV_X1 U9885 ( .A(n8072), .ZN(P1_U3534) );
  MUX2_X1 U9886 ( .A(n8073), .B(P1_REG0_REG_12__SCAN_IN), .S(n10072), .Z(n8074) );
  AOI21_X1 U9887 ( .B1(n6861), .B2(n9338), .A(n8074), .ZN(n8075) );
  INV_X1 U9888 ( .A(n8075), .ZN(P1_U3489) );
  XNOR2_X1 U9889 ( .A(n8076), .B(n8249), .ZN(n8077) );
  AOI22_X1 U9890 ( .A1(n9426), .A2(n9486), .B1(n9488), .B2(n9457), .ZN(n9407)
         );
  OAI21_X1 U9891 ( .B1(n8077), .B2(n9858), .A(n9407), .ZN(n8091) );
  INV_X1 U9892 ( .A(n8091), .ZN(n8087) );
  OAI21_X1 U9893 ( .B1(n8079), .B2(n5466), .A(n8078), .ZN(n8093) );
  AOI211_X1 U9894 ( .C1(n8082), .C2(n8081), .A(n9885), .B(n8080), .ZN(n8092)
         );
  NAND2_X1 U9895 ( .A1(n8092), .A2(n10057), .ZN(n8084) );
  AOI22_X1 U9896 ( .A1(n10063), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9409), .B2(
        n10052), .ZN(n8083) );
  OAI211_X1 U9897 ( .C1(n5135), .C2(n9891), .A(n8084), .B(n8083), .ZN(n8085)
         );
  AOI21_X1 U9898 ( .B1(n10049), .B2(n8093), .A(n8085), .ZN(n8086) );
  OAI21_X1 U9899 ( .B1(n10063), .B2(n8087), .A(n8086), .ZN(P1_U3280) );
  OAI222_X1 U9900 ( .A1(P1_U3086), .A2(n8090), .B1(n10029), .B2(n8089), .C1(
        n8088), .C2(n8378), .ZN(P1_U3330) );
  INV_X1 U9901 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8094) );
  AOI211_X1 U9902 ( .C1(n10071), .C2(n8093), .A(n8092), .B(n8091), .ZN(n8096)
         );
  MUX2_X1 U9903 ( .A(n8094), .B(n8096), .S(n10074), .Z(n8095) );
  OAI21_X1 U9904 ( .B1(n5135), .B2(n10017), .A(n8095), .ZN(P1_U3492) );
  MUX2_X1 U9905 ( .A(n8097), .B(n8096), .S(n10077), .Z(n8098) );
  OAI21_X1 U9906 ( .B1(n5135), .B2(n9961), .A(n8098), .ZN(P1_U3535) );
  INV_X1 U9907 ( .A(n8099), .ZN(n8102) );
  OAI222_X1 U9908 ( .A1(n9258), .A2(n8102), .B1(P2_U3151), .B2(n8100), .C1(
        n10429), .C2(n9246), .ZN(P2_U3269) );
  OAI222_X1 U9909 ( .A1(P1_U3086), .A2(n8103), .B1(n10029), .B2(n8102), .C1(
        n8101), .C2(n8378), .ZN(P1_U3329) );
  XNOR2_X1 U9910 ( .A(n9239), .B(n4460), .ZN(n8381) );
  XNOR2_X1 U9911 ( .A(n8381), .B(n8780), .ZN(n8383) );
  XOR2_X1 U9912 ( .A(n8384), .B(n8383), .Z(n8114) );
  NAND2_X1 U9913 ( .A1(n8565), .A2(n8108), .ZN(n8110) );
  AOI22_X1 U9914 ( .A1(n8561), .A2(n9091), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8109) );
  OAI211_X1 U9915 ( .C1(n8111), .C2(n8563), .A(n8110), .B(n8109), .ZN(n8112)
         );
  AOI21_X1 U9916 ( .B1(n9239), .B2(n8553), .A(n8112), .ZN(n8113) );
  OAI21_X1 U9917 ( .B1(n8114), .B2(n8555), .A(n8113), .ZN(P2_U3155) );
  AOI211_X1 U9918 ( .C1(n8225), .C2(n5780), .A(n8358), .B(n8296), .ZN(n8355)
         );
  INV_X1 U9919 ( .A(n9650), .ZN(n8212) );
  INV_X1 U9920 ( .A(n8290), .ZN(n8115) );
  INV_X1 U9921 ( .A(n8169), .ZN(n8117) );
  OAI21_X1 U9922 ( .B1(n8117), .B2(n8116), .A(n8168), .ZN(n8264) );
  INV_X1 U9923 ( .A(n8264), .ZN(n8120) );
  INV_X1 U9924 ( .A(n8118), .ZN(n8119) );
  NOR3_X1 U9925 ( .A1(n8120), .A2(n8119), .A3(n8297), .ZN(n8173) );
  OAI21_X1 U9926 ( .B1(n7739), .B2(n4797), .A(n8122), .ZN(n8124) );
  NAND2_X1 U9927 ( .A1(n8124), .A2(n8123), .ZN(n8128) );
  INV_X1 U9928 ( .A(n8129), .ZN(n8125) );
  AND2_X1 U9929 ( .A1(n8144), .A2(n8311), .ZN(n8131) );
  NAND2_X1 U9930 ( .A1(n9338), .A2(n8132), .ZN(n8318) );
  INV_X1 U9931 ( .A(n8318), .ZN(n8135) );
  INV_X1 U9932 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9933 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  NAND2_X1 U9934 ( .A1(n8138), .A2(n8145), .ZN(n8139) );
  NAND2_X1 U9935 ( .A1(n8141), .A2(n8140), .ZN(n8143) );
  INV_X1 U9936 ( .A(n8314), .ZN(n8142) );
  AOI21_X1 U9937 ( .B1(n8143), .B2(n8311), .A(n8142), .ZN(n8146) );
  NAND2_X1 U9938 ( .A1(n8145), .A2(n8144), .ZN(n8313) );
  OAI21_X1 U9939 ( .B1(n8146), .B2(n8313), .A(n8318), .ZN(n8147) );
  NAND2_X1 U9940 ( .A1(n8158), .A2(n8153), .ZN(n8150) );
  NAND4_X1 U9941 ( .A1(n8321), .A2(n8297), .A3(n9874), .A4(n8320), .ZN(n8148)
         );
  AOI21_X1 U9942 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8151) );
  INV_X1 U9943 ( .A(n8151), .ZN(n8162) );
  INV_X1 U9944 ( .A(n8154), .ZN(n8152) );
  INV_X1 U9945 ( .A(n9886), .ZN(n10018) );
  AOI22_X1 U9946 ( .A1(n8321), .A2(n8152), .B1(n10018), .B2(n8123), .ZN(n8161)
         );
  AOI21_X1 U9947 ( .B1(n8326), .B2(n9485), .A(n8297), .ZN(n8160) );
  NAND2_X1 U9948 ( .A1(n9874), .A2(n8153), .ZN(n8317) );
  OAI211_X1 U9949 ( .C1(n8317), .C2(n8156), .A(n8155), .B(n8154), .ZN(n8322)
         );
  NOR3_X1 U9950 ( .A1(n5807), .A2(n8322), .A3(n8297), .ZN(n8157) );
  MUX2_X1 U9951 ( .A(n8321), .B(n8326), .S(n8297), .Z(n8159) );
  NAND2_X1 U9952 ( .A1(n8177), .A2(n8163), .ZN(n8324) );
  OAI211_X1 U9953 ( .C1(n8174), .C2(n8324), .A(n8330), .B(n8176), .ZN(n8164)
         );
  NAND3_X1 U9954 ( .A1(n8164), .A2(n9771), .A3(n8178), .ZN(n8166) );
  INV_X1 U9955 ( .A(n8165), .ZN(n8228) );
  NAND3_X1 U9956 ( .A1(n8166), .A2(n8228), .A3(n8183), .ZN(n8172) );
  NAND2_X1 U9957 ( .A1(n8168), .A2(n8167), .ZN(n8267) );
  AND2_X1 U9958 ( .A1(n8267), .A2(n8169), .ZN(n8182) );
  OAI22_X1 U9959 ( .A1(n8264), .A2(n8297), .B1(n8227), .B2(n9749), .ZN(n8170)
         );
  AOI21_X1 U9960 ( .B1(n8182), .B2(n8297), .A(n8170), .ZN(n8171) );
  AOI211_X1 U9961 ( .C1(n8173), .C2(n8172), .A(n9729), .B(n8171), .ZN(n8190)
         );
  INV_X1 U9962 ( .A(n8174), .ZN(n8179) );
  AND2_X1 U9963 ( .A1(n8176), .A2(n8175), .ZN(n8327) );
  NAND2_X1 U9964 ( .A1(n8178), .A2(n8177), .ZN(n8331) );
  AOI21_X1 U9965 ( .B1(n8179), .B2(n8327), .A(n8331), .ZN(n8181) );
  NAND2_X1 U9966 ( .A1(n8228), .A2(n8330), .ZN(n8180) );
  OAI21_X1 U9967 ( .B1(n8181), .B2(n8180), .A(n8335), .ZN(n8185) );
  INV_X1 U9968 ( .A(n8182), .ZN(n8184) );
  NAND4_X1 U9969 ( .A1(n8185), .A2(n8297), .A3(n8184), .A4(n8183), .ZN(n8189)
         );
  INV_X1 U9970 ( .A(n8263), .ZN(n8187) );
  INV_X1 U9971 ( .A(n8270), .ZN(n8186) );
  MUX2_X1 U9972 ( .A(n8187), .B(n8186), .S(n8297), .Z(n8188) );
  NAND2_X1 U9973 ( .A1(n8192), .A2(n8191), .ZN(n8275) );
  NAND3_X1 U9974 ( .A1(n8272), .A2(n8123), .A3(n8273), .ZN(n8193) );
  INV_X1 U9975 ( .A(n8275), .ZN(n8197) );
  OAI21_X1 U9976 ( .B1(n8297), .B2(n8261), .A(n8262), .ZN(n8196) );
  NAND3_X1 U9977 ( .A1(n9706), .A2(n9359), .A3(n8297), .ZN(n8194) );
  NAND2_X1 U9978 ( .A1(n8280), .A2(n8194), .ZN(n8195) );
  NAND3_X1 U9979 ( .A1(n8261), .A2(n8297), .A3(n9698), .ZN(n8201) );
  AOI21_X1 U9980 ( .B1(n8202), .B2(n8273), .A(n8201), .ZN(n8203) );
  OAI21_X1 U9981 ( .B1(n8275), .B2(n8262), .A(n8280), .ZN(n8204) );
  NAND2_X1 U9982 ( .A1(n8290), .A2(n9470), .ZN(n8207) );
  INV_X1 U9983 ( .A(n9470), .ZN(n8226) );
  NOR3_X1 U9984 ( .A1(n9650), .A2(n9972), .A3(n8226), .ZN(n8209) );
  OAI21_X1 U9985 ( .B1(n9650), .B2(n8226), .A(n8211), .ZN(n8214) );
  INV_X1 U9986 ( .A(n8281), .ZN(n8213) );
  AND2_X1 U9987 ( .A1(n9972), .A2(n9470), .ZN(n8287) );
  NOR2_X1 U9988 ( .A1(n8215), .A2(n8123), .ZN(n8219) );
  AOI21_X1 U9989 ( .B1(n8216), .B2(n9654), .A(n8343), .ZN(n8217) );
  OAI21_X1 U9990 ( .B1(n8291), .B2(n7428), .A(n8221), .ZN(n8354) );
  INV_X1 U9991 ( .A(n8221), .ZN(n8224) );
  NAND2_X1 U9992 ( .A1(n5780), .A2(n8300), .ZN(n8298) );
  INV_X1 U9993 ( .A(n8298), .ZN(n8222) );
  NAND3_X1 U9994 ( .A1(n8224), .A2(n8223), .A3(n8222), .ZN(n8353) );
  INV_X1 U9995 ( .A(n8287), .ZN(n8340) );
  NAND2_X1 U9996 ( .A1(n9654), .A2(n8226), .ZN(n8286) );
  INV_X1 U9997 ( .A(n9686), .ZN(n8259) );
  INV_X1 U9998 ( .A(n9863), .ZN(n9855) );
  NOR2_X1 U9999 ( .A1(n8230), .A2(n8229), .ZN(n8233) );
  NAND4_X1 U10000 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8303), .ZN(n8238)
         );
  NAND2_X1 U10001 ( .A1(n8235), .A2(n8234), .ZN(n8237) );
  INV_X1 U10002 ( .A(n8239), .ZN(n8240) );
  NOR2_X1 U10003 ( .A1(n8241), .A2(n8240), .ZN(n8244) );
  NAND3_X1 U10004 ( .A1(n8249), .A2(n8248), .A3(n8247), .ZN(n8250) );
  OR3_X1 U10005 ( .A1(n9884), .A2(n8251), .A3(n8250), .ZN(n8252) );
  NOR2_X1 U10006 ( .A1(n9820), .A2(n8253), .ZN(n8254) );
  XNOR2_X1 U10007 ( .A(n9781), .B(n8255), .ZN(n9776) );
  NAND3_X1 U10008 ( .A1(n9717), .A2(n5817), .A3(n8256), .ZN(n8257) );
  NOR3_X1 U10009 ( .A1(n8295), .A2(n5780), .A3(n8260), .ZN(n8351) );
  AND2_X1 U10010 ( .A1(n8262), .A2(n8261), .ZN(n8336) );
  NAND2_X1 U10011 ( .A1(n8264), .A2(n8263), .ZN(n8266) );
  INV_X1 U10012 ( .A(n8267), .ZN(n8269) );
  NAND3_X1 U10013 ( .A1(n8270), .A2(n8269), .A3(n8268), .ZN(n8271) );
  NAND2_X1 U10014 ( .A1(n8334), .A2(n8271), .ZN(n8274) );
  NAND3_X1 U10015 ( .A1(n8274), .A2(n8273), .A3(n8272), .ZN(n8276) );
  AOI21_X1 U10016 ( .B1(n8336), .B2(n8276), .A(n8275), .ZN(n8339) );
  INV_X1 U10017 ( .A(n8339), .ZN(n8284) );
  INV_X1 U10018 ( .A(n8336), .ZN(n8279) );
  INV_X1 U10019 ( .A(n8334), .ZN(n8277) );
  NOR3_X1 U10020 ( .A1(n8279), .A2(n8278), .A3(n8277), .ZN(n8283) );
  NAND2_X1 U10021 ( .A1(n8281), .A2(n8280), .ZN(n8337) );
  INV_X1 U10022 ( .A(n8337), .ZN(n8282) );
  OAI21_X1 U10023 ( .B1(n8284), .B2(n8283), .A(n8282), .ZN(n8289) );
  NAND2_X1 U10024 ( .A1(n8286), .A2(n8285), .ZN(n8341) );
  INV_X1 U10025 ( .A(n8341), .ZN(n8288) );
  AOI22_X1 U10026 ( .A1(n8289), .A2(n8288), .B1(n8287), .B2(n8290), .ZN(n8294)
         );
  OAI21_X1 U10027 ( .B1(n9972), .B2(n8290), .A(n8208), .ZN(n8293) );
  OAI211_X1 U10028 ( .C1(n8294), .C2(n8293), .A(n8292), .B(n8291), .ZN(n8350)
         );
  INV_X1 U10029 ( .A(n8295), .ZN(n8299) );
  OAI22_X1 U10030 ( .A1(n8299), .A2(n8298), .B1(n8297), .B2(n8296), .ZN(n8349)
         );
  INV_X1 U10031 ( .A(n8356), .ZN(n8347) );
  NOR2_X1 U10032 ( .A1(n7428), .A2(n8300), .ZN(n8346) );
  OAI21_X1 U10033 ( .B1(n6124), .B2(n10055), .A(n8301), .ZN(n8302) );
  AOI211_X1 U10034 ( .C1(n8376), .C2(n9498), .A(n8303), .B(n8302), .ZN(n8306)
         );
  NAND4_X1 U10035 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n5793), .ZN(n8309)
         );
  INV_X1 U10036 ( .A(n8307), .ZN(n8308) );
  NAND2_X1 U10037 ( .A1(n8309), .A2(n8308), .ZN(n8312) );
  OAI211_X1 U10038 ( .C1(n7615), .C2(n8312), .A(n8311), .B(n8310), .ZN(n8315)
         );
  AOI21_X1 U10039 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8316) );
  INV_X1 U10040 ( .A(n8316), .ZN(n8319) );
  AOI21_X1 U10041 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(n8323) );
  OAI211_X1 U10042 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8320), .ZN(n8325)
         );
  AOI21_X1 U10043 ( .B1(n8326), .B2(n8325), .A(n8324), .ZN(n8329) );
  INV_X1 U10044 ( .A(n8327), .ZN(n8328) );
  NOR2_X1 U10045 ( .A1(n8329), .A2(n8328), .ZN(n8332) );
  OAI21_X1 U10046 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n8333) );
  NAND4_X1 U10047 ( .A1(n8336), .A2(n8335), .A3(n8334), .A4(n8333), .ZN(n8338)
         );
  OAI21_X1 U10048 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8344) );
  AOI21_X1 U10049 ( .B1(n8344), .B2(n8208), .A(n8343), .ZN(n8345) );
  MUX2_X1 U10050 ( .A(n8347), .B(n8346), .S(n8345), .Z(n8348) );
  AOI22_X1 U10051 ( .A1(n8355), .A2(n8354), .B1(n8353), .B2(n8352), .ZN(n8362)
         );
  NOR4_X1 U10052 ( .A1(n8357), .A2(n8356), .A3(n10031), .A4(n9369), .ZN(n8360)
         );
  OAI21_X1 U10053 ( .B1(n8361), .B2(n8358), .A(P1_B_REG_SCAN_IN), .ZN(n8359)
         );
  INV_X1 U10054 ( .A(n8363), .ZN(n8366) );
  OAI222_X1 U10055 ( .A1(n9258), .A2(n8366), .B1(n8365), .B2(P2_U3151), .C1(
        n8364), .C2(n9246), .ZN(P2_U3275) );
  INV_X1 U10056 ( .A(n8367), .ZN(n10028) );
  OAI222_X1 U10057 ( .A1(n9258), .A2(n10028), .B1(n8369), .B2(P2_U3151), .C1(
        n8368), .C2(n9246), .ZN(P2_U3266) );
  XNOR2_X1 U10058 ( .A(n8371), .B(n8370), .ZN(n8372) );
  NAND2_X1 U10059 ( .A1(n8372), .A2(n9434), .ZN(n8375) );
  AOI22_X1 U10060 ( .A1(n9460), .A2(n8373), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8440), .ZN(n8374) );
  OAI211_X1 U10061 ( .C1(n8376), .C2(n9412), .A(n8375), .B(n8374), .ZN(
        P1_U3237) );
  INV_X1 U10062 ( .A(n8575), .ZN(n8435) );
  OAI222_X1 U10063 ( .A1(n8378), .A2(n8377), .B1(n10029), .B2(n8435), .C1(
        P1_U3086), .C2(n4449), .ZN(P1_U3325) );
  INV_X1 U10064 ( .A(n8379), .ZN(n9254) );
  OAI222_X1 U10065 ( .A1(n8378), .A2(n8380), .B1(n10029), .B2(n9254), .C1(
        n5824), .C2(P1_U3086), .ZN(P1_U3327) );
  XNOR2_X1 U10066 ( .A(n9149), .B(n4460), .ZN(n8385) );
  XNOR2_X1 U10067 ( .A(n8385), .B(n9091), .ZN(n8559) );
  INV_X1 U10068 ( .A(n8385), .ZN(n8386) );
  NAND2_X1 U10069 ( .A1(n8386), .A2(n9091), .ZN(n8387) );
  XNOR2_X1 U10070 ( .A(n9231), .B(n8107), .ZN(n8388) );
  XNOR2_X1 U10071 ( .A(n8388), .B(n9081), .ZN(n8486) );
  INV_X1 U10072 ( .A(n8388), .ZN(n8389) );
  XNOR2_X1 U10073 ( .A(n9225), .B(n8107), .ZN(n8393) );
  XOR2_X1 U10074 ( .A(n9092), .B(n8393), .Z(n8496) );
  INV_X1 U10075 ( .A(n8496), .ZN(n8390) );
  NAND2_X1 U10076 ( .A1(n8391), .A2(n8390), .ZN(n8494) );
  NAND2_X1 U10077 ( .A1(n8393), .A2(n8392), .ZN(n8532) );
  NAND2_X1 U10078 ( .A1(n8494), .A2(n8532), .ZN(n8394) );
  XNOR2_X1 U10079 ( .A(n9219), .B(n8107), .ZN(n8395) );
  XNOR2_X1 U10080 ( .A(n8395), .B(n9082), .ZN(n8533) );
  NAND2_X1 U10081 ( .A1(n8395), .A2(n8466), .ZN(n8396) );
  XNOR2_X1 U10082 ( .A(n9060), .B(n4460), .ZN(n8397) );
  XOR2_X1 U10083 ( .A(n9067), .B(n8397), .Z(n8460) );
  INV_X1 U10084 ( .A(n8397), .ZN(n8398) );
  NAND2_X1 U10085 ( .A1(n8398), .A2(n9067), .ZN(n8399) );
  XNOR2_X1 U10086 ( .A(n6610), .B(n4460), .ZN(n8402) );
  XOR2_X1 U10087 ( .A(n9054), .B(n8402), .Z(n8516) );
  INV_X1 U10088 ( .A(n8516), .ZN(n8400) );
  NAND2_X1 U10089 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  XNOR2_X1 U10090 ( .A(n8472), .B(n4460), .ZN(n8404) );
  XNOR2_X1 U10091 ( .A(n8404), .B(n8527), .ZN(n8471) );
  INV_X1 U10092 ( .A(n8404), .ZN(n8405) );
  NAND2_X1 U10093 ( .A1(n8405), .A2(n8527), .ZN(n8406) );
  XNOR2_X1 U10094 ( .A(n9196), .B(n8107), .ZN(n8410) );
  XOR2_X1 U10095 ( .A(n9032), .B(n8410), .Z(n8522) );
  INV_X1 U10096 ( .A(n8522), .ZN(n8408) );
  INV_X1 U10097 ( .A(n8410), .ZN(n8411) );
  NAND2_X1 U10098 ( .A1(n8411), .A2(n9032), .ZN(n8412) );
  XNOR2_X1 U10099 ( .A(n8510), .B(n4460), .ZN(n8504) );
  XNOR2_X1 U10100 ( .A(n9190), .B(n8107), .ZN(n8413) );
  OAI22_X1 U10101 ( .A1(n8504), .A2(n9001), .B1(n8984), .B2(n8413), .ZN(n8417)
         );
  OAI21_X1 U10102 ( .B1(n8502), .B2(n9014), .A(n8779), .ZN(n8415) );
  NOR2_X1 U10103 ( .A1(n8779), .A2(n9014), .ZN(n8414) );
  AOI22_X1 U10104 ( .A1(n8415), .A2(n8504), .B1(n8414), .B2(n8413), .ZN(n8416)
         );
  XOR2_X1 U10105 ( .A(n4460), .B(n9180), .Z(n8419) );
  INV_X1 U10106 ( .A(n8419), .ZN(n8418) );
  XNOR2_X1 U10107 ( .A(n8418), .B(n8778), .ZN(n8479) );
  NOR2_X1 U10108 ( .A1(n8419), .A2(n8778), .ZN(n8420) );
  XNOR2_X1 U10109 ( .A(n8970), .B(n8107), .ZN(n8548) );
  NAND2_X1 U10110 ( .A1(n8548), .A2(n8975), .ZN(n8421) );
  NAND2_X1 U10111 ( .A1(n8547), .A2(n8421), .ZN(n8424) );
  INV_X1 U10112 ( .A(n8548), .ZN(n8422) );
  NAND2_X1 U10113 ( .A1(n8422), .A2(n8777), .ZN(n8423) );
  XNOR2_X1 U10114 ( .A(n8451), .B(n8107), .ZN(n8425) );
  XNOR2_X1 U10115 ( .A(n8425), .B(n8776), .ZN(n8446) );
  INV_X1 U10116 ( .A(n8425), .ZN(n8426) );
  XOR2_X1 U10117 ( .A(n4460), .B(n8610), .Z(n8427) );
  NAND2_X1 U10118 ( .A1(n8774), .A2(n8561), .ZN(n8430) );
  AOI22_X1 U10119 ( .A1(n8428), .A2(n8565), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8429) );
  OAI211_X1 U10120 ( .C1(n8966), .C2(n8563), .A(n8430), .B(n8429), .ZN(n8431)
         );
  AOI21_X1 U10121 ( .B1(n9169), .B2(n8553), .A(n8431), .ZN(n8432) );
  OAI222_X1 U10122 ( .A1(n9246), .A2(n8572), .B1(n9258), .B2(n8435), .C1(
        P2_U3151), .C2(n8433), .ZN(P2_U3265) );
  OAI21_X1 U10123 ( .B1(n8438), .B2(n8437), .A(n8436), .ZN(n8439) );
  NAND2_X1 U10124 ( .A1(n8439), .A2(n9434), .ZN(n8443) );
  AOI22_X1 U10125 ( .A1(n9460), .A2(n8441), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8440), .ZN(n8442) );
  OAI211_X1 U10126 ( .C1(n4588), .C2(n9412), .A(n8443), .B(n8442), .ZN(
        P1_U3222) );
  INV_X1 U10127 ( .A(n8445), .ZN(n9259) );
  OAI222_X1 U10128 ( .A1(n8378), .A2(n10285), .B1(P1_U3086), .B2(n10031), .C1(
        n9259), .C2(n10029), .ZN(P1_U3328) );
  XNOR2_X1 U10129 ( .A(n8447), .B(n8446), .ZN(n8453) );
  NAND2_X1 U10130 ( .A1(n8775), .A2(n8561), .ZN(n8449) );
  AOI22_X1 U10131 ( .A1(n8955), .A2(n8565), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8448) );
  OAI211_X1 U10132 ( .C1(n8975), .C2(n8563), .A(n8449), .B(n8448), .ZN(n8450)
         );
  AOI21_X1 U10133 ( .B1(n8451), .B2(n8553), .A(n8450), .ZN(n8452) );
  OAI21_X1 U10134 ( .B1(n8453), .B2(n8555), .A(n8452), .ZN(P2_U3154) );
  XNOR2_X1 U10135 ( .A(n8503), .B(n8984), .ZN(n8459) );
  NAND2_X1 U10136 ( .A1(n8779), .A2(n8561), .ZN(n8456) );
  AOI22_X1 U10137 ( .A1(n9005), .A2(n8565), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8455) );
  OAI211_X1 U10138 ( .C1(n9000), .C2(n8563), .A(n8456), .B(n8455), .ZN(n8457)
         );
  AOI21_X1 U10139 ( .B1(n9190), .B2(n8553), .A(n8457), .ZN(n8458) );
  OAI21_X1 U10140 ( .B1(n8459), .B2(n8555), .A(n8458), .ZN(P2_U3156) );
  INV_X1 U10141 ( .A(n9060), .ZN(n9212) );
  AOI21_X1 U10142 ( .B1(n8461), .B2(n8460), .A(n8555), .ZN(n8463) );
  NAND2_X1 U10143 ( .A1(n8463), .A2(n8462), .ZN(n8469) );
  NAND2_X1 U10144 ( .A1(n9054), .A2(n8561), .ZN(n8465) );
  OAI211_X1 U10145 ( .C1(n8466), .C2(n8563), .A(n8465), .B(n8464), .ZN(n8467)
         );
  AOI21_X1 U10146 ( .B1(n9059), .B2(n8565), .A(n8467), .ZN(n8468) );
  OAI211_X1 U10147 ( .C1(n9212), .C2(n8568), .A(n8469), .B(n8468), .ZN(
        P2_U3159) );
  XOR2_X1 U10148 ( .A(n8471), .B(n8470), .Z(n8477) );
  INV_X1 U10149 ( .A(n8472), .ZN(n9202) );
  AOI22_X1 U10150 ( .A1(n9054), .A2(n8539), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8474) );
  NAND2_X1 U10151 ( .A1(n9035), .A2(n8565), .ZN(n8473) );
  OAI211_X1 U10152 ( .C1(n9000), .C2(n8541), .A(n8474), .B(n8473), .ZN(n8475)
         );
  AOI21_X1 U10153 ( .B1(n9202), .B2(n8553), .A(n8475), .ZN(n8476) );
  OAI21_X1 U10154 ( .B1(n8477), .B2(n8555), .A(n8476), .ZN(P2_U3163) );
  XOR2_X1 U10155 ( .A(n8479), .B(n8478), .Z(n8484) );
  NAND2_X1 U10156 ( .A1(n8777), .A2(n8561), .ZN(n8481) );
  AOI22_X1 U10157 ( .A1(n8977), .A2(n8565), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8480) );
  OAI211_X1 U10158 ( .C1(n9001), .C2(n8563), .A(n8481), .B(n8480), .ZN(n8482)
         );
  AOI21_X1 U10159 ( .B1(n9180), .B2(n8553), .A(n8482), .ZN(n8483) );
  OAI21_X1 U10160 ( .B1(n8484), .B2(n8555), .A(n8483), .ZN(P2_U3165) );
  OAI211_X1 U10161 ( .C1(n8487), .C2(n8486), .A(n8485), .B(n8557), .ZN(n8492)
         );
  NAND2_X1 U10162 ( .A1(n9092), .A2(n8561), .ZN(n8488) );
  NAND2_X1 U10163 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8893) );
  OAI211_X1 U10164 ( .C1(n8489), .C2(n8563), .A(n8488), .B(n8893), .ZN(n8490)
         );
  AOI21_X1 U10165 ( .B1(n9095), .B2(n8565), .A(n8490), .ZN(n8491) );
  OAI211_X1 U10166 ( .C1(n8493), .C2(n8568), .A(n8492), .B(n8491), .ZN(
        P2_U3166) );
  INV_X1 U10167 ( .A(n8494), .ZN(n8535) );
  AOI21_X1 U10168 ( .B1(n8496), .B2(n8495), .A(n8535), .ZN(n8501) );
  NAND2_X1 U10169 ( .A1(n9082), .A2(n8561), .ZN(n8497) );
  NAND2_X1 U10170 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8905) );
  OAI211_X1 U10171 ( .C1(n9104), .C2(n8563), .A(n8497), .B(n8905), .ZN(n8498)
         );
  AOI21_X1 U10172 ( .B1(n9084), .B2(n8565), .A(n8498), .ZN(n8500) );
  NAND2_X1 U10173 ( .A1(n9225), .A2(n8553), .ZN(n8499) );
  OAI211_X1 U10174 ( .C1(n8501), .C2(n8555), .A(n8500), .B(n8499), .ZN(
        P2_U3168) );
  OAI22_X1 U10175 ( .A1(n8503), .A2(n9014), .B1(n8502), .B2(n8454), .ZN(n8506)
         );
  XNOR2_X1 U10176 ( .A(n8504), .B(n9001), .ZN(n8505) );
  XNOR2_X1 U10177 ( .A(n8506), .B(n8505), .ZN(n8512) );
  NAND2_X1 U10178 ( .A1(n8778), .A2(n8561), .ZN(n8508) );
  AOI22_X1 U10179 ( .A1(n8987), .A2(n8565), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8507) );
  OAI211_X1 U10180 ( .C1(n8984), .C2(n8563), .A(n8508), .B(n8507), .ZN(n8509)
         );
  AOI21_X1 U10181 ( .B1(n8510), .B2(n8553), .A(n8509), .ZN(n8511) );
  OAI21_X1 U10182 ( .B1(n8512), .B2(n8555), .A(n8511), .ZN(P2_U3169) );
  INV_X1 U10183 ( .A(n8513), .ZN(n8514) );
  AOI21_X1 U10184 ( .B1(n8516), .B2(n8515), .A(n8514), .ZN(n8521) );
  AOI22_X1 U10185 ( .A1(n9067), .A2(n8539), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8518) );
  NAND2_X1 U10186 ( .A1(n9046), .A2(n8565), .ZN(n8517) );
  OAI211_X1 U10187 ( .C1(n8527), .C2(n8541), .A(n8518), .B(n8517), .ZN(n8519)
         );
  AOI21_X1 U10188 ( .B1(n6610), .B2(n8553), .A(n8519), .ZN(n8520) );
  OAI21_X1 U10189 ( .B1(n8521), .B2(n8555), .A(n8520), .ZN(P2_U3173) );
  INV_X1 U10190 ( .A(n9196), .ZN(n8531) );
  AOI21_X1 U10191 ( .B1(n8523), .B2(n8522), .A(n8555), .ZN(n8525) );
  NAND2_X1 U10192 ( .A1(n8525), .A2(n8524), .ZN(n8530) );
  AOI22_X1 U10193 ( .A1(n9017), .A2(n8565), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8526) );
  OAI21_X1 U10194 ( .B1(n8527), .B2(n8563), .A(n8526), .ZN(n8528) );
  AOI21_X1 U10195 ( .B1(n9014), .B2(n8561), .A(n8528), .ZN(n8529) );
  OAI211_X1 U10196 ( .C1(n8531), .C2(n8568), .A(n8530), .B(n8529), .ZN(
        P2_U3175) );
  INV_X1 U10197 ( .A(n9219), .ZN(n8546) );
  INV_X1 U10198 ( .A(n8532), .ZN(n8534) );
  NOR3_X1 U10199 ( .A1(n8535), .A2(n8534), .A3(n8533), .ZN(n8538) );
  INV_X1 U10200 ( .A(n8536), .ZN(n8537) );
  OAI21_X1 U10201 ( .B1(n8538), .B2(n8537), .A(n8557), .ZN(n8545) );
  AND2_X1 U10202 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8936) );
  AOI21_X1 U10203 ( .B1(n9092), .B2(n8539), .A(n8936), .ZN(n8540) );
  OAI21_X1 U10204 ( .B1(n8542), .B2(n8541), .A(n8540), .ZN(n8543) );
  AOI21_X1 U10205 ( .B1(n9070), .B2(n8565), .A(n8543), .ZN(n8544) );
  OAI211_X1 U10206 ( .C1(n8546), .C2(n8568), .A(n8545), .B(n8544), .ZN(
        P2_U3178) );
  XNOR2_X1 U10207 ( .A(n8548), .B(n8777), .ZN(n8549) );
  XNOR2_X1 U10208 ( .A(n8547), .B(n8549), .ZN(n8556) );
  NAND2_X1 U10209 ( .A1(n8776), .A2(n8561), .ZN(n8551) );
  AOI22_X1 U10210 ( .A1(n8969), .A2(n8565), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8550) );
  OAI211_X1 U10211 ( .C1(n8985), .C2(n8563), .A(n8551), .B(n8550), .ZN(n8552)
         );
  AOI21_X1 U10212 ( .B1(n8970), .B2(n8553), .A(n8552), .ZN(n8554) );
  OAI21_X1 U10213 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(P2_U3180) );
  INV_X1 U10214 ( .A(n9149), .ZN(n8569) );
  OAI211_X1 U10215 ( .C1(n4599), .C2(n8559), .A(n8558), .B(n8557), .ZN(n8567)
         );
  NAND2_X1 U10216 ( .A1(n9081), .A2(n8561), .ZN(n8562) );
  NAND2_X1 U10217 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8874) );
  OAI211_X1 U10218 ( .C1(n9103), .C2(n8563), .A(n8562), .B(n8874), .ZN(n8564)
         );
  AOI21_X1 U10219 ( .B1(n9105), .B2(n8565), .A(n8564), .ZN(n8566) );
  OAI211_X1 U10220 ( .C1(n8569), .C2(n8568), .A(n8567), .B(n8566), .ZN(
        P2_U3181) );
  NAND2_X1 U10221 ( .A1(n9244), .A2(n6486), .ZN(n8571) );
  OR2_X1 U10222 ( .A1(n6430), .A2(n9247), .ZN(n8570) );
  INV_X1 U10223 ( .A(n9112), .ZN(n9161) );
  NOR2_X1 U10224 ( .A1(n6430), .A2(n8572), .ZN(n8574) );
  INV_X1 U10225 ( .A(n9164), .ZN(n8577) );
  OR2_X1 U10226 ( .A1(n9112), .A2(n8941), .ZN(n8580) );
  NAND2_X1 U10227 ( .A1(n8577), .A2(n8581), .ZN(n8745) );
  AND2_X1 U10228 ( .A1(n8745), .A2(n8578), .ZN(n8579) );
  INV_X1 U10229 ( .A(n8581), .ZN(n8773) );
  AND2_X1 U10230 ( .A1(n9164), .A2(n8773), .ZN(n8754) );
  INV_X1 U10231 ( .A(n8754), .ZN(n8746) );
  NAND2_X1 U10232 ( .A1(n8746), .A2(n8750), .ZN(n8582) );
  AND2_X1 U10233 ( .A1(n8582), .A2(n9112), .ZN(n8583) );
  XNOR2_X1 U10234 ( .A(n8585), .B(n8584), .ZN(n8616) );
  INV_X1 U10235 ( .A(n8737), .ZN(n8611) );
  AND2_X1 U10236 ( .A1(n9112), .A2(n8941), .ZN(n8755) );
  INV_X1 U10237 ( .A(n8729), .ZN(n8586) );
  INV_X1 U10238 ( .A(n8723), .ZN(n8587) );
  INV_X1 U10239 ( .A(n8718), .ZN(n8707) );
  NAND2_X1 U10240 ( .A1(n8707), .A2(n8588), .ZN(n8990) );
  INV_X1 U10241 ( .A(n8589), .ZN(n9030) );
  INV_X1 U10242 ( .A(n9077), .ZN(n9079) );
  NOR4_X1 U10243 ( .A1(n8593), .A2(n10119), .A3(n4620), .A4(n8592), .ZN(n8597)
         );
  NAND2_X1 U10244 ( .A1(n8595), .A2(n8594), .ZN(n10106) );
  NAND4_X1 U10245 ( .A1(n8597), .A2(n8596), .A3(n10106), .A4(n5087), .ZN(n8600) );
  NOR4_X1 U10246 ( .A1(n8601), .A2(n8600), .A3(n6476), .A4(n8599), .ZN(n8602)
         );
  NAND4_X1 U10247 ( .A1(n8604), .A2(n8603), .A3(n8670), .A4(n8602), .ZN(n8605)
         );
  NOR4_X1 U10248 ( .A1(n9089), .A2(n9101), .A3(n8674), .A4(n8605), .ZN(n8606)
         );
  NAND2_X1 U10249 ( .A1(n9079), .A2(n8606), .ZN(n8607) );
  NOR4_X1 U10250 ( .A1(n9041), .A2(n9065), .A3(n9052), .A4(n8607), .ZN(n8608)
         );
  NAND4_X1 U10251 ( .A1(n8996), .A2(n9012), .A3(n9030), .A4(n8608), .ZN(n8609)
         );
  OAI21_X1 U10252 ( .B1(n8614), .B2(n7011), .A(n8613), .ZN(n8615) );
  AOI21_X1 U10253 ( .B1(n8616), .B2(n7011), .A(n8615), .ZN(n8765) );
  OAI21_X1 U10254 ( .B1(n4889), .B2(n8617), .A(n8717), .ZN(n8709) );
  INV_X1 U10255 ( .A(n8618), .ZN(n8619) );
  AOI21_X1 U10256 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(n8673) );
  OAI211_X1 U10257 ( .C1(n8623), .C2(n7011), .A(n8622), .B(n6697), .ZN(n8630)
         );
  OAI22_X1 U10258 ( .A1(n8624), .A2(n4620), .B1(n8626), .B2(n4889), .ZN(n8629)
         );
  INV_X1 U10259 ( .A(n8625), .ZN(n8627) );
  MUX2_X1 U10260 ( .A(n8627), .B(n8626), .S(n4889), .Z(n8628) );
  NAND2_X1 U10261 ( .A1(n8631), .A2(n8637), .ZN(n8634) );
  NAND2_X1 U10262 ( .A1(n8632), .A2(n8651), .ZN(n8633) );
  MUX2_X1 U10263 ( .A(n8634), .B(n8633), .S(n4889), .Z(n8635) );
  OAI21_X1 U10264 ( .B1(n8636), .B2(n8635), .A(n5087), .ZN(n8654) );
  INV_X1 U10265 ( .A(n8637), .ZN(n8640) );
  NAND2_X1 U10266 ( .A1(n8790), .A2(n8638), .ZN(n8639) );
  OAI211_X1 U10267 ( .C1(n8654), .C2(n8640), .A(n8655), .B(n8639), .ZN(n8643)
         );
  NAND2_X1 U10268 ( .A1(n8662), .A2(n8661), .ZN(n8641) );
  NAND2_X1 U10269 ( .A1(n8646), .A2(n8645), .ZN(n8665) );
  AND2_X1 U10270 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  OAI211_X1 U10271 ( .C1(n8648), .C2(n8647), .A(n8666), .B(n8646), .ZN(n8649)
         );
  OAI21_X1 U10272 ( .B1(n8650), .B2(n8649), .A(n8663), .ZN(n8669) );
  INV_X1 U10273 ( .A(n8651), .ZN(n8653) );
  OAI211_X1 U10274 ( .C1(n8654), .C2(n8653), .A(n10102), .B(n8652), .ZN(n8657)
         );
  AND2_X1 U10275 ( .A1(n8661), .A2(n8660), .ZN(n8664) );
  OAI211_X1 U10276 ( .C1(n8665), .C2(n8664), .A(n8663), .B(n8662), .ZN(n8667)
         );
  MUX2_X1 U10277 ( .A(n8669), .B(n8668), .S(n6697), .Z(n8671) );
  INV_X1 U10278 ( .A(n8674), .ZN(n8678) );
  MUX2_X1 U10279 ( .A(n8676), .B(n8675), .S(n4889), .Z(n8677) );
  NAND2_X1 U10280 ( .A1(n8678), .A2(n8677), .ZN(n8683) );
  NAND2_X1 U10281 ( .A1(n8679), .A2(n8780), .ZN(n8680) );
  MUX2_X1 U10282 ( .A(n8681), .B(n8680), .S(n4889), .Z(n8682) );
  MUX2_X1 U10283 ( .A(n8685), .B(n8684), .S(n4889), .Z(n8686) );
  NOR2_X1 U10284 ( .A1(n9089), .A2(n8686), .ZN(n8690) );
  INV_X1 U10285 ( .A(n8687), .ZN(n9075) );
  MUX2_X1 U10286 ( .A(n9075), .B(n8688), .S(n6697), .Z(n8689) );
  NAND2_X1 U10287 ( .A1(n8695), .A2(n8691), .ZN(n8692) );
  OAI21_X1 U10288 ( .B1(n8698), .B2(n8692), .A(n8694), .ZN(n8699) );
  NAND2_X1 U10289 ( .A1(n8694), .A2(n8693), .ZN(n8697) );
  INV_X1 U10290 ( .A(n8700), .ZN(n8701) );
  INV_X1 U10291 ( .A(n8711), .ZN(n8703) );
  INV_X1 U10292 ( .A(n8710), .ZN(n9023) );
  AOI21_X1 U10293 ( .B1(n8713), .B2(n9024), .A(n8703), .ZN(n8705) );
  NAND3_X1 U10294 ( .A1(n9196), .A2(n9000), .A3(n4889), .ZN(n8706) );
  OAI211_X1 U10295 ( .C1(n8720), .C2(n6697), .A(n8707), .B(n8706), .ZN(n8708)
         );
  NAND3_X1 U10296 ( .A1(n8712), .A2(n8711), .A3(n8710), .ZN(n8714) );
  NAND2_X1 U10297 ( .A1(n8714), .A2(n8713), .ZN(n8716) );
  INV_X1 U10298 ( .A(n8717), .ZN(n8719) );
  AOI21_X1 U10299 ( .B1(n8720), .B2(n8719), .A(n8718), .ZN(n8721) );
  INV_X1 U10300 ( .A(n8722), .ZN(n8724) );
  MUX2_X1 U10301 ( .A(n8724), .B(n8723), .S(n6697), .Z(n8725) );
  INV_X1 U10302 ( .A(n8727), .ZN(n8728) );
  MUX2_X1 U10303 ( .A(n8729), .B(n8728), .S(n4889), .Z(n8730) );
  OAI21_X1 U10304 ( .B1(n8774), .B2(n6697), .A(n8752), .ZN(n8732) );
  OAI21_X1 U10305 ( .B1(n8733), .B2(n6697), .A(n8732), .ZN(n8739) );
  MUX2_X1 U10306 ( .A(n8735), .B(n8734), .S(n6697), .Z(n8736) );
  MUX2_X1 U10307 ( .A(n8775), .B(n9169), .S(n6697), .Z(n8738) );
  NAND2_X1 U10308 ( .A1(n8741), .A2(n8738), .ZN(n8756) );
  NAND2_X1 U10309 ( .A1(n8756), .A2(n8737), .ZN(n8744) );
  NOR2_X1 U10310 ( .A1(n8758), .A2(n8775), .ZN(n8743) );
  INV_X1 U10311 ( .A(n8745), .ZN(n8747) );
  OAI21_X1 U10312 ( .B1(n8747), .B2(n6697), .A(n8746), .ZN(n8748) );
  INV_X1 U10313 ( .A(n8748), .ZN(n8751) );
  OAI21_X1 U10314 ( .B1(n8748), .B2(n8941), .A(n9112), .ZN(n8749) );
  OAI21_X1 U10315 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(n8760) );
  INV_X1 U10316 ( .A(n8752), .ZN(n8753) );
  NOR4_X1 U10317 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n6697), .ZN(n8757)
         );
  OAI211_X1 U10318 ( .C1(n8758), .C2(n9169), .A(n8757), .B(n8756), .ZN(n8759)
         );
  NAND3_X1 U10319 ( .A1(n8768), .A2(n8767), .A3(n8766), .ZN(n8769) );
  OAI211_X1 U10320 ( .C1(n8771), .C2(n8770), .A(n8769), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8772) );
  MUX2_X1 U10321 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8773), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10322 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8774), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10323 ( .A(n8775), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8929), .Z(
        P2_U3519) );
  MUX2_X1 U10324 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8776), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10325 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8777), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10326 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8778), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10327 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8779), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10328 ( .A(n9014), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8929), .Z(
        P2_U3514) );
  MUX2_X1 U10329 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9032), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10330 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9043), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10331 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9054), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10332 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9067), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10333 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9082), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10334 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9092), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10335 ( .A(n9081), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8929), .Z(
        P2_U3507) );
  MUX2_X1 U10336 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9091), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10337 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8780), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10338 ( .A(n8781), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8929), .Z(
        P2_U3504) );
  MUX2_X1 U10339 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8782), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10340 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8783), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10341 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8784), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10342 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8785), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10343 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8786), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10344 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8787), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10345 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8788), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10346 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8789), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10347 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8790), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10348 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8791), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10349 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8792), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10350 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8793), .S(P2_U3893), .Z(
        P2_U3492) );
  OAI211_X1 U10351 ( .C1(n8796), .C2(n8795), .A(n8794), .B(n8883), .ZN(n8811)
         );
  OAI21_X1 U10352 ( .B1(n8928), .B2(n8798), .A(n8797), .ZN(n8799) );
  AOI21_X1 U10353 ( .B1(n10099), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8799), .ZN(
        n8810) );
  AND3_X1 U10354 ( .A1(n8801), .A2(n8800), .A3(n5941), .ZN(n8802) );
  OAI21_X1 U10355 ( .B1(n8803), .B2(n8802), .A(n8922), .ZN(n8809) );
  OAI21_X1 U10356 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n8807) );
  NAND2_X1 U10357 ( .A1(n10092), .A2(n8807), .ZN(n8808) );
  NAND4_X1 U10358 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(
        P2_U3186) );
  XNOR2_X1 U10359 ( .A(n8812), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n8824) );
  OAI21_X1 U10360 ( .B1(n8928), .B2(n4771), .A(n8813), .ZN(n8818) );
  NAND2_X1 U10361 ( .A1(n8815), .A2(n8814), .ZN(n8816) );
  AOI21_X1 U10362 ( .B1(n8832), .B2(n8816), .A(n10088), .ZN(n8817) );
  AOI211_X1 U10363 ( .C1(n10099), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8818), .B(
        n8817), .ZN(n8823) );
  XNOR2_X1 U10364 ( .A(n8820), .B(n8819), .ZN(n8821) );
  NAND2_X1 U10365 ( .A1(n8821), .A2(n8883), .ZN(n8822) );
  OAI211_X1 U10366 ( .C1(n8824), .C2(n8939), .A(n8823), .B(n8822), .ZN(
        P2_U3193) );
  XOR2_X1 U10367 ( .A(n8826), .B(n8825), .Z(n8842) );
  OAI21_X1 U10368 ( .B1(n8928), .B2(n8828), .A(n8827), .ZN(n8836) );
  INV_X1 U10369 ( .A(n8829), .ZN(n8831) );
  NAND3_X1 U10370 ( .A1(n8832), .A2(n8831), .A3(n8830), .ZN(n8833) );
  AOI21_X1 U10371 ( .B1(n8834), .B2(n8833), .A(n10088), .ZN(n8835) );
  AOI211_X1 U10372 ( .C1(n10099), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n8836), .B(
        n8835), .ZN(n8841) );
  XNOR2_X1 U10373 ( .A(n8838), .B(n8837), .ZN(n8839) );
  NAND2_X1 U10374 ( .A1(n8839), .A2(n8883), .ZN(n8840) );
  OAI211_X1 U10375 ( .C1(n8842), .C2(n8939), .A(n8841), .B(n8840), .ZN(
        P2_U3194) );
  XNOR2_X1 U10376 ( .A(n8843), .B(n10381), .ZN(n8855) );
  OAI21_X1 U10377 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8844), .A(n8863), .ZN(
        n8853) );
  XOR2_X1 U10378 ( .A(n8846), .B(n8845), .Z(n8851) );
  NAND2_X1 U10379 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n8847) );
  OAI21_X1 U10380 ( .B1(n8928), .B2(n8848), .A(n8847), .ZN(n8849) );
  AOI21_X1 U10381 ( .B1(n10099), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8849), .ZN(
        n8850) );
  OAI21_X1 U10382 ( .B1(n8851), .B2(n10095), .A(n8850), .ZN(n8852) );
  AOI21_X1 U10383 ( .B1(n8853), .B2(n8922), .A(n8852), .ZN(n8854) );
  OAI21_X1 U10384 ( .B1(n8855), .B2(n8939), .A(n8854), .ZN(P2_U3195) );
  XOR2_X1 U10385 ( .A(n8857), .B(n8856), .Z(n8870) );
  XNOR2_X1 U10386 ( .A(n8859), .B(n8858), .ZN(n8868) );
  NAND2_X1 U10387 ( .A1(n10099), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U10388 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8860) );
  OAI211_X1 U10389 ( .C1(n8928), .C2(n4785), .A(n8861), .B(n8860), .ZN(n8867)
         );
  NAND3_X1 U10390 ( .A1(n8863), .A2(n4562), .A3(n8862), .ZN(n8864) );
  AOI21_X1 U10391 ( .B1(n8865), .B2(n8864), .A(n10088), .ZN(n8866) );
  AOI211_X1 U10392 ( .C1(n8883), .C2(n8868), .A(n8867), .B(n8866), .ZN(n8869)
         );
  OAI21_X1 U10393 ( .B1(n8870), .B2(n8939), .A(n8869), .ZN(P2_U3196) );
  XOR2_X1 U10394 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8871), .Z(n8885) );
  XNOR2_X1 U10395 ( .A(n8873), .B(n8872), .ZN(n8882) );
  NAND2_X1 U10396 ( .A1(n10099), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8875) );
  OAI211_X1 U10397 ( .C1(n8928), .C2(n8876), .A(n8875), .B(n8874), .ZN(n8881)
         );
  NAND2_X1 U10398 ( .A1(n8877), .A2(n9107), .ZN(n8878) );
  AOI21_X1 U10399 ( .B1(n8879), .B2(n8878), .A(n10088), .ZN(n8880) );
  AOI211_X1 U10400 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(n8884)
         );
  OAI21_X1 U10401 ( .B1(n8885), .B2(n8939), .A(n8884), .ZN(P2_U3197) );
  XOR2_X1 U10402 ( .A(n8887), .B(n8886), .Z(n8900) );
  OAI21_X1 U10403 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8898) );
  XOR2_X1 U10404 ( .A(n8892), .B(n8891), .Z(n8896) );
  OAI21_X1 U10405 ( .B1(n8928), .B2(n5989), .A(n8893), .ZN(n8894) );
  AOI21_X1 U10406 ( .B1(n10099), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8894), .ZN(
        n8895) );
  OAI21_X1 U10407 ( .B1(n8896), .B2(n10095), .A(n8895), .ZN(n8897) );
  AOI21_X1 U10408 ( .B1(n8898), .B2(n8922), .A(n8897), .ZN(n8899) );
  OAI21_X1 U10409 ( .B1(n8939), .B2(n8900), .A(n8899), .ZN(P2_U3198) );
  XOR2_X1 U10410 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8901), .Z(n8913) );
  OAI21_X1 U10411 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8902), .A(n8916), .ZN(
        n8911) );
  XOR2_X1 U10412 ( .A(n8904), .B(n8903), .Z(n8909) );
  OAI21_X1 U10413 ( .B1(n8928), .B2(n8906), .A(n8905), .ZN(n8907) );
  AOI21_X1 U10414 ( .B1(n10099), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8907), .ZN(
        n8908) );
  OAI21_X1 U10415 ( .B1(n8909), .B2(n10095), .A(n8908), .ZN(n8910) );
  AOI21_X1 U10416 ( .B1(n8911), .B2(n8922), .A(n8910), .ZN(n8912) );
  OAI21_X1 U10417 ( .B1(n8913), .B2(n8939), .A(n8912), .ZN(P2_U3199) );
  INV_X1 U10418 ( .A(n8916), .ZN(n8920) );
  INV_X1 U10419 ( .A(n8917), .ZN(n8919) );
  INV_X1 U10420 ( .A(n8921), .ZN(n8923) );
  OAI21_X1 U10421 ( .B1(n8924), .B2(n8923), .A(n8922), .ZN(n8938) );
  INV_X1 U10422 ( .A(n8925), .ZN(n8926) );
  INV_X1 U10423 ( .A(n8931), .ZN(n8930) );
  OAI21_X1 U10424 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8934) );
  NOR2_X1 U10425 ( .A1(n8931), .A2(n10095), .ZN(n8933) );
  MUX2_X1 U10426 ( .A(n8934), .B(n8933), .S(n8932), .Z(n8935) );
  AOI211_X1 U10427 ( .C1(n10099), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8936), .B(
        n8935), .ZN(n8937) );
  NAND2_X1 U10428 ( .A1(n9112), .A2(n9109), .ZN(n8943) );
  NOR2_X1 U10429 ( .A1(n8942), .A2(n10123), .ZN(n8951) );
  AOI21_X1 U10430 ( .B1(n9159), .B2(n10141), .A(n8951), .ZN(n8946) );
  OAI211_X1 U10431 ( .C1(n10141), .C2(n8944), .A(n8943), .B(n8946), .ZN(
        P2_U3202) );
  NAND2_X1 U10432 ( .A1(n10144), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U10433 ( .C1(n9164), .C2(n10111), .A(n8946), .B(n8945), .ZN(
        P2_U3203) );
  NOR2_X1 U10434 ( .A1(n8948), .A2(n8947), .ZN(n8949) );
  AOI21_X1 U10435 ( .B1(n10144), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8951), .ZN(
        n8952) );
  INV_X1 U10436 ( .A(n8954), .ZN(n8961) );
  AOI22_X1 U10437 ( .A1(n8955), .A2(n9096), .B1(n10144), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8956) );
  OAI21_X1 U10438 ( .B1(n8957), .B2(n10111), .A(n8956), .ZN(n8958) );
  AOI21_X1 U10439 ( .B1(n8959), .B2(n8992), .A(n8958), .ZN(n8960) );
  OAI21_X1 U10440 ( .B1(n8961), .B2(n10144), .A(n8960), .ZN(P2_U3206) );
  XOR2_X1 U10441 ( .A(n8963), .B(n8962), .Z(n9174) );
  XNOR2_X1 U10442 ( .A(n8964), .B(n8963), .ZN(n8965) );
  OAI222_X1 U10443 ( .A1(n10127), .A2(n8966), .B1(n10125), .B2(n8985), .C1(
        n10132), .C2(n8965), .ZN(n9173) );
  INV_X1 U10444 ( .A(n9173), .ZN(n8967) );
  MUX2_X1 U10445 ( .A(n8968), .B(n8967), .S(n10141), .Z(n8972) );
  AOI22_X1 U10446 ( .A1(n8970), .A2(n9109), .B1(n9096), .B2(n8969), .ZN(n8971)
         );
  OAI211_X1 U10447 ( .C1(n9174), .C2(n10115), .A(n8972), .B(n8971), .ZN(
        P2_U3207) );
  NOR2_X1 U10448 ( .A1(n9118), .A2(n10122), .ZN(n8976) );
  XNOR2_X1 U10449 ( .A(n8973), .B(n4880), .ZN(n8974) );
  OAI222_X1 U10450 ( .A1(n10127), .A2(n8975), .B1(n10125), .B2(n9001), .C1(
        n8974), .C2(n10132), .ZN(n9177) );
  AOI211_X1 U10451 ( .C1(n9096), .C2(n8977), .A(n8976), .B(n9177), .ZN(n8981)
         );
  XNOR2_X1 U10452 ( .A(n8978), .B(n4880), .ZN(n9183) );
  INV_X1 U10453 ( .A(n9183), .ZN(n8979) );
  AOI22_X1 U10454 ( .A1(n8979), .A2(n8992), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10144), .ZN(n8980) );
  OAI21_X1 U10455 ( .B1(n8981), .B2(n10144), .A(n8980), .ZN(P2_U3208) );
  NOR2_X1 U10456 ( .A1(n9185), .A2(n10122), .ZN(n8986) );
  XNOR2_X1 U10457 ( .A(n8982), .B(n8990), .ZN(n8983) );
  OAI222_X1 U10458 ( .A1(n10127), .A2(n8985), .B1(n10125), .B2(n8984), .C1(
        n10132), .C2(n8983), .ZN(n9184) );
  AOI211_X1 U10459 ( .C1(n9096), .C2(n8987), .A(n8986), .B(n9184), .ZN(n8995)
         );
  NAND2_X1 U10460 ( .A1(n8989), .A2(n8988), .ZN(n8991) );
  XNOR2_X1 U10461 ( .A(n8991), .B(n8990), .ZN(n9186) );
  INV_X1 U10462 ( .A(n9186), .ZN(n8993) );
  AOI22_X1 U10463 ( .A1(n8993), .A2(n8992), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10144), .ZN(n8994) );
  OAI21_X1 U10464 ( .B1(n8995), .B2(n10144), .A(n8994), .ZN(P2_U3209) );
  XNOR2_X1 U10465 ( .A(n4614), .B(n8998), .ZN(n9193) );
  INV_X1 U10466 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9004) );
  XNOR2_X1 U10467 ( .A(n8999), .B(n8998), .ZN(n9003) );
  OAI22_X1 U10468 ( .A1(n9001), .A2(n10127), .B1(n9000), .B2(n10125), .ZN(
        n9002) );
  AOI21_X1 U10469 ( .B1(n9003), .B2(n9094), .A(n9002), .ZN(n9189) );
  MUX2_X1 U10470 ( .A(n9004), .B(n9189), .S(n10141), .Z(n9007) );
  AOI22_X1 U10471 ( .A1(n9190), .A2(n9109), .B1(n9096), .B2(n9005), .ZN(n9006)
         );
  OAI211_X1 U10472 ( .C1(n9193), .C2(n10115), .A(n9007), .B(n9006), .ZN(
        P2_U3210) );
  XNOR2_X1 U10473 ( .A(n9008), .B(n9012), .ZN(n9199) );
  INV_X1 U10474 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9016) );
  NAND3_X1 U10475 ( .A1(n9010), .A2(n9012), .A3(n9011), .ZN(n9013) );
  NAND2_X1 U10476 ( .A1(n9009), .A2(n9013), .ZN(n9015) );
  AOI222_X1 U10477 ( .A1(n9094), .A2(n9015), .B1(n9014), .B2(n6698), .C1(n9043), .C2(n9090), .ZN(n9194) );
  MUX2_X1 U10478 ( .A(n9016), .B(n9194), .S(n10141), .Z(n9019) );
  AOI22_X1 U10479 ( .A1(n9196), .A2(n9109), .B1(n9096), .B2(n9017), .ZN(n9018)
         );
  OAI211_X1 U10480 ( .C1(n9199), .C2(n10115), .A(n9019), .B(n9018), .ZN(
        P2_U3211) );
  INV_X1 U10481 ( .A(n9052), .ZN(n9049) );
  INV_X1 U10482 ( .A(n9021), .ZN(n9022) );
  AOI21_X1 U10483 ( .B1(n9050), .B2(n9049), .A(n9022), .ZN(n9038) );
  AOI21_X1 U10484 ( .B1(n9038), .B2(n9024), .A(n9023), .ZN(n9025) );
  XNOR2_X1 U10485 ( .A(n9025), .B(n9030), .ZN(n9205) );
  INV_X1 U10486 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U10487 ( .A1(n9066), .A2(n9065), .ZN(n9064) );
  INV_X1 U10488 ( .A(n9027), .ZN(n9028) );
  NAND2_X1 U10489 ( .A1(n9064), .A2(n9028), .ZN(n9051) );
  NAND3_X1 U10490 ( .A1(n9051), .A2(n9041), .A3(n9039), .ZN(n9040) );
  NAND3_X1 U10491 ( .A1(n9040), .A2(n9030), .A3(n9029), .ZN(n9031) );
  NAND2_X1 U10492 ( .A1(n9031), .A2(n9010), .ZN(n9033) );
  AOI222_X1 U10493 ( .A1(n9094), .A2(n9033), .B1(n9032), .B2(n6698), .C1(n9054), .C2(n9090), .ZN(n9200) );
  MUX2_X1 U10494 ( .A(n9034), .B(n9200), .S(n10141), .Z(n9037) );
  AOI22_X1 U10495 ( .A1(n9202), .A2(n9109), .B1(n9096), .B2(n9035), .ZN(n9036)
         );
  OAI211_X1 U10496 ( .C1(n9205), .C2(n10115), .A(n9037), .B(n9036), .ZN(
        P2_U3212) );
  XNOR2_X1 U10497 ( .A(n9038), .B(n9041), .ZN(n9210) );
  AND2_X1 U10498 ( .A1(n9051), .A2(n9039), .ZN(n9042) );
  OAI21_X1 U10499 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9044) );
  AOI222_X1 U10500 ( .A1(n9094), .A2(n9044), .B1(n9043), .B2(n6698), .C1(n9067), .C2(n9090), .ZN(n9206) );
  MUX2_X1 U10501 ( .A(n9045), .B(n9206), .S(n10141), .Z(n9048) );
  AOI22_X1 U10502 ( .A1(n6610), .A2(n9109), .B1(n9096), .B2(n9046), .ZN(n9047)
         );
  OAI211_X1 U10503 ( .C1(n9210), .C2(n10115), .A(n9048), .B(n9047), .ZN(
        P2_U3213) );
  XNOR2_X1 U10504 ( .A(n9050), .B(n9049), .ZN(n9213) );
  NAND2_X1 U10505 ( .A1(n9051), .A2(n9094), .ZN(n9057) );
  AOI21_X1 U10506 ( .B1(n9064), .B2(n9053), .A(n9052), .ZN(n9056) );
  AOI22_X1 U10507 ( .A1(n9054), .A2(n6698), .B1(n9090), .B2(n9082), .ZN(n9055)
         );
  OAI21_X1 U10508 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9214) );
  INV_X1 U10509 ( .A(n9214), .ZN(n9058) );
  MUX2_X1 U10510 ( .A(n10366), .B(n9058), .S(n10141), .Z(n9062) );
  AOI22_X1 U10511 ( .A1(n9060), .A2(n9109), .B1(n9096), .B2(n9059), .ZN(n9061)
         );
  OAI211_X1 U10512 ( .C1(n9213), .C2(n10115), .A(n9062), .B(n9061), .ZN(
        P2_U3214) );
  XNOR2_X1 U10513 ( .A(n9063), .B(n9065), .ZN(n9222) );
  OAI21_X1 U10514 ( .B1(n9066), .B2(n9065), .A(n9064), .ZN(n9068) );
  AOI222_X1 U10515 ( .A1(n9094), .A2(n9068), .B1(n9067), .B2(n6698), .C1(n9092), .C2(n9090), .ZN(n9217) );
  MUX2_X1 U10516 ( .A(n9069), .B(n9217), .S(n10141), .Z(n9072) );
  AOI22_X1 U10517 ( .A1(n9219), .A2(n9109), .B1(n9096), .B2(n9070), .ZN(n9071)
         );
  OAI211_X1 U10518 ( .C1(n9222), .C2(n10115), .A(n9072), .B(n9071), .ZN(
        P2_U3215) );
  NAND2_X1 U10519 ( .A1(n9074), .A2(n9073), .ZN(n9087) );
  AOI21_X1 U10520 ( .B1(n9087), .B2(n9076), .A(n9075), .ZN(n9078) );
  XNOR2_X1 U10521 ( .A(n9078), .B(n9077), .ZN(n9228) );
  XNOR2_X1 U10522 ( .A(n9080), .B(n9079), .ZN(n9083) );
  AOI222_X1 U10523 ( .A1(n9094), .A2(n9083), .B1(n9082), .B2(n6698), .C1(n9081), .C2(n9090), .ZN(n9223) );
  MUX2_X1 U10524 ( .A(n4917), .B(n9223), .S(n10141), .Z(n9086) );
  AOI22_X1 U10525 ( .A1(n9225), .A2(n9109), .B1(n9096), .B2(n9084), .ZN(n9085)
         );
  OAI211_X1 U10526 ( .C1(n9228), .C2(n10115), .A(n9086), .B(n9085), .ZN(
        P2_U3216) );
  XOR2_X1 U10527 ( .A(n9089), .B(n9087), .Z(n9235) );
  XOR2_X1 U10528 ( .A(n9088), .B(n9089), .Z(n9093) );
  AOI222_X1 U10529 ( .A1(n9094), .A2(n9093), .B1(n9092), .B2(n6698), .C1(n9091), .C2(n9090), .ZN(n9229) );
  MUX2_X1 U10530 ( .A(n10395), .B(n9229), .S(n10141), .Z(n9098) );
  AOI22_X1 U10531 ( .A1(n9231), .A2(n9109), .B1(n9096), .B2(n9095), .ZN(n9097)
         );
  OAI211_X1 U10532 ( .C1(n9235), .C2(n10115), .A(n9098), .B(n9097), .ZN(
        P2_U3217) );
  XNOR2_X1 U10533 ( .A(n9099), .B(n9101), .ZN(n9151) );
  XNOR2_X1 U10534 ( .A(n9100), .B(n9101), .ZN(n9102) );
  OAI222_X1 U10535 ( .A1(n10127), .A2(n9104), .B1(n10125), .B2(n9103), .C1(
        n9102), .C2(n10132), .ZN(n9148) );
  NAND2_X1 U10536 ( .A1(n9148), .A2(n10141), .ZN(n9111) );
  INV_X1 U10537 ( .A(n9105), .ZN(n9106) );
  OAI22_X1 U10538 ( .A1(n10141), .A2(n9107), .B1(n9106), .B2(n10123), .ZN(
        n9108) );
  AOI21_X1 U10539 ( .B1(n9149), .B2(n9109), .A(n9108), .ZN(n9110) );
  OAI211_X1 U10540 ( .C1(n9151), .C2(n10115), .A(n9111), .B(n9110), .ZN(
        P2_U3218) );
  NAND2_X1 U10541 ( .A1(n9112), .A2(n9154), .ZN(n9113) );
  NAND2_X1 U10542 ( .A1(n9159), .A2(n10189), .ZN(n9115) );
  OAI211_X1 U10543 ( .C1(n10189), .C2(n10498), .A(n9113), .B(n9115), .ZN(
        P2_U3490) );
  NAND2_X1 U10544 ( .A1(n10187), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9114) );
  OAI211_X1 U10545 ( .C1(n9164), .C2(n9135), .A(n9115), .B(n9114), .ZN(
        P2_U3489) );
  MUX2_X1 U10546 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9173), .S(n10189), .Z(
        n9117) );
  OAI22_X1 U10547 ( .A1(n9174), .A2(n9147), .B1(n6657), .B2(n9135), .ZN(n9116)
         );
  OR2_X1 U10548 ( .A1(n9117), .A2(n9116), .ZN(P2_U3485) );
  MUX2_X1 U10549 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9177), .S(n10189), .Z(
        n9120) );
  OAI22_X1 U10550 ( .A1(n9183), .A2(n9147), .B1(n9118), .B2(n9135), .ZN(n9119)
         );
  OR2_X1 U10551 ( .A1(n9120), .A2(n9119), .ZN(P2_U3484) );
  MUX2_X1 U10552 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9184), .S(n10189), .Z(
        n9122) );
  OAI22_X1 U10553 ( .A1(n9186), .A2(n9147), .B1(n9185), .B2(n9135), .ZN(n9121)
         );
  OR2_X1 U10554 ( .A1(n9122), .A2(n9121), .ZN(P2_U3483) );
  INV_X1 U10555 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9123) );
  MUX2_X1 U10556 ( .A(n9123), .B(n9189), .S(n10189), .Z(n9125) );
  NAND2_X1 U10557 ( .A1(n9190), .A2(n9154), .ZN(n9124) );
  OAI211_X1 U10558 ( .C1(n9193), .C2(n9147), .A(n9125), .B(n9124), .ZN(
        P2_U3482) );
  INV_X1 U10559 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9126) );
  MUX2_X1 U10560 ( .A(n9126), .B(n9194), .S(n10189), .Z(n9128) );
  NAND2_X1 U10561 ( .A1(n9196), .A2(n9154), .ZN(n9127) );
  OAI211_X1 U10562 ( .C1(n9199), .C2(n9147), .A(n9128), .B(n9127), .ZN(
        P2_U3481) );
  INV_X1 U10563 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10564 ( .A(n9129), .B(n9200), .S(n10189), .Z(n9131) );
  NAND2_X1 U10565 ( .A1(n9202), .A2(n9154), .ZN(n9130) );
  OAI211_X1 U10566 ( .C1(n9147), .C2(n9205), .A(n9131), .B(n9130), .ZN(
        P2_U3480) );
  INV_X1 U10567 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U10568 ( .A(n9132), .B(n9206), .S(n10189), .Z(n9134) );
  NAND2_X1 U10569 ( .A1(n6610), .A2(n9154), .ZN(n9133) );
  OAI211_X1 U10570 ( .C1(n9210), .C2(n9147), .A(n9134), .B(n9133), .ZN(
        P2_U3479) );
  OAI22_X1 U10571 ( .A1(n9213), .A2(n9147), .B1(n9212), .B2(n9135), .ZN(n9137)
         );
  MUX2_X1 U10572 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9214), .S(n10189), .Z(
        n9136) );
  OR2_X1 U10573 ( .A1(n9137), .A2(n9136), .ZN(P2_U3478) );
  MUX2_X1 U10574 ( .A(n9138), .B(n9217), .S(n10189), .Z(n9140) );
  NAND2_X1 U10575 ( .A1(n9219), .A2(n9154), .ZN(n9139) );
  OAI211_X1 U10576 ( .C1(n9147), .C2(n9222), .A(n9140), .B(n9139), .ZN(
        P2_U3477) );
  INV_X1 U10577 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10578 ( .A(n9141), .B(n9223), .S(n10189), .Z(n9143) );
  NAND2_X1 U10579 ( .A1(n9225), .A2(n9154), .ZN(n9142) );
  OAI211_X1 U10580 ( .C1(n9228), .C2(n9147), .A(n9143), .B(n9142), .ZN(
        P2_U3476) );
  MUX2_X1 U10581 ( .A(n9144), .B(n9229), .S(n10189), .Z(n9146) );
  NAND2_X1 U10582 ( .A1(n9231), .A2(n9154), .ZN(n9145) );
  OAI211_X1 U10583 ( .C1(n9235), .C2(n9147), .A(n9146), .B(n9145), .ZN(
        P2_U3475) );
  INV_X1 U10584 ( .A(n10162), .ZN(n10168) );
  AOI21_X1 U10585 ( .B1(n10161), .B2(n9149), .A(n9148), .ZN(n9150) );
  OAI21_X1 U10586 ( .B1(n10168), .B2(n9151), .A(n9150), .ZN(n9236) );
  MUX2_X1 U10587 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9236), .S(n10189), .Z(
        P2_U3474) );
  INV_X1 U10588 ( .A(n9152), .ZN(n9237) );
  MUX2_X1 U10589 ( .A(n9153), .B(n9237), .S(n10189), .Z(n9157) );
  AOI22_X1 U10590 ( .A1(n9241), .A2(n9155), .B1(n9154), .B2(n9239), .ZN(n9156)
         );
  NAND2_X1 U10591 ( .A1(n9157), .A2(n9156), .ZN(P2_U3473) );
  MUX2_X1 U10592 ( .A(n9158), .B(P2_REG1_REG_0__SCAN_IN), .S(n10187), .Z(
        P2_U3459) );
  NAND2_X1 U10593 ( .A1(n10180), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U10594 ( .A1(n9159), .A2(n10178), .ZN(n9163) );
  OAI211_X1 U10595 ( .C1(n9161), .C2(n9211), .A(n9160), .B(n9163), .ZN(
        P2_U3458) );
  NAND2_X1 U10596 ( .A1(n10180), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U10597 ( .C1(n9164), .C2(n9211), .A(n9163), .B(n9162), .ZN(
        P2_U3457) );
  NAND2_X1 U10598 ( .A1(n10180), .A2(n9166), .ZN(n9167) );
  NAND2_X1 U10599 ( .A1(n9169), .A2(n6799), .ZN(n9170) );
  MUX2_X1 U10600 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9173), .S(n10178), .Z(
        n9176) );
  OAI22_X1 U10601 ( .A1(n9174), .A2(n9234), .B1(n6657), .B2(n9211), .ZN(n9175)
         );
  OR2_X1 U10602 ( .A1(n9176), .A2(n9175), .ZN(P2_U3453) );
  INV_X1 U10603 ( .A(n9177), .ZN(n9178) );
  MUX2_X1 U10604 ( .A(n9179), .B(n9178), .S(n10178), .Z(n9182) );
  NAND2_X1 U10605 ( .A1(n9180), .A2(n6799), .ZN(n9181) );
  OAI211_X1 U10606 ( .C1(n9183), .C2(n9234), .A(n9182), .B(n9181), .ZN(
        P2_U3452) );
  MUX2_X1 U10607 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9184), .S(n10178), .Z(
        n9188) );
  OAI22_X1 U10608 ( .A1(n9186), .A2(n9234), .B1(n9185), .B2(n9211), .ZN(n9187)
         );
  OR2_X1 U10609 ( .A1(n9188), .A2(n9187), .ZN(P2_U3451) );
  MUX2_X1 U10610 ( .A(n10497), .B(n9189), .S(n10178), .Z(n9192) );
  NAND2_X1 U10611 ( .A1(n9190), .A2(n6799), .ZN(n9191) );
  OAI211_X1 U10612 ( .C1(n9193), .C2(n9234), .A(n9192), .B(n9191), .ZN(
        P2_U3450) );
  MUX2_X1 U10613 ( .A(n9195), .B(n9194), .S(n10178), .Z(n9198) );
  NAND2_X1 U10614 ( .A1(n9196), .A2(n6799), .ZN(n9197) );
  OAI211_X1 U10615 ( .C1(n9199), .C2(n9234), .A(n9198), .B(n9197), .ZN(
        P2_U3449) );
  MUX2_X1 U10616 ( .A(n9201), .B(n9200), .S(n10178), .Z(n9204) );
  NAND2_X1 U10617 ( .A1(n9202), .A2(n6799), .ZN(n9203) );
  OAI211_X1 U10618 ( .C1(n9205), .C2(n9234), .A(n9204), .B(n9203), .ZN(
        P2_U3448) );
  INV_X1 U10619 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9207) );
  MUX2_X1 U10620 ( .A(n9207), .B(n9206), .S(n10178), .Z(n9209) );
  NAND2_X1 U10621 ( .A1(n6610), .A2(n6799), .ZN(n9208) );
  OAI211_X1 U10622 ( .C1(n9210), .C2(n9234), .A(n9209), .B(n9208), .ZN(
        P2_U3447) );
  OAI22_X1 U10623 ( .A1(n9213), .A2(n9234), .B1(n9212), .B2(n9211), .ZN(n9216)
         );
  MUX2_X1 U10624 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9214), .S(n10178), .Z(
        n9215) );
  OR2_X1 U10625 ( .A1(n9216), .A2(n9215), .ZN(P2_U3446) );
  INV_X1 U10626 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9218) );
  MUX2_X1 U10627 ( .A(n9218), .B(n9217), .S(n10178), .Z(n9221) );
  NAND2_X1 U10628 ( .A1(n9219), .A2(n6799), .ZN(n9220) );
  OAI211_X1 U10629 ( .C1(n9222), .C2(n9234), .A(n9221), .B(n9220), .ZN(
        P2_U3444) );
  MUX2_X1 U10630 ( .A(n9224), .B(n9223), .S(n10178), .Z(n9227) );
  NAND2_X1 U10631 ( .A1(n9225), .A2(n6799), .ZN(n9226) );
  OAI211_X1 U10632 ( .C1(n9228), .C2(n9234), .A(n9227), .B(n9226), .ZN(
        P2_U3441) );
  INV_X1 U10633 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9230) );
  MUX2_X1 U10634 ( .A(n9230), .B(n9229), .S(n10178), .Z(n9233) );
  NAND2_X1 U10635 ( .A1(n9231), .A2(n6799), .ZN(n9232) );
  OAI211_X1 U10636 ( .C1(n9235), .C2(n9234), .A(n9233), .B(n9232), .ZN(
        P2_U3438) );
  MUX2_X1 U10637 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9236), .S(n10178), .Z(
        P2_U3435) );
  MUX2_X1 U10638 ( .A(n9238), .B(n9237), .S(n10178), .Z(n9243) );
  AOI22_X1 U10639 ( .A1(n9241), .A2(n9240), .B1(n6799), .B2(n9239), .ZN(n9242)
         );
  NAND2_X1 U10640 ( .A1(n9243), .A2(n9242), .ZN(P2_U3432) );
  INV_X1 U10641 ( .A(n9244), .ZN(n10026) );
  NAND3_X1 U10642 ( .A1(n4863), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9248) );
  OAI22_X1 U10643 ( .A1(n9249), .A2(n9248), .B1(n9247), .B2(n9246), .ZN(n9250)
         );
  INV_X1 U10644 ( .A(n9250), .ZN(n9251) );
  OAI21_X1 U10645 ( .B1(n10026), .B2(n9258), .A(n9251), .ZN(P2_U3264) );
  AOI21_X1 U10646 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9256), .A(n9252), .ZN(
        n9253) );
  OAI21_X1 U10647 ( .B1(n9254), .B2(n9258), .A(n9253), .ZN(P2_U3267) );
  AOI21_X1 U10648 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9256), .A(n9255), .ZN(
        n9257) );
  OAI21_X1 U10649 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(P2_U3268) );
  INV_X1 U10650 ( .A(n9260), .ZN(n9261) );
  MUX2_X1 U10651 ( .A(n9261), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10652 ( .B1(n9435), .B2(n9263), .A(n9262), .ZN(n9264) );
  OAI21_X1 U10653 ( .B1(n9265), .B2(n9264), .A(n9434), .ZN(n9274) );
  OR2_X1 U10654 ( .A1(n9266), .A2(n9455), .ZN(n9268) );
  NAND2_X1 U10655 ( .A1(n9474), .A2(n9457), .ZN(n9267) );
  AND2_X1 U10656 ( .A1(n9268), .A2(n9267), .ZN(n9685) );
  INV_X1 U10657 ( .A(n9685), .ZN(n9272) );
  INV_X1 U10658 ( .A(n9691), .ZN(n9270) );
  OAI22_X1 U10659 ( .A1(n9270), .A2(n9462), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9269), .ZN(n9271) );
  AOI21_X1 U10660 ( .B1(n9272), .B2(n9460), .A(n9271), .ZN(n9273) );
  OAI211_X1 U10661 ( .C1(n9975), .C2(n9412), .A(n9274), .B(n9273), .ZN(
        P1_U3214) );
  INV_X1 U10662 ( .A(n9275), .ZN(n9277) );
  NAND2_X1 U10663 ( .A1(n9277), .A2(n9276), .ZN(n9280) );
  NAND2_X1 U10664 ( .A1(n9280), .A2(n9279), .ZN(n9450) );
  INV_X1 U10665 ( .A(n9450), .ZN(n9282) );
  NAND2_X1 U10666 ( .A1(n9275), .A2(n9278), .ZN(n9449) );
  AOI21_X1 U10667 ( .B1(n9280), .B2(n9449), .A(n9279), .ZN(n9281) );
  AOI21_X1 U10668 ( .B1(n9282), .B2(n9449), .A(n9281), .ZN(n9291) );
  INV_X1 U10669 ( .A(n9283), .ZN(n9288) );
  NAND2_X1 U10670 ( .A1(n9460), .A2(n9284), .ZN(n9287) );
  INV_X1 U10671 ( .A(n9285), .ZN(n9286) );
  OAI211_X1 U10672 ( .C1(n9462), .C2(n9288), .A(n9287), .B(n9286), .ZN(n9289)
         );
  AOI21_X1 U10673 ( .B1(n9963), .B2(n9465), .A(n9289), .ZN(n9290) );
  OAI21_X1 U10674 ( .B1(n9291), .B2(n9467), .A(n9290), .ZN(P1_U3215) );
  INV_X1 U10675 ( .A(n9292), .ZN(n9293) );
  NOR2_X1 U10676 ( .A1(n9294), .A2(n9293), .ZN(n9295) );
  XNOR2_X1 U10677 ( .A(n9296), .B(n9295), .ZN(n9302) );
  AND2_X1 U10678 ( .A1(n9478), .A2(n9457), .ZN(n9297) );
  AOI21_X1 U10679 ( .B1(n9476), .B2(n9426), .A(n9297), .ZN(n9747) );
  INV_X1 U10680 ( .A(n9298), .ZN(n9753) );
  AOI22_X1 U10681 ( .A1(n9753), .A2(n9442), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9299) );
  OAI21_X1 U10682 ( .B1(n9747), .B2(n9444), .A(n9299), .ZN(n9300) );
  AOI21_X1 U10683 ( .B1(n9752), .B2(n9465), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10684 ( .B1(n9302), .B2(n9467), .A(n9301), .ZN(P1_U3216) );
  NOR2_X1 U10685 ( .A1(n9303), .A2(n9305), .ZN(n9421) );
  INV_X1 U10686 ( .A(n9304), .ZN(n9424) );
  NAND2_X1 U10687 ( .A1(n9303), .A2(n9305), .ZN(n9422) );
  OAI21_X1 U10688 ( .B1(n9421), .B2(n9424), .A(n9422), .ZN(n9309) );
  NAND2_X1 U10689 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  XNOR2_X1 U10690 ( .A(n9309), .B(n9308), .ZN(n9314) );
  NOR2_X1 U10691 ( .A1(n9462), .A2(n9811), .ZN(n9312) );
  AND2_X1 U10692 ( .A1(n9482), .A2(n9457), .ZN(n9310) );
  AOI21_X1 U10693 ( .B1(n9480), .B2(n9426), .A(n9310), .ZN(n9805) );
  NAND2_X1 U10694 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9641) );
  OAI21_X1 U10695 ( .B1(n9805), .B2(n9444), .A(n9641), .ZN(n9311) );
  AOI211_X1 U10696 ( .C1(n10006), .C2(n9465), .A(n9312), .B(n9311), .ZN(n9313)
         );
  OAI21_X1 U10697 ( .B1(n9314), .B2(n9467), .A(n9313), .ZN(P1_U3219) );
  NAND2_X1 U10698 ( .A1(n9460), .A2(n9315), .ZN(n9317) );
  OAI211_X1 U10699 ( .C1(n9462), .C2(n9318), .A(n9317), .B(n9316), .ZN(n9324)
         );
  AOI21_X1 U10700 ( .B1(n9321), .B2(n9320), .A(n9319), .ZN(n9322) );
  NOR2_X1 U10701 ( .A1(n9322), .A2(n9467), .ZN(n9323) );
  AOI211_X1 U10702 ( .C1(n9325), .C2(n9465), .A(n9324), .B(n9323), .ZN(n9326)
         );
  INV_X1 U10703 ( .A(n9326), .ZN(P1_U3221) );
  OAI211_X1 U10704 ( .C1(n9327), .C2(n9329), .A(n9328), .B(n9434), .ZN(n9337)
         );
  INV_X1 U10705 ( .A(n9330), .ZN(n9780) );
  NAND2_X1 U10706 ( .A1(n9478), .A2(n9426), .ZN(n9332) );
  NAND2_X1 U10707 ( .A1(n9480), .A2(n9457), .ZN(n9331) );
  NAND2_X1 U10708 ( .A1(n9332), .A2(n9331), .ZN(n9773) );
  INV_X1 U10709 ( .A(n9773), .ZN(n9334) );
  OAI22_X1 U10710 ( .A1(n9334), .A2(n9444), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9333), .ZN(n9335) );
  AOI21_X1 U10711 ( .B1(n9780), .B2(n9442), .A(n9335), .ZN(n9336) );
  OAI211_X1 U10712 ( .C1(n9999), .C2(n9412), .A(n9337), .B(n9336), .ZN(
        P1_U3223) );
  INV_X1 U10713 ( .A(n9338), .ZN(n9352) );
  INV_X1 U10714 ( .A(n9339), .ZN(n9341) );
  NOR3_X1 U10715 ( .A1(n9342), .A2(n9341), .A3(n9340), .ZN(n9345) );
  INV_X1 U10716 ( .A(n9343), .ZN(n9344) );
  OAI21_X1 U10717 ( .B1(n9345), .B2(n9344), .A(n9434), .ZN(n9351) );
  NOR2_X1 U10718 ( .A1(n9462), .A2(n9346), .ZN(n9347) );
  AOI211_X1 U10719 ( .C1(n9460), .C2(n9349), .A(n9348), .B(n9347), .ZN(n9350)
         );
  OAI211_X1 U10720 ( .C1(n9352), .C2(n9412), .A(n9351), .B(n9350), .ZN(
        P1_U3224) );
  OAI21_X1 U10721 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(n9356) );
  NAND2_X1 U10722 ( .A1(n9356), .A2(n9434), .ZN(n9363) );
  AOI22_X1 U10723 ( .A1(n9722), .A2(n9442), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9362) );
  NAND2_X1 U10724 ( .A1(n9357), .A2(n9465), .ZN(n9361) );
  OAI22_X1 U10725 ( .A1(n9359), .A2(n9455), .B1(n9358), .B2(n9369), .ZN(n9714)
         );
  NAND2_X1 U10726 ( .A1(n9714), .A2(n9460), .ZN(n9360) );
  NAND4_X1 U10727 ( .A1(n9363), .A2(n9362), .A3(n9361), .A4(n9360), .ZN(
        P1_U3225) );
  INV_X1 U10728 ( .A(n9365), .ZN(n9367) );
  NAND2_X1 U10729 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  XNOR2_X1 U10730 ( .A(n9364), .B(n9368), .ZN(n9376) );
  INV_X1 U10731 ( .A(n9868), .ZN(n9373) );
  OAI22_X1 U10732 ( .A1(n9371), .A2(n9455), .B1(n9370), .B2(n9369), .ZN(n9856)
         );
  AOI22_X1 U10733 ( .A1(n9460), .A2(n9856), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9372) );
  OAI21_X1 U10734 ( .B1(n9373), .B2(n9462), .A(n9372), .ZN(n9374) );
  AOI21_X1 U10735 ( .B1(n9867), .B2(n9465), .A(n9374), .ZN(n9375) );
  OAI21_X1 U10736 ( .B1(n9376), .B2(n9467), .A(n9375), .ZN(P1_U3226) );
  NOR2_X1 U10737 ( .A1(n9378), .A2(n4976), .ZN(n9379) );
  XNOR2_X1 U10738 ( .A(n9380), .B(n9379), .ZN(n9385) );
  AOI22_X1 U10739 ( .A1(n9484), .A2(n9457), .B1(n9426), .B2(n9482), .ZN(n9840)
         );
  NAND2_X1 U10740 ( .A1(n9442), .A2(n9846), .ZN(n9381) );
  OAI211_X1 U10741 ( .C1(n9444), .C2(n9840), .A(n9382), .B(n9381), .ZN(n9383)
         );
  AOI21_X1 U10742 ( .B1(n9842), .B2(n9465), .A(n9383), .ZN(n9384) );
  OAI21_X1 U10743 ( .B1(n9385), .B2(n9467), .A(n9384), .ZN(P1_U3228) );
  OAI21_X1 U10744 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9392) );
  AOI22_X1 U10745 ( .A1(n9475), .A2(n9426), .B1(n9457), .B2(n9477), .ZN(n9732)
         );
  NAND2_X1 U10746 ( .A1(n9736), .A2(n9465), .ZN(n9390) );
  AOI22_X1 U10747 ( .A1(n9737), .A2(n9442), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9389) );
  OAI211_X1 U10748 ( .C1(n9732), .C2(n9444), .A(n9390), .B(n9389), .ZN(n9391)
         );
  AOI21_X1 U10749 ( .B1(n9392), .B2(n9434), .A(n9391), .ZN(n9393) );
  INV_X1 U10750 ( .A(n9393), .ZN(P1_U3229) );
  NAND2_X1 U10751 ( .A1(n4557), .A2(n9395), .ZN(n9396) );
  XNOR2_X1 U10752 ( .A(n9394), .B(n9396), .ZN(n9401) );
  NOR2_X1 U10753 ( .A1(n9462), .A2(n9794), .ZN(n9399) );
  AOI22_X1 U10754 ( .A1(n9479), .A2(n9426), .B1(n9457), .B2(n9481), .ZN(n9787)
         );
  OAI22_X1 U10755 ( .A1(n9787), .A2(n9444), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9397), .ZN(n9398) );
  AOI211_X1 U10756 ( .C1(n9791), .C2(n9465), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OAI21_X1 U10757 ( .B1(n9401), .B2(n9467), .A(n9400), .ZN(P1_U3233) );
  OAI21_X1 U10758 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n9405) );
  NAND2_X1 U10759 ( .A1(n9405), .A2(n9434), .ZN(n9411) );
  OAI21_X1 U10760 ( .B1(n9444), .B2(n9407), .A(n9406), .ZN(n9408) );
  AOI21_X1 U10761 ( .B1(n9409), .B2(n9442), .A(n9408), .ZN(n9410) );
  OAI211_X1 U10762 ( .C1(n5135), .C2(n9412), .A(n9411), .B(n9410), .ZN(
        P1_U3234) );
  NAND2_X1 U10763 ( .A1(n4534), .A2(n9413), .ZN(n9415) );
  XNOR2_X1 U10764 ( .A(n9415), .B(n9414), .ZN(n9420) );
  AOI22_X1 U10765 ( .A1(n9477), .A2(n9426), .B1(n9457), .B2(n9479), .ZN(n9761)
         );
  AOI22_X1 U10766 ( .A1(n9442), .A2(n9764), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9416) );
  OAI21_X1 U10767 ( .B1(n9761), .B2(n9444), .A(n9416), .ZN(n9417) );
  AOI21_X1 U10768 ( .B1(n9418), .B2(n9465), .A(n9417), .ZN(n9419) );
  OAI21_X1 U10769 ( .B1(n9420), .B2(n9467), .A(n9419), .ZN(P1_U3235) );
  INV_X1 U10770 ( .A(n9421), .ZN(n9423) );
  NAND2_X1 U10771 ( .A1(n9423), .A2(n9422), .ZN(n9425) );
  XNOR2_X1 U10772 ( .A(n9425), .B(n9424), .ZN(n9432) );
  NAND2_X1 U10773 ( .A1(n9943), .A2(n9465), .ZN(n9430) );
  NAND2_X1 U10774 ( .A1(n9481), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U10775 ( .A1(n9483), .A2(n9457), .ZN(n9427) );
  NAND2_X1 U10776 ( .A1(n9428), .A2(n9427), .ZN(n9825) );
  AOI22_X1 U10777 ( .A1(n9460), .A2(n9825), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9429) );
  OAI211_X1 U10778 ( .C1(n9462), .C2(n9828), .A(n9430), .B(n9429), .ZN(n9431)
         );
  AOI21_X1 U10779 ( .B1(n9432), .B2(n9434), .A(n9431), .ZN(n9433) );
  INV_X1 U10780 ( .A(n9433), .ZN(P1_U3238) );
  NAND2_X1 U10781 ( .A1(n9435), .A2(n9434), .ZN(n9448) );
  AOI21_X1 U10782 ( .B1(n9353), .B2(n9437), .A(n9436), .ZN(n9447) );
  OR2_X1 U10783 ( .A1(n9438), .A2(n9455), .ZN(n9440) );
  NAND2_X1 U10784 ( .A1(n9475), .A2(n9457), .ZN(n9439) );
  AND2_X1 U10785 ( .A1(n9440), .A2(n9439), .ZN(n9701) );
  INV_X1 U10786 ( .A(n9441), .ZN(n9707) );
  AOI22_X1 U10787 ( .A1(n9707), .A2(n9442), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9443) );
  OAI21_X1 U10788 ( .B1(n9701), .B2(n9444), .A(n9443), .ZN(n9445) );
  AOI21_X1 U10789 ( .B1(n9706), .B2(n9465), .A(n9445), .ZN(n9446) );
  OAI21_X1 U10790 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(P1_U3240) );
  NAND2_X1 U10791 ( .A1(n9450), .A2(n9449), .ZN(n9454) );
  XNOR2_X1 U10792 ( .A(n9452), .B(n9451), .ZN(n9453) );
  XNOR2_X1 U10793 ( .A(n9454), .B(n9453), .ZN(n9468) );
  INV_X1 U10794 ( .A(n9888), .ZN(n9463) );
  OR2_X1 U10795 ( .A1(n9456), .A2(n9455), .ZN(n9459) );
  NAND2_X1 U10796 ( .A1(n9486), .A2(n9457), .ZN(n9458) );
  NAND2_X1 U10797 ( .A1(n9459), .A2(n9458), .ZN(n9880) );
  AOI22_X1 U10798 ( .A1(n9460), .A2(n9880), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9461) );
  OAI21_X1 U10799 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  AOI21_X1 U10800 ( .B1(n9886), .B2(n9465), .A(n9464), .ZN(n9466) );
  OAI21_X1 U10801 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(P1_U3241) );
  MUX2_X1 U10802 ( .A(n9470), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9469), .Z(
        P1_U3584) );
  MUX2_X1 U10803 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9471), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10804 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9472), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10805 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9473), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10806 ( .A(n9474), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9469), .Z(
        P1_U3580) );
  MUX2_X1 U10807 ( .A(n9475), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9469), .Z(
        P1_U3579) );
  MUX2_X1 U10808 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9476), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10809 ( .A(n9477), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9469), .Z(
        P1_U3577) );
  MUX2_X1 U10810 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9478), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10811 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9479), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10812 ( .A(n9480), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9469), .Z(
        P1_U3574) );
  MUX2_X1 U10813 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9481), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10814 ( .A(n9482), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9469), .Z(
        P1_U3572) );
  MUX2_X1 U10815 ( .A(n9483), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9469), .Z(
        P1_U3571) );
  MUX2_X1 U10816 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9484), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10817 ( .A(n9485), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9469), .Z(
        P1_U3569) );
  MUX2_X1 U10818 ( .A(n9486), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9469), .Z(
        P1_U3568) );
  MUX2_X1 U10819 ( .A(n9487), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9469), .Z(
        P1_U3567) );
  MUX2_X1 U10820 ( .A(n9488), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9469), .Z(
        P1_U3566) );
  MUX2_X1 U10821 ( .A(n9489), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9469), .Z(
        P1_U3565) );
  MUX2_X1 U10822 ( .A(n9490), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9469), .Z(
        P1_U3564) );
  MUX2_X1 U10823 ( .A(n9491), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9469), .Z(
        P1_U3563) );
  MUX2_X1 U10824 ( .A(n9492), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9469), .Z(
        P1_U3562) );
  MUX2_X1 U10825 ( .A(n9493), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9469), .Z(
        P1_U3561) );
  MUX2_X1 U10826 ( .A(n9494), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9469), .Z(
        P1_U3560) );
  MUX2_X1 U10827 ( .A(n9495), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9469), .Z(
        P1_U3559) );
  MUX2_X1 U10828 ( .A(n9496), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9469), .Z(
        P1_U3558) );
  MUX2_X1 U10829 ( .A(n9497), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9469), .Z(
        P1_U3557) );
  MUX2_X1 U10830 ( .A(n9498), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9469), .Z(
        P1_U3556) );
  MUX2_X1 U10831 ( .A(n5317), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9469), .Z(
        P1_U3555) );
  INV_X1 U10832 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9515) );
  MUX2_X1 U10833 ( .A(n9499), .B(P1_REG1_REG_1__SCAN_IN), .S(n9502), .Z(n9500)
         );
  OAI21_X1 U10834 ( .B1(n6127), .B2(n9515), .A(n9500), .ZN(n9501) );
  NAND3_X1 U10835 ( .A1(n9632), .A2(n9523), .A3(n9501), .ZN(n9509) );
  AOI22_X1 U10836 ( .A1(n10038), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9508) );
  NAND2_X1 U10837 ( .A1(n9636), .A2(n9502), .ZN(n9507) );
  OAI211_X1 U10838 ( .C1(n9505), .C2(n9504), .A(n9638), .B(n9503), .ZN(n9506)
         );
  NAND4_X1 U10839 ( .A1(n9509), .A2(n9508), .A3(n9507), .A4(n9506), .ZN(
        P1_U3244) );
  INV_X1 U10840 ( .A(n9510), .ZN(n9511) );
  MUX2_X1 U10841 ( .A(n9512), .B(n9511), .S(n10031), .Z(n9516) );
  OR2_X1 U10842 ( .A1(n10031), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U10843 ( .A1(n9514), .A2(n9513), .ZN(n10032) );
  NAND2_X1 U10844 ( .A1(n10032), .A2(n9515), .ZN(n10035) );
  OAI211_X1 U10845 ( .C1(n9516), .C2(n5824), .A(P1_U3973), .B(n10035), .ZN(
        n9559) );
  INV_X1 U10846 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9518) );
  INV_X1 U10847 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9517) );
  OAI22_X1 U10848 ( .A1(n9643), .A2(n9518), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9517), .ZN(n9519) );
  AOI21_X1 U10849 ( .B1(n9636), .B2(n9520), .A(n9519), .ZN(n9532) );
  MUX2_X1 U10850 ( .A(n9521), .B(P1_REG1_REG_2__SCAN_IN), .S(n9520), .Z(n9524)
         );
  NAND3_X1 U10851 ( .A1(n9524), .A2(n9523), .A3(n9522), .ZN(n9525) );
  NAND3_X1 U10852 ( .A1(n9632), .A2(n9526), .A3(n9525), .ZN(n9531) );
  OAI211_X1 U10853 ( .C1(n9529), .C2(n9528), .A(n9638), .B(n9527), .ZN(n9530)
         );
  NAND4_X1 U10854 ( .A1(n9559), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(
        P1_U3245) );
  OAI211_X1 U10855 ( .C1(n9534), .C2(n9533), .A(n9632), .B(n9554), .ZN(n9543)
         );
  INV_X1 U10856 ( .A(n9535), .ZN(n9537) );
  INV_X1 U10857 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10226) );
  OAI22_X1 U10858 ( .A1(n9643), .A2(n10226), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10043), .ZN(n9536) );
  AOI21_X1 U10859 ( .B1(n9636), .B2(n9537), .A(n9536), .ZN(n9542) );
  OAI211_X1 U10860 ( .C1(n9540), .C2(n9539), .A(n9638), .B(n9538), .ZN(n9541)
         );
  NAND3_X1 U10861 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(P1_U3246) );
  INV_X1 U10862 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9545) );
  OAI21_X1 U10863 ( .B1(n9643), .B2(n9545), .A(n9544), .ZN(n9546) );
  AOI21_X1 U10864 ( .B1(n9636), .B2(n9547), .A(n9546), .ZN(n9558) );
  OAI211_X1 U10865 ( .C1(n9550), .C2(n9549), .A(n9638), .B(n9548), .ZN(n9557)
         );
  INV_X1 U10866 ( .A(n9551), .ZN(n9564) );
  NAND3_X1 U10867 ( .A1(n9554), .A2(n9553), .A3(n9552), .ZN(n9555) );
  NAND3_X1 U10868 ( .A1(n9632), .A2(n9564), .A3(n9555), .ZN(n9556) );
  NAND4_X1 U10869 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(
        P1_U3247) );
  INV_X1 U10870 ( .A(n9560), .ZN(n9563) );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6930), .S(n9561), .Z(n9562)
         );
  NAND3_X1 U10872 ( .A1(n9564), .A2(n9563), .A3(n9562), .ZN(n9565) );
  NAND3_X1 U10873 ( .A1(n9632), .A2(n9584), .A3(n9565), .ZN(n9575) );
  INV_X1 U10874 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9567) );
  OAI21_X1 U10875 ( .B1(n9643), .B2(n9567), .A(n9566), .ZN(n9568) );
  AOI21_X1 U10876 ( .B1(n9636), .B2(n9569), .A(n9568), .ZN(n9574) );
  OAI211_X1 U10877 ( .C1(n9572), .C2(n9571), .A(n9638), .B(n9570), .ZN(n9573)
         );
  NAND3_X1 U10878 ( .A1(n9575), .A2(n9574), .A3(n9573), .ZN(P1_U3248) );
  AND2_X1 U10879 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9578) );
  NOR2_X1 U10880 ( .A1(n9592), .A2(n9576), .ZN(n9577) );
  AOI211_X1 U10881 ( .C1(n10038), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9578), .B(
        n9577), .ZN(n9589) );
  OAI211_X1 U10882 ( .C1(n9581), .C2(n9580), .A(n9638), .B(n9579), .ZN(n9588)
         );
  INV_X1 U10883 ( .A(n9604), .ZN(n9586) );
  NAND3_X1 U10884 ( .A1(n9584), .A2(n9583), .A3(n9582), .ZN(n9585) );
  NAND3_X1 U10885 ( .A1(n9632), .A2(n9586), .A3(n9585), .ZN(n9587) );
  NAND3_X1 U10886 ( .A1(n9589), .A2(n9588), .A3(n9587), .ZN(P1_U3249) );
  INV_X1 U10887 ( .A(n9590), .ZN(n9594) );
  NOR2_X1 U10888 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  AOI211_X1 U10889 ( .C1(n10038), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n9594), .B(
        n9593), .ZN(n9607) );
  OAI211_X1 U10890 ( .C1(n9597), .C2(n9596), .A(n9638), .B(n9595), .ZN(n9606)
         );
  MUX2_X1 U10891 ( .A(n6933), .B(P1_REG1_REG_7__SCAN_IN), .S(n9598), .Z(n9601)
         );
  INV_X1 U10892 ( .A(n9599), .ZN(n9600) );
  NAND2_X1 U10893 ( .A1(n9601), .A2(n9600), .ZN(n9603) );
  OAI211_X1 U10894 ( .C1(n9604), .C2(n9603), .A(n9632), .B(n9602), .ZN(n9605)
         );
  NAND3_X1 U10895 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(P1_U3250) );
  NOR2_X1 U10896 ( .A1(n9614), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9609) );
  XNOR2_X1 U10897 ( .A(n9627), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9608) );
  NOR3_X1 U10898 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(n9625) );
  INV_X1 U10899 ( .A(n9625), .ZN(n9612) );
  OAI21_X1 U10900 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9611) );
  NAND3_X1 U10901 ( .A1(n9612), .A2(n9632), .A3(n9611), .ZN(n9624) );
  NOR2_X1 U10902 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5570), .ZN(n9613) );
  AOI21_X1 U10903 ( .B1(n10038), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9613), .ZN(
        n9623) );
  OR2_X1 U10904 ( .A1(n9614), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U10905 ( .A1(n9616), .A2(n9615), .ZN(n9619) );
  MUX2_X1 U10906 ( .A(n9617), .B(P1_REG2_REG_18__SCAN_IN), .S(n9627), .Z(n9618) );
  NAND2_X1 U10907 ( .A1(n9619), .A2(n9618), .ZN(n9620) );
  NAND3_X1 U10908 ( .A1(n9629), .A2(n9638), .A3(n9620), .ZN(n9622) );
  NAND2_X1 U10909 ( .A1(n9636), .A2(n9627), .ZN(n9621) );
  NAND4_X1 U10910 ( .A1(n9624), .A2(n9623), .A3(n9622), .A4(n9621), .ZN(
        P1_U3261) );
  INV_X1 U10911 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9644) );
  XNOR2_X1 U10912 ( .A(n9626), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U10913 ( .A1(n9627), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U10914 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  XNOR2_X1 U10915 ( .A(n9630), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9637) );
  INV_X1 U10916 ( .A(n9637), .ZN(n9631) );
  AOI22_X1 U10917 ( .A1(n9634), .A2(n9632), .B1(n9638), .B2(n9631), .ZN(n9640)
         );
  NOR2_X1 U10918 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  AOI211_X1 U10919 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9639)
         );
  MUX2_X1 U10920 ( .A(n9640), .B(n9639), .S(n5780), .Z(n9642) );
  OAI211_X1 U10921 ( .C1(n9644), .C2(n9643), .A(n9642), .B(n9641), .ZN(
        P1_U3262) );
  NAND2_X1 U10922 ( .A1(n9646), .A2(n9645), .ZN(n9649) );
  INV_X1 U10923 ( .A(n9895), .ZN(n9647) );
  NOR2_X1 U10924 ( .A1(n10063), .A2(n9647), .ZN(n9655) );
  AOI21_X1 U10925 ( .B1(n10063), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9655), .ZN(
        n9648) );
  OAI211_X1 U10926 ( .C1(n9650), .C2(n9891), .A(n9649), .B(n9648), .ZN(
        P1_U3263) );
  INV_X1 U10927 ( .A(n9652), .ZN(n9653) );
  NAND2_X1 U10928 ( .A1(n9896), .A2(n10057), .ZN(n9657) );
  AOI21_X1 U10929 ( .B1(n10063), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9655), .ZN(
        n9656) );
  OAI211_X1 U10930 ( .C1(n9972), .C2(n9891), .A(n9657), .B(n9656), .ZN(
        P1_U3264) );
  AOI21_X1 U10931 ( .B1(n9660), .B2(n10052), .A(n9659), .ZN(n9672) );
  XNOR2_X1 U10932 ( .A(n9664), .B(n9663), .ZN(n9670) );
  AOI22_X1 U10933 ( .A1(n9665), .A2(n10054), .B1(n10063), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9666) );
  OAI21_X1 U10934 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9669) );
  AOI21_X1 U10935 ( .B1(n9670), .B2(n10049), .A(n9669), .ZN(n9671) );
  OAI21_X1 U10936 ( .B1(n9672), .B2(n10063), .A(n9671), .ZN(P1_U3356) );
  NAND2_X1 U10937 ( .A1(n9673), .A2(n10049), .ZN(n9681) );
  INV_X1 U10938 ( .A(n9674), .ZN(n9679) );
  AOI22_X1 U10939 ( .A1(n9675), .A2(n10052), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10063), .ZN(n9676) );
  OAI21_X1 U10940 ( .B1(n9677), .B2(n9891), .A(n9676), .ZN(n9678) );
  AOI21_X1 U10941 ( .B1(n9679), .B2(n10057), .A(n9678), .ZN(n9680) );
  OAI211_X1 U10942 ( .C1(n9682), .C2(n10063), .A(n9681), .B(n9680), .ZN(
        P1_U3265) );
  XNOR2_X1 U10943 ( .A(n9683), .B(n9686), .ZN(n9684) );
  INV_X1 U10944 ( .A(n9899), .ZN(n9696) );
  XNOR2_X1 U10945 ( .A(n9687), .B(n9686), .ZN(n9901) );
  NAND2_X1 U10946 ( .A1(n9901), .A2(n10049), .ZN(n9695) );
  AOI211_X1 U10947 ( .C1(n9690), .C2(n9688), .A(n9885), .B(n5127), .ZN(n9900)
         );
  AOI22_X1 U10948 ( .A1(n9691), .A2(n10052), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10063), .ZN(n9692) );
  OAI21_X1 U10949 ( .B1(n9975), .B2(n9891), .A(n9692), .ZN(n9693) );
  AOI21_X1 U10950 ( .B1(n9900), .B2(n10057), .A(n9693), .ZN(n9694) );
  OAI211_X1 U10951 ( .C1(n9696), .C2(n10063), .A(n9695), .B(n9694), .ZN(
        P1_U3266) );
  NAND2_X1 U10952 ( .A1(n9697), .A2(n9698), .ZN(n9699) );
  XNOR2_X1 U10953 ( .A(n9699), .B(n9704), .ZN(n9700) );
  NAND2_X1 U10954 ( .A1(n9700), .A2(n9878), .ZN(n9702) );
  NAND2_X1 U10955 ( .A1(n9702), .A2(n9701), .ZN(n9902) );
  INV_X1 U10956 ( .A(n9902), .ZN(n9712) );
  XOR2_X1 U10957 ( .A(n9704), .B(n9703), .Z(n9904) );
  NAND2_X1 U10958 ( .A1(n9904), .A2(n10049), .ZN(n9711) );
  INV_X1 U10959 ( .A(n9720), .ZN(n9705) );
  AOI211_X1 U10960 ( .C1(n9706), .C2(n9705), .A(n9885), .B(n5131), .ZN(n9903)
         );
  AOI22_X1 U10961 ( .A1(n9707), .A2(n10052), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10063), .ZN(n9708) );
  OAI21_X1 U10962 ( .B1(n9979), .B2(n9891), .A(n9708), .ZN(n9709) );
  AOI21_X1 U10963 ( .B1(n9903), .B2(n10057), .A(n9709), .ZN(n9710) );
  OAI211_X1 U10964 ( .C1(n10063), .C2(n9712), .A(n9711), .B(n9710), .ZN(
        P1_U3267) );
  OAI211_X1 U10965 ( .C1(n9717), .C2(n9713), .A(n9697), .B(n9878), .ZN(n9716)
         );
  INV_X1 U10966 ( .A(n9714), .ZN(n9715) );
  NAND2_X1 U10967 ( .A1(n9716), .A2(n9715), .ZN(n9906) );
  INV_X1 U10968 ( .A(n9906), .ZN(n9727) );
  XOR2_X1 U10969 ( .A(n9718), .B(n9717), .Z(n9908) );
  NAND2_X1 U10970 ( .A1(n9908), .A2(n10049), .ZN(n9726) );
  OAI21_X1 U10971 ( .B1(n9719), .B2(n9983), .A(n9843), .ZN(n9721) );
  NOR2_X1 U10972 ( .A1(n9721), .A2(n9720), .ZN(n9907) );
  AOI22_X1 U10973 ( .A1(n9722), .A2(n10052), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10063), .ZN(n9723) );
  OAI21_X1 U10974 ( .B1(n9983), .B2(n9891), .A(n9723), .ZN(n9724) );
  AOI21_X1 U10975 ( .B1(n9907), .B2(n10057), .A(n9724), .ZN(n9725) );
  OAI211_X1 U10976 ( .C1(n10063), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        P1_U3268) );
  NAND2_X1 U10977 ( .A1(n9728), .A2(n9729), .ZN(n9730) );
  NAND3_X1 U10978 ( .A1(n9731), .A2(n9878), .A3(n9730), .ZN(n9733) );
  NAND2_X1 U10979 ( .A1(n9733), .A2(n9732), .ZN(n9911) );
  INV_X1 U10980 ( .A(n9911), .ZN(n9742) );
  XNOR2_X1 U10981 ( .A(n9734), .B(n5817), .ZN(n9913) );
  NAND2_X1 U10982 ( .A1(n9913), .A2(n10049), .ZN(n9741) );
  AOI211_X1 U10983 ( .C1(n9736), .C2(n9735), .A(n9885), .B(n9719), .ZN(n9912)
         );
  AOI22_X1 U10984 ( .A1(n9737), .A2(n10052), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10063), .ZN(n9738) );
  OAI21_X1 U10985 ( .B1(n9987), .B2(n9891), .A(n9738), .ZN(n9739) );
  AOI21_X1 U10986 ( .B1(n9912), .B2(n10057), .A(n9739), .ZN(n9740) );
  OAI211_X1 U10987 ( .C1(n10063), .C2(n9742), .A(n9741), .B(n9740), .ZN(
        P1_U3269) );
  NAND2_X1 U10988 ( .A1(n9743), .A2(n9744), .ZN(n9745) );
  XNOR2_X1 U10989 ( .A(n9745), .B(n9749), .ZN(n9746) );
  NAND2_X1 U10990 ( .A1(n9746), .A2(n9878), .ZN(n9748) );
  NAND2_X1 U10991 ( .A1(n9748), .A2(n9747), .ZN(n9916) );
  INV_X1 U10992 ( .A(n9916), .ZN(n9758) );
  XNOR2_X1 U10993 ( .A(n9750), .B(n9749), .ZN(n9918) );
  NAND2_X1 U10994 ( .A1(n9918), .A2(n10049), .ZN(n9757) );
  AOI21_X1 U10995 ( .B1(n4536), .B2(n9752), .A(n9885), .ZN(n9751) );
  AND2_X1 U10996 ( .A1(n9751), .A2(n9735), .ZN(n9915) );
  INV_X1 U10997 ( .A(n9752), .ZN(n9991) );
  AOI22_X1 U10998 ( .A1(n9753), .A2(n10052), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10063), .ZN(n9754) );
  OAI21_X1 U10999 ( .B1(n9991), .B2(n9891), .A(n9754), .ZN(n9755) );
  AOI21_X1 U11000 ( .B1(n9915), .B2(n10057), .A(n9755), .ZN(n9756) );
  OAI211_X1 U11001 ( .C1(n10063), .C2(n9758), .A(n9757), .B(n9756), .ZN(
        P1_U3270) );
  XNOR2_X1 U11002 ( .A(n9759), .B(n5814), .ZN(n9923) );
  INV_X1 U11003 ( .A(n9923), .ZN(n9769) );
  OAI211_X1 U11004 ( .C1(n9760), .C2(n5814), .A(n9743), .B(n9878), .ZN(n9762)
         );
  NAND2_X1 U11005 ( .A1(n9762), .A2(n9761), .ZN(n9921) );
  OR2_X1 U11006 ( .A1(n9778), .A2(n9995), .ZN(n9763) );
  AND3_X1 U11007 ( .A1(n4536), .A2(n9763), .A3(n9843), .ZN(n9922) );
  NAND2_X1 U11008 ( .A1(n9922), .A2(n10057), .ZN(n9766) );
  AOI22_X1 U11009 ( .A1(n9764), .A2(n10052), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10063), .ZN(n9765) );
  OAI211_X1 U11010 ( .C1(n9995), .C2(n9891), .A(n9766), .B(n9765), .ZN(n9767)
         );
  AOI21_X1 U11011 ( .B1(n9921), .B2(n9850), .A(n9767), .ZN(n9768) );
  OAI21_X1 U11012 ( .B1(n9769), .B2(n9852), .A(n9768), .ZN(P1_U3271) );
  OAI21_X1 U11013 ( .B1(n9770), .B2(n9786), .A(n9771), .ZN(n9772) );
  XNOR2_X1 U11014 ( .A(n9772), .B(n9776), .ZN(n9774) );
  AOI21_X1 U11015 ( .B1(n9774), .B2(n9878), .A(n9773), .ZN(n9928) );
  XNOR2_X1 U11016 ( .A(n9775), .B(n9776), .ZN(n9926) );
  OAI21_X1 U11017 ( .B1(n9999), .B2(n9777), .A(n9843), .ZN(n9779) );
  OR2_X1 U11018 ( .A1(n9779), .A2(n9778), .ZN(n9927) );
  AOI22_X1 U11019 ( .A1(n9780), .A2(n10052), .B1(n10063), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U11020 ( .A1(n9781), .A2(n10054), .ZN(n9782) );
  OAI211_X1 U11021 ( .C1(n9927), .C2(n9814), .A(n9783), .B(n9782), .ZN(n9784)
         );
  AOI21_X1 U11022 ( .B1(n9926), .B2(n10049), .A(n9784), .ZN(n9785) );
  OAI21_X1 U11023 ( .B1(n10063), .B2(n9928), .A(n9785), .ZN(P1_U3272) );
  XNOR2_X1 U11024 ( .A(n9770), .B(n9786), .ZN(n9788) );
  OAI21_X1 U11025 ( .B1(n9788), .B2(n9858), .A(n9787), .ZN(n9932) );
  INV_X1 U11026 ( .A(n9932), .ZN(n9800) );
  XNOR2_X1 U11027 ( .A(n9790), .B(n9789), .ZN(n9934) );
  NAND2_X1 U11028 ( .A1(n4473), .A2(n9791), .ZN(n9792) );
  NAND2_X1 U11029 ( .A1(n9792), .A2(n9843), .ZN(n9793) );
  NOR2_X1 U11030 ( .A1(n9777), .A2(n9793), .ZN(n9933) );
  NAND2_X1 U11031 ( .A1(n9933), .A2(n10057), .ZN(n9797) );
  INV_X1 U11032 ( .A(n9794), .ZN(n9795) );
  AOI22_X1 U11033 ( .A1(n10063), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9795), 
        .B2(n10052), .ZN(n9796) );
  OAI211_X1 U11034 ( .C1(n10003), .C2(n9891), .A(n9797), .B(n9796), .ZN(n9798)
         );
  AOI21_X1 U11035 ( .B1(n9934), .B2(n10049), .A(n9798), .ZN(n9799) );
  OAI21_X1 U11036 ( .B1(n9800), .B2(n10063), .A(n9799), .ZN(P1_U3273) );
  XNOR2_X1 U11037 ( .A(n9801), .B(n9804), .ZN(n9938) );
  OAI21_X1 U11038 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9807) );
  INV_X1 U11039 ( .A(n9805), .ZN(n9806) );
  AOI21_X1 U11040 ( .B1(n9807), .B2(n9878), .A(n9806), .ZN(n9937) );
  INV_X1 U11041 ( .A(n9937), .ZN(n9816) );
  AOI21_X1 U11042 ( .B1(n9808), .B2(n10006), .A(n9885), .ZN(n9809) );
  NAND2_X1 U11043 ( .A1(n9809), .A2(n4473), .ZN(n9936) );
  NAND2_X1 U11044 ( .A1(n10063), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9810) );
  OAI21_X1 U11045 ( .B1(n9829), .B2(n9811), .A(n9810), .ZN(n9812) );
  AOI21_X1 U11046 ( .B1(n10006), .B2(n10054), .A(n9812), .ZN(n9813) );
  OAI21_X1 U11047 ( .B1(n9936), .B2(n9814), .A(n9813), .ZN(n9815) );
  AOI21_X1 U11048 ( .B1(n9816), .B2(n9850), .A(n9815), .ZN(n9817) );
  OAI21_X1 U11049 ( .B1(n9852), .B2(n9938), .A(n9817), .ZN(P1_U3274) );
  XNOR2_X1 U11050 ( .A(n9818), .B(n9820), .ZN(n9946) );
  INV_X1 U11051 ( .A(n9819), .ZN(n9822) );
  OAI21_X1 U11052 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9824) );
  AOI21_X1 U11053 ( .B1(n9824), .B2(n9823), .A(n9858), .ZN(n9826) );
  NOR2_X1 U11054 ( .A1(n9826), .A2(n9825), .ZN(n9945) );
  NAND2_X1 U11055 ( .A1(n10063), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9827) );
  OAI21_X1 U11056 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(n9830) );
  AOI21_X1 U11057 ( .B1(n9943), .B2(n10054), .A(n9830), .ZN(n9834) );
  OR2_X1 U11058 ( .A1(n4556), .A2(n9831), .ZN(n9832) );
  AND3_X1 U11059 ( .A1(n9808), .A2(n9843), .A3(n9832), .ZN(n9942) );
  NAND2_X1 U11060 ( .A1(n9942), .A2(n10057), .ZN(n9833) );
  OAI211_X1 U11061 ( .C1(n9945), .C2(n10063), .A(n9834), .B(n9833), .ZN(n9835)
         );
  INV_X1 U11062 ( .A(n9835), .ZN(n9836) );
  OAI21_X1 U11063 ( .B1(n9852), .B2(n9946), .A(n9836), .ZN(P1_U3275) );
  XOR2_X1 U11064 ( .A(n9837), .B(n9838), .Z(n9949) );
  INV_X1 U11065 ( .A(n9949), .ZN(n9853) );
  OAI211_X1 U11066 ( .C1(n9839), .C2(n5808), .A(n9878), .B(n9819), .ZN(n9841)
         );
  NAND2_X1 U11067 ( .A1(n9841), .A2(n9840), .ZN(n9947) );
  INV_X1 U11068 ( .A(n9842), .ZN(n10011) );
  NAND2_X1 U11069 ( .A1(n9865), .A2(n9842), .ZN(n9844) );
  NAND2_X1 U11070 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  NOR2_X1 U11071 ( .A1(n4556), .A2(n9845), .ZN(n9948) );
  NAND2_X1 U11072 ( .A1(n9948), .A2(n10057), .ZN(n9848) );
  AOI22_X1 U11073 ( .A1(n10063), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9846), 
        .B2(n10052), .ZN(n9847) );
  OAI211_X1 U11074 ( .C1(n10011), .C2(n9891), .A(n9848), .B(n9847), .ZN(n9849)
         );
  AOI21_X1 U11075 ( .B1(n9947), .B2(n9850), .A(n9849), .ZN(n9851) );
  OAI21_X1 U11076 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(P1_U3276) );
  XNOR2_X1 U11077 ( .A(n9854), .B(n9855), .ZN(n9859) );
  INV_X1 U11078 ( .A(n9856), .ZN(n9857) );
  OAI21_X1 U11079 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9951) );
  INV_X1 U11080 ( .A(n9951), .ZN(n9873) );
  INV_X1 U11081 ( .A(n9860), .ZN(n9861) );
  AOI21_X1 U11082 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(n9953) );
  INV_X1 U11083 ( .A(n9865), .ZN(n9866) );
  AOI211_X1 U11084 ( .C1(n9867), .C2(n9864), .A(n9885), .B(n9866), .ZN(n9952)
         );
  NAND2_X1 U11085 ( .A1(n9952), .A2(n10057), .ZN(n9870) );
  AOI22_X1 U11086 ( .A1(n10063), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9868), 
        .B2(n10052), .ZN(n9869) );
  OAI211_X1 U11087 ( .C1(n5126), .C2(n9891), .A(n9870), .B(n9869), .ZN(n9871)
         );
  AOI21_X1 U11088 ( .B1(n9953), .B2(n10049), .A(n9871), .ZN(n9872) );
  OAI21_X1 U11089 ( .B1(n10063), .B2(n9873), .A(n9872), .ZN(P1_U3277) );
  NAND2_X1 U11090 ( .A1(n8010), .A2(n9874), .ZN(n9875) );
  NAND2_X1 U11091 ( .A1(n9875), .A2(n9884), .ZN(n9877) );
  NAND2_X1 U11092 ( .A1(n9877), .A2(n9876), .ZN(n9879) );
  NAND2_X1 U11093 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  INV_X1 U11094 ( .A(n9880), .ZN(n9881) );
  NAND2_X1 U11095 ( .A1(n9882), .A2(n9881), .ZN(n9959) );
  INV_X1 U11096 ( .A(n9959), .ZN(n9894) );
  XNOR2_X1 U11097 ( .A(n9883), .B(n9884), .ZN(n9956) );
  AOI21_X1 U11098 ( .B1(n8017), .B2(n9886), .A(n9885), .ZN(n9887) );
  AND2_X1 U11099 ( .A1(n9887), .A2(n9864), .ZN(n9957) );
  NAND2_X1 U11100 ( .A1(n9957), .A2(n10057), .ZN(n9890) );
  AOI22_X1 U11101 ( .A1(n10063), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9888), 
        .B2(n10052), .ZN(n9889) );
  OAI211_X1 U11102 ( .C1(n10018), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9892)
         );
  AOI21_X1 U11103 ( .B1(n9956), .B2(n10049), .A(n9892), .ZN(n9893) );
  OAI21_X1 U11104 ( .B1(n9894), .B2(n10063), .A(n9893), .ZN(P1_U3278) );
  INV_X1 U11105 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9897) );
  MUX2_X1 U11106 ( .A(n9897), .B(n9969), .S(n10077), .Z(n9898) );
  OAI21_X1 U11107 ( .B1(n9972), .B2(n9961), .A(n9898), .ZN(P1_U3552) );
  AOI211_X1 U11108 ( .C1(n9904), .C2(n10071), .A(n9903), .B(n9902), .ZN(n9976)
         );
  MUX2_X1 U11109 ( .A(n10437), .B(n9976), .S(n10077), .Z(n9905) );
  OAI21_X1 U11110 ( .B1(n9979), .B2(n9961), .A(n9905), .ZN(P1_U3548) );
  AOI211_X1 U11111 ( .C1(n9908), .C2(n10071), .A(n9907), .B(n9906), .ZN(n9980)
         );
  MUX2_X1 U11112 ( .A(n9909), .B(n9980), .S(n10077), .Z(n9910) );
  OAI21_X1 U11113 ( .B1(n9983), .B2(n9961), .A(n9910), .ZN(P1_U3547) );
  AOI211_X1 U11114 ( .C1(n9913), .C2(n10071), .A(n9912), .B(n9911), .ZN(n9984)
         );
  MUX2_X1 U11115 ( .A(n10341), .B(n9984), .S(n10077), .Z(n9914) );
  OAI21_X1 U11116 ( .B1(n9987), .B2(n9961), .A(n9914), .ZN(P1_U3546) );
  OR2_X1 U11117 ( .A1(n9916), .A2(n9915), .ZN(n9917) );
  AOI21_X1 U11118 ( .B1(n9918), .B2(n10071), .A(n9917), .ZN(n9988) );
  MUX2_X1 U11119 ( .A(n9919), .B(n9988), .S(n10077), .Z(n9920) );
  OAI21_X1 U11120 ( .B1(n9991), .B2(n9961), .A(n9920), .ZN(P1_U3545) );
  AOI211_X1 U11121 ( .C1(n9923), .C2(n10071), .A(n9922), .B(n9921), .ZN(n9992)
         );
  MUX2_X1 U11122 ( .A(n9924), .B(n9992), .S(n10077), .Z(n9925) );
  OAI21_X1 U11123 ( .B1(n9995), .B2(n9961), .A(n9925), .ZN(P1_U3544) );
  NAND2_X1 U11124 ( .A1(n9926), .A2(n10071), .ZN(n9929) );
  AND3_X1 U11125 ( .A1(n9929), .A2(n9928), .A3(n9927), .ZN(n9996) );
  MUX2_X1 U11126 ( .A(n9930), .B(n9996), .S(n10077), .Z(n9931) );
  OAI21_X1 U11127 ( .B1(n9999), .B2(n9961), .A(n9931), .ZN(P1_U3543) );
  INV_X1 U11128 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10483) );
  AOI211_X1 U11129 ( .C1(n9934), .C2(n10071), .A(n9933), .B(n9932), .ZN(n10000) );
  MUX2_X1 U11130 ( .A(n10483), .B(n10000), .S(n10077), .Z(n9935) );
  OAI21_X1 U11131 ( .B1(n10003), .B2(n9961), .A(n9935), .ZN(P1_U3542) );
  OAI211_X1 U11132 ( .C1(n9938), .C2(n9968), .A(n9937), .B(n9936), .ZN(n10004)
         );
  MUX2_X1 U11133 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10004), .S(n10077), .Z(
        n9939) );
  AOI21_X1 U11134 ( .B1(n9940), .B2(n10006), .A(n9939), .ZN(n9941) );
  INV_X1 U11135 ( .A(n9941), .ZN(P1_U3541) );
  AOI21_X1 U11136 ( .B1(n9964), .B2(n9943), .A(n9942), .ZN(n9944) );
  OAI211_X1 U11137 ( .C1(n9968), .C2(n9946), .A(n9945), .B(n9944), .ZN(n10008)
         );
  MUX2_X1 U11138 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10008), .S(n10077), .Z(
        P1_U3540) );
  INV_X1 U11139 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10426) );
  AOI211_X1 U11140 ( .C1(n9949), .C2(n10071), .A(n9948), .B(n9947), .ZN(n10009) );
  MUX2_X1 U11141 ( .A(n10426), .B(n10009), .S(n10077), .Z(n9950) );
  OAI21_X1 U11142 ( .B1(n10011), .B2(n9961), .A(n9950), .ZN(P1_U3539) );
  AOI211_X1 U11143 ( .C1(n9953), .C2(n10071), .A(n9952), .B(n9951), .ZN(n10012) );
  MUX2_X1 U11144 ( .A(n9954), .B(n10012), .S(n10077), .Z(n9955) );
  OAI21_X1 U11145 ( .B1(n5126), .B2(n9961), .A(n9955), .ZN(P1_U3538) );
  AND2_X1 U11146 ( .A1(n9956), .A2(n10071), .ZN(n9958) );
  NOR3_X1 U11147 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n10015) );
  MUX2_X1 U11148 ( .A(n10015), .B(n10353), .S(n4655), .Z(n9960) );
  OAI21_X1 U11149 ( .B1(n10018), .B2(n9961), .A(n9960), .ZN(P1_U3537) );
  AOI21_X1 U11150 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9965) );
  OAI211_X1 U11151 ( .C1(n9968), .C2(n9967), .A(n9966), .B(n9965), .ZN(n10019)
         );
  MUX2_X1 U11152 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10019), .S(n10077), .Z(
        P1_U3536) );
  INV_X1 U11153 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U11154 ( .A(n9970), .B(n9969), .S(n10074), .Z(n9971) );
  OAI21_X1 U11155 ( .B1(n9972), .B2(n10017), .A(n9971), .ZN(P1_U3520) );
  OAI21_X1 U11156 ( .B1(n9975), .B2(n10017), .A(n9974), .ZN(P1_U3517) );
  INV_X1 U11157 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9977) );
  MUX2_X1 U11158 ( .A(n9977), .B(n9976), .S(n10074), .Z(n9978) );
  OAI21_X1 U11159 ( .B1(n9979), .B2(n10017), .A(n9978), .ZN(P1_U3516) );
  INV_X1 U11160 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9981) );
  MUX2_X1 U11161 ( .A(n9981), .B(n9980), .S(n10074), .Z(n9982) );
  OAI21_X1 U11162 ( .B1(n9983), .B2(n10017), .A(n9982), .ZN(P1_U3515) );
  INV_X1 U11163 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9985) );
  MUX2_X1 U11164 ( .A(n9985), .B(n9984), .S(n10074), .Z(n9986) );
  OAI21_X1 U11165 ( .B1(n9987), .B2(n10017), .A(n9986), .ZN(P1_U3514) );
  INV_X1 U11166 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9989) );
  MUX2_X1 U11167 ( .A(n9989), .B(n9988), .S(n10074), .Z(n9990) );
  OAI21_X1 U11168 ( .B1(n9991), .B2(n10017), .A(n9990), .ZN(P1_U3513) );
  INV_X1 U11169 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9993) );
  MUX2_X1 U11170 ( .A(n9993), .B(n9992), .S(n10074), .Z(n9994) );
  OAI21_X1 U11171 ( .B1(n9995), .B2(n10017), .A(n9994), .ZN(P1_U3512) );
  INV_X1 U11172 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9997) );
  MUX2_X1 U11173 ( .A(n9997), .B(n9996), .S(n10074), .Z(n9998) );
  OAI21_X1 U11174 ( .B1(n9999), .B2(n10017), .A(n9998), .ZN(P1_U3511) );
  INV_X1 U11175 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10001) );
  MUX2_X1 U11176 ( .A(n10001), .B(n10000), .S(n10074), .Z(n10002) );
  OAI21_X1 U11177 ( .B1(n10003), .B2(n10017), .A(n10002), .ZN(P1_U3510) );
  MUX2_X1 U11178 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10004), .S(n10074), .Z(
        n10005) );
  AOI21_X1 U11179 ( .B1(n6861), .B2(n10006), .A(n10005), .ZN(n10007) );
  INV_X1 U11180 ( .A(n10007), .ZN(P1_U3509) );
  MUX2_X1 U11181 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10008), .S(n10074), .Z(
        P1_U3507) );
  INV_X1 U11182 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10495) );
  MUX2_X1 U11183 ( .A(n10495), .B(n10009), .S(n10074), .Z(n10010) );
  OAI21_X1 U11184 ( .B1(n10011), .B2(n10017), .A(n10010), .ZN(P1_U3504) );
  INV_X1 U11185 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10013) );
  MUX2_X1 U11186 ( .A(n10013), .B(n10012), .S(n10074), .Z(n10014) );
  OAI21_X1 U11187 ( .B1(n5126), .B2(n10017), .A(n10014), .ZN(P1_U3501) );
  INV_X1 U11188 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10398) );
  MUX2_X1 U11189 ( .A(n10398), .B(n10015), .S(n10074), .Z(n10016) );
  OAI21_X1 U11190 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(P1_U3498) );
  MUX2_X1 U11191 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10019), .S(n10074), .Z(
        P1_U3495) );
  MUX2_X1 U11192 ( .A(P1_D_REG_0__SCAN_IN), .B(n10021), .S(n10020), .Z(
        P1_U3439) );
  NOR4_X1 U11193 ( .A1(n4809), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10022), .A4(
        P1_U3086), .ZN(n10023) );
  AOI21_X1 U11194 ( .B1(n10024), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10023), 
        .ZN(n10025) );
  OAI21_X1 U11195 ( .B1(n10026), .B2(n10029), .A(n10025), .ZN(P1_U3324) );
  OAI222_X1 U11196 ( .A1(n8378), .A2(n10287), .B1(n10029), .B2(n10028), .C1(
        n10027), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U11197 ( .A(n10030), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11198 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X1 U11199 ( .A1(n10031), .A2(n6127), .ZN(n10034) );
  NOR2_X1 U11200 ( .A1(n10032), .A2(n10034), .ZN(n10033) );
  MUX2_X1 U11201 ( .A(n10034), .B(n10033), .S(P1_IR_REG_0__SCAN_IN), .Z(n10037) );
  INV_X1 U11202 ( .A(n10035), .ZN(n10036) );
  OR2_X1 U11203 ( .A1(n10037), .A2(n10036), .ZN(n10040) );
  AOI22_X1 U11204 ( .A1(n10038), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10039) );
  OAI21_X1 U11205 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(P1_U3243) );
  NAND2_X1 U11206 ( .A1(n10042), .A2(n10057), .ZN(n10045) );
  AOI22_X1 U11207 ( .A1(n10063), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10052), 
        .B2(n10043), .ZN(n10044) );
  OAI211_X1 U11208 ( .C1(n10046), .C2(n9891), .A(n10045), .B(n10044), .ZN(
        n10047) );
  AOI21_X1 U11209 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n10050) );
  OAI21_X1 U11210 ( .B1(n10063), .B2(n10051), .A(n10050), .ZN(P1_U3290) );
  AOI22_X1 U11211 ( .A1(n10052), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n10063), .ZN(n10061) );
  INV_X1 U11212 ( .A(n10053), .ZN(n10058) );
  AOI222_X1 U11213 ( .A1(n10059), .A2(n10058), .B1(n10057), .B2(n10056), .C1(
        n10055), .C2(n10054), .ZN(n10060) );
  OAI211_X1 U11214 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        P1_U3292) );
  INV_X1 U11215 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10352) );
  NOR2_X1 U11216 ( .A1(n10064), .A2(n10352), .ZN(P1_U3294) );
  AND2_X1 U11217 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10223), .ZN(P1_U3295) );
  AND2_X1 U11218 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10223), .ZN(P1_U3296) );
  AND2_X1 U11219 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10223), .ZN(P1_U3297) );
  AND2_X1 U11220 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10223), .ZN(P1_U3298) );
  AND2_X1 U11221 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10223), .ZN(P1_U3299) );
  AND2_X1 U11222 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10223), .ZN(P1_U3300) );
  AND2_X1 U11223 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10223), .ZN(P1_U3301) );
  AND2_X1 U11224 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10223), .ZN(P1_U3302) );
  AND2_X1 U11225 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10223), .ZN(P1_U3303) );
  AND2_X1 U11226 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10223), .ZN(P1_U3304) );
  AND2_X1 U11227 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10223), .ZN(P1_U3305) );
  AND2_X1 U11228 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10223), .ZN(P1_U3306) );
  AND2_X1 U11229 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10223), .ZN(P1_U3307) );
  AND2_X1 U11230 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10223), .ZN(P1_U3308) );
  INV_X1 U11231 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U11232 ( .A1(n10064), .A2(n10397), .ZN(P1_U3309) );
  AND2_X1 U11233 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10223), .ZN(P1_U3310) );
  AND2_X1 U11234 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10223), .ZN(P1_U3312) );
  INV_X1 U11235 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10484) );
  NOR2_X1 U11236 ( .A1(n10064), .A2(n10484), .ZN(P1_U3313) );
  AND2_X1 U11237 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10223), .ZN(P1_U3314) );
  AND2_X1 U11238 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10223), .ZN(P1_U3315) );
  AND2_X1 U11239 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10223), .ZN(P1_U3316) );
  INV_X1 U11240 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10480) );
  NOR2_X1 U11241 ( .A1(n10064), .A2(n10480), .ZN(P1_U3317) );
  AND2_X1 U11242 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10223), .ZN(P1_U3318) );
  AND2_X1 U11243 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10223), .ZN(P1_U3319) );
  INV_X1 U11244 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10326) );
  NOR2_X1 U11245 ( .A1(n10064), .A2(n10326), .ZN(P1_U3320) );
  AND2_X1 U11246 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10223), .ZN(P1_U3321) );
  AND2_X1 U11247 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10223), .ZN(P1_U3322) );
  AND2_X1 U11248 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10223), .ZN(P1_U3323) );
  OAI21_X1 U11249 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10069) );
  AOI211_X1 U11250 ( .C1(n10071), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10076) );
  INV_X1 U11251 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11252 ( .A1(n10074), .A2(n10076), .B1(n10073), .B2(n10072), .ZN(
        P1_U3465) );
  AOI22_X1 U11253 ( .A1(n10077), .A2(n10076), .B1(n10075), .B2(n4655), .ZN(
        P1_U3526) );
  OAI21_X1 U11254 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10091) );
  AOI21_X1 U11255 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10089) );
  NAND2_X1 U11256 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  OAI211_X1 U11257 ( .C1(n10089), .C2(n10088), .A(n10087), .B(n10086), .ZN(
        n10090) );
  AOI21_X1 U11258 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10101) );
  NAND2_X1 U11259 ( .A1(n10094), .A2(n10093), .ZN(n10096) );
  AOI21_X1 U11260 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10098) );
  AOI21_X1 U11261 ( .B1(n10099), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10098), .ZN(
        n10100) );
  NAND2_X1 U11262 ( .A1(n10101), .A2(n10100), .ZN(P2_U3188) );
  NAND2_X1 U11263 ( .A1(n4450), .A2(n10102), .ZN(n10104) );
  XOR2_X1 U11264 ( .A(n10106), .B(n10104), .Z(n10169) );
  XOR2_X1 U11265 ( .A(n10105), .B(n10106), .Z(n10107) );
  OAI222_X1 U11266 ( .A1(n10127), .A2(n10109), .B1(n10125), .B2(n10108), .C1(
        n10132), .C2(n10107), .ZN(n10171) );
  MUX2_X1 U11267 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10171), .S(n10141), .Z(
        n10113) );
  OAI22_X1 U11268 ( .A1(n10111), .A2(n10167), .B1(n10110), .B2(n10123), .ZN(
        n10112) );
  NOR2_X1 U11269 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  OAI21_X1 U11270 ( .B1(n10169), .B2(n10115), .A(n10114), .ZN(P2_U3227) );
  OAI21_X1 U11271 ( .B1(n4620), .B2(n10117), .A(n10116), .ZN(n10121) );
  INV_X1 U11272 ( .A(n10119), .ZN(n10130) );
  NAND2_X1 U11273 ( .A1(n10121), .A2(n10130), .ZN(n10120) );
  OAI21_X1 U11274 ( .B1(n10121), .B2(n10130), .A(n10120), .ZN(n10152) );
  OAI22_X1 U11275 ( .A1(n10123), .A2(n7184), .B1(n4567), .B2(n10122), .ZN(
        n10139) );
  INV_X1 U11276 ( .A(n10124), .ZN(n10137) );
  OAI22_X1 U11277 ( .A1(n10128), .A2(n10127), .B1(n10126), .B2(n10125), .ZN(
        n10136) );
  NAND3_X1 U11278 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(n10133) );
  AOI21_X1 U11279 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10135) );
  AOI211_X1 U11280 ( .C1(n10137), .C2(n10152), .A(n10136), .B(n10135), .ZN(
        n10154) );
  INV_X1 U11281 ( .A(n10154), .ZN(n10138) );
  AOI211_X1 U11282 ( .C1(n10140), .C2(n10152), .A(n10139), .B(n10138), .ZN(
        n10142) );
  AOI22_X1 U11283 ( .A1(n10144), .A2(n10143), .B1(n10142), .B2(n10141), .ZN(
        P2_U3231) );
  INV_X1 U11284 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10149) );
  INV_X1 U11285 ( .A(n10145), .ZN(n10148) );
  OAI21_X1 U11286 ( .B1(n7016), .B2(n10172), .A(n10146), .ZN(n10147) );
  AOI21_X1 U11287 ( .B1(n10162), .B2(n10148), .A(n10147), .ZN(n10181) );
  AOI22_X1 U11288 ( .A1(n10180), .A2(n10149), .B1(n10181), .B2(n10178), .ZN(
        P2_U3393) );
  INV_X1 U11289 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11290 ( .A1(n10152), .A2(n10151), .B1(n10161), .B2(n10150), .ZN(
        n10153) );
  AND2_X1 U11291 ( .A1(n10154), .A2(n10153), .ZN(n10182) );
  AOI22_X1 U11292 ( .A1(n10180), .A2(n10155), .B1(n10182), .B2(n10178), .ZN(
        P2_U3396) );
  INV_X1 U11293 ( .A(n10156), .ZN(n10160) );
  OAI22_X1 U11294 ( .A1(n10158), .A2(n10168), .B1(n10157), .B2(n10172), .ZN(
        n10159) );
  NOR2_X1 U11295 ( .A1(n10160), .A2(n10159), .ZN(n10183) );
  AOI22_X1 U11296 ( .A1(n10180), .A2(n6423), .B1(n10183), .B2(n10178), .ZN(
        P2_U3399) );
  INV_X1 U11297 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U11298 ( .A1(n10163), .A2(n10162), .B1(n10161), .B2(n6739), .ZN(
        n10164) );
  AND2_X1 U11299 ( .A1(n10165), .A2(n10164), .ZN(n10184) );
  AOI22_X1 U11300 ( .A1(n10180), .A2(n10166), .B1(n10184), .B2(n10178), .ZN(
        P2_U3405) );
  OAI22_X1 U11301 ( .A1(n10169), .A2(n10168), .B1(n10167), .B2(n10172), .ZN(
        n10170) );
  NOR2_X1 U11302 ( .A1(n10171), .A2(n10170), .ZN(n10186) );
  AOI22_X1 U11303 ( .A1(n10180), .A2(n6459), .B1(n10186), .B2(n10178), .ZN(
        P2_U3408) );
  INV_X1 U11304 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10179) );
  OAI22_X1 U11305 ( .A1(n10175), .A2(n10174), .B1(n10173), .B2(n10172), .ZN(
        n10176) );
  NOR2_X1 U11306 ( .A1(n10177), .A2(n10176), .ZN(n10188) );
  AOI22_X1 U11307 ( .A1(n10180), .A2(n10179), .B1(n10188), .B2(n10178), .ZN(
        P2_U3411) );
  AOI22_X1 U11308 ( .A1(n10189), .A2(n10181), .B1(n6394), .B2(n10187), .ZN(
        P2_U3460) );
  AOI22_X1 U11309 ( .A1(n10189), .A2(n10182), .B1(n6413), .B2(n10187), .ZN(
        P2_U3461) );
  AOI22_X1 U11310 ( .A1(n10189), .A2(n10183), .B1(n6425), .B2(n10187), .ZN(
        P2_U3462) );
  AOI22_X1 U11311 ( .A1(n10189), .A2(n10184), .B1(n6448), .B2(n10187), .ZN(
        P2_U3464) );
  INV_X1 U11312 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U11313 ( .A1(n10189), .A2(n10186), .B1(n10185), .B2(n10187), .ZN(
        P2_U3465) );
  AOI22_X1 U11314 ( .A1(n10189), .A2(n10188), .B1(n6471), .B2(n10187), .ZN(
        P2_U3466) );
  OAI222_X1 U11315 ( .A1(n10194), .A2(n10193), .B1(n10194), .B2(n10192), .C1(
        n10191), .C2(n10190), .ZN(ADD_1068_U5) );
  XOR2_X1 U11316 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11317 ( .B1(n10197), .B2(n10196), .A(n10195), .ZN(n10198) );
  XNOR2_X1 U11318 ( .A(n10198), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11319 ( .B1(n10201), .B2(n10200), .A(n10199), .ZN(ADD_1068_U56) );
  OAI21_X1 U11320 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(ADD_1068_U57) );
  OAI21_X1 U11321 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(ADD_1068_U58) );
  OAI21_X1 U11322 ( .B1(n10210), .B2(n10209), .A(n10208), .ZN(ADD_1068_U59) );
  OAI21_X1 U11323 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(ADD_1068_U60) );
  OAI21_X1 U11324 ( .B1(n10216), .B2(n10215), .A(n10214), .ZN(ADD_1068_U61) );
  OAI21_X1 U11325 ( .B1(n10219), .B2(n10218), .A(n10217), .ZN(ADD_1068_U62) );
  OAI21_X1 U11326 ( .B1(n10222), .B2(n10221), .A(n10220), .ZN(ADD_1068_U63) );
  NAND2_X1 U11327 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10223), .ZN(n10516) );
  INV_X1 U11328 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10224) );
  NOR3_X1 U11329 ( .A1(n10225), .A2(n10224), .A3(n9567), .ZN(n10227) );
  NAND4_X1 U11330 ( .A1(n10228), .A2(P1_IR_REG_7__SCAN_IN), .A3(n10227), .A4(
        n10226), .ZN(n10239) );
  NAND4_X1 U11331 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(P2_REG3_REG_1__SCAN_IN), 
        .A3(P1_REG3_REG_16__SCAN_IN), .A4(n10453), .ZN(n10238) );
  NAND4_X1 U11332 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), 
        .A3(P2_D_REG_12__SCAN_IN), .A4(P1_REG2_REG_3__SCAN_IN), .ZN(n10237) );
  INV_X1 U11333 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10229) );
  NAND4_X1 U11334 ( .A1(n10229), .A2(n10493), .A3(P1_B_REG_SCAN_IN), .A4(
        P1_REG3_REG_3__SCAN_IN), .ZN(n10235) );
  INV_X1 U11335 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10232) );
  NOR4_X1 U11336 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P1_REG1_REG_5__SCAN_IN), 
        .A3(P1_REG2_REG_5__SCAN_IN), .A4(n10472), .ZN(n10231) );
  NOR4_X1 U11337 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_REG0_REG_23__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(n10495), .ZN(n10230) );
  NAND4_X1 U11338 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(
        P2_IR_REG_30__SCAN_IN), .ZN(n10234) );
  INV_X1 U11339 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10233) );
  OR4_X1 U11340 ( .A1(n10235), .A2(n10234), .A3(P1_IR_REG_22__SCAN_IN), .A4(
        n10233), .ZN(n10236) );
  NOR4_X1 U11341 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10282) );
  NAND4_X1 U11342 ( .A1(n10285), .A2(n10288), .A3(n10284), .A4(n10426), .ZN(
        n10280) );
  INV_X1 U11343 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10427) );
  NAND4_X1 U11344 ( .A1(SI_17_), .A2(P1_REG0_REG_2__SCAN_IN), .A3(n10429), 
        .A4(n10427), .ZN(n10279) );
  NAND4_X1 U11345 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n10312), .A4(n6848), .ZN(n10240) );
  NOR3_X1 U11346 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .A3(n10240), .ZN(n10246) );
  NAND4_X1 U11347 ( .A1(n6813), .A2(n10292), .A3(n5608), .A4(
        P1_REG2_REG_4__SCAN_IN), .ZN(n10244) );
  NAND4_X1 U11348 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), .A3(n10303), .A4(n10302), .ZN(n10243) );
  NAND4_X1 U11349 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(P1_REG1_REG_9__SCAN_IN), .A4(P1_REG2_REG_6__SCAN_IN), .ZN(n10242)
         );
  NAND4_X1 U11350 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P1_DATAO_REG_4__SCAN_IN), 
        .A3(n10300), .A4(n10316), .ZN(n10241) );
  NOR4_X1 U11351 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  NAND4_X1 U11352 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10246), .A3(n10245), .A4(
        n6663), .ZN(n10278) );
  INV_X1 U11353 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10424) );
  INV_X1 U11354 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10422) );
  NAND4_X1 U11355 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_DATAO_REG_31__SCAN_IN), 
        .A3(n10424), .A4(n10422), .ZN(n10250) );
  NAND4_X1 U11356 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P1_REG0_REG_0__SCAN_IN), .A4(n10394), .ZN(n10249) );
  NAND4_X1 U11357 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), 
        .A3(n10400), .A4(n10398), .ZN(n10248) );
  NAND4_X1 U11358 ( .A1(n5056), .A2(n10437), .A3(P2_DATAO_REG_16__SCAN_IN), 
        .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n10247) );
  NOR4_X1 U11359 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10276) );
  NAND4_X1 U11360 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(P1_REG1_REG_20__SCAN_IN), .A3(n10487), .A4(n10410), .ZN(n10254) );
  NAND4_X1 U11361 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P2_REG1_REG_12__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10253) );
  INV_X1 U11362 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10401) );
  NAND4_X1 U11363 ( .A1(n10401), .A2(n8968), .A3(n8944), .A4(
        P2_REG1_REG_8__SCAN_IN), .ZN(n10252) );
  NAND4_X1 U11364 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(P2_DATAO_REG_2__SCAN_IN), 
        .A3(P1_REG2_REG_11__SCAN_IN), .A4(n6933), .ZN(n10251) );
  NOR4_X1 U11365 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10275) );
  INV_X1 U11366 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U11367 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n6684), .A3(n10255), .A4(
        n10366), .ZN(n10261) );
  NAND4_X1 U11368 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .A3(n10381), .A4(n10256), .ZN(n10259) );
  NAND4_X1 U11369 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(n6409), .A4(n10257), .ZN(n10258) );
  OR4_X1 U11370 ( .A1(n10371), .A2(n10259), .A3(n10258), .A4(
        P1_REG3_REG_18__SCAN_IN), .ZN(n10260) );
  NOR4_X1 U11371 ( .A1(n10261), .A2(n10260), .A3(P1_DATAO_REG_7__SCAN_IN), 
        .A4(P1_REG1_REG_19__SCAN_IN), .ZN(n10274) );
  INV_X1 U11372 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10262) );
  NAND4_X1 U11373 ( .A1(n10263), .A2(n10262), .A3(n10342), .A4(n6448), .ZN(
        n10272) );
  NAND4_X1 U11374 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(SI_11_), .ZN(
        n10271) );
  NAND4_X1 U11375 ( .A1(n10268), .A2(n10267), .A3(P2_REG0_REG_18__SCAN_IN), 
        .A4(P1_REG3_REG_14__SCAN_IN), .ZN(n10270) );
  NAND4_X1 U11376 ( .A1(n10353), .A2(P1_REG2_REG_8__SCAN_IN), .A3(
        P1_REG0_REG_9__SCAN_IN), .A4(P1_REG1_REG_24__SCAN_IN), .ZN(n10269) );
  NOR4_X1 U11377 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  NAND4_X1 U11378 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n10277) );
  NOR4_X1 U11379 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        n10281) );
  AOI21_X1 U11380 ( .B1(n10282), .B2(n10281), .A(P2_IR_REG_26__SCAN_IN), .ZN(
        n10514) );
  AOI22_X1 U11381 ( .A1(n10285), .A2(keyinput74), .B1(keyinput81), .B2(n10284), 
        .ZN(n10283) );
  OAI221_X1 U11382 ( .B1(n10285), .B2(keyinput74), .C1(n10284), .C2(keyinput81), .A(n10283), .ZN(n10297) );
  AOI22_X1 U11383 ( .A1(n10288), .A2(keyinput46), .B1(n10287), .B2(keyinput124), .ZN(n10286) );
  OAI221_X1 U11384 ( .B1(n10288), .B2(keyinput46), .C1(n10287), .C2(
        keyinput124), .A(n10286), .ZN(n10296) );
  INV_X1 U11385 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U11386 ( .A1(n10290), .A2(keyinput31), .B1(n5608), .B2(keyinput85), 
        .ZN(n10289) );
  OAI221_X1 U11387 ( .B1(n10290), .B2(keyinput31), .C1(n5608), .C2(keyinput85), 
        .A(n10289), .ZN(n10295) );
  AOI22_X1 U11388 ( .A1(n10293), .A2(keyinput82), .B1(n10292), .B2(keyinput116), .ZN(n10291) );
  OAI221_X1 U11389 ( .B1(n10293), .B2(keyinput82), .C1(n10292), .C2(
        keyinput116), .A(n10291), .ZN(n10294) );
  NOR4_X1 U11390 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10339) );
  AOI22_X1 U11391 ( .A1(n6813), .A2(keyinput99), .B1(keyinput26), .B2(n10224), 
        .ZN(n10298) );
  OAI221_X1 U11392 ( .B1(n6813), .B2(keyinput99), .C1(n10224), .C2(keyinput26), 
        .A(n10298), .ZN(n10310) );
  AOI22_X1 U11393 ( .A1(n10300), .A2(keyinput77), .B1(keyinput13), .B2(n5868), 
        .ZN(n10299) );
  OAI221_X1 U11394 ( .B1(n10300), .B2(keyinput77), .C1(n5868), .C2(keyinput13), 
        .A(n10299), .ZN(n10309) );
  AOI22_X1 U11395 ( .A1(n10303), .A2(keyinput80), .B1(n10302), .B2(keyinput38), 
        .ZN(n10301) );
  OAI221_X1 U11396 ( .B1(n10303), .B2(keyinput80), .C1(n10302), .C2(keyinput38), .A(n10301), .ZN(n10308) );
  XOR2_X1 U11397 ( .A(n10304), .B(keyinput104), .Z(n10306) );
  XNOR2_X1 U11398 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput33), .ZN(n10305)
         );
  NAND2_X1 U11399 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NOR4_X1 U11400 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10338) );
  AOI22_X1 U11401 ( .A1(n10313), .A2(keyinput90), .B1(keyinput1), .B2(n10312), 
        .ZN(n10311) );
  OAI221_X1 U11402 ( .B1(n10313), .B2(keyinput90), .C1(n10312), .C2(keyinput1), 
        .A(n10311), .ZN(n10324) );
  AOI22_X1 U11403 ( .A1(n10316), .A2(keyinput6), .B1(keyinput56), .B2(n10315), 
        .ZN(n10314) );
  OAI221_X1 U11404 ( .B1(n10316), .B2(keyinput6), .C1(n10315), .C2(keyinput56), 
        .A(n10314), .ZN(n10323) );
  XOR2_X1 U11405 ( .A(n10317), .B(keyinput65), .Z(n10321) );
  XNOR2_X1 U11406 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput111), .ZN(n10320) );
  XNOR2_X1 U11407 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput121), .ZN(n10319)
         );
  XNOR2_X1 U11408 ( .A(P2_REG1_REG_18__SCAN_IN), .B(keyinput76), .ZN(n10318)
         );
  NAND4_X1 U11409 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10322) );
  NOR3_X1 U11410 ( .A1(n10324), .A2(n10323), .A3(n10322), .ZN(n10337) );
  AOI22_X1 U11411 ( .A1(n6663), .A2(keyinput93), .B1(keyinput126), .B2(n10326), 
        .ZN(n10325) );
  OAI221_X1 U11412 ( .B1(n6663), .B2(keyinput93), .C1(n10326), .C2(keyinput126), .A(n10325), .ZN(n10335) );
  AOI22_X1 U11413 ( .A1(n10328), .A2(keyinput97), .B1(keyinput61), .B2(n7220), 
        .ZN(n10327) );
  OAI221_X1 U11414 ( .B1(n10328), .B2(keyinput97), .C1(n7220), .C2(keyinput61), 
        .A(n10327), .ZN(n10334) );
  XOR2_X1 U11415 ( .A(n6848), .B(keyinput28), .Z(n10332) );
  XNOR2_X1 U11416 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput58), .ZN(n10331)
         );
  XNOR2_X1 U11417 ( .A(SI_20_), .B(keyinput30), .ZN(n10330) );
  XNOR2_X1 U11418 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput49), .ZN(n10329) );
  NAND4_X1 U11419 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10333) );
  NOR3_X1 U11420 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10336) );
  NAND4_X1 U11421 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10512) );
  AOI22_X1 U11422 ( .A1(n10341), .A2(keyinput94), .B1(n5481), .B2(keyinput48), 
        .ZN(n10340) );
  OAI221_X1 U11423 ( .B1(n10341), .B2(keyinput94), .C1(n5481), .C2(keyinput48), 
        .A(n10340), .ZN(n10350) );
  XNOR2_X1 U11424 ( .A(keyinput47), .B(n10342), .ZN(n10349) );
  XNOR2_X1 U11425 ( .A(keyinput114), .B(n6448), .ZN(n10348) );
  XNOR2_X1 U11426 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput12), .ZN(n10346) );
  XNOR2_X1 U11427 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput92), .ZN(n10345)
         );
  XNOR2_X1 U11428 ( .A(P2_REG0_REG_18__SCAN_IN), .B(keyinput115), .ZN(n10344)
         );
  XNOR2_X1 U11429 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput4), .ZN(n10343) );
  NAND4_X1 U11430 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10347) );
  NOR4_X1 U11431 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10392) );
  AOI22_X1 U11432 ( .A1(n10353), .A2(keyinput57), .B1(n10352), .B2(keyinput84), 
        .ZN(n10351) );
  OAI221_X1 U11433 ( .B1(n10353), .B2(keyinput57), .C1(n10352), .C2(keyinput84), .A(n10351), .ZN(n10364) );
  INV_X1 U11434 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U11435 ( .A1(n10356), .A2(keyinput36), .B1(keyinput37), .B2(n10355), 
        .ZN(n10354) );
  OAI221_X1 U11436 ( .B1(n10356), .B2(keyinput36), .C1(n10355), .C2(keyinput37), .A(n10354), .ZN(n10363) );
  XOR2_X1 U11437 ( .A(n10357), .B(keyinput35), .Z(n10361) );
  XNOR2_X1 U11438 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput17), .ZN(n10360)
         );
  XNOR2_X1 U11439 ( .A(P1_REG2_REG_31__SCAN_IN), .B(keyinput18), .ZN(n10359)
         );
  XNOR2_X1 U11440 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput20), .ZN(n10358)
         );
  NAND4_X1 U11441 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10362) );
  NOR3_X1 U11442 ( .A1(n10364), .A2(n10363), .A3(n10362), .ZN(n10391) );
  AOI22_X1 U11443 ( .A1(n6409), .A2(keyinput55), .B1(keyinput91), .B2(n10366), 
        .ZN(n10365) );
  OAI221_X1 U11444 ( .B1(n6409), .B2(keyinput55), .C1(n10366), .C2(keyinput91), 
        .A(n10365), .ZN(n10377) );
  AOI22_X1 U11445 ( .A1(n5570), .A2(keyinput70), .B1(keyinput66), .B2(n10368), 
        .ZN(n10367) );
  OAI221_X1 U11446 ( .B1(n5570), .B2(keyinput70), .C1(n10368), .C2(keyinput66), 
        .A(n10367), .ZN(n10376) );
  AOI22_X1 U11447 ( .A1(n10371), .A2(keyinput21), .B1(keyinput106), .B2(n10370), .ZN(n10369) );
  OAI221_X1 U11448 ( .B1(n10371), .B2(keyinput21), .C1(n10370), .C2(
        keyinput106), .A(n10369), .ZN(n10375) );
  XNOR2_X1 U11449 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput112), .ZN(n10373)
         );
  XNOR2_X1 U11450 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput64), .ZN(n10372) );
  NAND2_X1 U11451 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  NOR4_X1 U11452 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10390) );
  AOI22_X1 U11453 ( .A1(n6684), .A2(keyinput96), .B1(keyinput10), .B2(n10379), 
        .ZN(n10378) );
  OAI221_X1 U11454 ( .B1(n6684), .B2(keyinput96), .C1(n10379), .C2(keyinput10), 
        .A(n10378), .ZN(n10388) );
  AOI22_X1 U11455 ( .A1(n10381), .A2(keyinput101), .B1(n9045), .B2(keyinput5), 
        .ZN(n10380) );
  OAI221_X1 U11456 ( .B1(n10381), .B2(keyinput101), .C1(n9045), .C2(keyinput5), 
        .A(n10380), .ZN(n10387) );
  XNOR2_X1 U11457 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput88), .ZN(n10385) );
  XNOR2_X1 U11458 ( .A(P2_REG0_REG_30__SCAN_IN), .B(keyinput44), .ZN(n10384)
         );
  XNOR2_X1 U11459 ( .A(P1_REG1_REG_12__SCAN_IN), .B(keyinput29), .ZN(n10383)
         );
  XNOR2_X1 U11460 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput100), .ZN(n10382)
         );
  NAND4_X1 U11461 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10386) );
  NOR3_X1 U11462 ( .A1(n10388), .A2(n10387), .A3(n10386), .ZN(n10389) );
  NAND4_X1 U11463 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10511) );
  AOI22_X1 U11464 ( .A1(n10395), .A2(keyinput120), .B1(keyinput52), .B2(n10394), .ZN(n10393) );
  OAI221_X1 U11465 ( .B1(n10395), .B2(keyinput120), .C1(n10394), .C2(
        keyinput52), .A(n10393), .ZN(n10408) );
  AOI22_X1 U11466 ( .A1(n10398), .A2(keyinput87), .B1(n10397), .B2(keyinput14), 
        .ZN(n10396) );
  OAI221_X1 U11467 ( .B1(n10398), .B2(keyinput87), .C1(n10397), .C2(keyinput14), .A(n10396), .ZN(n10407) );
  AOI22_X1 U11468 ( .A1(n10401), .A2(keyinput122), .B1(keyinput119), .B2(
        n10400), .ZN(n10399) );
  OAI221_X1 U11469 ( .B1(n10401), .B2(keyinput122), .C1(n10400), .C2(
        keyinput119), .A(n10399), .ZN(n10406) );
  XOR2_X1 U11470 ( .A(n10402), .B(keyinput34), .Z(n10404) );
  XNOR2_X1 U11471 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput41), .ZN(n10403) );
  NAND2_X1 U11472 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  NOR4_X1 U11473 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10451) );
  AOI22_X1 U11474 ( .A1(n10410), .A2(keyinput75), .B1(keyinput27), .B2(n7034), 
        .ZN(n10409) );
  OAI221_X1 U11475 ( .B1(n10410), .B2(keyinput75), .C1(n7034), .C2(keyinput27), 
        .A(n10409), .ZN(n10419) );
  AOI22_X1 U11476 ( .A1(n10412), .A2(keyinput22), .B1(keyinput24), .B2(n8944), 
        .ZN(n10411) );
  OAI221_X1 U11477 ( .B1(n10412), .B2(keyinput22), .C1(n8944), .C2(keyinput24), 
        .A(n10411), .ZN(n10418) );
  AOI22_X1 U11478 ( .A1(n6933), .A2(keyinput63), .B1(n8968), .B2(keyinput117), 
        .ZN(n10413) );
  OAI221_X1 U11479 ( .B1(n6933), .B2(keyinput63), .C1(n8968), .C2(keyinput117), 
        .A(n10413), .ZN(n10417) );
  XNOR2_X1 U11480 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput7), .ZN(n10415) );
  XNOR2_X1 U11481 ( .A(P2_REG1_REG_8__SCAN_IN), .B(keyinput60), .ZN(n10414) );
  NAND2_X1 U11482 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  NOR4_X1 U11483 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10450) );
  AOI22_X1 U11484 ( .A1(n10422), .A2(keyinput45), .B1(n10421), .B2(keyinput71), 
        .ZN(n10420) );
  OAI221_X1 U11485 ( .B1(n10422), .B2(keyinput45), .C1(n10421), .C2(keyinput71), .A(n10420), .ZN(n10434) );
  AOI22_X1 U11486 ( .A1(n10424), .A2(keyinput50), .B1(keyinput51), .B2(n6127), 
        .ZN(n10423) );
  OAI221_X1 U11487 ( .B1(n10424), .B2(keyinput50), .C1(n6127), .C2(keyinput51), 
        .A(n10423), .ZN(n10433) );
  AOI22_X1 U11488 ( .A1(n10427), .A2(keyinput107), .B1(n10426), .B2(keyinput86), .ZN(n10425) );
  OAI221_X1 U11489 ( .B1(n10427), .B2(keyinput107), .C1(n10426), .C2(
        keyinput86), .A(n10425), .ZN(n10432) );
  INV_X1 U11490 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U11491 ( .A1(n10430), .A2(keyinput59), .B1(n10429), .B2(keyinput67), 
        .ZN(n10428) );
  OAI221_X1 U11492 ( .B1(n10430), .B2(keyinput59), .C1(n10429), .C2(keyinput67), .A(n10428), .ZN(n10431) );
  NOR4_X1 U11493 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10449) );
  INV_X1 U11494 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U11495 ( .A1(n10437), .A2(keyinput32), .B1(keyinput53), .B2(n10436), 
        .ZN(n10435) );
  OAI221_X1 U11496 ( .B1(n10437), .B2(keyinput32), .C1(n10436), .C2(keyinput53), .A(n10435), .ZN(n10447) );
  AOI22_X1 U11497 ( .A1(n9567), .A2(keyinput42), .B1(n9247), .B2(keyinput72), 
        .ZN(n10438) );
  OAI221_X1 U11498 ( .B1(n9567), .B2(keyinput42), .C1(n9247), .C2(keyinput72), 
        .A(n10438), .ZN(n10446) );
  AOI22_X1 U11499 ( .A1(n10441), .A2(keyinput11), .B1(keyinput19), .B2(n10440), 
        .ZN(n10439) );
  OAI221_X1 U11500 ( .B1(n10441), .B2(keyinput11), .C1(n10440), .C2(keyinput19), .A(n10439), .ZN(n10445) );
  XOR2_X1 U11501 ( .A(n10226), .B(keyinput89), .Z(n10443) );
  XNOR2_X1 U11502 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput108), .ZN(n10442) );
  NAND2_X1 U11503 ( .A1(n10443), .A2(n10442), .ZN(n10444) );
  NOR4_X1 U11504 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  NAND4_X1 U11505 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10510) );
  AOI22_X1 U11506 ( .A1(n10454), .A2(keyinput105), .B1(keyinput39), .B2(n10453), .ZN(n10452) );
  OAI221_X1 U11507 ( .B1(n10454), .B2(keyinput105), .C1(n10453), .C2(
        keyinput39), .A(n10452), .ZN(n10463) );
  AOI22_X1 U11508 ( .A1(n5988), .A2(keyinput16), .B1(keyinput125), .B2(n5877), 
        .ZN(n10455) );
  OAI221_X1 U11509 ( .B1(n5988), .B2(keyinput16), .C1(n5877), .C2(keyinput125), 
        .A(n10455), .ZN(n10462) );
  AOI22_X1 U11510 ( .A1(n5524), .A2(keyinput15), .B1(n10457), .B2(keyinput25), 
        .ZN(n10456) );
  OAI221_X1 U11511 ( .B1(n5524), .B2(keyinput15), .C1(n10457), .C2(keyinput25), 
        .A(n10456), .ZN(n10461) );
  AOI22_X1 U11512 ( .A1(n10459), .A2(keyinput102), .B1(n7170), .B2(keyinput54), 
        .ZN(n10458) );
  OAI221_X1 U11513 ( .B1(n10459), .B2(keyinput102), .C1(n7170), .C2(keyinput54), .A(n10458), .ZN(n10460) );
  NOR4_X1 U11514 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10508) );
  XNOR2_X1 U11515 ( .A(n10464), .B(keyinput43), .ZN(n10465) );
  AOI21_X1 U11516 ( .B1(keyinput3), .B2(n10466), .A(n10465), .ZN(n10469) );
  XOR2_X1 U11517 ( .A(n4863), .B(keyinput123), .Z(n10468) );
  XNOR2_X1 U11518 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput83), .ZN(n10467) );
  NAND3_X1 U11519 ( .A1(n10469), .A2(n10468), .A3(n10467), .ZN(n10476) );
  AOI22_X1 U11520 ( .A1(n10472), .A2(keyinput69), .B1(keyinput109), .B2(n10471), .ZN(n10470) );
  OAI221_X1 U11521 ( .B1(n10472), .B2(keyinput69), .C1(n10471), .C2(
        keyinput109), .A(n10470), .ZN(n10475) );
  AOI22_X1 U11522 ( .A1(n6930), .A2(keyinput9), .B1(keyinput79), .B2(n6944), 
        .ZN(n10473) );
  OAI221_X1 U11523 ( .B1(n6930), .B2(keyinput9), .C1(n6944), .C2(keyinput79), 
        .A(n10473), .ZN(n10474) );
  NOR3_X1 U11524 ( .A1(n10476), .A2(n10475), .A3(n10474), .ZN(n10507) );
  AOI22_X1 U11525 ( .A1(n5921), .A2(keyinput98), .B1(keyinput78), .B2(n10478), 
        .ZN(n10477) );
  OAI221_X1 U11526 ( .B1(n5921), .B2(keyinput98), .C1(n10478), .C2(keyinput78), 
        .A(n10477), .ZN(n10491) );
  INV_X1 U11527 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11528 ( .A1(n10481), .A2(keyinput73), .B1(keyinput68), .B2(n10480), 
        .ZN(n10479) );
  OAI221_X1 U11529 ( .B1(n10481), .B2(keyinput73), .C1(n10480), .C2(keyinput68), .A(n10479), .ZN(n10490) );
  AOI22_X1 U11530 ( .A1(n10484), .A2(keyinput0), .B1(keyinput118), .B2(n10483), 
        .ZN(n10482) );
  OAI221_X1 U11531 ( .B1(n10484), .B2(keyinput0), .C1(n10483), .C2(keyinput118), .A(n10482), .ZN(n10489) );
  AOI22_X1 U11532 ( .A1(n10487), .A2(keyinput113), .B1(keyinput103), .B2(
        n10486), .ZN(n10485) );
  OAI221_X1 U11533 ( .B1(n10487), .B2(keyinput113), .C1(n10486), .C2(
        keyinput103), .A(n10485), .ZN(n10488) );
  NOR4_X1 U11534 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10506) );
  AOI22_X1 U11535 ( .A1(n10493), .A2(keyinput127), .B1(n10232), .B2(
        keyinput110), .ZN(n10492) );
  OAI221_X1 U11536 ( .B1(n10493), .B2(keyinput127), .C1(n10232), .C2(
        keyinput110), .A(n10492), .ZN(n10504) );
  AOI22_X1 U11537 ( .A1(n5886), .A2(keyinput2), .B1(keyinput8), .B2(n10495), 
        .ZN(n10494) );
  OAI221_X1 U11538 ( .B1(n5886), .B2(keyinput2), .C1(n10495), .C2(keyinput8), 
        .A(n10494), .ZN(n10503) );
  AOI22_X1 U11539 ( .A1(n10498), .A2(keyinput23), .B1(n10497), .B2(keyinput95), 
        .ZN(n10496) );
  OAI221_X1 U11540 ( .B1(n10498), .B2(keyinput23), .C1(n10497), .C2(keyinput95), .A(n10496), .ZN(n10502) );
  XNOR2_X1 U11541 ( .A(P1_REG3_REG_3__SCAN_IN), .B(keyinput62), .ZN(n10500) );
  XNOR2_X1 U11542 ( .A(keyinput40), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n10499)
         );
  NAND2_X1 U11543 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  NOR4_X1 U11544 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10505) );
  NAND4_X1 U11545 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  NOR4_X1 U11546 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10513) );
  OAI21_X1 U11547 ( .B1(keyinput3), .B2(n10514), .A(n10513), .ZN(n10515) );
  XOR2_X1 U11548 ( .A(n10516), .B(n10515), .Z(P1_U3311) );
  OAI21_X1 U11549 ( .B1(n10519), .B2(n10518), .A(n10517), .ZN(ADD_1068_U51) );
  OAI21_X1 U11550 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(ADD_1068_U47) );
  OAI21_X1 U11551 ( .B1(n10525), .B2(n10524), .A(n10523), .ZN(ADD_1068_U49) );
  OAI21_X1 U11552 ( .B1(n10528), .B2(n10527), .A(n10526), .ZN(ADD_1068_U48) );
  OAI21_X1 U11553 ( .B1(n10531), .B2(n10530), .A(n10529), .ZN(ADD_1068_U50) );
  AOI21_X1 U11554 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(ADD_1068_U54) );
  AOI21_X1 U11555 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(ADD_1068_U53) );
  OAI21_X1 U11556 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(ADD_1068_U52) );
  XNOR2_X1 U7301 ( .A(n5613), .B(n5612), .ZN(n7751) );
  CLKBUF_X1 U4976 ( .A(n6555), .Z(n4447) );
  CLKBUF_X1 U4995 ( .A(n6412), .Z(n4612) );
endmodule

