

module b20_C_gen_AntiSAT_k_256_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608;

  MUX2_X1 U5020 ( .A(n6895), .B(n6909), .S(n10570), .Z(n6897) );
  NAND2_X1 U5021 ( .A1(n6371), .A2(n6370), .ZN(n9601) );
  NAND2_X1 U5022 ( .A1(n6234), .A2(n6233), .ZN(n9627) );
  INV_X2 U5023 ( .A(n6451), .ZN(n6446) );
  AND2_X2 U5024 ( .A1(n6464), .A2(n6469), .ZN(n6461) );
  INV_X1 U5025 ( .A(n5336), .ZN(n5730) );
  INV_X1 U5026 ( .A(n7144), .ZN(n10479) );
  INV_X2 U5027 ( .A(n4519), .ZN(n4523) );
  INV_X1 U5028 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U5029 ( .A1(n5886), .A2(n4517), .ZN(n4514) );
  AND2_X1 U5030 ( .A1(n4514), .A2(n4515), .ZN(n5889) );
  OR2_X1 U5031 ( .A1(n4516), .A2(n6884), .ZN(n4515) );
  INV_X1 U5032 ( .A(n4742), .ZN(n4516) );
  AND2_X1 U5033 ( .A1(n4743), .A2(n4742), .ZN(n4517) );
  OAI22_X1 U5034 ( .A1(n5937), .A2(n5936), .B1(n9096), .B2(n8849), .ZN(n4518)
         );
  OAI22_X1 U5035 ( .A1(n5937), .A2(n5936), .B1(n9096), .B2(n8849), .ZN(n5939)
         );
  INV_X1 U5036 ( .A(n8523), .ZN(n5123) );
  INV_X1 U5037 ( .A(n6461), .ZN(n6781) );
  NOR2_X1 U5038 ( .A1(n10276), .A2(n6440), .ZN(n10257) );
  INV_X1 U5039 ( .A(n8351), .ZN(n8508) );
  INV_X1 U5040 ( .A(n8569), .ZN(n8556) );
  INV_X1 U5041 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8146) );
  AND2_X1 U5042 ( .A1(n9535), .A2(n8403), .ZN(n9520) );
  NOR2_X2 U5043 ( .A1(n8024), .A2(n9222), .ZN(n8023) );
  NAND2_X1 U5044 ( .A1(n4843), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4842) );
  NOR2_X1 U5045 ( .A1(n4755), .A2(n4573), .ZN(n4754) );
  AND3_X1 U5046 ( .A1(n6006), .A2(n6005), .A3(n6004), .ZN(n10298) );
  NOR2_X1 U5047 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6002) );
  INV_X1 U5048 ( .A(n6929), .ZN(n4993) );
  OAI211_X2 U5049 ( .C1(n6936), .C2(n6071), .A(n4842), .B(n5150), .ZN(n10276)
         );
  NAND2_X1 U5050 ( .A1(n5421), .A2(n5420), .ZN(n5419) );
  NAND4_X2 U5051 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n8738)
         );
  MUX2_X1 U5052 ( .A(n6910), .B(n6909), .S(n10545), .Z(n6911) );
  NAND2_X1 U5053 ( .A1(n5303), .A2(n9165), .ZN(n4519) );
  NAND2_X1 U5054 ( .A1(n5304), .A2(n5303), .ZN(n4520) );
  INV_X2 U5055 ( .A(n9568), .ZN(n9197) );
  INV_X1 U5056 ( .A(n6461), .ZN(n4521) );
  NAND2_X4 U5057 ( .A1(n6437), .A2(n7469), .ZN(n6451) );
  OAI21_X2 U5058 ( .B1(n8921), .B2(n6854), .A(n6853), .ZN(n8906) );
  AOI21_X2 U5059 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7841), .A(n7828), .ZN(
        n6681) );
  AOI21_X2 U5060 ( .B1(n8690), .B2(n8613), .A(n8612), .ZN(n8672) );
  AND2_X1 U5061 ( .A1(n8580), .A2(n5304), .ZN(n4522) );
  AOI21_X2 U5062 ( .B1(n8056), .B2(n4765), .A(n4762), .ZN(n9599) );
  XNOR2_X2 U5063 ( .A(n6687), .B(n8822), .ZN(n8809) );
  OAI21_X2 U5064 ( .B1(n5591), .B2(n5590), .A(n5232), .ZN(n5609) );
  XNOR2_X2 U5065 ( .A(n5990), .B(n5989), .ZN(n6326) );
  BUF_X2 U5066 ( .A(n6324), .Z(n4524) );
  XNOR2_X1 U5067 ( .A(n5991), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6324) );
  XNOR2_X2 U5068 ( .A(n5437), .B(n5436), .ZN(n6955) );
  OAI21_X2 U5069 ( .B1(n5426), .B2(n5427), .A(n5193), .ZN(n5437) );
  INV_X4 U5070 ( .A(n6864), .ZN(n6773) );
  INV_X1 U5071 ( .A(n4520), .ZN(n4525) );
  INV_X1 U5072 ( .A(n4520), .ZN(n4526) );
  NAND3_X1 U5073 ( .A1(n5073), .A2(n5339), .A3(n5365), .ZN(n5400) );
  NOR2_X4 U5074 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5339) );
  INV_X1 U5075 ( .A(n8236), .ZN(n10318) );
  NAND2_X2 U5076 ( .A1(n5806), .A2(n5804), .ZN(n10440) );
  INV_X1 U5077 ( .A(n10428), .ZN(n7330) );
  INV_X1 U5078 ( .A(n10303), .ZN(n7609) );
  INV_X1 U5079 ( .A(n10426), .ZN(n10455) );
  AND2_X1 U5081 ( .A1(n9756), .A2(n5984), .ZN(n8162) );
  NAND2_X1 U5082 ( .A1(n4810), .A2(n4808), .ZN(n8856) );
  NAND2_X1 U5083 ( .A1(n9520), .A2(n9523), .ZN(n9519) );
  OAI21_X1 U5084 ( .B1(n9193), .B2(n4645), .A(n4939), .ZN(n6801) );
  NAND2_X1 U5085 ( .A1(n5114), .A2(n5130), .ZN(n6804) );
  NAND2_X1 U5086 ( .A1(n5117), .A2(n4564), .ZN(n5114) );
  NAND2_X1 U5087 ( .A1(n6593), .A2(n6592), .ZN(n9259) );
  NAND2_X1 U5088 ( .A1(n8158), .A2(n8157), .ZN(n9713) );
  NAND2_X1 U5089 ( .A1(n6368), .A2(n8300), .ZN(n4852) );
  NAND2_X1 U5090 ( .A1(n9103), .A2(n8727), .ZN(n5130) );
  NOR2_X1 U5091 ( .A1(n4557), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U5092 ( .A1(n6125), .A2(n7594), .ZN(n7598) );
  OR2_X1 U5093 ( .A1(n7747), .A2(n4612), .ZN(n4999) );
  AND2_X1 U5094 ( .A1(n6143), .A2(n6142), .ZN(n10383) );
  OR2_X1 U5095 ( .A1(n6271), .A2(n6270), .ZN(n9568) );
  NOR2_X1 U5096 ( .A1(n7064), .A2(n6460), .ZN(n7175) );
  AND2_X1 U5097 ( .A1(n6060), .A2(n6059), .ZN(n10332) );
  NAND2_X1 U5098 ( .A1(n6818), .A2(n5374), .ZN(n7374) );
  OAI21_X1 U5099 ( .B1(n5426), .B2(n4672), .A(n4670), .ZN(n5456) );
  NAND2_X1 U5100 ( .A1(n6335), .A2(n6334), .ZN(n10246) );
  OAI21_X2 U5101 ( .B1(n6645), .B2(n6636), .A(n9603), .ZN(n6637) );
  NAND2_X1 U5102 ( .A1(n4761), .A2(n4760), .ZN(n10268) );
  OR2_X1 U5103 ( .A1(n6067), .A2(n6066), .ZN(n10322) );
  OR2_X1 U5104 ( .A1(n6026), .A2(n6025), .ZN(n9306) );
  OR2_X1 U5105 ( .A1(n6080), .A2(n6079), .ZN(n9305) );
  OR2_X1 U5106 ( .A1(n6057), .A2(n6056), .ZN(n10341) );
  OR2_X1 U5107 ( .A1(n6039), .A2(n6038), .ZN(n10323) );
  NAND4_X1 U5108 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n10426)
         );
  NAND2_X1 U5109 ( .A1(n6703), .A2(n6932), .ZN(n7302) );
  NAND2_X1 U5110 ( .A1(n5351), .A2(n5350), .ZN(n5349) );
  AND2_X1 U5111 ( .A1(n5984), .A2(n5986), .ZN(n6008) );
  NAND2_X1 U5112 ( .A1(n5959), .A2(n5958), .ZN(n7996) );
  XNOR2_X1 U5113 ( .A(n5594), .B(n5752), .ZN(n7660) );
  NAND2_X1 U5114 ( .A1(n5024), .A2(n5022), .ZN(n7805) );
  NAND2_X1 U5115 ( .A1(n5593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5594) );
  OR2_X1 U5116 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U5117 ( .A1(n4703), .A2(n5318), .ZN(n6936) );
  OR2_X1 U5118 ( .A1(n6392), .A2(n6390), .ZN(n6434) );
  NAND2_X1 U5119 ( .A1(n5445), .A2(n5444), .ZN(n5480) );
  INV_X1 U5120 ( .A(n5304), .ZN(n9165) );
  XNOR2_X1 U5121 ( .A(n6408), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8082) );
  INV_X1 U5122 ( .A(n5446), .ZN(n5445) );
  OAI211_X1 U5123 ( .C1(n7284), .C2(n4993), .A(n4991), .B(n4988), .ZN(n7250)
         );
  XNOR2_X1 U5124 ( .A(n5295), .B(n5294), .ZN(n5963) );
  NAND2_X1 U5125 ( .A1(n5298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  AND2_X1 U5126 ( .A1(n5171), .A2(n5172), .ZN(n5350) );
  AND2_X1 U5128 ( .A1(n4768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  AND2_X1 U5129 ( .A1(n4769), .A2(n4812), .ZN(n6311) );
  AND3_X1 U5130 ( .A1(n5288), .A2(n4546), .A3(n5782), .ZN(n5082) );
  OAI21_X1 U5131 ( .B1(n6166), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U5132 ( .A1(n5341), .A2(n5353), .ZN(n6949) );
  NOR2_X1 U5133 ( .A1(n4791), .A2(n5287), .ZN(n5288) );
  NAND2_X1 U5134 ( .A1(n5311), .A2(n5310), .ZN(n7263) );
  AND2_X1 U5135 ( .A1(n4813), .A2(n4554), .ZN(n4769) );
  NAND2_X1 U5136 ( .A1(n4729), .A2(n4728), .ZN(n5161) );
  AND4_X1 U5137 ( .A1(n6154), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4813)
         );
  NAND2_X1 U5138 ( .A1(n5339), .A2(n5340), .ZN(n5353) );
  INV_X1 U5139 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5753) );
  NOR2_X1 U5140 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4793) );
  INV_X1 U5141 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6316) );
  NOR2_X1 U5142 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4710) );
  NOR2_X1 U5143 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6027) );
  NOR2_X1 U5144 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4711) );
  NOR2_X1 U5145 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4712) );
  INV_X1 U5146 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5525) );
  INV_X4 U5147 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5148 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10083) );
  INV_X1 U5149 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9899) );
  INV_X1 U5150 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5470) );
  NOR2_X1 U5151 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10191) );
  INV_X4 U5152 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AND2_X1 U5153 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10190) );
  NOR2_X1 U5154 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6154) );
  NOR2_X1 U5155 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6153) );
  NOR2_X1 U5156 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6152) );
  NOR2_X1 U5157 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5966) );
  INV_X1 U5158 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5475) );
  AOI21_X2 U5159 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6935), .A(n7297), .ZN(
        n6673) );
  NAND2_X1 U5160 ( .A1(n6866), .A2(n6914), .ZN(n4527) );
  OAI21_X1 U5161 ( .B1(n8229), .B2(n4706), .A(n4704), .ZN(n8251) );
  NAND2_X1 U5162 ( .A1(n8508), .A2(n8231), .ZN(n4706) );
  NAND2_X1 U5163 ( .A1(n8229), .A2(n4705), .ZN(n4704) );
  NOR2_X1 U5164 ( .A1(n8508), .A2(n8228), .ZN(n4705) );
  AND2_X1 U5165 ( .A1(n5882), .A2(n5890), .ZN(n4743) );
  OR2_X1 U5166 ( .A1(n9106), .A2(n8526), .ZN(n5905) );
  INV_X1 U5167 ( .A(n4970), .ZN(n4969) );
  CLKBUF_X3 U5168 ( .A(n5344), .Z(n5733) );
  AND2_X1 U5169 ( .A1(n8580), .A2(n9165), .ZN(n5344) );
  NAND2_X1 U5170 ( .A1(n8254), .A2(n8255), .ZN(n4687) );
  INV_X1 U5171 ( .A(n6827), .ZN(n4785) );
  NAND2_X1 U5172 ( .A1(n4923), .A2(n4925), .ZN(n4631) );
  AND2_X1 U5173 ( .A1(n9728), .A2(n9658), .ZN(n8324) );
  NOR2_X1 U5174 ( .A1(n7377), .A2(n7103), .ZN(n7108) );
  NAND2_X1 U5175 ( .A1(n7106), .A2(n7105), .ZN(n7107) );
  NAND2_X1 U5176 ( .A1(n4878), .A2(n4567), .ZN(n4877) );
  NAND2_X1 U5177 ( .A1(n6896), .A2(n8862), .ZN(n5916) );
  OR2_X1 U5178 ( .A1(n6896), .A2(n8862), .ZN(n5917) );
  NOR2_X1 U5179 ( .A1(n4775), .A2(n4774), .ZN(n4773) );
  INV_X1 U5180 ( .A(n6857), .ZN(n4774) );
  OR2_X1 U5181 ( .A1(n8940), .A2(n8951), .ZN(n5898) );
  OAI21_X1 U5182 ( .B1(n4786), .B2(n4785), .A(n7700), .ZN(n4784) );
  AND2_X1 U5183 ( .A1(n5655), .A2(n8908), .ZN(n5903) );
  AND2_X1 U5184 ( .A1(n8961), .A2(n6847), .ZN(n4799) );
  OR2_X1 U5185 ( .A1(n8984), .A2(n8697), .ZN(n5890) );
  AND3_X1 U5186 ( .A1(n5376), .A2(n5283), .A3(n5284), .ZN(n5073) );
  INV_X1 U5187 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5284) );
  INV_X1 U5188 ( .A(n6574), .ZN(n4926) );
  INV_X1 U5189 ( .A(n8086), .ZN(n4922) );
  INV_X1 U5190 ( .A(n8087), .ZN(n4921) );
  OR2_X1 U5191 ( .A1(n9724), .A2(n6451), .ZN(n6616) );
  INV_X1 U5192 ( .A(n8324), .ZN(n8403) );
  NOR2_X1 U5193 ( .A1(n9557), .A2(n4759), .ZN(n4758) );
  INV_X1 U5194 ( .A(n8397), .ZN(n4759) );
  NOR2_X1 U5195 ( .A1(n10326), .A2(n9305), .ZN(n8449) );
  NAND2_X1 U5196 ( .A1(n9310), .A2(n10290), .ZN(n8441) );
  XNOR2_X1 U5197 ( .A(n5273), .B(n5272), .ZN(n5719) );
  NAND2_X1 U5198 ( .A1(n4951), .A2(n4949), .ZN(n5694) );
  AOI21_X1 U5199 ( .B1(n4953), .B2(n4955), .A(n4950), .ZN(n4949) );
  INV_X1 U5200 ( .A(n5262), .ZN(n4950) );
  OAI21_X1 U5201 ( .B1(n5609), .B2(n9918), .A(n5233), .ZN(n5235) );
  NOR2_X1 U5202 ( .A1(n5467), .A2(n4948), .ZN(n4947) );
  INV_X1 U5203 ( .A(n5198), .ZN(n4948) );
  XNOR2_X1 U5204 ( .A(n5199), .B(SI_11_), .ZN(n5467) );
  INV_X1 U5205 ( .A(n5456), .ZN(n5454) );
  XNOR2_X1 U5206 ( .A(n5194), .B(n9886), .ZN(n5436) );
  NAND2_X1 U5207 ( .A1(n5419), .A2(n5190), .ZN(n5426) );
  XNOR2_X1 U5208 ( .A(n5191), .B(SI_8_), .ZN(n5427) );
  NAND2_X1 U5209 ( .A1(n10190), .A2(n5154), .ZN(n4728) );
  INV_X1 U5210 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5153) );
  NAND2_X1 U5211 ( .A1(n5041), .A2(n5038), .ZN(n5037) );
  OAI21_X1 U5212 ( .B1(n8570), .B2(n4528), .A(n5043), .ZN(n5041) );
  NAND2_X1 U5213 ( .A1(n5040), .A2(n5039), .ZN(n5038) );
  INV_X1 U5214 ( .A(n8570), .ZN(n5040) );
  AND2_X1 U5215 ( .A1(n5054), .A2(n5052), .ZN(n5051) );
  INV_X1 U5216 ( .A(n8645), .ZN(n5052) );
  AND2_X1 U5217 ( .A1(n7324), .A2(n7321), .ZN(n8658) );
  AOI21_X1 U5218 ( .B1(n7535), .B2(n7390), .A(n5027), .ZN(n5026) );
  XNOR2_X1 U5219 ( .A(n6949), .B(n10550), .ZN(n7286) );
  AND2_X1 U5220 ( .A1(n6706), .A2(n7363), .ZN(n6708) );
  OAI22_X1 U5221 ( .A1(n6859), .A2(n6858), .B1(n5706), .B2(n8728), .ZN(n8861)
         );
  AND2_X1 U5222 ( .A1(n5121), .A2(n5120), .ZN(n5119) );
  NAND2_X1 U5223 ( .A1(n5123), .A2(n5131), .ZN(n5120) );
  INV_X1 U5224 ( .A(n5127), .ZN(n5124) );
  NAND2_X1 U5225 ( .A1(n5115), .A2(n5118), .ZN(n5117) );
  AND2_X1 U5226 ( .A1(n5125), .A2(n5131), .ZN(n5118) );
  AND2_X1 U5227 ( .A1(n5692), .A2(n5691), .ZN(n8526) );
  AND2_X1 U5228 ( .A1(n5681), .A2(n5680), .ZN(n8885) );
  NAND2_X1 U5229 ( .A1(n6866), .A2(n6914), .ZN(n5319) );
  AND4_X1 U5230 ( .A1(n5589), .A2(n5588), .A3(n5587), .A4(n5586), .ZN(n8977)
         );
  INV_X1 U5231 ( .A(n5319), .ZN(n5596) );
  INV_X1 U5232 ( .A(n6866), .ZN(n5595) );
  OR2_X1 U5233 ( .A1(n8145), .A2(n8146), .ZN(n5299) );
  NAND2_X1 U5234 ( .A1(n4905), .A2(n4904), .ZN(n8100) );
  AOI21_X1 U5235 ( .B1(n4907), .B2(n4910), .A(n4541), .ZN(n4904) );
  NAND2_X1 U5236 ( .A1(n9227), .A2(n6611), .ZN(n9193) );
  AND2_X1 U5237 ( .A1(n5985), .A2(n9756), .ZN(n8163) );
  AND2_X1 U5238 ( .A1(n5986), .A2(n5985), .ZN(n6171) );
  OR2_X1 U5239 ( .A1(n9576), .A2(n9683), .ZN(n4832) );
  NOR2_X1 U5240 ( .A1(n4848), .A2(n4576), .ZN(n4847) );
  NAND2_X1 U5241 ( .A1(n7962), .A2(n8381), .ZN(n4849) );
  INV_X1 U5242 ( .A(n8278), .ZN(n8464) );
  INV_X1 U5243 ( .A(n6013), .ZN(n6224) );
  INV_X1 U5244 ( .A(n8141), .ZN(n5979) );
  NAND4_X1 U5245 ( .A1(n4769), .A2(n4814), .A3(n4812), .A4(n4722), .ZN(n4723)
         );
  INV_X1 U5246 ( .A(n5974), .ZN(n4722) );
  NAND2_X1 U5247 ( .A1(n4957), .A2(n5217), .ZN(n5565) );
  AOI21_X1 U5248 ( .B1(n5403), .B2(n4979), .A(n4978), .ZN(n4976) );
  INV_X1 U5249 ( .A(n5186), .ZN(n4978) );
  NAND2_X1 U5250 ( .A1(n5178), .A2(SI_5_), .ZN(n5181) );
  NAND2_X2 U5251 ( .A1(n5962), .A2(n5963), .ZN(n6866) );
  INV_X1 U5252 ( .A(n9658), .ZN(n9559) );
  NAND2_X1 U5253 ( .A1(n5833), .A2(n5873), .ZN(n4741) );
  NAND2_X1 U5254 ( .A1(n4740), .A2(n6884), .ZN(n4739) );
  NOR2_X1 U5255 ( .A1(n8449), .A2(n8351), .ZN(n4689) );
  NAND2_X1 U5256 ( .A1(n5852), .A2(n5851), .ZN(n4749) );
  AND2_X1 U5257 ( .A1(n5853), .A2(n6884), .ZN(n4748) );
  NAND2_X1 U5258 ( .A1(n4683), .A2(n8259), .ZN(n8272) );
  NAND2_X1 U5259 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  INV_X1 U5260 ( .A(n8260), .ZN(n4684) );
  NAND2_X1 U5261 ( .A1(n5876), .A2(n5870), .ZN(n4679) );
  NAND2_X1 U5262 ( .A1(n8287), .A2(n4692), .ZN(n4691) );
  NAND2_X1 U5263 ( .A1(n8474), .A2(n8351), .ZN(n4692) );
  OAI21_X1 U5264 ( .B1(n8283), .B2(n4695), .A(n4694), .ZN(n4693) );
  NAND2_X1 U5265 ( .A1(n8285), .A2(n4696), .ZN(n4695) );
  NOR2_X1 U5266 ( .A1(n8286), .A2(n8289), .ZN(n4694) );
  OAI21_X1 U5267 ( .B1(n4702), .B2(n4701), .A(n8397), .ZN(n4700) );
  NOR2_X1 U5268 ( .A1(n8396), .A2(n8508), .ZN(n4701) );
  NOR2_X1 U5269 ( .A1(n8314), .A2(n9582), .ZN(n4702) );
  NAND2_X1 U5270 ( .A1(n8404), .A2(n8508), .ZN(n4699) );
  NAND2_X1 U5271 ( .A1(n5787), .A2(n8523), .ZN(n5914) );
  INV_X1 U5272 ( .A(n5902), .ZN(n4731) );
  AOI21_X1 U5273 ( .B1(n8496), .B2(n8333), .A(n8332), .ZN(n8335) );
  OR2_X1 U5274 ( .A1(n9048), .A2(n5746), .ZN(n5932) );
  AND2_X1 U5275 ( .A1(n9720), .A2(n9659), .ZN(n8333) );
  NOR2_X1 U5276 ( .A1(n9513), .A2(n9532), .ZN(n4727) );
  NOR2_X1 U5277 ( .A1(n9627), .A2(n4719), .ZN(n4718) );
  INV_X1 U5278 ( .A(n4720), .ZN(n4719) );
  NOR2_X1 U5279 ( .A1(n5227), .A2(n4964), .ZN(n4961) );
  NAND2_X1 U5280 ( .A1(n4980), .A2(n4606), .ZN(n5213) );
  NAND2_X1 U5281 ( .A1(n5070), .A2(n7981), .ZN(n5069) );
  INV_X1 U5282 ( .A(n5069), .ZN(n5065) );
  INV_X1 U5283 ( .A(n7936), .ZN(n5071) );
  XNOR2_X1 U5284 ( .A(n8940), .B(n8569), .ZN(n8553) );
  AOI21_X1 U5285 ( .B1(n5051), .B2(n8636), .A(n8692), .ZN(n5049) );
  INV_X1 U5286 ( .A(n5051), .ZN(n5050) );
  INV_X1 U5287 ( .A(n5929), .ZN(n5930) );
  INV_X1 U5288 ( .A(n5922), .ZN(n4745) );
  AND2_X1 U5289 ( .A1(n4882), .A2(n6932), .ZN(n6672) );
  INV_X1 U5290 ( .A(n8834), .ZN(n5007) );
  INV_X1 U5291 ( .A(n6719), .ZN(n5006) );
  NOR2_X1 U5292 ( .A1(n5839), .A2(n5095), .ZN(n5094) );
  INV_X1 U5293 ( .A(n5843), .ZN(n5095) );
  INV_X1 U5294 ( .A(n5849), .ZN(n5839) );
  AND2_X1 U5295 ( .A1(n6824), .A2(n4781), .ZN(n4780) );
  NOR2_X1 U5296 ( .A1(n6826), .A2(n4785), .ZN(n4781) );
  AND2_X1 U5297 ( .A1(n10428), .A2(n8663), .ZN(n6820) );
  OR2_X1 U5298 ( .A1(n9118), .A2(n8560), .ZN(n5910) );
  OR2_X1 U5299 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  NOR2_X1 U5300 ( .A1(n9010), .A2(n6840), .ZN(n6841) );
  OR2_X1 U5301 ( .A1(n9158), .A2(n8718), .ZN(n5879) );
  AND2_X1 U5302 ( .A1(n5861), .A2(n5109), .ZN(n5108) );
  NAND2_X1 U5303 ( .A1(n5518), .A2(n5517), .ZN(n5109) );
  NAND2_X1 U5304 ( .A1(n10519), .A2(n8735), .ZN(n5843) );
  AOI21_X1 U5305 ( .B1(n5088), .B2(n7649), .A(n5087), .ZN(n5086) );
  INV_X1 U5306 ( .A(n5841), .ZN(n5087) );
  NOR2_X1 U5307 ( .A1(n7722), .A2(n5021), .ZN(n7105) );
  INV_X1 U5308 ( .A(n4935), .ZN(n4934) );
  OAI22_X1 U5309 ( .A1(n7580), .A2(n4936), .B1(n6495), .B2(n6496), .ZN(n4935)
         );
  NOR2_X1 U5310 ( .A1(n7580), .A2(n4938), .ZN(n4937) );
  INV_X1 U5311 ( .A(n7456), .ZN(n4938) );
  NOR2_X1 U5312 ( .A1(n4916), .A2(n4914), .ZN(n4913) );
  INV_X1 U5313 ( .A(n7808), .ZN(n4914) );
  OAI21_X1 U5314 ( .B1(n4627), .B2(n4930), .A(n4927), .ZN(n6514) );
  AOI21_X1 U5315 ( .B1(n4931), .B2(n4929), .A(n4928), .ZN(n4927) );
  INV_X1 U5316 ( .A(n4931), .ZN(n4930) );
  NAND2_X1 U5317 ( .A1(n4628), .A2(n6484), .ZN(n4627) );
  OAI22_X1 U5318 ( .A1(n7175), .A2(n4647), .B1(n5151), .B2(n4548), .ZN(n6482)
         );
  NAND2_X1 U5319 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  INV_X1 U5320 ( .A(n5151), .ZN(n4648) );
  AOI21_X1 U5321 ( .B1(n8351), .B2(n8350), .A(n8341), .ZN(n8349) );
  AND2_X1 U5322 ( .A1(n9713), .A2(n8351), .ZN(n8343) );
  NOR3_X1 U5323 ( .A1(n8352), .A2(n8351), .A3(n9713), .ZN(n8353) );
  AND2_X1 U5324 ( .A1(n8434), .A2(n6391), .ZN(n8351) );
  NOR2_X1 U5325 ( .A1(n9371), .A2(n4616), .ZN(n4855) );
  NOR2_X1 U5326 ( .A1(n4855), .A2(n9373), .ZN(n9396) );
  INV_X1 U5327 ( .A(n8333), .ZN(n8492) );
  NOR2_X1 U5328 ( .A1(n10210), .A2(n8048), .ZN(n4715) );
  AND2_X1 U5329 ( .A1(n6139), .A2(n8460), .ZN(n8376) );
  OR2_X1 U5330 ( .A1(n10342), .A2(n7811), .ZN(n8261) );
  NAND2_X1 U5331 ( .A1(n6393), .A2(n7479), .ZN(n6435) );
  NAND2_X1 U5332 ( .A1(n5237), .A2(n4975), .ZN(n4974) );
  INV_X1 U5333 ( .A(n5631), .ZN(n4975) );
  NAND2_X1 U5334 ( .A1(n4610), .A2(n5223), .ZN(n4962) );
  INV_X1 U5335 ( .A(n5217), .ZN(n4965) );
  INV_X1 U5336 ( .A(n5213), .ZN(n5538) );
  INV_X1 U5337 ( .A(n5427), .ZN(n4673) );
  INV_X1 U5338 ( .A(n5193), .ZN(n4671) );
  OAI21_X1 U5339 ( .B1(n8151), .B2(n4668), .A(n4667), .ZN(n5175) );
  OAI21_X1 U5340 ( .B1(n5161), .B2(n5156), .A(n5155), .ZN(n5159) );
  NAND2_X1 U5341 ( .A1(n5063), .A2(n5060), .ZN(n5059) );
  INV_X1 U5342 ( .A(n5061), .ZN(n5060) );
  AOI21_X1 U5343 ( .B1(n8670), .B2(n8671), .A(n5062), .ZN(n5061) );
  INV_X1 U5344 ( .A(n8620), .ZN(n5062) );
  AOI21_X1 U5345 ( .B1(n5055), .B2(n4529), .A(n4574), .ZN(n5054) );
  AND2_X1 U5346 ( .A1(n8658), .A2(n7317), .ZN(n5029) );
  NAND2_X1 U5347 ( .A1(n7766), .A2(n7765), .ZN(n7791) );
  AND2_X1 U5348 ( .A1(n8613), .A2(n8544), .ZN(n8691) );
  NAND2_X1 U5349 ( .A1(n7660), .A2(n7722), .ZN(n7102) );
  AND4_X1 U5350 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n7394)
         );
  NAND2_X1 U5351 ( .A1(n4522), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5308) );
  XNOR2_X1 U5352 ( .A(n6949), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7283) );
  NAND2_X1 U5353 ( .A1(n7284), .A2(n4985), .ZN(n4991) );
  NAND2_X1 U5354 ( .A1(n4880), .A2(n4883), .ZN(n4878) );
  INV_X1 U5355 ( .A(n7253), .ZN(n4880) );
  NAND2_X1 U5356 ( .A1(n6702), .A2(n7233), .ZN(n6704) );
  INV_X1 U5357 ( .A(n6708), .ZN(n5015) );
  OAI21_X1 U5358 ( .B1(n6708), .B2(P2_REG1_REG_7__SCAN_IN), .A(n5014), .ZN(
        n5013) );
  INV_X1 U5359 ( .A(n7402), .ZN(n5014) );
  OR2_X1 U5360 ( .A1(n6708), .A2(n6707), .ZN(n7357) );
  NAND2_X1 U5361 ( .A1(n5012), .A2(n5010), .ZN(n6709) );
  NAND2_X1 U5362 ( .A1(n5013), .A2(n4547), .ZN(n5012) );
  NAND2_X1 U5363 ( .A1(n7357), .A2(n5011), .ZN(n5010) );
  AND2_X1 U5364 ( .A1(n5015), .A2(n4547), .ZN(n5011) );
  XNOR2_X1 U5365 ( .A(n6711), .B(n7745), .ZN(n7747) );
  NOR2_X1 U5366 ( .A1(n7672), .A2(n7671), .ZN(n7670) );
  NAND2_X1 U5367 ( .A1(n6712), .A2(n4998), .ZN(n4997) );
  INV_X1 U5368 ( .A(n7837), .ZN(n4998) );
  OR2_X1 U5369 ( .A1(n7747), .A2(n10566), .ZN(n5001) );
  NOR2_X1 U5370 ( .A1(n8822), .A2(n6718), .ZN(n6720) );
  NOR2_X1 U5371 ( .A1(n6720), .A2(n6719), .ZN(n8811) );
  NAND2_X1 U5372 ( .A1(n5006), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5005) );
  INV_X1 U5373 ( .A(n5963), .ZN(n6864) );
  AND2_X1 U5374 ( .A1(n8574), .A2(n8727), .ZN(n6860) );
  NAND2_X1 U5375 ( .A1(n5917), .A2(n5916), .ZN(n6862) );
  OAI21_X1 U5376 ( .B1(n8854), .B2(n10451), .A(n6867), .ZN(n4809) );
  NOR2_X1 U5377 ( .A1(n5772), .A2(n5128), .ZN(n5127) );
  NAND2_X1 U5378 ( .A1(n5905), .A2(n5904), .ZN(n5126) );
  OAI21_X1 U5379 ( .B1(n8975), .B2(n4796), .A(n4794), .ZN(n6850) );
  INV_X1 U5380 ( .A(n4795), .ZN(n4794) );
  OR2_X1 U5381 ( .A1(n9072), .A2(n8932), .ZN(n8936) );
  AND3_X1 U5382 ( .A1(n5639), .A2(n5638), .A3(n5637), .ZN(n8951) );
  NOR2_X1 U5383 ( .A1(n6828), .A2(n4790), .ZN(n4786) );
  OR2_X1 U5384 ( .A1(n7421), .A2(n7394), .ZN(n6825) );
  OAI21_X1 U5385 ( .B1(n10424), .B2(n6817), .A(n6816), .ZN(n7369) );
  OAI211_X1 U5386 ( .C1(n5319), .C2(n5156), .A(n5342), .B(n5152), .ZN(n7144)
         );
  NOR2_X1 U5387 ( .A1(n7805), .A2(n6900), .ZN(n7377) );
  AND2_X1 U5388 ( .A1(n5685), .A2(n5684), .ZN(n8566) );
  NAND2_X1 U5389 ( .A1(n4584), .A2(n4530), .ZN(n4775) );
  NAND2_X1 U5390 ( .A1(n6856), .A2(n6855), .ZN(n4777) );
  NAND2_X1 U5391 ( .A1(n8906), .A2(n4604), .ZN(n4772) );
  AND2_X1 U5392 ( .A1(n5787), .A2(n5905), .ZN(n8883) );
  OR2_X1 U5393 ( .A1(n8920), .A2(n5903), .ZN(n8914) );
  NAND2_X1 U5394 ( .A1(n8975), .A2(n4799), .ZN(n8960) );
  INV_X1 U5395 ( .A(n8975), .ZN(n4798) );
  NAND2_X1 U5396 ( .A1(n5077), .A2(n5078), .ZN(n8971) );
  INV_X1 U5397 ( .A(n5079), .ZN(n5078) );
  OAI21_X1 U5398 ( .B1(n6844), .B2(n5080), .A(n8973), .ZN(n5079) );
  NAND2_X1 U5399 ( .A1(n5100), .A2(n5097), .ZN(n9011) );
  INV_X1 U5400 ( .A(n5098), .ZN(n5097) );
  OAI21_X1 U5401 ( .B1(n5880), .B2(n5099), .A(n5865), .ZN(n5098) );
  AOI21_X1 U5402 ( .B1(n5108), .B2(n5105), .A(n5104), .ZN(n5103) );
  INV_X1 U5403 ( .A(n5517), .ZN(n5105) );
  INV_X1 U5404 ( .A(n5862), .ZN(n5104) );
  INV_X1 U5405 ( .A(n5108), .ZN(n5106) );
  NAND2_X1 U5406 ( .A1(n5509), .A2(n5508), .ZN(n7930) );
  AND2_X1 U5407 ( .A1(n7095), .A2(n6884), .ZN(n10425) );
  INV_X1 U5408 ( .A(n10454), .ZN(n10427) );
  INV_X1 U5409 ( .A(n7788), .ZN(n10526) );
  NAND2_X1 U5410 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U5411 ( .A1(n5957), .A2(n5956), .ZN(n5959) );
  NAND2_X1 U5412 ( .A1(n5288), .A2(n4546), .ZN(n5084) );
  NAND2_X1 U5413 ( .A1(n5754), .A2(n5139), .ZN(n5756) );
  INV_X1 U5414 ( .A(n5554), .ZN(n5032) );
  AND2_X1 U5415 ( .A1(n5376), .A2(n5283), .ZN(n5072) );
  NOR2_X1 U5416 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5365) );
  NOR2_X1 U5417 ( .A1(n6088), .A2(n6087), .ZN(n6111) );
  OR2_X1 U5418 ( .A1(n9249), .A2(n9250), .ZN(n6580) );
  AND2_X1 U5419 ( .A1(n8043), .A2(n6533), .ZN(n7946) );
  NAND2_X1 U5420 ( .A1(n9204), .A2(n4639), .ZN(n4637) );
  AND2_X1 U5421 ( .A1(n9204), .A2(n4556), .ZN(n4635) );
  NAND2_X1 U5422 ( .A1(n4919), .A2(n4568), .ZN(n9227) );
  OR2_X1 U5423 ( .A1(n9171), .A2(n9225), .ZN(n4920) );
  NAND2_X1 U5424 ( .A1(n8162), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4845) );
  INV_X2 U5425 ( .A(n6469), .ZN(n6786) );
  XNOR2_X1 U5426 ( .A(n6456), .B(n6546), .ZN(n6457) );
  NAND2_X1 U5427 ( .A1(n6411), .A2(n8082), .ZN(n6437) );
  AND2_X1 U5428 ( .A1(n8036), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U5429 ( .A1(n7044), .A2(n7045), .ZN(n4866) );
  NOR2_X1 U5430 ( .A1(n8216), .A2(n4609), .ZN(n7058) );
  OR2_X1 U5431 ( .A1(n9331), .A2(n9330), .ZN(n4862) );
  AND2_X1 U5432 ( .A1(n4862), .A2(n4861), .ZN(n9341) );
  NAND2_X1 U5433 ( .A1(n7006), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4861) );
  OR2_X1 U5434 ( .A1(n9341), .A2(n9340), .ZN(n4860) );
  AND2_X1 U5435 ( .A1(n4860), .A2(n4859), .ZN(n6999) );
  NAND2_X1 U5436 ( .A1(n9344), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4859) );
  NOR2_X1 U5437 ( .A1(n8191), .A2(n8190), .ZN(n9371) );
  NAND2_X1 U5438 ( .A1(n4858), .A2(n4857), .ZN(n9457) );
  AOI21_X1 U5439 ( .B1(n4542), .B2(n9421), .A(n4617), .ZN(n4857) );
  NAND2_X1 U5440 ( .A1(n8160), .A2(n8159), .ZN(n9472) );
  NAND2_X1 U5441 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  INV_X1 U5442 ( .A(n6385), .ZN(n4835) );
  NOR2_X1 U5443 ( .A1(n6382), .A2(n4841), .ZN(n4840) );
  INV_X1 U5444 ( .A(n6380), .ZN(n4841) );
  AND2_X1 U5445 ( .A1(n8492), .A2(n8330), .ZN(n9514) );
  INV_X1 U5446 ( .A(n4757), .ZN(n4756) );
  OAI21_X1 U5447 ( .B1(n4758), .B2(n8318), .A(n9546), .ZN(n4757) );
  AND2_X1 U5448 ( .A1(n8403), .A2(n8410), .ZN(n9546) );
  NAND2_X1 U5449 ( .A1(n6261), .A2(n4758), .ZN(n9561) );
  INV_X1 U5450 ( .A(n9575), .ZN(n4831) );
  AND2_X1 U5451 ( .A1(n8313), .A2(n8397), .ZN(n9574) );
  OR2_X2 U5452 ( .A1(n4716), .A2(n7961), .ZN(n8024) );
  NAND2_X1 U5453 ( .A1(n7897), .A2(n6361), .ZN(n4625) );
  NAND2_X1 U5454 ( .A1(n8464), .A2(n8267), .ZN(n8379) );
  NAND2_X1 U5455 ( .A1(n6132), .A2(n6131), .ZN(n7944) );
  OR2_X1 U5456 ( .A1(n7024), .A2(n6071), .ZN(n6132) );
  INV_X1 U5457 ( .A(n8376), .ZN(n7681) );
  INV_X1 U5458 ( .A(n10352), .ZN(n7484) );
  AOI21_X1 U5459 ( .B1(n4818), .B2(n4820), .A(n4571), .ZN(n4816) );
  NAND2_X1 U5460 ( .A1(n10247), .A2(n8445), .ZN(n6007) );
  AND4_X1 U5461 ( .A1(n6331), .A2(n6332), .A3(n6333), .A4(n6330), .ZN(n10265)
         );
  NAND2_X1 U5462 ( .A1(n6256), .A2(n6255), .ZN(n9576) );
  NAND2_X1 U5463 ( .A1(n6226), .A2(n6225), .ZN(n8129) );
  OR2_X1 U5464 ( .A1(n7074), .A2(n6071), .ZN(n6143) );
  AND2_X1 U5465 ( .A1(n6073), .A2(n6072), .ZN(n10326) );
  OAI211_X1 U5466 ( .C1(n6013), .C2(n4709), .A(n6018), .B(n6017), .ZN(n10303)
         );
  OAI21_X1 U5467 ( .B1(n5719), .B2(n5275), .A(n5274), .ZN(n5729) );
  OR2_X1 U5468 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  XNOR2_X1 U5469 ( .A(n5729), .B(n5728), .ZN(n8532) );
  INV_X1 U5470 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U5471 ( .A1(n6402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5472 ( .A1(n6311), .A2(n4814), .ZN(n6402) );
  OAI21_X1 U5473 ( .B1(n4974), .B2(n4972), .A(n5242), .ZN(n4971) );
  INV_X1 U5474 ( .A(n5238), .ZN(n4972) );
  INV_X1 U5475 ( .A(n4974), .ZN(n4973) );
  NAND2_X1 U5476 ( .A1(n6313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U5477 ( .B1(n5622), .B2(n5238), .A(n5237), .ZN(n5632) );
  NAND2_X1 U5478 ( .A1(n5505), .A2(n5209), .ZN(n5519) );
  AOI21_X1 U5479 ( .B1(n4945), .B2(n4947), .A(n4579), .ZN(n4944) );
  OR2_X1 U5480 ( .A1(n5454), .A2(n4946), .ZN(n4943) );
  INV_X1 U5481 ( .A(n4947), .ZN(n4946) );
  NAND2_X1 U5482 ( .A1(n4943), .A2(n4941), .ZN(n5489) );
  AND2_X1 U5483 ( .A1(n4944), .A2(n4942), .ZN(n4941) );
  INV_X1 U5484 ( .A(n5486), .ZN(n4942) );
  NAND2_X1 U5485 ( .A1(n5458), .A2(n5198), .ZN(n5468) );
  AND2_X1 U5486 ( .A1(n5190), .A2(n5189), .ZN(n5420) );
  AND2_X1 U5487 ( .A1(n5181), .A2(n5180), .ZN(n5378) );
  AND2_X1 U5488 ( .A1(n6040), .A2(n6032), .ZN(n7013) );
  NAND2_X1 U5489 ( .A1(n5330), .A2(n5331), .ZN(n5335) );
  OR2_X1 U5490 ( .A1(n6002), .A2(n6103), .ZN(n6029) );
  OAI21_X1 U5491 ( .B1(n4666), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4669), .ZN(
        n5314) );
  NAND2_X1 U5492 ( .A1(n8151), .A2(n6937), .ZN(n4669) );
  NAND2_X1 U5493 ( .A1(n5697), .A2(n5696), .ZN(n5706) );
  AND3_X1 U5494 ( .A1(n5618), .A2(n5617), .A3(n5616), .ZN(n8978) );
  NOR2_X1 U5495 ( .A1(n4534), .A2(n8711), .ZN(n5034) );
  NAND2_X1 U5496 ( .A1(n5037), .A2(n5042), .ZN(n5036) );
  NAND2_X1 U5497 ( .A1(n8570), .A2(n4528), .ZN(n5042) );
  AND4_X1 U5498 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n7714)
         );
  AND4_X1 U5499 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n8697)
         );
  NAND2_X1 U5500 ( .A1(n8565), .A2(n8564), .ZN(n8701) );
  AND2_X1 U5501 ( .A1(n5946), .A2(n5945), .ZN(n4736) );
  AND2_X1 U5502 ( .A1(n5745), .A2(n5726), .ZN(n8862) );
  INV_X1 U5503 ( .A(n8526), .ZN(n8895) );
  XNOR2_X1 U5504 ( .A(n6709), .B(n7563), .ZN(n7551) );
  NOR2_X1 U5505 ( .A1(n7551), .A2(n10562), .ZN(n7550) );
  OAI211_X1 U5506 ( .C1(n7672), .C2(n4888), .A(n4887), .B(n4884), .ZN(n7736)
         );
  INV_X1 U5507 ( .A(n4889), .ZN(n4888) );
  NOR2_X1 U5508 ( .A1(n4885), .A2(n4531), .ZN(n4884) );
  NOR2_X1 U5509 ( .A1(n7736), .A2(n7824), .ZN(n7735) );
  XNOR2_X1 U5510 ( .A(n6681), .B(n8754), .ZN(n8741) );
  NAND2_X1 U5511 ( .A1(n5598), .A2(n5597), .ZN(n8984) );
  NAND2_X1 U5512 ( .A1(n5081), .A2(n6844), .ZN(n9082) );
  INV_X1 U5513 ( .A(n8995), .ZN(n5081) );
  NAND2_X1 U5514 ( .A1(n5583), .A2(n5582), .ZN(n8994) );
  OAI211_X1 U5515 ( .C1(n6866), .C2(n6935), .A(n5407), .B(n5406), .ZN(n10505)
         );
  NAND2_X1 U5516 ( .A1(n5647), .A2(n5646), .ZN(n9124) );
  NAND2_X1 U5517 ( .A1(n5569), .A2(n5568), .ZN(n9151) );
  INV_X1 U5518 ( .A(n6801), .ZN(n6796) );
  NAND2_X2 U5519 ( .A1(n6263), .A2(n6262), .ZN(n6378) );
  OR2_X1 U5520 ( .A1(n6284), .A2(n6283), .ZN(n9649) );
  OR2_X1 U5521 ( .A1(n6276), .A2(n6275), .ZN(n9658) );
  OR2_X1 U5522 ( .A1(n9422), .A2(n9421), .ZN(n9440) );
  NAND2_X1 U5523 ( .A1(n7726), .A2(n8464), .ZN(n10203) );
  INV_X1 U5524 ( .A(n6013), .ZN(n4843) );
  INV_X1 U5525 ( .A(n8154), .ZN(n8155) );
  NOR2_X1 U5526 ( .A1(n5976), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5977) );
  INV_X1 U5527 ( .A(n4723), .ZN(n5988) );
  NAND2_X1 U5528 ( .A1(n5832), .A2(n5843), .ZN(n4740) );
  NAND2_X1 U5529 ( .A1(n5845), .A2(n4661), .ZN(n5850) );
  OAI21_X1 U5530 ( .B1(n4561), .B2(n6884), .A(n4663), .ZN(n4662) );
  OAI211_X1 U5531 ( .C1(n8252), .C2(n4688), .A(n4687), .B(n4686), .ZN(n4685)
         );
  NAND2_X1 U5532 ( .A1(n4569), .A2(n4689), .ZN(n4688) );
  INV_X1 U5533 ( .A(n8253), .ZN(n4686) );
  NAND2_X1 U5534 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  AOI21_X1 U5535 ( .B1(n8272), .B2(n8453), .A(n8271), .ZN(n8277) );
  NOR2_X1 U5536 ( .A1(n8282), .A2(n8468), .ZN(n4696) );
  NAND2_X1 U5537 ( .A1(n5877), .A2(n5873), .ZN(n4742) );
  OAI21_X1 U5538 ( .B1(n4678), .B2(n5873), .A(n5875), .ZN(n5886) );
  OAI21_X1 U5539 ( .B1(n8288), .B2(n8289), .A(n4690), .ZN(n8293) );
  AOI21_X1 U5540 ( .B1(n4693), .B2(n8508), .A(n4691), .ZN(n4690) );
  INV_X1 U5541 ( .A(n5894), .ZN(n4659) );
  NAND2_X1 U5542 ( .A1(n5897), .A2(n6884), .ZN(n4733) );
  INV_X1 U5543 ( .A(n8938), .ZN(n4734) );
  AOI21_X1 U5544 ( .B1(n4698), .B2(n4697), .A(n4580), .ZN(n8325) );
  AOI21_X1 U5545 ( .B1(n8316), .B2(n8508), .A(n9557), .ZN(n4697) );
  NAND2_X1 U5546 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  AND2_X1 U5547 ( .A1(n8326), .A2(n8322), .ZN(n8323) );
  NOR2_X1 U5548 ( .A1(n5128), .A2(n4983), .ZN(n4982) );
  INV_X1 U5549 ( .A(n5914), .ZN(n4984) );
  OR2_X1 U5550 ( .A1(n5913), .A2(n6884), .ZN(n4983) );
  NAND2_X1 U5551 ( .A1(n5917), .A2(n5790), .ZN(n5791) );
  OR2_X1 U5552 ( .A1(n5786), .A2(n5785), .ZN(n5792) );
  INV_X1 U5553 ( .A(n5916), .ZN(n5793) );
  INV_X1 U5554 ( .A(n5907), .ZN(n4682) );
  NAND2_X1 U5555 ( .A1(n5520), .A2(SI_14_), .ZN(n4981) );
  NOR2_X1 U5556 ( .A1(n5706), .A2(n8886), .ZN(n5788) );
  NAND2_X1 U5557 ( .A1(n10526), .A2(n8734), .ZN(n5849) );
  INV_X1 U5558 ( .A(n9013), .ZN(n4806) );
  AOI21_X1 U5559 ( .B1(n7643), .B2(n5089), .A(n4578), .ZN(n5088) );
  INV_X1 U5560 ( .A(n5826), .ZN(n5089) );
  INV_X1 U5561 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4792) );
  INV_X1 U5562 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5286) );
  AND2_X1 U5563 ( .A1(n4934), .A2(n4932), .ZN(n4931) );
  INV_X1 U5564 ( .A(n6511), .ZN(n4932) );
  INV_X1 U5565 ( .A(n4937), .ZN(n4929) );
  INV_X1 U5566 ( .A(n6510), .ZN(n4928) );
  OAI21_X1 U5567 ( .B1(n8339), .B2(n8338), .A(n8419), .ZN(n8342) );
  AOI21_X1 U5568 ( .B1(n8337), .B2(n8496), .A(n8336), .ZN(n8339) );
  NOR2_X1 U5569 ( .A1(n8423), .A2(n8422), .ZN(n8497) );
  OR2_X1 U5570 ( .A1(n9480), .A2(n9496), .ZN(n8419) );
  AND2_X1 U5571 ( .A1(n9532), .A2(n9196), .ZN(n8321) );
  AND2_X1 U5572 ( .A1(n9541), .A2(n9559), .ZN(n8320) );
  AND2_X1 U5573 ( .A1(n7961), .A2(n8092), .ZN(n8289) );
  INV_X1 U5574 ( .A(n4954), .ZN(n4953) );
  OAI21_X1 U5575 ( .B1(n5670), .B2(n4955), .A(n5682), .ZN(n4954) );
  INV_X1 U5576 ( .A(n5258), .ZN(n4955) );
  INV_X1 U5577 ( .A(n4971), .ZN(n4967) );
  OAI21_X1 U5578 ( .B1(n4971), .B2(n4973), .A(n5644), .ZN(n4970) );
  INV_X1 U5579 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5967) );
  AOI21_X1 U5580 ( .B1(n4528), .B2(n5044), .A(n4583), .ZN(n5043) );
  INV_X1 U5581 ( .A(n8702), .ZN(n5044) );
  INV_X1 U5582 ( .A(n8621), .ZN(n5063) );
  XNOR2_X1 U5583 ( .A(n8556), .B(n10489), .ZN(n7319) );
  XNOR2_X1 U5584 ( .A(n8556), .B(n10485), .ZN(n7315) );
  INV_X1 U5585 ( .A(n7254), .ZN(n4883) );
  AOI21_X1 U5586 ( .B1(n7227), .B2(n7298), .A(n7299), .ZN(n7297) );
  AOI21_X1 U5587 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6959), .A(n7661), .ZN(
        n6711) );
  AOI21_X1 U5588 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6952), .A(n7410), .ZN(
        n6676) );
  AND3_X1 U5589 ( .A1(n4999), .A2(n4997), .A3(n4613), .ZN(n6714) );
  AOI21_X1 U5590 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7238), .A(n8763), .ZN(
        n6716) );
  INV_X1 U5591 ( .A(n5788), .ZN(n5131) );
  NAND2_X1 U5592 ( .A1(n5698), .A2(n9846), .ZN(n5712) );
  INV_X1 U5593 ( .A(n6848), .ZN(n4796) );
  OAI21_X1 U5594 ( .B1(n4799), .B2(n4796), .A(n8948), .ZN(n4795) );
  NAND2_X1 U5595 ( .A1(n10441), .A2(n7168), .ZN(n5819) );
  AND2_X1 U5596 ( .A1(n5911), .A2(n8913), .ZN(n5907) );
  NAND2_X1 U5597 ( .A1(n5133), .A2(n4806), .ZN(n4804) );
  NAND2_X1 U5598 ( .A1(n4806), .A2(n5134), .ZN(n4805) );
  NAND2_X1 U5599 ( .A1(n5103), .A2(n5106), .ZN(n5099) );
  NOR2_X1 U5600 ( .A1(n5880), .A2(n5102), .ZN(n5101) );
  INV_X1 U5601 ( .A(n5103), .ZN(n5102) );
  NAND2_X1 U5602 ( .A1(n5292), .A2(n5110), .ZN(n5954) );
  AND2_X1 U5603 ( .A1(n5291), .A2(n5111), .ZN(n5110) );
  INV_X1 U5604 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5111) );
  INV_X1 U5605 ( .A(n5292), .ZN(n5777) );
  NAND2_X1 U5606 ( .A1(n5032), .A2(n5031), .ZN(n5751) );
  AND2_X1 U5607 ( .A1(n5566), .A2(n5581), .ZN(n5031) );
  INV_X1 U5608 ( .A(n7174), .ZN(n4649) );
  NAND2_X1 U5609 ( .A1(n8439), .A2(n8512), .ZN(n6433) );
  AOI21_X1 U5610 ( .B1(n8042), .B2(n4909), .A(n4908), .ZN(n4907) );
  INV_X1 U5611 ( .A(n8043), .ZN(n4909) );
  INV_X1 U5612 ( .A(n6539), .ZN(n4908) );
  AND2_X1 U5613 ( .A1(n8331), .A2(n8330), .ZN(n8496) );
  NOR2_X1 U5614 ( .A1(n6387), .A2(n4726), .ZN(n4725) );
  INV_X1 U5615 ( .A(n4727), .ZN(n4726) );
  NAND2_X1 U5616 ( .A1(n8419), .A2(n8421), .ZN(n8338) );
  NOR2_X1 U5617 ( .A1(n4839), .A2(n6385), .ZN(n4838) );
  INV_X1 U5618 ( .A(n4840), .ZN(n4839) );
  NAND2_X1 U5619 ( .A1(n6386), .A2(n6383), .ZN(n4836) );
  INV_X1 U5620 ( .A(n8321), .ZN(n8488) );
  OR2_X1 U5621 ( .A1(n9576), .A2(n9590), .ZN(n8313) );
  AND2_X1 U5622 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n6241), .ZN(n6248) );
  NOR2_X1 U5623 ( .A1(n4766), .A2(n9620), .ZN(n4765) );
  NOR2_X1 U5624 ( .A1(n4767), .A2(n6232), .ZN(n4766) );
  INV_X1 U5625 ( .A(n6369), .ZN(n4851) );
  AND2_X1 U5626 ( .A1(n8385), .A2(n8294), .ZN(n4767) );
  NOR2_X1 U5627 ( .A1(n9275), .A2(n8129), .ZN(n4720) );
  INV_X1 U5628 ( .A(n6362), .ZN(n4848) );
  INV_X1 U5629 ( .A(n8289), .ZN(n8476) );
  AND2_X1 U5630 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(n6182), .ZN(n6195) );
  OR2_X1 U5631 ( .A1(n6094), .A2(n6093), .ZN(n8452) );
  INV_X1 U5632 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U5633 ( .B1(n10225), .B2(n4820), .A(n7639), .ZN(n4819) );
  INV_X1 U5634 ( .A(n6350), .ZN(n4820) );
  AND2_X1 U5635 ( .A1(n6346), .A2(n6344), .ZN(n4824) );
  NOR2_X1 U5636 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  INV_X1 U5637 ( .A(n9306), .ZN(n6470) );
  NAND2_X1 U5638 ( .A1(n9539), .A2(n9724), .ZN(n9529) );
  AND2_X1 U5639 ( .A1(n4718), .A2(n9740), .ZN(n4717) );
  NAND2_X1 U5640 ( .A1(n7730), .A2(n10383), .ZN(n10212) );
  NAND2_X1 U5641 ( .A1(n5271), .A2(n5270), .ZN(n5273) );
  INV_X1 U5642 ( .A(n4960), .ZN(n4959) );
  OAI21_X1 U5643 ( .B1(n4962), .B2(n5227), .A(n5226), .ZN(n4960) );
  INV_X1 U5644 ( .A(n5181), .ZN(n4979) );
  CLKBUF_X1 U5645 ( .A(n6046), .Z(n6047) );
  OAI21_X1 U5646 ( .B1(n8151), .B2(n4665), .A(n4664), .ZN(n5182) );
  INV_X1 U5647 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5648 ( .A1(n8151), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4664) );
  OR2_X1 U5649 ( .A1(n5161), .A2(n5169), .ZN(n4708) );
  NAND2_X1 U5650 ( .A1(n5170), .A2(SI_3_), .ZN(n5172) );
  INV_X1 U5651 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5384) );
  INV_X1 U5652 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9941) );
  INV_X1 U5653 ( .A(n5068), .ZN(n5067) );
  OAI21_X1 U5654 ( .B1(n4545), .B2(n5069), .A(n7982), .ZN(n5068) );
  INV_X1 U5655 ( .A(n5043), .ZN(n5039) );
  NAND2_X1 U5656 ( .A1(n5625), .A2(n9786), .ZN(n5635) );
  INV_X1 U5657 ( .A(n5626), .ZN(n5625) );
  NAND2_X1 U5658 ( .A1(n8710), .A2(n5055), .ZN(n5053) );
  AND2_X1 U5659 ( .A1(n4537), .A2(n8682), .ZN(n5057) );
  NAND2_X1 U5660 ( .A1(n9833), .A2(n9941), .ZN(n5386) );
  OAI21_X1 U5661 ( .B1(n8672), .B2(n8671), .A(n8670), .ZN(n8669) );
  NAND2_X1 U5662 ( .A1(n5071), .A2(n7929), .ZN(n5070) );
  XNOR2_X1 U5663 ( .A(n7791), .B(n7820), .ZN(n7768) );
  NAND2_X1 U5664 ( .A1(n5048), .A2(n5046), .ZN(n8690) );
  AOI21_X1 U5665 ( .B1(n5049), .B2(n5050), .A(n5047), .ZN(n5046) );
  INV_X1 U5666 ( .A(n8691), .ZN(n5047) );
  OR2_X1 U5667 ( .A1(n5934), .A2(n5146), .ZN(n5137) );
  NAND2_X1 U5668 ( .A1(n5928), .A2(n8602), .ZN(n5935) );
  AND4_X1 U5669 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(n8638)
         );
  CLKBUF_X3 U5670 ( .A(n4523), .Z(n5734) );
  OR2_X1 U5671 ( .A1(n7266), .A2(n10548), .ZN(n7264) );
  NOR2_X1 U5672 ( .A1(n6672), .A2(n4881), .ZN(n7228) );
  NAND2_X1 U5673 ( .A1(n4622), .A2(n6704), .ZN(n7303) );
  OAI21_X1 U5674 ( .B1(n4996), .B2(n6704), .A(n4994), .ZN(n7305) );
  AOI21_X1 U5675 ( .B1(n7302), .B2(n4995), .A(n4623), .ZN(n4994) );
  NAND2_X1 U5676 ( .A1(n4900), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4899) );
  AND2_X1 U5677 ( .A1(n4899), .A2(n4898), .ZN(n7412) );
  NOR2_X1 U5678 ( .A1(n7412), .A2(n7411), .ZN(n7410) );
  NOR2_X1 U5679 ( .A1(n7357), .A2(n10558), .ZN(n7358) );
  XNOR2_X1 U5680 ( .A(n6676), .B(n7563), .ZN(n7559) );
  INV_X1 U5681 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5469) );
  NOR2_X1 U5682 ( .A1(n4891), .A2(n4886), .ZN(n4885) );
  INV_X1 U5683 ( .A(n7671), .ZN(n4886) );
  AOI21_X1 U5684 ( .B1(n7671), .B2(n4890), .A(n7745), .ZN(n4889) );
  INV_X1 U5685 ( .A(n5019), .ZN(n8780) );
  INV_X1 U5686 ( .A(n6720), .ZN(n5004) );
  NAND2_X1 U5687 ( .A1(n5003), .A2(n5002), .ZN(n8833) );
  NAND2_X1 U5688 ( .A1(n5006), .A2(n4620), .ZN(n5003) );
  OR2_X1 U5689 ( .A1(n5712), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8850) );
  NOR2_X1 U5690 ( .A1(n8862), .A2(n10454), .ZN(n8863) );
  NAND2_X1 U5691 ( .A1(n4771), .A2(n4770), .ZN(n6859) );
  NOR2_X1 U5692 ( .A1(n4773), .A2(n4558), .ZN(n4770) );
  OR2_X1 U5693 ( .A1(n5686), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U5694 ( .A1(n5674), .A2(n5673), .ZN(n5686) );
  INV_X1 U5695 ( .A(n5675), .ZN(n5674) );
  NAND2_X1 U5696 ( .A1(n5660), .A2(n9920), .ZN(n5675) );
  INV_X1 U5697 ( .A(n5661), .ZN(n5660) );
  NAND2_X1 U5698 ( .A1(n5600), .A2(n5599), .ZN(n5614) );
  INV_X1 U5699 ( .A(n5601), .ZN(n5600) );
  NAND2_X1 U5700 ( .A1(n5570), .A2(n9974), .ZN(n5584) );
  INV_X1 U5701 ( .A(n5571), .ZN(n5570) );
  OR2_X1 U5702 ( .A1(n5558), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U5703 ( .A1(n5543), .A2(n10098), .ZN(n5558) );
  INV_X1 U5704 ( .A(n5544), .ZN(n5543) );
  OR2_X1 U5705 ( .A1(n5530), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U5706 ( .A1(n5494), .A2(n5493), .ZN(n5511) );
  INV_X1 U5707 ( .A(n5495), .ZN(n5494) );
  NAND2_X1 U5708 ( .A1(n5510), .A2(n9950), .ZN(n5530) );
  INV_X1 U5709 ( .A(n5511), .ZN(n5510) );
  AND2_X1 U5710 ( .A1(n5856), .A2(n5855), .ZN(n7922) );
  NAND2_X1 U5711 ( .A1(n5090), .A2(n5091), .ZN(n7923) );
  AOI21_X1 U5712 ( .B1(n5092), .B2(n4533), .A(n5847), .ZN(n5091) );
  AOI21_X1 U5713 ( .B1(n7711), .B2(n5094), .A(n5764), .ZN(n5092) );
  INV_X1 U5714 ( .A(n5094), .ZN(n5093) );
  INV_X1 U5715 ( .A(n4784), .ZN(n4783) );
  NAND2_X1 U5716 ( .A1(n5410), .A2(n5409), .ZN(n5430) );
  INV_X1 U5717 ( .A(n5411), .ZN(n5410) );
  NAND2_X1 U5718 ( .A1(n10500), .A2(n5826), .ZN(n7647) );
  NAND2_X1 U5719 ( .A1(n7647), .A2(n7643), .ZN(n7699) );
  OAI21_X1 U5720 ( .B1(n7369), .B2(n6820), .A(n6819), .ZN(n6823) );
  AND2_X1 U5721 ( .A1(n5828), .A2(n5826), .ZN(n9042) );
  OR2_X1 U5722 ( .A1(n5392), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U5723 ( .A1(n5385), .A2(n5384), .ZN(n5392) );
  INV_X1 U5724 ( .A(n5386), .ZN(n5385) );
  NAND2_X1 U5725 ( .A1(n6815), .A2(n6814), .ZN(n10424) );
  NAND2_X1 U5726 ( .A1(n5721), .A2(n5720), .ZN(n6896) );
  OR2_X1 U5727 ( .A1(n5903), .A2(n5759), .ZN(n8922) );
  NAND2_X1 U5728 ( .A1(n5640), .A2(n5619), .ZN(n5075) );
  INV_X1 U5729 ( .A(n9010), .ZN(n9015) );
  AND2_X1 U5730 ( .A1(n5879), .A2(n5871), .ZN(n9010) );
  INV_X1 U5731 ( .A(n4802), .ZN(n9014) );
  OAI21_X1 U5732 ( .B1(n7919), .B2(n4803), .A(n4807), .ZN(n4802) );
  INV_X1 U5733 ( .A(n5134), .ZN(n4803) );
  AND4_X1 U5734 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(n8718)
         );
  NAND2_X1 U5735 ( .A1(n7709), .A2(n5843), .ZN(n7777) );
  AND2_X1 U5736 ( .A1(n7081), .A2(n6979), .ZN(n7097) );
  AND2_X1 U5737 ( .A1(n5291), .A2(n5113), .ZN(n5112) );
  NOR2_X1 U5738 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5113) );
  OR2_X1 U5739 ( .A1(n5400), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U5740 ( .A1(n6228), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6235) );
  AND2_X1 U5741 ( .A1(n6625), .A2(n6624), .ZN(n6798) );
  NOR2_X1 U5742 ( .A1(n6235), .A2(n9252), .ZN(n6241) );
  AOI21_X1 U5743 ( .B1(n4924), .B2(n4926), .A(n4552), .ZN(n4923) );
  NOR2_X1 U5744 ( .A1(n4633), .A2(n6552), .ZN(n4632) );
  INV_X1 U5745 ( .A(n4637), .ZN(n4633) );
  AND2_X1 U5746 ( .A1(n6611), .A2(n6610), .ZN(n9226) );
  INV_X1 U5747 ( .A(n9236), .ZN(n6474) );
  INV_X1 U5748 ( .A(n9235), .ZN(n6475) );
  NAND2_X1 U5749 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  INV_X1 U5750 ( .A(n7175), .ZN(n4650) );
  NAND2_X1 U5751 ( .A1(n7458), .A2(n4937), .ZN(n4933) );
  NAND2_X1 U5752 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  NAND2_X1 U5753 ( .A1(n6516), .A2(n7879), .ZN(n4911) );
  INV_X1 U5754 ( .A(n6591), .ZN(n6592) );
  AND2_X1 U5755 ( .A1(n6450), .A2(n6449), .ZN(n7025) );
  NAND2_X1 U5756 ( .A1(n6457), .A2(n6458), .ZN(n6459) );
  AND2_X1 U5757 ( .A1(n6213), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U5758 ( .A1(n8358), .A2(n8357), .ZN(n8509) );
  NAND2_X1 U5759 ( .A1(n8162), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U5760 ( .A1(n6171), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U5761 ( .A1(n4866), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U5762 ( .A1(n6990), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4865) );
  NOR2_X1 U5763 ( .A1(n7126), .A2(n4600), .ZN(n7130) );
  NOR2_X1 U5764 ( .A1(n7130), .A2(n7129), .ZN(n7215) );
  NOR2_X1 U5765 ( .A1(n7215), .A2(n4863), .ZN(n7217) );
  AND2_X1 U5766 ( .A1(n7216), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5767 ( .A1(n7217), .A2(n7218), .ZN(n7336) );
  NOR2_X1 U5768 ( .A1(n8186), .A2(n4867), .ZN(n8199) );
  AND2_X1 U5769 ( .A1(n8187), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5770 ( .A1(n8199), .A2(n8200), .ZN(n8198) );
  NOR2_X1 U5771 ( .A1(n9359), .A2(n4856), .ZN(n8191) );
  AND2_X1 U5772 ( .A1(n8189), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4856) );
  AOI21_X1 U5773 ( .B1(n4855), .B2(n9373), .A(n9396), .ZN(n9374) );
  NAND2_X1 U5774 ( .A1(n9539), .A2(n4725), .ZN(n9498) );
  INV_X1 U5775 ( .A(n9488), .ZN(n9501) );
  AOI21_X1 U5776 ( .B1(n6377), .B2(n4829), .A(n4535), .ZN(n4828) );
  NOR2_X1 U5777 ( .A1(n6378), .A2(n9572), .ZN(n9552) );
  NAND2_X1 U5778 ( .A1(n9591), .A2(n6396), .ZN(n9592) );
  OR2_X1 U5779 ( .A1(n9592), .A2(n9576), .ZN(n9572) );
  INV_X1 U5780 ( .A(n4763), .ZN(n4762) );
  AOI21_X1 U5781 ( .B1(n4765), .B2(n6232), .A(n4764), .ZN(n4763) );
  INV_X1 U5782 ( .A(n8305), .ZN(n4764) );
  AOI21_X1 U5783 ( .B1(n8056), .B2(n4767), .A(n6232), .ZN(n9621) );
  AND2_X1 U5784 ( .A1(n8296), .A2(n8484), .ZN(n8385) );
  NAND2_X1 U5785 ( .A1(n8023), .A2(n6395), .ZN(n8128) );
  NAND2_X1 U5786 ( .A1(n7730), .A2(n4715), .ZN(n10213) );
  AND2_X1 U5787 ( .A1(n4715), .A2(n4714), .ZN(n4713) );
  OR2_X1 U5788 ( .A1(n6144), .A2(n9352), .ZN(n6160) );
  NAND2_X1 U5789 ( .A1(n6150), .A2(n6149), .ZN(n7726) );
  INV_X1 U5790 ( .A(n8379), .ZN(n6149) );
  NOR2_X1 U5791 ( .A1(n7685), .A2(n7944), .ZN(n7730) );
  OR2_X1 U5792 ( .A1(n7588), .A2(n10362), .ZN(n7685) );
  AND2_X1 U5793 ( .A1(n10226), .A2(n10338), .ZN(n10228) );
  OR2_X1 U5794 ( .A1(n6064), .A2(n6053), .ZN(n6088) );
  INV_X1 U5795 ( .A(n10332), .ZN(n7497) );
  NOR2_X1 U5796 ( .A1(n7520), .A2(n7497), .ZN(n10226) );
  OR2_X1 U5797 ( .A1(n10239), .A2(n8236), .ZN(n7519) );
  OR2_X1 U5798 ( .A1(n7519), .A2(n8240), .ZN(n7520) );
  NAND2_X1 U5799 ( .A1(n10257), .A2(n10298), .ZN(n10256) );
  NOR2_X1 U5800 ( .A1(n10256), .A2(n10303), .ZN(n10240) );
  INV_X1 U5801 ( .A(n10266), .ZN(n4760) );
  INV_X1 U5802 ( .A(n8361), .ZN(n4761) );
  OR2_X1 U5803 ( .A1(n10366), .A2(n8439), .ZN(n6635) );
  OR2_X1 U5804 ( .A1(n8508), .A2(n6390), .ZN(n10366) );
  AND3_X1 U5805 ( .A1(n6035), .A2(n6034), .A3(n6033), .ZN(n10311) );
  NAND2_X1 U5806 ( .A1(n7471), .A2(n10366), .ZN(n10385) );
  XNOR2_X1 U5807 ( .A(n5719), .B(SI_29_), .ZN(n9163) );
  NAND2_X1 U5808 ( .A1(n4952), .A2(n5258), .ZN(n5683) );
  NAND2_X1 U5809 ( .A1(n6318), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6317) );
  AND2_X1 U5810 ( .A1(n4958), .A2(n4962), .ZN(n5579) );
  AOI21_X1 U5811 ( .B1(n5436), .B2(n4671), .A(n4581), .ZN(n4670) );
  NAND2_X1 U5812 ( .A1(n4673), .A2(n5436), .ZN(n4672) );
  AND2_X1 U5813 ( .A1(n5176), .A2(n5177), .ZN(n5369) );
  NAND2_X1 U5814 ( .A1(n5335), .A2(n5168), .ZN(n5351) );
  NAND2_X1 U5815 ( .A1(n5167), .A2(n4746), .ZN(n5331) );
  NAND2_X1 U5816 ( .A1(n4707), .A2(n5166), .ZN(n5167) );
  AND2_X1 U5817 ( .A1(n5160), .A2(n5168), .ZN(n5330) );
  AND2_X1 U5818 ( .A1(n7112), .A2(n7145), .ZN(n7116) );
  NAND2_X1 U5819 ( .A1(n5058), .A2(n5059), .ZN(n8623) );
  NAND2_X1 U5820 ( .A1(n5053), .A2(n5054), .ZN(n8644) );
  AND2_X1 U5821 ( .A1(n7318), .A2(n7317), .ZN(n8659) );
  NAND2_X1 U5822 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  NAND2_X1 U5823 ( .A1(n5066), .A2(n5070), .ZN(n7984) );
  NAND2_X1 U5824 ( .A1(n7866), .A2(n4545), .ZN(n5066) );
  NAND2_X1 U5825 ( .A1(n5634), .A2(n5633), .ZN(n8940) );
  AND2_X1 U5826 ( .A1(n7100), .A2(n7095), .ZN(n8715) );
  OR2_X1 U5827 ( .A1(n7157), .A2(n7156), .ZN(n8720) );
  INV_X1 U5828 ( .A(n8885), .ZN(n8907) );
  INV_X1 U5829 ( .A(n7714), .ZN(n8736) );
  INV_X1 U5830 ( .A(n7394), .ZN(n9035) );
  NAND2_X1 U5831 ( .A1(n5733), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5346) );
  OR2_X1 U5832 ( .A1(n7081), .A2(n7092), .ZN(n8831) );
  NAND2_X1 U5833 ( .A1(n4992), .A2(n4991), .ZN(n7184) );
  NAND2_X1 U5834 ( .A1(n4987), .A2(n6929), .ZN(n4992) );
  NOR2_X1 U5835 ( .A1(n7358), .A2(n6708), .ZN(n7403) );
  NAND2_X1 U5836 ( .A1(n7357), .A2(n5015), .ZN(n5008) );
  INV_X1 U5837 ( .A(n5013), .ZN(n5009) );
  NOR2_X1 U5838 ( .A1(n7550), .A2(n6710), .ZN(n7663) );
  NOR2_X1 U5839 ( .A1(n7663), .A2(n7662), .ZN(n7661) );
  NOR2_X1 U5840 ( .A1(n6679), .A2(n7735), .ZN(n7830) );
  NOR2_X1 U5841 ( .A1(n7670), .A2(n4894), .ZN(n6678) );
  AND2_X1 U5842 ( .A1(n5001), .A2(n5000), .ZN(n7838) );
  NAND2_X1 U5843 ( .A1(n4999), .A2(n4997), .ZN(n7836) );
  NOR2_X1 U5844 ( .A1(n8741), .A2(n8742), .ZN(n8740) );
  OAI21_X1 U5845 ( .B1(n8741), .B2(n4902), .A(n4901), .ZN(n8758) );
  NAND2_X1 U5846 ( .A1(n4903), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4902) );
  INV_X1 U5847 ( .A(n8759), .ZN(n4903) );
  OR2_X1 U5848 ( .A1(n8782), .A2(n8781), .ZN(n5019) );
  INV_X1 U5849 ( .A(n6717), .ZN(n5018) );
  OAI21_X1 U5850 ( .B1(n8782), .B2(n5017), .A(n5016), .ZN(n8792) );
  NAND2_X1 U5851 ( .A1(n5020), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U5852 ( .A1(n6717), .A2(n5020), .ZN(n5016) );
  INV_X1 U5853 ( .A(n8793), .ZN(n5020) );
  NOR2_X1 U5854 ( .A1(n5005), .A2(n6720), .ZN(n8813) );
  NOR2_X1 U5855 ( .A1(n8809), .A2(n8810), .ZN(n8808) );
  NAND2_X1 U5856 ( .A1(n4897), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U5857 ( .A1(n6688), .A2(n4897), .ZN(n4895) );
  INV_X1 U5858 ( .A(n8826), .ZN(n4897) );
  INV_X1 U5859 ( .A(n4809), .ZN(n4808) );
  OAI21_X1 U5860 ( .B1(n8866), .B2(n10459), .A(n8865), .ZN(n9051) );
  NOR2_X1 U5861 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  XNOR2_X1 U5862 ( .A(n8861), .B(n5116), .ZN(n8866) );
  NOR2_X1 U5863 ( .A1(n8886), .A2(n10456), .ZN(n8864) );
  NAND2_X1 U5864 ( .A1(n5117), .A2(n5119), .ZN(n8868) );
  NAND2_X1 U5865 ( .A1(n5122), .A2(n5125), .ZN(n8522) );
  NAND2_X1 U5866 ( .A1(n8900), .A2(n5127), .ZN(n5122) );
  NAND2_X1 U5867 ( .A1(n8960), .A2(n6848), .ZN(n8949) );
  NAND2_X1 U5868 ( .A1(n5624), .A2(n5623), .ZN(n9072) );
  NAND2_X1 U5869 ( .A1(n5462), .A2(n5461), .ZN(n7788) );
  NAND2_X1 U5870 ( .A1(n5443), .A2(n5442), .ZN(n10518) );
  NAND2_X1 U5871 ( .A1(n4782), .A2(n6827), .ZN(n7696) );
  NAND2_X1 U5872 ( .A1(n4787), .A2(n4786), .ZN(n4782) );
  NAND2_X1 U5873 ( .A1(n4787), .A2(n4789), .ZN(n7644) );
  AND2_X1 U5874 ( .A1(n10471), .A2(n7378), .ZN(n10433) );
  INV_X1 U5875 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U5876 ( .A1(n5732), .A2(n5731), .ZN(n9048) );
  INV_X1 U5877 ( .A(n5926), .ZN(n9096) );
  NAND2_X1 U5878 ( .A1(n4772), .A2(n4775), .ZN(n8884) );
  NAND2_X1 U5879 ( .A1(n8900), .A2(n5912), .ZN(n5129) );
  NAND2_X1 U5880 ( .A1(n5672), .A2(n5671), .ZN(n9112) );
  NAND2_X1 U5881 ( .A1(n4776), .A2(n6855), .ZN(n8894) );
  OR2_X1 U5882 ( .A1(n8906), .A2(n6856), .ZN(n4776) );
  NAND2_X1 U5883 ( .A1(n5659), .A2(n5658), .ZN(n9118) );
  NAND2_X1 U5884 ( .A1(n5611), .A2(n5610), .ZN(n9138) );
  NOR2_X1 U5885 ( .A1(n4798), .A2(n4797), .ZN(n8962) );
  INV_X1 U5886 ( .A(n6847), .ZN(n4797) );
  NAND2_X1 U5887 ( .A1(n9082), .A2(n5882), .ZN(n8969) );
  NAND2_X1 U5888 ( .A1(n5557), .A2(n5556), .ZN(n9158) );
  NAND2_X1 U5889 ( .A1(n5542), .A2(n5541), .ZN(n9012) );
  OR2_X1 U5890 ( .A1(n7966), .A2(n5106), .ZN(n5096) );
  NAND2_X1 U5891 ( .A1(n5529), .A2(n5528), .ZN(n8078) );
  NAND2_X1 U5892 ( .A1(n5107), .A2(n5517), .ZN(n8066) );
  OR2_X1 U5893 ( .A1(n7966), .A2(n5518), .ZN(n5107) );
  AND2_X1 U5894 ( .A1(n6908), .A2(n6907), .ZN(n10547) );
  INV_X1 U5895 ( .A(n6871), .ZN(n8099) );
  XNOR2_X1 U5896 ( .A(n5951), .B(n5950), .ZN(n6885) );
  NAND2_X1 U5897 ( .A1(n5959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  NOR2_X1 U5898 ( .A1(n5755), .A2(n5023), .ZN(n5022) );
  OAI21_X1 U5899 ( .B1(n5756), .B2(P2_IR_REG_20__SCAN_IN), .A(n4551), .ZN(
        n5024) );
  NOR2_X1 U5900 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5023) );
  NAND2_X1 U5901 ( .A1(n5756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5902 ( .A1(n5032), .A2(n5566), .ZN(n5580) );
  OR2_X1 U5903 ( .A1(n5401), .A2(n5083), .ZN(n6935) );
  AND3_X1 U5904 ( .A1(n5339), .A2(n5283), .A3(n5365), .ZN(n5375) );
  XNOR2_X1 U5905 ( .A(n5367), .B(n5283), .ZN(n7261) );
  OAI21_X1 U5906 ( .B1(n5338), .B2(n5340), .A(n5337), .ZN(n5341) );
  NAND2_X1 U5907 ( .A1(n5340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5337) );
  INV_X1 U5908 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5156) );
  MUX2_X1 U5909 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5309), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5311) );
  AOI21_X1 U5910 ( .B1(n9193), .B2(n4643), .A(n4641), .ZN(n4640) );
  INV_X1 U5911 ( .A(n4642), .ZN(n4641) );
  AOI21_X1 U5912 ( .B1(n4643), .B2(n4645), .A(n6631), .ZN(n4642) );
  AOI21_X1 U5913 ( .B1(n6619), .B2(n4644), .A(n4553), .ZN(n4643) );
  AND2_X1 U5914 ( .A1(n6109), .A2(n6108), .ZN(n10352) );
  NAND2_X1 U5915 ( .A1(n9179), .A2(n9178), .ZN(n9177) );
  NAND2_X1 U5916 ( .A1(n6567), .A2(n9268), .ZN(n9179) );
  AND2_X1 U5917 ( .A1(n6797), .A2(n9285), .ZN(n6795) );
  AND2_X1 U5918 ( .A1(n6630), .A2(n4940), .ZN(n4939) );
  NAND2_X1 U5919 ( .A1(n6619), .A2(n4644), .ZN(n4940) );
  OAI211_X1 U5920 ( .C1(n9268), .C2(n4925), .A(n4630), .B(n4923), .ZN(n9185)
         );
  OR2_X1 U5921 ( .A1(n6567), .A2(n4925), .ZN(n4630) );
  NAND2_X1 U5922 ( .A1(n4636), .A2(n4638), .ZN(n9203) );
  AND2_X1 U5923 ( .A1(n6483), .A2(n6484), .ZN(n4918) );
  NAND2_X1 U5924 ( .A1(n4608), .A2(n6483), .ZN(n7449) );
  NAND2_X1 U5925 ( .A1(n6192), .A2(n6191), .ZN(n9222) );
  NAND2_X2 U5926 ( .A1(n6085), .A2(n6084), .ZN(n10342) );
  AND4_X1 U5927 ( .A1(n5987), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n7068)
         );
  NAND2_X1 U5928 ( .A1(n6008), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U5929 ( .A1(n6171), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U5930 ( .A1(n9177), .A2(n6574), .ZN(n9248) );
  NAND2_X1 U5931 ( .A1(n4906), .A2(n8042), .ZN(n8045) );
  NAND2_X1 U5932 ( .A1(n7948), .A2(n8043), .ZN(n4906) );
  INV_X1 U5933 ( .A(n6516), .ZN(n4917) );
  OAI22_X1 U5934 ( .A1(n6395), .A2(n6451), .B1(n9181), .B2(n6469), .ZN(n9270)
         );
  NAND2_X1 U5935 ( .A1(n7449), .A2(n6484), .ZN(n7458) );
  NAND2_X1 U5936 ( .A1(n9281), .A2(n6619), .ZN(n9284) );
  OR2_X1 U5937 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  OR2_X1 U5938 ( .A1(n6294), .A2(n6293), .ZN(n9659) );
  OR2_X1 U5939 ( .A1(n6124), .A2(n6123), .ZN(n10373) );
  OR2_X1 U5940 ( .A1(n6115), .A2(n6114), .ZN(n9304) );
  OR2_X1 U5941 ( .A1(n6092), .A2(n6091), .ZN(n10349) );
  NAND4_X1 U5942 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n9308)
         );
  NAND4_X1 U5943 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n7032)
         );
  INV_X1 U5944 ( .A(n4866), .ZN(n7047) );
  AND2_X1 U5945 ( .A1(n6992), .A2(n4864), .ZN(n8216) );
  INV_X1 U5946 ( .A(n4864), .ZN(n8218) );
  INV_X1 U5947 ( .A(n4862), .ZN(n9329) );
  INV_X1 U5948 ( .A(n4860), .ZN(n9339) );
  NOR2_X1 U5949 ( .A1(n7432), .A2(n4868), .ZN(n7436) );
  AND2_X1 U5950 ( .A1(n7433), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U5951 ( .A1(n7436), .A2(n7435), .ZN(n8186) );
  NAND2_X1 U5952 ( .A1(n9440), .A2(n4542), .ZN(n9456) );
  AND2_X1 U5953 ( .A1(n9440), .A2(n9439), .ZN(n9445) );
  AOI21_X1 U5954 ( .B1(n9467), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9466), .ZN(
        n4873) );
  NAND2_X1 U5955 ( .A1(n9463), .A2(n4555), .ZN(n4870) );
  OAI22_X1 U5956 ( .A1(n9461), .A2(n9458), .B1(n9464), .B2(n9459), .ZN(n4874)
         );
  NAND2_X1 U5957 ( .A1(n9491), .A2(n9490), .ZN(n9646) );
  AOI21_X1 U5958 ( .B1(n6381), .B2(n4840), .A(n6384), .ZN(n9505) );
  NAND2_X1 U5959 ( .A1(n6287), .A2(n6286), .ZN(n9513) );
  NAND2_X1 U5960 ( .A1(n6381), .A2(n6380), .ZN(n9522) );
  NAND2_X1 U5961 ( .A1(n9561), .A2(n8399), .ZN(n9536) );
  NAND2_X1 U5962 ( .A1(n6261), .A2(n8397), .ZN(n9558) );
  NAND2_X1 U5963 ( .A1(n4830), .A2(n4832), .ZN(n9551) );
  NAND2_X1 U5964 ( .A1(n4831), .A2(n4833), .ZN(n4830) );
  NAND2_X1 U5965 ( .A1(n6247), .A2(n6246), .ZN(n9595) );
  NAND2_X1 U5966 ( .A1(n4852), .A2(n6369), .ZN(n9619) );
  NAND2_X1 U5967 ( .A1(n4849), .A2(n6362), .ZN(n8027) );
  NAND2_X1 U5968 ( .A1(n4854), .A2(n6358), .ZN(n10201) );
  NAND2_X1 U5969 ( .A1(n6157), .A2(n6156), .ZN(n10210) );
  NAND2_X1 U5970 ( .A1(n7598), .A2(n8373), .ZN(n7682) );
  AND2_X1 U5971 ( .A1(n6119), .A2(n6118), .ZN(n7887) );
  NAND2_X1 U5972 ( .A1(n10224), .A2(n10225), .ZN(n4817) );
  NAND2_X1 U5973 ( .A1(n7515), .A2(n7516), .ZN(n4825) );
  INV_X1 U5974 ( .A(n10271), .ZN(n9603) );
  INV_X1 U5975 ( .A(n10257), .ZN(n10272) );
  INV_X2 U5976 ( .A(n10282), .ZN(n10261) );
  INV_X1 U5977 ( .A(n9612), .ZN(n10278) );
  INV_X1 U5978 ( .A(n7068), .ZN(n9310) );
  AND2_X1 U5979 ( .A1(n9470), .A2(n9636), .ZN(n8169) );
  NAND2_X1 U5980 ( .A1(n8532), .A2(n8156), .ZN(n8158) );
  INV_X1 U5981 ( .A(n9513), .ZN(n9720) );
  AND2_X1 U5982 ( .A1(n6273), .A2(n6272), .ZN(n9728) );
  INV_X1 U5983 ( .A(n9595), .ZN(n6396) );
  XNOR2_X1 U5984 ( .A(n5282), .B(n5281), .ZN(n8153) );
  OAI21_X1 U5985 ( .B1(n5729), .B2(n5728), .A(n5279), .ZN(n5282) );
  XNOR2_X1 U5986 ( .A(n5983), .B(n5982), .ZN(n5985) );
  NAND2_X1 U5987 ( .A1(n8141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5988 ( .A1(n5981), .A2(n5980), .ZN(n9756) );
  NOR2_X1 U5989 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NOR2_X1 U5990 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5978) );
  NAND2_X1 U5991 ( .A1(n4723), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U5992 ( .A1(n6407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  INV_X1 U5993 ( .A(n4968), .ZN(n5645) );
  AOI21_X1 U5994 ( .B1(n5622), .B2(n4973), .A(n4971), .ZN(n4968) );
  OR2_X1 U5995 ( .A1(n6314), .A2(n9899), .ZN(n6315) );
  NAND2_X1 U5996 ( .A1(n6319), .A2(n6318), .ZN(n8512) );
  NAND2_X1 U5997 ( .A1(n4653), .A2(n4652), .ZN(n6319) );
  NAND2_X1 U5998 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6312), .ZN(n4652) );
  OAI21_X1 U5999 ( .B1(n6311), .B2(n6103), .A(P1_IR_REG_20__SCAN_IN), .ZN(
        n4653) );
  NAND2_X1 U6000 ( .A1(n4943), .A2(n4944), .ZN(n5487) );
  NAND2_X1 U6001 ( .A1(n5404), .A2(n5403), .ZN(n5402) );
  NAND2_X1 U6002 ( .A1(n5381), .A2(n5181), .ZN(n5404) );
  XNOR2_X1 U6003 ( .A(n6016), .B(n6015), .ZN(n8224) );
  OAI21_X1 U6004 ( .B1(n6029), .B2(n6003), .A(n6014), .ZN(n7043) );
  NAND2_X1 U6005 ( .A1(n5315), .A2(SI_1_), .ZN(n4703) );
  XNOR2_X1 U6006 ( .A(n5993), .B(n5992), .ZN(n9315) );
  NAND2_X1 U6007 ( .A1(n5036), .A2(n8693), .ZN(n5035) );
  OR2_X1 U6008 ( .A1(n6778), .A2(n8839), .ZN(n5145) );
  AOI211_X1 U6009 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n10414), .A(n6731), .B(
        n6730), .ZN(n6779) );
  NAND2_X1 U6010 ( .A1(n4871), .A2(n4869), .ZN(P1_U3262) );
  AOI21_X1 U6011 ( .B1(n4874), .B2(n7479), .A(n4872), .ZN(n4871) );
  NAND2_X1 U6012 ( .A1(n4870), .A2(n8434), .ZN(n4869) );
  INV_X1 U6013 ( .A(n4873), .ZN(n4872) );
  NOR2_X1 U6014 ( .A1(n6429), .A2(n6431), .ZN(n6432) );
  NAND2_X1 U6015 ( .A1(n4753), .A2(n4751), .ZN(P1_U3518) );
  INV_X1 U6016 ( .A(n4752), .ZN(n4751) );
  NAND2_X1 U6017 ( .A1(n9715), .A2(n10395), .ZN(n4753) );
  OAI22_X1 U6018 ( .A1(n9716), .A2(n9747), .B1(n10395), .B2(n6298), .ZN(n4752)
         );
  AND2_X1 U6019 ( .A1(n8598), .A2(n4605), .ZN(n4528) );
  NOR2_X1 U6020 ( .A1(n4894), .A2(n4893), .ZN(n4892) );
  NAND2_X1 U6021 ( .A1(n6297), .A2(n6296), .ZN(n6387) );
  NAND2_X1 U6022 ( .A1(n8155), .A2(n6045), .ZN(n8359) );
  INV_X1 U6023 ( .A(n6619), .ZN(n4645) );
  XNOR2_X1 U6024 ( .A(n5355), .B(n5354), .ZN(n6929) );
  NOR2_X1 U6025 ( .A1(n5400), .A2(n5084), .ZN(n5755) );
  INV_X1 U6026 ( .A(n9194), .ZN(n4644) );
  INV_X1 U6027 ( .A(n6844), .ZN(n8996) );
  AND2_X1 U6028 ( .A1(n5882), .A2(n5876), .ZN(n6844) );
  AND2_X1 U6029 ( .A1(n8538), .A2(n9017), .ZN(n4529) );
  XNOR2_X1 U6030 ( .A(n8574), .B(n8602), .ZN(n8867) );
  INV_X1 U6031 ( .A(n8867), .ZN(n5116) );
  OR2_X1 U6032 ( .A1(n9112), .A2(n8907), .ZN(n4530) );
  AND2_X1 U6033 ( .A1(n4889), .A2(n4894), .ZN(n4531) );
  NAND2_X1 U6034 ( .A1(n9112), .A2(n8885), .ZN(n5912) );
  INV_X1 U6035 ( .A(n5912), .ZN(n5128) );
  NOR2_X1 U6036 ( .A1(n6490), .A2(n6489), .ZN(n4532) );
  NOR2_X1 U6037 ( .A1(n6600), .A2(n6599), .ZN(n9225) );
  AND2_X1 U6038 ( .A1(n5093), .A2(n5851), .ZN(n4533) );
  NAND2_X1 U6039 ( .A1(n6170), .A2(n6169), .ZN(n8284) );
  INV_X1 U6040 ( .A(n8284), .ZN(n4714) );
  AND2_X1 U6041 ( .A1(n5037), .A2(n4550), .ZN(n4534) );
  INV_X1 U6042 ( .A(n5455), .ZN(n4945) );
  AND2_X1 U6043 ( .A1(n6378), .A2(n9568), .ZN(n4535) );
  NAND2_X1 U6044 ( .A1(n5910), .A2(n5909), .ZN(n4536) );
  AND2_X1 U6045 ( .A1(n5059), .A2(n4566), .ZN(n4537) );
  AND2_X1 U6046 ( .A1(n4724), .A2(n4725), .ZN(n4538) );
  AND2_X1 U6047 ( .A1(n4883), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4539) );
  AND2_X1 U6048 ( .A1(n8023), .A2(n4718), .ZN(n4540) );
  INV_X1 U6049 ( .A(n6377), .ZN(n4833) );
  INV_X1 U6050 ( .A(n4892), .ZN(n4891) );
  XOR2_X1 U6051 ( .A(n6540), .B(n6612), .Z(n4541) );
  OR2_X1 U6052 ( .A1(n9138), .A2(n8978), .ZN(n5895) );
  XNOR2_X1 U6053 ( .A(n6317), .B(n6316), .ZN(n6325) );
  INV_X1 U6054 ( .A(n8711), .ZN(n8693) );
  AND2_X1 U6055 ( .A1(n9444), .A2(n9439), .ZN(n4542) );
  INV_X1 U6056 ( .A(n8359), .ZN(n8358) );
  NAND3_X1 U6057 ( .A1(n6435), .A2(n6437), .A3(n6433), .ZN(n6464) );
  INV_X1 U6058 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U6059 ( .A1(n6438), .A2(n6437), .ZN(n6469) );
  INV_X1 U6060 ( .A(n4925), .ZN(n4924) );
  OAI21_X1 U6061 ( .B1(n9178), .B2(n4926), .A(n6580), .ZN(n4925) );
  INV_X1 U6062 ( .A(n7416), .ZN(n6952) );
  INV_X1 U6063 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6064 ( .A1(n9169), .A2(n9171), .ZN(n9170) );
  NAND2_X1 U6065 ( .A1(n5076), .A2(n5895), .ZN(n8934) );
  AND2_X1 U6066 ( .A1(n9000), .A2(n6843), .ZN(n4543) );
  NAND2_X1 U6067 ( .A1(n9539), .A2(n4727), .ZN(n4544) );
  OR2_X1 U6068 ( .A1(n9112), .A2(n8885), .ZN(n5904) );
  AND2_X1 U6069 ( .A1(n5071), .A2(n7865), .ZN(n4545) );
  NAND3_X1 U6070 ( .A1(n5357), .A2(n5143), .A3(n5356), .ZN(n7168) );
  INV_X1 U6071 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5340) );
  AND4_X1 U6072 ( .A1(n5290), .A2(n5289), .A3(n5753), .A4(n5581), .ZN(n4546)
         );
  INV_X1 U6073 ( .A(n7722), .ZN(n6900) );
  OR2_X1 U6074 ( .A1(n7416), .A2(n10560), .ZN(n4547) );
  AND2_X1 U6075 ( .A1(n6475), .A2(n6474), .ZN(n4548) );
  AND2_X1 U6076 ( .A1(n5129), .A2(n5904), .ZN(n4549) );
  OR2_X1 U6077 ( .A1(n5039), .A2(n8570), .ZN(n4550) );
  AND2_X1 U6078 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4551) );
  AND2_X1 U6079 ( .A1(n9249), .A2(n9250), .ZN(n4552) );
  AND3_X1 U6080 ( .A1(n5339), .A2(n5365), .A3(n5072), .ZN(n5398) );
  INV_X1 U6081 ( .A(n8735), .ZN(n7780) );
  AND2_X1 U6082 ( .A1(n6629), .A2(n6628), .ZN(n4553) );
  INV_X1 U6083 ( .A(n8636), .ZN(n5055) );
  AND3_X1 U6084 ( .A1(n6153), .A2(n6152), .A3(n6167), .ZN(n4554) );
  OR2_X1 U6085 ( .A1(n9465), .A2(n9464), .ZN(n4555) );
  NOR2_X1 U6086 ( .A1(n9307), .A2(n7609), .ZN(n8444) );
  NAND2_X2 U6087 ( .A1(n6045), .A2(n8151), .ZN(n6013) );
  AND2_X1 U6088 ( .A1(n5836), .A2(n7698), .ZN(n7643) );
  OR2_X1 U6089 ( .A1(n4922), .A2(n4921), .ZN(n4556) );
  AND2_X1 U6090 ( .A1(n9627), .A2(n9693), .ZN(n4557) );
  AND2_X1 U6091 ( .A1(n9106), .A2(n8895), .ZN(n4558) );
  INV_X1 U6092 ( .A(n9275), .ZN(n6395) );
  NAND2_X1 U6093 ( .A1(n6212), .A2(n6211), .ZN(n9275) );
  AND2_X1 U6094 ( .A1(n6181), .A2(n6180), .ZN(n10196) );
  NOR2_X1 U6095 ( .A1(n8808), .A2(n6688), .ZN(n4559) );
  NOR2_X1 U6096 ( .A1(n5974), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4560) );
  AND3_X1 U6097 ( .A1(n5849), .A2(n5843), .A3(n5842), .ZN(n4561) );
  NAND2_X1 U6098 ( .A1(n8284), .A2(n9301), .ZN(n4562) );
  AND2_X1 U6099 ( .A1(n8472), .A2(n8477), .ZN(n8384) );
  AND2_X1 U6100 ( .A1(n5005), .A2(n5004), .ZN(n4563) );
  INV_X1 U6101 ( .A(n4639), .ZN(n4638) );
  NOR2_X1 U6102 ( .A1(n8086), .A2(n8087), .ZN(n4639) );
  INV_X1 U6103 ( .A(n4790), .ZN(n4789) );
  AND2_X1 U6104 ( .A1(n5119), .A2(n5116), .ZN(n4564) );
  AND2_X1 U6105 ( .A1(n6278), .A2(n6277), .ZN(n9724) );
  INV_X1 U6106 ( .A(n9724), .ZN(n9532) );
  INV_X1 U6107 ( .A(n6387), .ZN(n9716) );
  AND2_X1 U6108 ( .A1(n5297), .A2(n5293), .ZN(n4565) );
  XNOR2_X1 U6109 ( .A(n5299), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6110 ( .A1(n8552), .A2(n8932), .ZN(n4566) );
  NAND2_X1 U6111 ( .A1(n7261), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4567) );
  AND2_X1 U6112 ( .A1(n9106), .A2(n8526), .ZN(n5772) );
  AND2_X1 U6113 ( .A1(n4920), .A2(n9226), .ZN(n4568) );
  AND2_X1 U6114 ( .A1(n8230), .A2(n6343), .ZN(n4569) );
  OR2_X1 U6115 ( .A1(n10536), .A2(n7921), .ZN(n5853) );
  AND2_X1 U6116 ( .A1(n5643), .A2(n5075), .ZN(n4570) );
  NOR2_X1 U6117 ( .A1(n10342), .A2(n10349), .ZN(n4571) );
  OR2_X1 U6118 ( .A1(n6866), .A2(n7263), .ZN(n4572) );
  NAND2_X1 U6119 ( .A1(n9644), .A2(n9643), .ZN(n4573) );
  NOR2_X1 U6120 ( .A1(n8539), .A2(n8718), .ZN(n4574) );
  NAND2_X1 U6121 ( .A1(n6311), .A2(n5968), .ZN(n4575) );
  AND2_X1 U6122 ( .A1(n9222), .A2(n9299), .ZN(n4576) );
  AND2_X1 U6123 ( .A1(n4984), .A2(n4982), .ZN(n4577) );
  NAND2_X1 U6124 ( .A1(n5832), .A2(n7698), .ZN(n4578) );
  AND2_X1 U6125 ( .A1(n5200), .A2(n10104), .ZN(n4579) );
  OR2_X1 U6126 ( .A1(n8490), .A2(n8319), .ZN(n4580) );
  NOR2_X1 U6127 ( .A1(n5194), .A2(SI_9_), .ZN(n4581) );
  AND2_X1 U6128 ( .A1(n10196), .A2(n9300), .ZN(n8474) );
  OR2_X1 U6129 ( .A1(n5123), .A2(n5906), .ZN(n4582) );
  AND2_X1 U6130 ( .A1(n8568), .A2(n8728), .ZN(n4583) );
  NAND2_X1 U6131 ( .A1(n8901), .A2(n4777), .ZN(n4584) );
  OR2_X1 U6132 ( .A1(n8935), .A2(n6884), .ZN(n4585) );
  INV_X1 U6133 ( .A(n9103), .ZN(n8574) );
  AND2_X1 U6134 ( .A1(n5711), .A2(n5710), .ZN(n9103) );
  AND2_X1 U6135 ( .A1(n8056), .A2(n8294), .ZN(n4586) );
  AND2_X1 U6136 ( .A1(n5058), .A2(n4537), .ZN(n4587) );
  AND2_X1 U6137 ( .A1(n9186), .A2(n4631), .ZN(n4588) );
  OR2_X1 U6138 ( .A1(n6378), .A2(n9197), .ZN(n8399) );
  AND3_X1 U6139 ( .A1(n4530), .A2(n6857), .A3(n6855), .ZN(n4589) );
  AND2_X1 U6140 ( .A1(n5092), .A2(n5851), .ZN(n4590) );
  OR2_X1 U6141 ( .A1(n6378), .A2(n9568), .ZN(n4591) );
  AND2_X1 U6142 ( .A1(n5209), .A2(n4981), .ZN(n4592) );
  AND2_X1 U6143 ( .A1(n5063), .A2(n8670), .ZN(n4593) );
  AND2_X1 U6144 ( .A1(n8376), .A2(n8373), .ZN(n4594) );
  INV_X1 U6145 ( .A(n6346), .ZN(n4826) );
  INV_X1 U6146 ( .A(n5882), .ZN(n5080) );
  OR2_X1 U6147 ( .A1(n8994), .A2(n8977), .ZN(n5882) );
  AND2_X1 U6148 ( .A1(n6165), .A2(n8464), .ZN(n4595) );
  NAND2_X1 U6149 ( .A1(n5163), .A2(n5162), .ZN(n4596) );
  AND2_X1 U6150 ( .A1(n5112), .A2(n4565), .ZN(n4597) );
  AND2_X1 U6151 ( .A1(n7619), .A2(n7615), .ZN(n4598) );
  NAND2_X1 U6152 ( .A1(n5126), .A2(n5787), .ZN(n5125) );
  AND2_X1 U6153 ( .A1(n4734), .A2(n4733), .ZN(n4599) );
  AND2_X1 U6154 ( .A1(n4832), .A2(n4591), .ZN(n4829) );
  INV_X2 U6155 ( .A(n8163), .ZN(n6305) );
  INV_X1 U6156 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U6157 ( .A1(n4933), .A2(n4934), .ZN(n7752) );
  AND2_X1 U6158 ( .A1(n5053), .A2(n5051), .ZN(n8643) );
  NAND2_X1 U6159 ( .A1(n7794), .A2(n7793), .ZN(n7866) );
  NAND2_X1 U6160 ( .A1(n7866), .A2(n7865), .ZN(n7935) );
  INV_X1 U6161 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U6162 ( .A1(n4625), .A2(n4562), .ZN(n7962) );
  NAND2_X1 U6163 ( .A1(n8101), .A2(n6544), .ZN(n8085) );
  NAND2_X1 U6164 ( .A1(n5074), .A2(n4570), .ZN(n8920) );
  AND2_X1 U6165 ( .A1(n7127), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U6166 ( .A1(n5216), .A2(n5550), .ZN(n4601) );
  NAND2_X1 U6167 ( .A1(n6304), .A2(n6303), .ZN(n9480) );
  INV_X1 U6168 ( .A(n9480), .ZN(n4724) );
  AND2_X1 U6169 ( .A1(n4915), .A2(n7879), .ZN(n4602) );
  AND2_X1 U6170 ( .A1(n4634), .A2(n4637), .ZN(n9202) );
  INV_X1 U6171 ( .A(n7745), .ZN(n4893) );
  INV_X1 U6172 ( .A(n4894), .ZN(n4890) );
  NOR2_X1 U6173 ( .A1(n7676), .A2(n7786), .ZN(n4894) );
  NOR2_X1 U6174 ( .A1(n8740), .A2(n6682), .ZN(n4603) );
  AND2_X1 U6175 ( .A1(n4530), .A2(n6855), .ZN(n4604) );
  NAND2_X1 U6176 ( .A1(n8023), .A2(n4720), .ZN(n4721) );
  OR2_X1 U6177 ( .A1(n8567), .A2(n8895), .ZN(n4605) );
  OR2_X1 U6178 ( .A1(n5520), .A2(SI_14_), .ZN(n4606) );
  AND2_X1 U6179 ( .A1(n5019), .A2(n5018), .ZN(n4607) );
  AND2_X1 U6180 ( .A1(n6484), .A2(n7450), .ZN(n4608) );
  AND2_X1 U6181 ( .A1(n6993), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4609) );
  INV_X1 U6182 ( .A(n4964), .ZN(n4963) );
  NAND2_X1 U6183 ( .A1(n4601), .A2(n5223), .ZN(n4964) );
  INV_X1 U6184 ( .A(n5133), .ZN(n4807) );
  OR2_X1 U6185 ( .A1(n5564), .A2(n4965), .ZN(n4610) );
  INV_X1 U6186 ( .A(n9591), .ZN(n9611) );
  AND2_X1 U6187 ( .A1(n8023), .A2(n4717), .ZN(n9591) );
  NOR2_X1 U6188 ( .A1(n8710), .A2(n4529), .ZN(n4611) );
  OR2_X1 U6189 ( .A1(n7837), .A2(n10566), .ZN(n4612) );
  OR2_X1 U6190 ( .A1(n6763), .A2(n6713), .ZN(n4613) );
  INV_X1 U6191 ( .A(n4605), .ZN(n5045) );
  XNOR2_X1 U6192 ( .A(n5301), .B(n5293), .ZN(n5962) );
  NAND2_X1 U6193 ( .A1(n7536), .A2(n7535), .ZN(n7539) );
  NAND2_X1 U6194 ( .A1(n5028), .A2(n7391), .ZN(n7536) );
  AOI21_X1 U6195 ( .B1(n7458), .B2(n7456), .A(n4532), .ZN(n7579) );
  NAND2_X1 U6196 ( .A1(n6345), .A2(n6344), .ZN(n7515) );
  OAI21_X1 U6197 ( .B1(n5453), .B2(n5093), .A(n5092), .ZN(n7816) );
  NAND2_X1 U6198 ( .A1(n4825), .A2(n6346), .ZN(n7493) );
  NAND2_X1 U6199 ( .A1(n4817), .A2(n6350), .ZN(n7626) );
  NAND2_X1 U6200 ( .A1(n5096), .A2(n5103), .ZN(n8004) );
  INV_X1 U6201 ( .A(n8042), .ZN(n4910) );
  NAND2_X1 U6202 ( .A1(n5453), .A2(n5452), .ZN(n7709) );
  NAND2_X1 U6203 ( .A1(n4651), .A2(n4548), .ZN(n4614) );
  AND2_X1 U6204 ( .A1(n6824), .A2(n4788), .ZN(n4615) );
  NAND2_X1 U6205 ( .A1(n6315), .A2(n6412), .ZN(n6391) );
  INV_X1 U6206 ( .A(n6391), .ZN(n6393) );
  INV_X1 U6207 ( .A(n6045), .ZN(n6920) );
  AND2_X1 U6208 ( .A1(n9372), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4616) );
  INV_X1 U6209 ( .A(n7805), .ZN(n5021) );
  INV_X1 U6210 ( .A(n7538), .ZN(n5027) );
  AND2_X1 U6211 ( .A1(n9455), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4617) );
  INV_X1 U6212 ( .A(n4532), .ZN(n4936) );
  NAND2_X1 U6213 ( .A1(n6704), .A2(n7302), .ZN(n4618) );
  NOR2_X1 U6214 ( .A1(n6673), .A2(n6745), .ZN(n6674) );
  INV_X1 U6215 ( .A(n6674), .ZN(n4898) );
  AND2_X1 U6216 ( .A1(n4879), .A2(n4878), .ZN(n4619) );
  AND2_X1 U6217 ( .A1(n5007), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4620) );
  AND2_X1 U6218 ( .A1(n5009), .A2(n5008), .ZN(n4621) );
  AND2_X1 U6219 ( .A1(n7302), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4622) );
  XOR2_X1 U6220 ( .A(n6935), .B(n6742), .Z(n4623) );
  AND2_X1 U6221 ( .A1(n5292), .A2(n4597), .ZN(n8145) );
  INV_X1 U6222 ( .A(n6325), .ZN(n8439) );
  INV_X1 U6223 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U6224 ( .A1(n4624), .A2(n6901), .ZN(n10443) );
  NAND2_X1 U6225 ( .A1(n6900), .A2(n5021), .ZN(n4624) );
  XNOR2_X1 U6226 ( .A(n5758), .B(n5757), .ZN(n7722) );
  XNOR2_X1 U6227 ( .A(n6716), .B(n8785), .ZN(n8782) );
  AOI21_X1 U6228 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n7385), .A(n8792), .ZN(
        n6718) );
  AND2_X1 U6229 ( .A1(n6718), .A2(n8822), .ZN(n6719) );
  INV_X2 U6230 ( .A(n8149), .ZN(n9167) );
  INV_X2 U6231 ( .A(n8143), .ZN(n9754) );
  INV_X1 U6232 ( .A(n4662), .ZN(n4661) );
  NAND2_X1 U6233 ( .A1(n4741), .A2(n4739), .ZN(n5838) );
  OR2_X1 U6234 ( .A1(n5170), .A2(SI_3_), .ZN(n5171) );
  NAND2_X1 U6235 ( .A1(n5858), .A2(n5857), .ZN(n4677) );
  AOI21_X1 U6236 ( .B1(n5908), .B2(n5909), .A(n4682), .ZN(n4681) );
  AOI21_X1 U6237 ( .B1(n5935), .B2(n4744), .A(n5137), .ZN(n5936) );
  AOI21_X1 U6238 ( .B1(n5850), .B2(n5848), .A(n5847), .ZN(n5854) );
  AOI21_X1 U6239 ( .B1(n5869), .B2(n5868), .A(n4679), .ZN(n4678) );
  NAND2_X1 U6240 ( .A1(n5844), .A2(n6884), .ZN(n4663) );
  NAND2_X1 U6241 ( .A1(n7728), .A2(n8379), .ZN(n4854) );
  NOR2_X1 U6242 ( .A1(n9646), .A2(n10307), .ZN(n4755) );
  NAND2_X1 U6243 ( .A1(n10191), .A2(n5153), .ZN(n4729) );
  NAND2_X1 U6244 ( .A1(n4837), .A2(n4834), .ZN(n9489) );
  NAND2_X1 U6245 ( .A1(n9645), .A2(n4754), .ZN(n9715) );
  NAND2_X1 U6246 ( .A1(n4626), .A2(n9259), .ZN(n9169) );
  NAND3_X1 U6247 ( .A1(n9259), .A2(n4626), .A3(n6601), .ZN(n4919) );
  NAND2_X1 U6248 ( .A1(n9258), .A2(n9260), .ZN(n4626) );
  NAND2_X1 U6249 ( .A1(n6483), .A2(n7450), .ZN(n4628) );
  NOR2_X1 U6250 ( .A1(n6514), .A2(n6513), .ZN(n6516) );
  NAND2_X1 U6251 ( .A1(n4629), .A2(n4588), .ZN(n6588) );
  NAND3_X1 U6252 ( .A1(n6567), .A2(n4923), .A3(n9268), .ZN(n4629) );
  NAND2_X1 U6253 ( .A1(n4634), .A2(n4632), .ZN(n9213) );
  NAND3_X1 U6254 ( .A1(n8101), .A2(n4635), .A3(n6544), .ZN(n4634) );
  NAND3_X1 U6255 ( .A1(n8101), .A2(n6544), .A3(n4556), .ZN(n4636) );
  OAI21_X1 U6256 ( .B1(n6796), .B2(n4640), .A(n9285), .ZN(n6654) );
  NAND2_X1 U6257 ( .A1(n9193), .A2(n9194), .ZN(n9281) );
  INV_X1 U6258 ( .A(n6631), .ZN(n4646) );
  INV_X1 U6259 ( .A(n4651), .ZN(n7173) );
  NAND2_X1 U6260 ( .A1(n4654), .A2(n4599), .ZN(n4732) );
  NAND2_X1 U6261 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  INV_X1 U6262 ( .A(n5896), .ZN(n4655) );
  NAND2_X1 U6263 ( .A1(n4657), .A2(n8936), .ZN(n4656) );
  NAND2_X1 U6264 ( .A1(n4658), .A2(n4585), .ZN(n4657) );
  NAND2_X1 U6265 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  OR3_X1 U6266 ( .A1(n5889), .A2(n5888), .A3(n5887), .ZN(n4660) );
  NAND2_X1 U6267 ( .A1(n8151), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4667) );
  MUX2_X1 U6268 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8151), .Z(n5178) );
  MUX2_X1 U6269 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8151), .Z(n5187) );
  MUX2_X1 U6270 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n4666), .Z(n5191) );
  MUX2_X1 U6271 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n4666), .Z(n5194) );
  MUX2_X1 U6272 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n4666), .Z(n5201) );
  MUX2_X1 U6273 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n4666), .Z(n5520) );
  MUX2_X1 U6274 ( .A(n9970), .B(n5218), .S(n4666), .Z(n5220) );
  MUX2_X1 U6275 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n4666), .Z(n5551) );
  MUX2_X1 U6276 ( .A(n7657), .B(n7658), .S(n4666), .Z(n5229) );
  MUX2_X1 U6277 ( .A(n10072), .B(n7877), .S(n4666), .Z(n5239) );
  MUX2_X1 U6278 ( .A(n7992), .B(n7994), .S(n4666), .Z(n5249) );
  MUX2_X1 U6279 ( .A(n8576), .B(n5709), .S(n4666), .Z(n5269) );
  MUX2_X1 U6280 ( .A(n9755), .B(n9166), .S(n4666), .Z(n5272) );
  NAND2_X2 U6281 ( .A1(n6045), .A2(n6914), .ZN(n6071) );
  INV_X2 U6282 ( .A(n4666), .ZN(n6914) );
  NAND2_X1 U6283 ( .A1(n4674), .A2(n8071), .ZN(n4730) );
  NAND2_X1 U6284 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U6285 ( .A1(n4677), .A2(n5147), .ZN(n4675) );
  OAI21_X1 U6286 ( .B1(n4677), .B2(n6836), .A(n5860), .ZN(n4676) );
  OAI211_X2 U6287 ( .C1(n4681), .C2(n4582), .A(n5915), .B(n4680), .ZN(n5921)
         );
  OAI21_X2 U6288 ( .B1(n5908), .B2(n4536), .A(n4577), .ZN(n4680) );
  NAND2_X2 U6289 ( .A1(n6007), .A2(n5135), .ZN(n8229) );
  INV_X1 U6290 ( .A(n8151), .ZN(n4707) );
  OAI21_X1 U6291 ( .B1(n8151), .B2(n4709), .A(n4708), .ZN(n5170) );
  MUX2_X1 U6292 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n8151), .Z(n5312) );
  NAND2_X1 U6293 ( .A1(n7730), .A2(n4713), .ZN(n4716) );
  INV_X1 U6294 ( .A(n4716), .ZN(n7958) );
  INV_X1 U6295 ( .A(n4721), .ZN(n9625) );
  NAND2_X1 U6296 ( .A1(n9539), .A2(n4538), .ZN(n9471) );
  NAND2_X1 U6297 ( .A1(n4730), .A2(n5863), .ZN(n5864) );
  AND2_X2 U6298 ( .A1(n4732), .A2(n4731), .ZN(n5908) );
  NAND2_X1 U6299 ( .A1(n4735), .A2(n5965), .ZN(P2_U3296) );
  NAND2_X1 U6300 ( .A1(n4737), .A2(n4736), .ZN(n4735) );
  OAI21_X1 U6301 ( .B1(n4518), .B2(n5938), .A(n4738), .ZN(n4737) );
  NAND2_X1 U6302 ( .A1(n5939), .A2(n7102), .ZN(n4738) );
  AND2_X2 U6303 ( .A1(n5931), .A2(n5930), .ZN(n4744) );
  OR2_X2 U6304 ( .A1(n5921), .A2(n4745), .ZN(n5931) );
  NAND2_X1 U6305 ( .A1(n8151), .A2(n4596), .ZN(n4746) );
  NAND3_X1 U6306 ( .A1(n4750), .A2(n7922), .A3(n4747), .ZN(n5858) );
  OR2_X2 U6307 ( .A1(n5854), .A2(n6884), .ZN(n4750) );
  NAND4_X1 U6308 ( .A1(n6027), .A2(n6002), .A3(n5966), .A4(n5967), .ZN(n6046)
         );
  OAI21_X2 U6309 ( .B1(n6261), .B2(n8318), .A(n4756), .ZN(n9535) );
  NAND2_X2 U6310 ( .A1(n10268), .A2(n5997), .ZN(n10247) );
  NAND2_X2 U6311 ( .A1(n8441), .A2(n5997), .ZN(n8361) );
  NAND2_X1 U6312 ( .A1(n7726), .A2(n4595), .ZN(n10205) );
  NAND2_X1 U6313 ( .A1(n7598), .A2(n4594), .ZN(n7684) );
  NAND4_X1 U6314 ( .A1(n4769), .A2(n4814), .A3(n4560), .A4(n4812), .ZN(n4768)
         );
  NAND2_X1 U6315 ( .A1(n8906), .A2(n4589), .ZN(n4771) );
  INV_X1 U6316 ( .A(n6859), .ZN(n8524) );
  INV_X1 U6317 ( .A(n10473), .ZN(n6811) );
  OAI211_X1 U6318 ( .C1(n5336), .C2(n6936), .A(n4572), .B(n4778), .ZN(n10473)
         );
  OR2_X1 U6319 ( .A1(n4527), .A2(n6937), .ZN(n4778) );
  NAND2_X1 U6320 ( .A1(n6811), .A2(n7109), .ZN(n5796) );
  NAND2_X1 U6321 ( .A1(n4615), .A2(n6825), .ZN(n4787) );
  NAND2_X1 U6322 ( .A1(n4779), .A2(n4783), .ZN(n6830) );
  NAND2_X1 U6323 ( .A1(n6825), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U6324 ( .A1(n6825), .A2(n6824), .ZN(n9034) );
  INV_X1 U6325 ( .A(n6826), .ZN(n4788) );
  NOR2_X1 U6326 ( .A1(n10505), .A2(n8737), .ZN(n4790) );
  NAND4_X1 U6327 ( .A1(n4793), .A2(n5285), .A3(n5286), .A4(n4792), .ZN(n4791)
         );
  NAND3_X1 U6328 ( .A1(n4801), .A2(n6842), .A3(n4800), .ZN(n9002) );
  NAND3_X1 U6329 ( .A1(n4804), .A2(n6841), .A3(n4805), .ZN(n4800) );
  NAND3_X1 U6330 ( .A1(n7919), .A2(n6841), .A3(n4804), .ZN(n4801) );
  NOR2_X1 U6331 ( .A1(n8856), .A2(n6869), .ZN(n6909) );
  NAND2_X1 U6332 ( .A1(n4811), .A2(n10443), .ZN(n4810) );
  XNOR2_X1 U6333 ( .A(n6863), .B(n6862), .ZN(n4811) );
  AND2_X2 U6334 ( .A1(n5082), .A2(n5083), .ZN(n5292) );
  INV_X1 U6335 ( .A(n6046), .ZN(n4812) );
  AND3_X1 U6336 ( .A1(n5966), .A2(n6002), .A3(n6027), .ZN(n6068) );
  AND2_X2 U6337 ( .A1(n5968), .A2(n5969), .ZN(n4814) );
  AND4_X2 U6338 ( .A1(n6312), .A2(n6316), .A3(n9899), .A4(n10083), .ZN(n5968)
         );
  NAND2_X1 U6339 ( .A1(n4815), .A2(n4816), .ZN(n7463) );
  NAND2_X1 U6340 ( .A1(n10224), .A2(n4818), .ZN(n4815) );
  NAND2_X1 U6341 ( .A1(n4823), .A2(n4821), .ZN(n6349) );
  INV_X1 U6342 ( .A(n4822), .ZN(n4821) );
  OAI21_X1 U6343 ( .B1(n7516), .B2(n4826), .A(n7634), .ZN(n4822) );
  NAND2_X1 U6344 ( .A1(n6345), .A2(n4824), .ZN(n4823) );
  NAND2_X1 U6345 ( .A1(n9575), .A2(n4829), .ZN(n4827) );
  NAND2_X1 U6346 ( .A1(n4827), .A2(n4828), .ZN(n9547) );
  INV_X1 U6347 ( .A(n9547), .ZN(n6379) );
  NAND2_X1 U6348 ( .A1(n6381), .A2(n4838), .ZN(n4837) );
  INV_X1 U6349 ( .A(n10276), .ZN(n10290) );
  NAND2_X1 U6350 ( .A1(n7068), .A2(n10276), .ZN(n5997) );
  NAND2_X1 U6351 ( .A1(n4849), .A2(n4847), .ZN(n6364) );
  NAND2_X1 U6352 ( .A1(n4852), .A2(n4850), .ZN(n6371) );
  NAND2_X1 U6353 ( .A1(n4854), .A2(n4853), .ZN(n6360) );
  AND2_X1 U6354 ( .A1(n5132), .A2(n6358), .ZN(n4853) );
  NAND2_X1 U6355 ( .A1(n9422), .A2(n4542), .ZN(n4858) );
  NAND2_X1 U6356 ( .A1(n4879), .A2(n7233), .ZN(n4876) );
  NAND2_X1 U6357 ( .A1(n7186), .A2(n4539), .ZN(n4879) );
  NAND2_X1 U6358 ( .A1(n4875), .A2(n4879), .ZN(n4882) );
  INV_X1 U6359 ( .A(n4877), .ZN(n4875) );
  NOR2_X1 U6360 ( .A1(n4876), .A2(n4877), .ZN(n4881) );
  NAND2_X1 U6361 ( .A1(n7186), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U6362 ( .A1(n7672), .A2(n4892), .ZN(n4887) );
  OAI21_X1 U6363 ( .B1(n8809), .B2(n4896), .A(n4895), .ZN(n8825) );
  NAND2_X1 U6364 ( .A1(n6673), .A2(n6745), .ZN(n4900) );
  NOR2_X1 U6365 ( .A1(n6674), .A2(n4899), .ZN(n7350) );
  NAND2_X1 U6366 ( .A1(n4898), .A2(n4900), .ZN(n7351) );
  NAND2_X1 U6367 ( .A1(n6682), .A2(n4903), .ZN(n4901) );
  NOR2_X1 U6368 ( .A1(n7559), .A2(n7716), .ZN(n7558) );
  NOR2_X1 U6369 ( .A1(n7830), .A2(n7829), .ZN(n7828) );
  OAI21_X1 U6370 ( .B1(n7948), .B2(n4910), .A(n4907), .ZN(n6542) );
  NAND2_X1 U6371 ( .A1(n7948), .A2(n4907), .ZN(n4905) );
  NAND2_X1 U6372 ( .A1(n7807), .A2(n7808), .ZN(n7806) );
  NAND3_X1 U6373 ( .A1(n4912), .A2(n4911), .A3(n7945), .ZN(n6534) );
  NAND2_X1 U6374 ( .A1(n7807), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U6375 ( .A1(n7806), .A2(n4917), .ZN(n4915) );
  INV_X1 U6376 ( .A(n7879), .ZN(n4916) );
  OAI21_X1 U6377 ( .B1(n7450), .B2(n4918), .A(n7449), .ZN(n7451) );
  NAND2_X1 U6378 ( .A1(n5454), .A2(n5455), .ZN(n5458) );
  NAND2_X1 U6379 ( .A1(n5669), .A2(n4953), .ZN(n4951) );
  NAND2_X1 U6380 ( .A1(n5669), .A2(n5670), .ZN(n4952) );
  NAND3_X1 U6381 ( .A1(n5215), .A2(n5214), .A3(n4961), .ZN(n4956) );
  NAND2_X1 U6382 ( .A1(n4956), .A2(n4959), .ZN(n5591) );
  NAND3_X1 U6383 ( .A1(n5215), .A2(n4601), .A3(n5214), .ZN(n4957) );
  NAND2_X1 U6384 ( .A1(n5215), .A2(n5214), .ZN(n5553) );
  NAND3_X1 U6385 ( .A1(n5215), .A2(n5214), .A3(n4963), .ZN(n4958) );
  NAND2_X1 U6386 ( .A1(n5235), .A2(n5234), .ZN(n5622) );
  NAND2_X1 U6387 ( .A1(n4966), .A2(n4969), .ZN(n5248) );
  NAND3_X1 U6388 ( .A1(n5235), .A2(n4967), .A3(n5234), .ZN(n4966) );
  NAND2_X1 U6389 ( .A1(n4977), .A2(n4976), .ZN(n5421) );
  NAND3_X1 U6390 ( .A1(n5379), .A2(n5403), .A3(n5378), .ZN(n4977) );
  NAND2_X1 U6391 ( .A1(n5379), .A2(n5378), .ZN(n5381) );
  NAND2_X1 U6392 ( .A1(n5505), .A2(n4592), .ZN(n4980) );
  XNOR2_X2 U6393 ( .A(n5706), .B(n8728), .ZN(n8523) );
  NOR2_X1 U6394 ( .A1(n6929), .A2(n4986), .ZN(n4985) );
  INV_X1 U6395 ( .A(n6699), .ZN(n4986) );
  NAND2_X1 U6396 ( .A1(n7284), .A2(n6699), .ZN(n4987) );
  INV_X1 U6397 ( .A(n4989), .ZN(n4988) );
  OAI21_X1 U6398 ( .B1(n4993), .B2(n6699), .A(P2_REG1_REG_3__SCAN_IN), .ZN(
        n4989) );
  NAND2_X1 U6399 ( .A1(n4990), .A2(n6929), .ZN(n7245) );
  NAND2_X1 U6400 ( .A1(n7284), .A2(n6699), .ZN(n4990) );
  INV_X1 U6401 ( .A(n7302), .ZN(n4996) );
  INV_X1 U6402 ( .A(n5001), .ZN(n7746) );
  INV_X1 U6403 ( .A(n6712), .ZN(n5000) );
  NAND2_X1 U6404 ( .A1(n6720), .A2(n5007), .ZN(n5002) );
  NAND2_X1 U6405 ( .A1(n7389), .A2(n7535), .ZN(n5025) );
  INV_X1 U6406 ( .A(n7389), .ZN(n5028) );
  NAND2_X1 U6407 ( .A1(n5025), .A2(n5026), .ZN(n7541) );
  NAND2_X1 U6408 ( .A1(n7318), .A2(n5029), .ZN(n7325) );
  NAND2_X1 U6409 ( .A1(n7325), .A2(n7324), .ZN(n5030) );
  NAND2_X1 U6410 ( .A1(n5030), .A2(n7326), .ZN(n7388) );
  NAND2_X1 U6411 ( .A1(n7616), .A2(n4598), .ZN(n7766) );
  NAND2_X1 U6412 ( .A1(n8701), .A2(n5034), .ZN(n5033) );
  AOI21_X1 U6413 ( .B1(n8701), .B2(n8702), .A(n5045), .ZN(n8599) );
  OAI211_X1 U6414 ( .C1(n8701), .C2(n5035), .A(n8575), .B(n5033), .ZN(P2_U3160) );
  NAND2_X1 U6415 ( .A1(n8710), .A2(n5049), .ZN(n5048) );
  NAND2_X1 U6416 ( .A1(n8672), .A2(n4593), .ZN(n5058) );
  NAND2_X1 U6417 ( .A1(n5058), .A2(n5057), .ZN(n8555) );
  NAND2_X1 U6419 ( .A1(n5064), .A2(n5067), .ZN(n8535) );
  NAND3_X1 U6420 ( .A1(n7793), .A2(n7794), .A3(n5065), .ZN(n5064) );
  INV_X1 U6421 ( .A(n8959), .ZN(n5076) );
  NAND2_X1 U6422 ( .A1(n8959), .A2(n5640), .ZN(n5074) );
  NAND2_X1 U6423 ( .A1(n8995), .A2(n5882), .ZN(n5077) );
  INV_X1 U6424 ( .A(n5400), .ZN(n5083) );
  NAND2_X1 U6425 ( .A1(n5083), .A2(n5288), .ZN(n5554) );
  NAND2_X1 U6426 ( .A1(n10500), .A2(n5088), .ZN(n5085) );
  NAND2_X1 U6427 ( .A1(n5085), .A2(n5086), .ZN(n7708) );
  NAND2_X1 U6428 ( .A1(n5453), .A2(n4590), .ZN(n5090) );
  NAND2_X1 U6429 ( .A1(n7966), .A2(n5101), .ZN(n5100) );
  NAND2_X1 U6430 ( .A1(n5292), .A2(n5112), .ZN(n5298) );
  NAND2_X1 U6431 ( .A1(n5292), .A2(n5291), .ZN(n5952) );
  INV_X1 U6432 ( .A(n8900), .ZN(n5115) );
  NAND3_X1 U6433 ( .A1(n5124), .A2(n5125), .A3(n5131), .ZN(n5121) );
  AOI211_X1 U6434 ( .C1(n10342), .C2(n6637), .A(n7858), .B(n7857), .ZN(n7859)
         );
  OAI21_X1 U6435 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8329) );
  XNOR2_X1 U6436 ( .A(n5707), .B(n5708), .ZN(n8137) );
  AOI21_X1 U6437 ( .B1(n9480), .B2(n6660), .A(n6659), .ZN(n6661) );
  AOI21_X2 U6438 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n7385), .A(n8799), .ZN(
        n6687) );
  NAND2_X1 U6439 ( .A1(n5159), .A2(SI_2_), .ZN(n5168) );
  INV_X1 U6440 ( .A(n6590), .ZN(n6593) );
  AND2_X1 U6441 ( .A1(n8515), .A2(n8514), .ZN(n8521) );
  NAND2_X1 U6442 ( .A1(n5988), .A2(n5977), .ZN(n8141) );
  INV_X1 U6443 ( .A(n5985), .ZN(n5984) );
  NAND2_X2 U6444 ( .A1(n6326), .A2(n6324), .ZN(n6045) );
  AND2_X1 U6445 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  AND2_X1 U6446 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U6447 ( .A1(n10452), .A2(n5800), .ZN(n10436) );
  INV_X1 U6448 ( .A(n5303), .ZN(n8580) );
  AND2_X1 U6449 ( .A1(n6868), .A2(n10474), .ZN(n6869) );
  NOR2_X1 U6450 ( .A1(n6804), .A2(n5727), .ZN(n5747) );
  OR2_X1 U6451 ( .A1(n10210), .A2(n9302), .ZN(n5132) );
  INV_X1 U6452 ( .A(n10202), .ZN(n6165) );
  NOR2_X1 U6453 ( .A1(n6839), .A2(n6838), .ZN(n5133) );
  NOR2_X1 U6454 ( .A1(n8068), .A2(n6839), .ZN(n5134) );
  OR2_X1 U6455 ( .A1(n9308), .A2(n10298), .ZN(n5135) );
  OR2_X1 U6456 ( .A1(n8860), .A2(n9078), .ZN(n5136) );
  AND2_X1 U6457 ( .A1(n6442), .A2(n6546), .ZN(n5138) );
  AND2_X1 U6458 ( .A1(n5753), .A2(n5752), .ZN(n5139) );
  OR2_X1 U6459 ( .A1(n8860), .A2(n9143), .ZN(n5140) );
  NOR2_X1 U6460 ( .A1(n6938), .A2(n4524), .ZN(n5141) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5169) );
  OR2_X1 U6462 ( .A1(n9728), .A2(n9559), .ZN(n5142) );
  OR2_X1 U6463 ( .A1(n6866), .A2(n6929), .ZN(n5143) );
  INV_X1 U6464 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5173) );
  AND4_X1 U6465 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n5144)
         );
  OAI21_X1 U6466 ( .B1(n9601), .B2(n6373), .A(n6372), .ZN(n9584) );
  INV_X1 U6467 ( .A(n7479), .ZN(n8434) );
  XNOR2_X1 U6468 ( .A(n6223), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6392) );
  INV_X1 U6469 ( .A(n8383), .ZN(n8053) );
  AND2_X1 U6470 ( .A1(n8295), .A2(n8294), .ZN(n8383) );
  INV_X1 U6471 ( .A(n5706), .ZN(n8877) );
  AND2_X1 U6472 ( .A1(n5933), .A2(n6884), .ZN(n5146) );
  AND2_X1 U6473 ( .A1(n7930), .A2(n8731), .ZN(n5147) );
  INV_X1 U6474 ( .A(n9747), .ZN(n6660) );
  INV_X1 U6475 ( .A(n10395), .ZN(n6662) );
  AND2_X1 U6476 ( .A1(n6653), .A2(n6652), .ZN(n5148) );
  AND3_X1 U6477 ( .A1(n6800), .A2(n9285), .A3(n6799), .ZN(n5149) );
  OR2_X1 U6478 ( .A1(n6045), .A2(n9315), .ZN(n5150) );
  AND2_X1 U6479 ( .A1(n6477), .A2(n6476), .ZN(n5151) );
  INV_X1 U6480 ( .A(n9295), .ZN(n8357) );
  OR2_X1 U6481 ( .A1(n6866), .A2(n6949), .ZN(n5152) );
  MUX2_X1 U6482 ( .A(n5873), .B(n5797), .S(n5796), .Z(n5798) );
  NAND2_X1 U6483 ( .A1(n5807), .A2(n5873), .ZN(n5808) );
  NAND2_X1 U6484 ( .A1(n5874), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U6485 ( .A1(n8324), .A2(n8351), .ZN(n8322) );
  NAND2_X1 U6486 ( .A1(n5784), .A2(n6884), .ZN(n5785) );
  NAND2_X1 U6487 ( .A1(n5918), .A2(n5922), .ZN(n5919) );
  AND2_X1 U6488 ( .A1(n8261), .A2(n7637), .ZN(n8257) );
  NOR2_X1 U6489 ( .A1(n9012), .A2(n9017), .ZN(n6840) );
  INV_X1 U6490 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5285) );
  INV_X1 U6491 ( .A(n8923), .ZN(n8560) );
  NOR2_X1 U6492 ( .A1(n8877), .A2(n8886), .ZN(n6858) );
  INV_X1 U6493 ( .A(n7711), .ZN(n5452) );
  INV_X1 U6494 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5522) );
  INV_X1 U6495 ( .A(n6571), .ZN(n6572) );
  NAND2_X1 U6496 ( .A1(n10276), .A2(n4521), .ZN(n6444) );
  INV_X1 U6497 ( .A(n8512), .ZN(n6390) );
  NAND2_X1 U6498 ( .A1(n8559), .A2(n8560), .ZN(n8561) );
  AND2_X1 U6499 ( .A1(n7795), .A2(n7861), .ZN(n7793) );
  NAND2_X1 U6500 ( .A1(n7264), .A2(n6698), .ZN(n7285) );
  INV_X1 U6501 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5154) );
  AOI21_X1 U6502 ( .B1(n6378), .B2(n6446), .A(n6605), .ZN(n6607) );
  INV_X1 U6503 ( .A(n6464), .ZN(n6546) );
  OR2_X1 U6504 ( .A1(n10298), .A2(n6461), .ZN(n6454) );
  INV_X1 U6505 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6074) );
  AND2_X1 U6506 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n6274), .ZN(n6279) );
  AND2_X1 U6507 ( .A1(n6195), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6213) );
  INV_X1 U6508 ( .A(SI_5_), .ZN(n9975) );
  AND2_X1 U6509 ( .A1(n7868), .A2(n7867), .ZN(n7865) );
  NOR2_X1 U6510 ( .A1(n7282), .A2(n7283), .ZN(n7281) );
  NOR2_X1 U6511 ( .A1(n6715), .A2(n8747), .ZN(n8765) );
  NAND2_X1 U6512 ( .A1(n5954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5295) );
  INV_X1 U6513 ( .A(n8837), .ZN(n6725) );
  NAND2_X1 U6514 ( .A1(n7373), .A2(n5814), .ZN(n7425) );
  INV_X1 U6515 ( .A(n6449), .ZN(n6447) );
  OR2_X1 U6516 ( .A1(n6135), .A2(n6134), .ZN(n6144) );
  AND2_X1 U6517 ( .A1(n6111), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6121) );
  NOR2_X1 U6518 ( .A1(n6266), .A2(n9230), .ZN(n6274) );
  AND2_X1 U6519 ( .A1(n6248), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6258) );
  NOR2_X1 U6520 ( .A1(n6160), .A2(n6159), .ZN(n6172) );
  NAND2_X1 U6521 ( .A1(n8229), .A2(n7607), .ZN(n7606) );
  NOR2_X1 U6522 ( .A1(n4724), .A2(n9710), .ZN(n6429) );
  NAND2_X1 U6523 ( .A1(n6044), .A2(n8450), .ZN(n7517) );
  NAND2_X1 U6524 ( .A1(n6206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6209) );
  INV_X1 U6525 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U6526 ( .A1(n5192), .A2(n10073), .ZN(n5193) );
  NAND2_X1 U6527 ( .A1(n5175), .A2(SI_4_), .ZN(n5177) );
  AND2_X1 U6528 ( .A1(n8620), .A2(n8551), .ZN(n8670) );
  INV_X1 U6529 ( .A(n8734), .ZN(n7820) );
  NAND2_X1 U6530 ( .A1(n6872), .A2(n6871), .ZN(n6889) );
  INV_X1 U6531 ( .A(n8338), .ZN(n8393) );
  INV_X1 U6532 ( .A(n10372), .ZN(n8104) );
  INV_X1 U6533 ( .A(n8381), .ZN(n7963) );
  NAND2_X1 U6534 ( .A1(n6116), .A2(n6351), .ZN(n7594) );
  INV_X1 U6535 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6312) );
  AND2_X1 U6536 ( .A1(n5209), .A2(n5208), .ZN(n5502) );
  AND2_X1 U6537 ( .A1(n5198), .A2(n5197), .ZN(n5455) );
  AND2_X1 U6538 ( .A1(n5186), .A2(n5185), .ZN(n5403) );
  INV_X1 U6539 ( .A(n7109), .ZN(n6810) );
  AND2_X1 U6540 ( .A1(n5718), .A2(n5717), .ZN(n8602) );
  AND3_X1 U6541 ( .A1(n5630), .A2(n5629), .A3(n5628), .ZN(n8932) );
  AND4_X1 U6542 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n7921)
         );
  INV_X1 U6543 ( .A(n10466), .ZN(n9041) );
  NAND2_X1 U6544 ( .A1(n5904), .A2(n5912), .ZN(n8901) );
  AND2_X1 U6545 ( .A1(n9006), .A2(n9005), .ZN(n9150) );
  INV_X1 U6546 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6547 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  AND2_X1 U6548 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6037) );
  OAI21_X1 U6549 ( .B1(n6458), .B2(n6457), .A(n6459), .ZN(n7065) );
  AOI22_X1 U6550 ( .A1(n8513), .A2(n8512), .B1(n8511), .B2(n8510), .ZN(n8514)
         );
  OR3_X1 U6551 ( .A1(n9389), .A2(n9387), .A3(n9386), .ZN(n9412) );
  NOR2_X1 U6552 ( .A1(n10413), .A2(n6430), .ZN(n6431) );
  XNOR2_X1 U6553 ( .A(n5683), .B(n5682), .ZN(n8081) );
  INV_X1 U6554 ( .A(n6392), .ZN(n7479) );
  AND2_X1 U6555 ( .A1(n7122), .A2(n7121), .ZN(n8711) );
  INV_X1 U6556 ( .A(n5927), .ZN(n8849) );
  INV_X1 U6557 ( .A(n6896), .ZN(n8860) );
  INV_X1 U6558 ( .A(n10433), .ZN(n9024) );
  INV_X1 U6559 ( .A(n10570), .ZN(n10568) );
  INV_X1 U6560 ( .A(n9243), .ZN(n9288) );
  INV_X1 U6561 ( .A(n6637), .ZN(n9294) );
  OR2_X1 U6562 ( .A1(n6301), .A2(n6300), .ZN(n9650) );
  INV_X1 U6563 ( .A(n10242), .ZN(n9635) );
  INV_X1 U6564 ( .A(n10413), .ZN(n10411) );
  NAND2_X1 U6565 ( .A1(n5161), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5155) );
  INV_X1 U6566 ( .A(n5159), .ZN(n5158) );
  INV_X1 U6567 ( .A(SI_2_), .ZN(n5157) );
  NAND2_X1 U6568 ( .A1(n5158), .A2(n5157), .ZN(n5160) );
  INV_X4 U6569 ( .A(n5161), .ZN(n8151) );
  OAI211_X1 U6570 ( .C1(SI_1_), .C2(P1_DATAO_REG_1__SCAN_IN), .A(SI_0_), .B(
        P1_DATAO_REG_0__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6571 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5162) );
  OAI211_X1 U6572 ( .C1(SI_1_), .C2(P2_DATAO_REG_1__SCAN_IN), .A(SI_0_), .B(
        P2_DATAO_REG_0__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6573 ( .A1(SI_1_), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6574 ( .A1(n5165), .A2(n5164), .ZN(n5166) );
  NAND2_X1 U6575 ( .A1(n5349), .A2(n5172), .ZN(n5370) );
  INV_X1 U6576 ( .A(n5175), .ZN(n5174) );
  INV_X1 U6577 ( .A(SI_4_), .ZN(n10127) );
  NAND2_X1 U6578 ( .A1(n5174), .A2(n10127), .ZN(n5176) );
  NAND2_X1 U6579 ( .A1(n5370), .A2(n5369), .ZN(n5368) );
  NAND2_X1 U6580 ( .A1(n5368), .A2(n5177), .ZN(n5379) );
  INV_X1 U6581 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6582 ( .A1(n5179), .A2(n9975), .ZN(n5180) );
  NAND2_X1 U6583 ( .A1(n5182), .A2(SI_6_), .ZN(n5186) );
  INV_X1 U6584 ( .A(n5182), .ZN(n5184) );
  INV_X1 U6585 ( .A(SI_6_), .ZN(n5183) );
  NAND2_X1 U6586 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  NAND2_X1 U6587 ( .A1(n5187), .A2(SI_7_), .ZN(n5190) );
  INV_X1 U6588 ( .A(n5187), .ZN(n5188) );
  INV_X1 U6589 ( .A(SI_7_), .ZN(n9940) );
  NAND2_X1 U6590 ( .A1(n5188), .A2(n9940), .ZN(n5189) );
  INV_X1 U6591 ( .A(n5191), .ZN(n5192) );
  INV_X1 U6592 ( .A(SI_8_), .ZN(n10073) );
  INV_X1 U6593 ( .A(SI_9_), .ZN(n9886) );
  MUX2_X1 U6594 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6914), .Z(n5195) );
  NAND2_X1 U6595 ( .A1(n5195), .A2(SI_10_), .ZN(n5198) );
  INV_X1 U6596 ( .A(n5195), .ZN(n5196) );
  INV_X1 U6597 ( .A(SI_10_), .ZN(n10085) );
  NAND2_X1 U6598 ( .A1(n5196), .A2(n10085), .ZN(n5197) );
  MUX2_X1 U6599 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6914), .Z(n5199) );
  INV_X1 U6600 ( .A(n5199), .ZN(n5200) );
  INV_X1 U6601 ( .A(SI_11_), .ZN(n10104) );
  NAND2_X1 U6602 ( .A1(n5201), .A2(SI_12_), .ZN(n5205) );
  INV_X1 U6603 ( .A(n5201), .ZN(n5203) );
  INV_X1 U6604 ( .A(SI_12_), .ZN(n5202) );
  NAND2_X1 U6605 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U6606 ( .A1(n5205), .A2(n5204), .ZN(n5486) );
  NAND2_X1 U6607 ( .A1(n5489), .A2(n5205), .ZN(n5503) );
  MUX2_X1 U6608 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6914), .Z(n5206) );
  NAND2_X1 U6609 ( .A1(n5206), .A2(SI_13_), .ZN(n5209) );
  INV_X1 U6610 ( .A(n5206), .ZN(n5207) );
  INV_X1 U6611 ( .A(SI_13_), .ZN(n9857) );
  NAND2_X1 U6612 ( .A1(n5207), .A2(n9857), .ZN(n5208) );
  NAND2_X1 U6613 ( .A1(n5503), .A2(n5502), .ZN(n5505) );
  NAND2_X1 U6614 ( .A1(n5538), .A2(SI_15_), .ZN(n5211) );
  MUX2_X1 U6615 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6914), .Z(n5536) );
  INV_X1 U6616 ( .A(n5536), .ZN(n5210) );
  NAND2_X1 U6617 ( .A1(n5211), .A2(n5210), .ZN(n5215) );
  INV_X1 U6618 ( .A(SI_15_), .ZN(n5212) );
  NAND2_X1 U6619 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  INV_X1 U6620 ( .A(n5551), .ZN(n5216) );
  INV_X1 U6621 ( .A(SI_16_), .ZN(n5550) );
  NAND2_X1 U6622 ( .A1(n5551), .A2(SI_16_), .ZN(n5217) );
  INV_X1 U6623 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5218) );
  INV_X1 U6624 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9970) );
  INV_X1 U6625 ( .A(SI_17_), .ZN(n5219) );
  NAND2_X1 U6626 ( .A1(n5220), .A2(n5219), .ZN(n5223) );
  INV_X1 U6627 ( .A(n5220), .ZN(n5221) );
  NAND2_X1 U6628 ( .A1(n5221), .A2(SI_17_), .ZN(n5222) );
  NAND2_X1 U6629 ( .A1(n5223), .A2(n5222), .ZN(n5564) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7569) );
  INV_X1 U6631 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9837) );
  MUX2_X1 U6632 ( .A(n7569), .B(n9837), .S(n6914), .Z(n5224) );
  XNOR2_X1 U6633 ( .A(n5224), .B(SI_18_), .ZN(n5578) );
  INV_X1 U6634 ( .A(n5578), .ZN(n5227) );
  INV_X1 U6635 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6636 ( .A1(n5225), .A2(SI_18_), .ZN(n5226) );
  INV_X1 U6637 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7658) );
  INV_X1 U6638 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7657) );
  INV_X1 U6639 ( .A(SI_19_), .ZN(n5228) );
  NAND2_X1 U6640 ( .A1(n5229), .A2(n5228), .ZN(n5232) );
  INV_X1 U6641 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6642 ( .A1(n5230), .A2(SI_19_), .ZN(n5231) );
  NAND2_X1 U6643 ( .A1(n5232), .A2(n5231), .ZN(n5590) );
  INV_X1 U6644 ( .A(SI_20_), .ZN(n9918) );
  MUX2_X1 U6645 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6914), .Z(n5607) );
  INV_X1 U6646 ( .A(n5607), .ZN(n5233) );
  NAND2_X1 U6647 ( .A1(n5609), .A2(n9918), .ZN(n5234) );
  INV_X1 U6648 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7803) );
  INV_X1 U6649 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7761) );
  MUX2_X1 U6650 ( .A(n7803), .B(n7761), .S(n6914), .Z(n5620) );
  AND2_X1 U6651 ( .A1(n5620), .A2(n10075), .ZN(n5238) );
  INV_X1 U6652 ( .A(n5620), .ZN(n5236) );
  NAND2_X1 U6653 ( .A1(n5236), .A2(SI_21_), .ZN(n5237) );
  INV_X1 U6654 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7877) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10072) );
  INV_X1 U6656 ( .A(SI_22_), .ZN(n9906) );
  NAND2_X1 U6657 ( .A1(n5239), .A2(n9906), .ZN(n5242) );
  INV_X1 U6658 ( .A(n5239), .ZN(n5240) );
  NAND2_X1 U6659 ( .A1(n5240), .A2(SI_22_), .ZN(n5241) );
  NAND2_X1 U6660 ( .A1(n5242), .A2(n5241), .ZN(n5631) );
  INV_X1 U6661 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7896) );
  INV_X1 U6662 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7891) );
  MUX2_X1 U6663 ( .A(n7896), .B(n7891), .S(n6914), .Z(n5244) );
  INV_X1 U6664 ( .A(SI_23_), .ZN(n5243) );
  NAND2_X1 U6665 ( .A1(n5244), .A2(n5243), .ZN(n5247) );
  INV_X1 U6666 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6667 ( .A1(n5245), .A2(SI_23_), .ZN(n5246) );
  AND2_X1 U6668 ( .A1(n5247), .A2(n5246), .ZN(n5644) );
  NAND2_X1 U6669 ( .A1(n5248), .A2(n5247), .ZN(n5656) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7994) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U6672 ( .A1(n5249), .A2(n9937), .ZN(n5252) );
  INV_X1 U6673 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6674 ( .A1(n5250), .A2(SI_24_), .ZN(n5251) );
  AND2_X1 U6675 ( .A1(n5252), .A2(n5251), .ZN(n5657) );
  NAND2_X1 U6676 ( .A1(n5656), .A2(n5657), .ZN(n5253) );
  NAND2_X1 U6677 ( .A1(n5253), .A2(n5252), .ZN(n5669) );
  INV_X1 U6678 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8050) );
  INV_X1 U6679 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8037) );
  MUX2_X1 U6680 ( .A(n8050), .B(n8037), .S(n6914), .Z(n5255) );
  INV_X1 U6681 ( .A(SI_25_), .ZN(n5254) );
  NAND2_X1 U6682 ( .A1(n5255), .A2(n5254), .ZN(n5258) );
  INV_X1 U6683 ( .A(n5255), .ZN(n5256) );
  NAND2_X1 U6684 ( .A1(n5256), .A2(SI_25_), .ZN(n5257) );
  AND2_X1 U6685 ( .A1(n5258), .A2(n5257), .ZN(n5670) );
  INV_X1 U6686 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8096) );
  INV_X1 U6687 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8083) );
  MUX2_X1 U6688 ( .A(n8096), .B(n8083), .S(n6914), .Z(n5259) );
  INV_X1 U6689 ( .A(SI_26_), .ZN(n9845) );
  NAND2_X1 U6690 ( .A1(n5259), .A2(n9845), .ZN(n5262) );
  INV_X1 U6691 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6692 ( .A1(n5260), .A2(SI_26_), .ZN(n5261) );
  AND2_X1 U6693 ( .A1(n5262), .A2(n5261), .ZN(n5682) );
  INV_X1 U6694 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5695) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10101) );
  MUX2_X1 U6696 ( .A(n5695), .B(n10101), .S(n6914), .Z(n5264) );
  INV_X1 U6697 ( .A(SI_27_), .ZN(n5263) );
  NAND2_X1 U6698 ( .A1(n5264), .A2(n5263), .ZN(n5267) );
  INV_X1 U6699 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6700 ( .A1(n5265), .A2(SI_27_), .ZN(n5266) );
  AND2_X1 U6701 ( .A1(n5267), .A2(n5266), .ZN(n5693) );
  NAND2_X1 U6702 ( .A1(n5694), .A2(n5693), .ZN(n5268) );
  NAND2_X1 U6703 ( .A1(n5268), .A2(n5267), .ZN(n5707) );
  INV_X1 U6704 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5709) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8576) );
  XNOR2_X1 U6706 ( .A(n5269), .B(SI_28_), .ZN(n5708) );
  NAND2_X1 U6707 ( .A1(n5707), .A2(n5708), .ZN(n5271) );
  INV_X1 U6708 ( .A(SI_28_), .ZN(n10070) );
  NAND2_X1 U6709 ( .A1(n5269), .A2(n10070), .ZN(n5270) );
  INV_X1 U6710 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9166) );
  INV_X1 U6711 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9755) );
  INV_X1 U6712 ( .A(SI_29_), .ZN(n5275) );
  INV_X1 U6713 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9951) );
  INV_X1 U6714 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8578) );
  MUX2_X1 U6715 ( .A(n9951), .B(n8578), .S(n8151), .Z(n5276) );
  INV_X1 U6716 ( .A(SI_30_), .ZN(n10088) );
  NAND2_X1 U6717 ( .A1(n5276), .A2(n10088), .ZN(n5279) );
  INV_X1 U6718 ( .A(n5276), .ZN(n5277) );
  NAND2_X1 U6719 ( .A1(n5277), .A2(SI_30_), .ZN(n5278) );
  NAND2_X1 U6720 ( .A1(n5279), .A2(n5278), .ZN(n5728) );
  MUX2_X1 U6721 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8151), .Z(n5280) );
  XNOR2_X1 U6722 ( .A(n5280), .B(SI_31_), .ZN(n5281) );
  NAND4_X1 U6723 ( .A1(n5522), .A2(n5525), .A3(n5470), .A4(n5475), .ZN(n5287)
         );
  NOR2_X1 U6724 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5290) );
  NOR2_X1 U6725 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5289) );
  INV_X1 U6726 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5581) );
  INV_X1 U6727 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5782) );
  NOR3_X1 U6728 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5291) );
  INV_X1 U6729 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5294) );
  INV_X1 U6730 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6731 ( .A1(n6866), .A2(n8151), .ZN(n5336) );
  INV_X1 U6732 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5296) );
  OAI22_X1 U6733 ( .A1(n8153), .A2(n5336), .B1(n5319), .B2(n5296), .ZN(n5926)
         );
  INV_X1 U6734 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6735 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5300) );
  NAND2_X1 U6736 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  XNOR2_X2 U6737 ( .A(n5302), .B(n5297), .ZN(n5304) );
  AND2_X2 U6738 ( .A1(n8580), .A2(n5304), .ZN(n5359) );
  NAND2_X1 U6739 ( .A1(n4525), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6740 ( .A1(n5344), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6741 ( .A1(n4523), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5305) );
  NAND4_X1 U6742 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n7109)
         );
  NAND2_X1 U6743 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5309) );
  INV_X1 U6744 ( .A(n5339), .ZN(n5310) );
  INV_X1 U6745 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6937) );
  INV_X1 U6746 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U6747 ( .A1(n5312), .A2(SI_0_), .ZN(n5313) );
  XNOR2_X1 U6748 ( .A(n5314), .B(n5313), .ZN(n5317) );
  INV_X1 U6749 ( .A(n5317), .ZN(n5315) );
  INV_X1 U6750 ( .A(SI_1_), .ZN(n5316) );
  NAND2_X1 U6751 ( .A1(n5317), .A2(n5316), .ZN(n5318) );
  NAND2_X1 U6752 ( .A1(n6810), .A2(n10473), .ZN(n5800) );
  NAND2_X1 U6753 ( .A1(n5796), .A2(n5800), .ZN(n6809) );
  INV_X1 U6754 ( .A(n6809), .ZN(n5325) );
  NAND2_X1 U6755 ( .A1(n4525), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6756 ( .A1(n4523), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6757 ( .A1(n5344), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6758 ( .A1(n5359), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5320) );
  NAND4_X1 U6759 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n8739)
         );
  INV_X1 U6760 ( .A(n8739), .ZN(n10457) );
  NAND2_X1 U6761 ( .A1(n8151), .A2(SI_0_), .ZN(n5324) );
  XNOR2_X1 U6762 ( .A(n5324), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9168) );
  MUX2_X1 U6763 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9168), .S(n6866), .Z(n8583) );
  NAND2_X1 U6764 ( .A1(n10457), .A2(n8583), .ZN(n7114) );
  INV_X1 U6765 ( .A(n7114), .ZN(n10453) );
  NAND2_X1 U6766 ( .A1(n5325), .A2(n10453), .ZN(n10452) );
  NAND2_X1 U6767 ( .A1(n4525), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6768 ( .A1(n4523), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6769 ( .A1(n5359), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6770 ( .A1(n5344), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5326) );
  INV_X1 U6771 ( .A(n5330), .ZN(n5333) );
  INV_X1 U6772 ( .A(n5331), .ZN(n5332) );
  NAND2_X1 U6773 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  NAND2_X1 U6774 ( .A1(n5335), .A2(n5334), .ZN(n6948) );
  OR2_X1 U6775 ( .A1(n5336), .A2(n6948), .ZN(n5342) );
  NOR2_X1 U6776 ( .A1(n5339), .A2(n8146), .ZN(n5338) );
  NAND2_X1 U6777 ( .A1(n10455), .A2(n7144), .ZN(n5806) );
  NAND2_X1 U6778 ( .A1(n10479), .A2(n10426), .ZN(n5804) );
  INV_X1 U6779 ( .A(n10440), .ZN(n5761) );
  NAND2_X1 U6780 ( .A1(n10436), .A2(n5761), .ZN(n5343) );
  NAND2_X1 U6781 ( .A1(n5343), .A2(n5806), .ZN(n10430) );
  NAND2_X1 U6782 ( .A1(n4526), .A2(n9833), .ZN(n5348) );
  NAND2_X1 U6783 ( .A1(n5734), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6784 ( .A1(n5359), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6785 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  NAND2_X1 U6786 ( .A1(n5349), .A2(n5352), .ZN(n6928) );
  OR2_X1 U6787 ( .A1(n5336), .A2(n6928), .ZN(n5357) );
  NAND2_X1 U6788 ( .A1(n5353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5355) );
  INV_X1 U6789 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5354) );
  OR2_X1 U6790 ( .A1(n5319), .A2(n5169), .ZN(n5356) );
  XNOR2_X1 U6791 ( .A(n8738), .B(n7168), .ZN(n10431) );
  NAND2_X1 U6792 ( .A1(n10430), .A2(n10431), .ZN(n5358) );
  INV_X1 U6793 ( .A(n8738), .ZN(n10441) );
  NAND2_X1 U6794 ( .A1(n5358), .A2(n5819), .ZN(n7375) );
  NAND2_X1 U6795 ( .A1(n5359), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6796 ( .A1(n4523), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6797 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5360) );
  NAND2_X1 U6798 ( .A1(n5386), .A2(n5360), .ZN(n8664) );
  NAND2_X1 U6799 ( .A1(n4526), .A2(n8664), .ZN(n5362) );
  NAND2_X1 U6800 ( .A1(n5733), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5361) );
  NAND4_X1 U6801 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), .ZN(n10428)
         );
  NAND2_X1 U6802 ( .A1(n5365), .A2(n5339), .ZN(n5366) );
  NAND2_X1 U6803 ( .A1(n5366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5367) );
  OR2_X1 U6804 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6805 ( .A1(n5368), .A2(n5371), .ZN(n6927) );
  OR2_X1 U6806 ( .A1(n5336), .A2(n6927), .ZN(n5373) );
  OR2_X1 U6807 ( .A1(n5319), .A2(n5173), .ZN(n5372) );
  OAI211_X1 U6808 ( .C1(n6866), .C2(n7261), .A(n5373), .B(n5372), .ZN(n8663)
         );
  INV_X1 U6809 ( .A(n8663), .ZN(n10489) );
  NAND2_X1 U6810 ( .A1(n7330), .A2(n10489), .ZN(n6818) );
  INV_X1 U6811 ( .A(n6820), .ZN(n5374) );
  NAND2_X1 U6812 ( .A1(n7375), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U6813 ( .A1(n7330), .A2(n8663), .ZN(n5814) );
  OR2_X1 U6814 ( .A1(n5375), .A2(n8146), .ZN(n5377) );
  XNOR2_X1 U6815 ( .A(n5377), .B(n5376), .ZN(n6932) );
  OR2_X1 U6816 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND2_X1 U6817 ( .A1(n5381), .A2(n5380), .ZN(n6931) );
  OR2_X1 U6818 ( .A1(n5336), .A2(n6931), .ZN(n5383) );
  INV_X1 U6819 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6930) );
  OR2_X1 U6820 ( .A1(n5319), .A2(n6930), .ZN(n5382) );
  OAI211_X1 U6821 ( .C1(n6866), .C2(n6932), .A(n5383), .B(n5382), .ZN(n10495)
         );
  INV_X1 U6822 ( .A(n10495), .ZN(n6821) );
  NAND2_X1 U6823 ( .A1(n5359), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6824 ( .A1(n4523), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6825 ( .A1(n5386), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6826 ( .A1(n5392), .A2(n5387), .ZN(n7427) );
  NAND2_X1 U6827 ( .A1(n4526), .A2(n7427), .ZN(n5389) );
  NAND2_X1 U6828 ( .A1(n5733), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5388) );
  NOR2_X1 U6829 ( .A1(n6821), .A2(n9035), .ZN(n5813) );
  NAND2_X1 U6830 ( .A1(n6821), .A2(n9035), .ZN(n5821) );
  OAI21_X1 U6831 ( .B1(n7425), .B2(n5813), .A(n5821), .ZN(n9043) );
  NAND2_X1 U6832 ( .A1(n5359), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6833 ( .A1(n4523), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6834 ( .A1(n5392), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6835 ( .A1(n5411), .A2(n5393), .ZN(n9039) );
  NAND2_X1 U6836 ( .A1(n4526), .A2(n9039), .ZN(n5395) );
  NAND2_X1 U6837 ( .A1(n5733), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5394) );
  NAND4_X1 U6838 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n8737)
         );
  INV_X1 U6839 ( .A(n8737), .ZN(n7646) );
  NOR2_X1 U6840 ( .A1(n5398), .A2(n8146), .ZN(n5399) );
  MUX2_X1 U6841 ( .A(n8146), .B(n5399), .S(P2_IR_REG_6__SCAN_IN), .Z(n5401) );
  OR2_X1 U6842 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U6843 ( .A1(n5402), .A2(n5405), .ZN(n6934) );
  OR2_X1 U6844 ( .A1(n5336), .A2(n6934), .ZN(n5407) );
  INV_X1 U6845 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6933) );
  OR2_X1 U6846 ( .A1(n5319), .A2(n6933), .ZN(n5406) );
  NAND2_X1 U6847 ( .A1(n7646), .A2(n10505), .ZN(n5828) );
  INV_X1 U6848 ( .A(n10505), .ZN(n5408) );
  NAND2_X1 U6849 ( .A1(n5408), .A2(n8737), .ZN(n5826) );
  NAND2_X1 U6850 ( .A1(n9043), .A2(n9042), .ZN(n10500) );
  NAND2_X1 U6851 ( .A1(n5359), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6852 ( .A1(n5734), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5415) );
  INV_X1 U6853 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6854 ( .A1(n5411), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6855 ( .A1(n5430), .A2(n5412), .ZN(n8593) );
  NAND2_X1 U6856 ( .A1(n4526), .A2(n8593), .ZN(n5414) );
  NAND2_X1 U6857 ( .A1(n5733), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5413) );
  NAND4_X1 U6858 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n9036)
         );
  INV_X1 U6859 ( .A(n9036), .ZN(n7544) );
  NAND2_X1 U6860 ( .A1(n5400), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5417) );
  MUX2_X1 U6861 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5417), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5418) );
  NAND2_X1 U6862 ( .A1(n5418), .A2(n5438), .ZN(n7363) );
  OR2_X1 U6863 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U6864 ( .A1(n5419), .A2(n5422), .ZN(n6926) );
  OR2_X1 U6865 ( .A1(n5336), .A2(n6926), .ZN(n5424) );
  INV_X1 U6866 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6925) );
  OR2_X1 U6867 ( .A1(n5319), .A2(n6925), .ZN(n5423) );
  OAI211_X1 U6868 ( .C1(n6866), .C2(n7363), .A(n5424), .B(n5423), .ZN(n8592)
         );
  NAND2_X1 U6869 ( .A1(n7544), .A2(n8592), .ZN(n5836) );
  INV_X1 U6870 ( .A(n8592), .ZN(n10507) );
  NAND2_X1 U6871 ( .A1(n10507), .A2(n9036), .ZN(n7698) );
  NAND2_X1 U6872 ( .A1(n5438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U6873 ( .A(n5425), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7416) );
  XNOR2_X1 U6874 ( .A(n5426), .B(n5427), .ZN(n6950) );
  NAND2_X1 U6875 ( .A1(n6950), .A2(n5730), .ZN(n5429) );
  INV_X1 U6876 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6951) );
  OR2_X1 U6877 ( .A1(n5319), .A2(n6951), .ZN(n5428) );
  OAI211_X1 U6878 ( .C1(n6866), .C2(n6952), .A(n5429), .B(n5428), .ZN(n10513)
         );
  INV_X1 U6879 ( .A(n10513), .ZN(n7704) );
  NAND2_X1 U6880 ( .A1(n5359), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6881 ( .A1(n4523), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5434) );
  OR2_X2 U6882 ( .A1(n5430), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6883 ( .A1(n5430), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6884 ( .A1(n5446), .A2(n5431), .ZN(n7702) );
  NAND2_X1 U6885 ( .A1(n4526), .A2(n7702), .ZN(n5433) );
  NAND2_X1 U6886 ( .A1(n5733), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6887 ( .A1(n7704), .A2(n8736), .ZN(n5832) );
  NAND2_X1 U6888 ( .A1(n7714), .A2(n10513), .ZN(n5841) );
  INV_X1 U6889 ( .A(n7708), .ZN(n5453) );
  NAND2_X1 U6890 ( .A1(n6955), .A2(n5730), .ZN(n5443) );
  OR2_X1 U6891 ( .A1(n5438), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6892 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5440) );
  INV_X1 U6893 ( .A(n5440), .ZN(n5439) );
  NAND2_X1 U6894 ( .A1(n5439), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6895 ( .A1(n5440), .A2(n5470), .ZN(n5459) );
  AND2_X1 U6896 ( .A1(n5441), .A2(n5459), .ZN(n7563) );
  AOI22_X1 U6897 ( .A1(n5596), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5595), .B2(
        n7563), .ZN(n5442) );
  NAND2_X1 U6898 ( .A1(n5359), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6899 ( .A1(n5734), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5450) );
  INV_X1 U6900 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6901 ( .A1(n5446), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6902 ( .A1(n5480), .A2(n5447), .ZN(n7613) );
  NAND2_X1 U6903 ( .A1(n4526), .A2(n7613), .ZN(n5449) );
  NAND2_X1 U6904 ( .A1(n5733), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5448) );
  NAND4_X1 U6905 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n8735)
         );
  NAND2_X1 U6906 ( .A1(n10518), .A2(n7780), .ZN(n5840) );
  NAND2_X1 U6907 ( .A1(n5843), .A2(n5840), .ZN(n7711) );
  NAND2_X1 U6908 ( .A1(n5456), .A2(n4945), .ZN(n5457) );
  NAND2_X1 U6909 ( .A1(n5458), .A2(n5457), .ZN(n6958) );
  OR2_X1 U6910 ( .A1(n6958), .A2(n5336), .ZN(n5462) );
  NAND2_X1 U6911 ( .A1(n5459), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6912 ( .A(n5460), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7676) );
  AOI22_X1 U6913 ( .A1(n5596), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5595), .B2(
        n7676), .ZN(n5461) );
  NAND2_X1 U6914 ( .A1(n5359), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6915 ( .A1(n5734), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U6916 ( .A(n5480), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U6917 ( .A1(n4526), .A2(n7762), .ZN(n5464) );
  NAND2_X1 U6918 ( .A1(n5733), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5463) );
  NAND4_X1 U6919 ( .A1(n5466), .A2(n5465), .A3(n5464), .A4(n5463), .ZN(n8734)
         );
  NAND2_X1 U6920 ( .A1(n7788), .A2(n7820), .ZN(n5846) );
  XNOR2_X1 U6921 ( .A(n5468), .B(n5467), .ZN(n6963) );
  NAND2_X1 U6922 ( .A1(n6963), .A2(n5730), .ZN(n5479) );
  NAND2_X1 U6923 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NOR2_X1 U6924 ( .A1(n5472), .A2(n5471), .ZN(n5476) );
  NOR2_X1 U6925 ( .A1(n5476), .A2(n8146), .ZN(n5473) );
  MUX2_X1 U6926 ( .A(n8146), .B(n5473), .S(P2_IR_REG_11__SCAN_IN), .Z(n5474)
         );
  INV_X1 U6927 ( .A(n5474), .ZN(n5477) );
  NAND2_X1 U6928 ( .A1(n5476), .A2(n5475), .ZN(n5506) );
  AND2_X1 U6929 ( .A1(n5477), .A2(n5506), .ZN(n7745) );
  AOI22_X1 U6930 ( .A1(n5596), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5595), .B2(
        n7745), .ZN(n5478) );
  NAND2_X1 U6931 ( .A1(n5479), .A2(n5478), .ZN(n10536) );
  NAND2_X1 U6932 ( .A1(n5359), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6933 ( .A1(n5734), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5484) );
  OAI21_X1 U6934 ( .B1(n5480), .B2(P2_REG3_REG_10__SCAN_IN), .A(
        P2_REG3_REG_11__SCAN_IN), .ZN(n5481) );
  OR3_X2 U6935 ( .A1(n5480), .A2(P2_REG3_REG_11__SCAN_IN), .A3(
        P2_REG3_REG_10__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6936 ( .A1(n5481), .A2(n5495), .ZN(n7822) );
  NAND2_X1 U6937 ( .A1(n4526), .A2(n7822), .ZN(n5483) );
  NAND2_X1 U6938 ( .A1(n5733), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6939 ( .A1(n10536), .A2(n7921), .ZN(n5851) );
  NAND2_X1 U6940 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  NAND2_X1 U6941 ( .A1(n5489), .A2(n5488), .ZN(n7024) );
  OR2_X1 U6942 ( .A1(n7024), .A2(n5336), .ZN(n5492) );
  NAND2_X1 U6943 ( .A1(n5506), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5490) );
  XNOR2_X1 U6944 ( .A(n5490), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U6945 ( .A1(n5596), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5595), .B2(
        n6763), .ZN(n5491) );
  NAND2_X1 U6946 ( .A1(n5492), .A2(n5491), .ZN(n7863) );
  NAND2_X1 U6947 ( .A1(n4522), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6948 ( .A1(n5734), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5499) );
  INV_X1 U6949 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6950 ( .A1(n5495), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6951 ( .A1(n5511), .A2(n5496), .ZN(n7924) );
  NAND2_X1 U6952 ( .A1(n4525), .A2(n7924), .ZN(n5498) );
  NAND2_X1 U6953 ( .A1(n5733), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5497) );
  NAND4_X1 U6954 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n8732)
         );
  INV_X1 U6955 ( .A(n8732), .ZN(n7821) );
  OR2_X1 U6956 ( .A1(n7863), .A2(n7821), .ZN(n5856) );
  NAND2_X1 U6957 ( .A1(n7863), .A2(n7821), .ZN(n5855) );
  NAND2_X1 U6958 ( .A1(n7923), .A2(n7922), .ZN(n5501) );
  NAND2_X1 U6959 ( .A1(n5501), .A2(n5856), .ZN(n7966) );
  OR2_X1 U6960 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  NAND2_X1 U6961 ( .A1(n5505), .A2(n5504), .ZN(n7074) );
  OR2_X1 U6962 ( .A1(n7074), .A2(n5336), .ZN(n5509) );
  OR2_X1 U6963 ( .A1(n5506), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6964 ( .A1(n5507), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5523) );
  XNOR2_X1 U6965 ( .A(n5523), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8754) );
  AOI22_X1 U6966 ( .A1(n5596), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5595), .B2(
        n8754), .ZN(n5508) );
  NAND2_X1 U6967 ( .A1(n4522), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6968 ( .A1(n4523), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5515) );
  INV_X1 U6969 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U6970 ( .A1(n5511), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6971 ( .A1(n5530), .A2(n5512), .ZN(n7978) );
  NAND2_X1 U6972 ( .A1(n4525), .A2(n7978), .ZN(n5514) );
  NAND2_X1 U6973 ( .A1(n5733), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5513) );
  NAND4_X1 U6974 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n8731)
         );
  INV_X1 U6975 ( .A(n8731), .ZN(n7931) );
  NOR2_X1 U6976 ( .A1(n7930), .A2(n7931), .ZN(n5518) );
  NAND2_X1 U6977 ( .A1(n7930), .A2(n7931), .ZN(n5517) );
  XNOR2_X1 U6978 ( .A(n5520), .B(SI_14_), .ZN(n5521) );
  XNOR2_X1 U6979 ( .A(n5519), .B(n5521), .ZN(n7171) );
  NAND2_X1 U6980 ( .A1(n7171), .A2(n5730), .ZN(n5529) );
  NAND2_X1 U6981 ( .A1(n5523), .A2(n5522), .ZN(n5524) );
  NAND2_X1 U6982 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5526) );
  OR2_X1 U6983 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U6984 ( .A1(n5526), .A2(n5525), .ZN(n5539) );
  AND2_X1 U6985 ( .A1(n5527), .A2(n5539), .ZN(n8767) );
  AOI22_X1 U6986 ( .A1(n5596), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5595), .B2(
        n8767), .ZN(n5528) );
  NAND2_X1 U6987 ( .A1(n4522), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6988 ( .A1(n4523), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U6989 ( .A1(n5530), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6990 ( .A1(n5544), .A2(n5531), .ZN(n9029) );
  NAND2_X1 U6991 ( .A1(n4526), .A2(n9029), .ZN(n5533) );
  NAND2_X1 U6992 ( .A1(n5733), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5532) );
  NAND4_X1 U6993 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n8730)
         );
  INV_X1 U6994 ( .A(n8730), .ZN(n7940) );
  OR2_X1 U6995 ( .A1(n8078), .A2(n7940), .ZN(n5861) );
  NAND2_X1 U6996 ( .A1(n8078), .A2(n7940), .ZN(n5862) );
  XNOR2_X1 U6997 ( .A(n5536), .B(SI_15_), .ZN(n5537) );
  XNOR2_X1 U6998 ( .A(n5538), .B(n5537), .ZN(n7277) );
  NAND2_X1 U6999 ( .A1(n7277), .A2(n5730), .ZN(n5542) );
  NAND2_X1 U7000 ( .A1(n5539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5540) );
  XNOR2_X1 U7001 ( .A(n5540), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8785) );
  AOI22_X1 U7002 ( .A1(n5596), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5595), .B2(
        n8785), .ZN(n5541) );
  NAND2_X1 U7003 ( .A1(n4522), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7004 ( .A1(n5734), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5548) );
  INV_X1 U7005 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U7006 ( .A1(n5544), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7007 ( .A1(n5558), .A2(n5545), .ZN(n8721) );
  NAND2_X1 U7008 ( .A1(n4525), .A2(n8721), .ZN(n5547) );
  NAND2_X1 U7009 ( .A1(n5733), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5546) );
  NAND4_X1 U7010 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n9017)
         );
  INV_X1 U7011 ( .A(n9017), .ZN(n8536) );
  AND2_X1 U7012 ( .A1(n9012), .A2(n8536), .ZN(n5880) );
  OR2_X1 U7013 ( .A1(n9012), .A2(n8536), .ZN(n5865) );
  XNOR2_X1 U7014 ( .A(n5551), .B(n5550), .ZN(n5552) );
  XNOR2_X1 U7015 ( .A(n5553), .B(n5552), .ZN(n7348) );
  NAND2_X1 U7016 ( .A1(n7348), .A2(n5730), .ZN(n5557) );
  NAND2_X1 U7017 ( .A1(n5554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5555) );
  INV_X1 U7018 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5566) );
  XNOR2_X1 U7019 ( .A(n5555), .B(n5566), .ZN(n7385) );
  INV_X1 U7020 ( .A(n7385), .ZN(n8796) );
  AOI22_X1 U7021 ( .A1(n5596), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5595), .B2(
        n8796), .ZN(n5556) );
  NAND2_X1 U7022 ( .A1(n4522), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7023 ( .A1(n4523), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7024 ( .A1(n5558), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7025 ( .A1(n5571), .A2(n5559), .ZN(n9021) );
  NAND2_X1 U7026 ( .A1(n4526), .A2(n9021), .ZN(n5561) );
  NAND2_X1 U7027 ( .A1(n5733), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7028 ( .A1(n9158), .A2(n8718), .ZN(n5871) );
  OAI21_X1 U7029 ( .B1(n9011), .B2(n9015), .A(n5871), .ZN(n8999) );
  XNOR2_X1 U7030 ( .A(n5565), .B(n5564), .ZN(n7400) );
  NAND2_X1 U7031 ( .A1(n7400), .A2(n5730), .ZN(n5569) );
  NAND2_X1 U7032 ( .A1(n5580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7033 ( .A(n5567), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8822) );
  AOI22_X1 U7034 ( .A1(n5596), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5595), .B2(
        n8822), .ZN(n5568) );
  NAND2_X1 U7035 ( .A1(n5734), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7036 ( .A1(n5359), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5575) );
  INV_X1 U7037 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U7038 ( .A1(n5571), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7039 ( .A1(n5584), .A2(n5572), .ZN(n9007) );
  NAND2_X1 U7040 ( .A1(n4525), .A2(n9007), .ZN(n5574) );
  NAND2_X1 U7041 ( .A1(n5733), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5573) );
  OR2_X1 U7042 ( .A1(n9151), .A2(n8638), .ZN(n5883) );
  NAND2_X1 U7043 ( .A1(n9151), .A2(n8638), .ZN(n5870) );
  NAND2_X1 U7044 ( .A1(n5883), .A2(n5870), .ZN(n9001) );
  INV_X1 U7045 ( .A(n9001), .ZN(n5868) );
  NAND2_X1 U7046 ( .A1(n8999), .A2(n5868), .ZN(n5577) );
  NAND2_X1 U7047 ( .A1(n5577), .A2(n5870), .ZN(n8995) );
  XNOR2_X1 U7048 ( .A(n5579), .B(n5578), .ZN(n7567) );
  NAND2_X1 U7049 ( .A1(n7567), .A2(n5730), .ZN(n5583) );
  NAND2_X1 U7050 ( .A1(n5751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5592) );
  XNOR2_X1 U7051 ( .A(n5592), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8844) );
  AOI22_X1 U7052 ( .A1(n5596), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5595), .B2(
        n8844), .ZN(n5582) );
  NAND2_X1 U7053 ( .A1(n4522), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7054 ( .A1(n5734), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5588) );
  OR2_X2 U7055 ( .A1(n5584), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7056 ( .A1(n5584), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7057 ( .A1(n5601), .A2(n5585), .ZN(n8990) );
  NAND2_X1 U7058 ( .A1(n4526), .A2(n8990), .ZN(n5587) );
  NAND2_X1 U7059 ( .A1(n5733), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7060 ( .A1(n8994), .A2(n8977), .ZN(n5876) );
  XNOR2_X1 U7061 ( .A(n5591), .B(n5590), .ZN(n7656) );
  NAND2_X1 U7062 ( .A1(n7656), .A2(n5730), .ZN(n5598) );
  NAND2_X1 U7063 ( .A1(n5592), .A2(n5753), .ZN(n5593) );
  INV_X1 U7064 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5752) );
  INV_X1 U7065 ( .A(n7660), .ZN(n7376) );
  AOI22_X1 U7066 ( .A1(n5596), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7376), .B2(
        n5595), .ZN(n5597) );
  NAND2_X1 U7067 ( .A1(n5734), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7068 ( .A1(n5733), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5605) );
  INV_X1 U7069 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7070 ( .A1(n5601), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7071 ( .A1(n5614), .A2(n5602), .ZN(n8983) );
  NAND2_X1 U7072 ( .A1(n4526), .A2(n8983), .ZN(n5604) );
  NAND2_X1 U7073 ( .A1(n4522), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7074 ( .A1(n8984), .A2(n8697), .ZN(n5891) );
  NAND2_X1 U7075 ( .A1(n5890), .A2(n5891), .ZN(n6845) );
  INV_X1 U7076 ( .A(n6845), .ZN(n8973) );
  NAND2_X1 U7077 ( .A1(n8971), .A2(n5890), .ZN(n8959) );
  XNOR2_X1 U7078 ( .A(n5607), .B(n9918), .ZN(n5608) );
  XNOR2_X1 U7079 ( .A(n5609), .B(n5608), .ZN(n7707) );
  NAND2_X1 U7080 ( .A1(n7707), .A2(n5730), .ZN(n5611) );
  INV_X1 U7081 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7720) );
  OR2_X1 U7082 ( .A1(n4527), .A2(n7720), .ZN(n5610) );
  NAND2_X1 U7083 ( .A1(n4522), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7084 ( .A1(n4523), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5612) );
  AND2_X1 U7085 ( .A1(n5613), .A2(n5612), .ZN(n5618) );
  OR2_X2 U7086 ( .A1(n5614), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7087 ( .A1(n5614), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7088 ( .A1(n5626), .A2(n5615), .ZN(n8966) );
  NAND2_X1 U7089 ( .A1(n8966), .A2(n4526), .ZN(n5617) );
  NAND2_X1 U7090 ( .A1(n5733), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5616) );
  INV_X1 U7091 ( .A(n5895), .ZN(n5619) );
  XNOR2_X1 U7092 ( .A(n5620), .B(SI_21_), .ZN(n5621) );
  XNOR2_X1 U7093 ( .A(n5622), .B(n5621), .ZN(n7760) );
  NAND2_X1 U7094 ( .A1(n7760), .A2(n5730), .ZN(n5624) );
  OR2_X1 U7095 ( .A1(n5319), .A2(n7803), .ZN(n5623) );
  INV_X1 U7096 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U7097 ( .A1(n5626), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7098 ( .A1(n5635), .A2(n5627), .ZN(n8952) );
  NAND2_X1 U7099 ( .A1(n8952), .A2(n4526), .ZN(n5630) );
  AOI22_X1 U7100 ( .A1(n4522), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5734), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7101 ( .A1(n5733), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7102 ( .A1(n9072), .A2(n8932), .ZN(n5794) );
  NAND2_X1 U7103 ( .A1(n9138), .A2(n8978), .ZN(n8946) );
  AND2_X1 U7104 ( .A1(n5794), .A2(n8946), .ZN(n8935) );
  XNOR2_X1 U7105 ( .A(n5632), .B(n5631), .ZN(n7876) );
  NAND2_X1 U7106 ( .A1(n7876), .A2(n5730), .ZN(n5634) );
  OR2_X1 U7107 ( .A1(n5319), .A2(n7877), .ZN(n5633) );
  OR2_X2 U7108 ( .A1(n5635), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7109 ( .A1(n5635), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7110 ( .A1(n5648), .A2(n5636), .ZN(n8941) );
  NAND2_X1 U7111 ( .A1(n8941), .A2(n4525), .ZN(n5639) );
  AOI22_X1 U7112 ( .A1(n5359), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n4523), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7113 ( .A1(n5733), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7114 ( .A1(n8940), .A2(n8951), .ZN(n5899) );
  AND2_X1 U7115 ( .A1(n8935), .A2(n5899), .ZN(n5640) );
  INV_X1 U7116 ( .A(n5899), .ZN(n5642) );
  AND2_X1 U7117 ( .A1(n8936), .A2(n5898), .ZN(n5641) );
  XNOR2_X1 U7118 ( .A(n5645), .B(n5644), .ZN(n7893) );
  NAND2_X1 U7119 ( .A1(n7893), .A2(n5730), .ZN(n5647) );
  OR2_X1 U7120 ( .A1(n4527), .A2(n7896), .ZN(n5646) );
  INV_X1 U7121 ( .A(n9124), .ZN(n5655) );
  OR2_X2 U7122 ( .A1(n5648), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7123 ( .A1(n5648), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7124 ( .A1(n5661), .A2(n5649), .ZN(n8927) );
  NAND2_X1 U7125 ( .A1(n8927), .A2(n4526), .ZN(n5654) );
  INV_X1 U7126 ( .A(n5359), .ZN(n5738) );
  INV_X1 U7127 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U7128 ( .A1(n5733), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7129 ( .A1(n4523), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5650) );
  OAI211_X1 U7130 ( .C1(n5738), .C2(n9064), .A(n5651), .B(n5650), .ZN(n5652)
         );
  INV_X1 U7131 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7132 ( .A1(n5654), .A2(n5653), .ZN(n8908) );
  XNOR2_X1 U7133 ( .A(n5656), .B(n5657), .ZN(n7991) );
  NAND2_X1 U7134 ( .A1(n7991), .A2(n5730), .ZN(n5659) );
  OR2_X1 U7135 ( .A1(n5319), .A2(n7994), .ZN(n5658) );
  INV_X1 U7136 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U7137 ( .A1(n5661), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7138 ( .A1(n5675), .A2(n5662), .ZN(n8912) );
  NAND2_X1 U7139 ( .A1(n8912), .A2(n4526), .ZN(n5667) );
  INV_X1 U7140 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U7141 ( .A1(n4523), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U7142 ( .A1(n5733), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5663) );
  OAI211_X1 U7143 ( .C1(n5738), .C2(n9061), .A(n5664), .B(n5663), .ZN(n5665)
         );
  INV_X1 U7144 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7145 ( .A1(n5667), .A2(n5666), .ZN(n8923) );
  NAND2_X1 U7146 ( .A1(n9118), .A2(n8560), .ZN(n5911) );
  INV_X1 U7147 ( .A(n8908), .ZN(n8933) );
  NAND2_X1 U7148 ( .A1(n9124), .A2(n8933), .ZN(n8913) );
  NAND2_X1 U7149 ( .A1(n8914), .A2(n5907), .ZN(n5668) );
  NAND2_X1 U7150 ( .A1(n5668), .A2(n5910), .ZN(n8900) );
  XNOR2_X1 U7151 ( .A(n5669), .B(n5670), .ZN(n8035) );
  NAND2_X1 U7152 ( .A1(n8035), .A2(n5730), .ZN(n5672) );
  OR2_X1 U7153 ( .A1(n5319), .A2(n8050), .ZN(n5671) );
  INV_X1 U7154 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7155 ( .A1(n5675), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7156 ( .A1(n5686), .A2(n5676), .ZN(n8899) );
  NAND2_X1 U7157 ( .A1(n8899), .A2(n4525), .ZN(n5681) );
  INV_X1 U7158 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U7159 ( .A1(n5734), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7160 ( .A1(n5733), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5677) );
  OAI211_X1 U7161 ( .C1(n9058), .C2(n5738), .A(n5678), .B(n5677), .ZN(n5679)
         );
  INV_X1 U7162 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7163 ( .A1(n8081), .A2(n5730), .ZN(n5685) );
  OR2_X1 U7164 ( .A1(n4527), .A2(n8096), .ZN(n5684) );
  INV_X1 U7165 ( .A(n8566), .ZN(n9106) );
  NAND2_X1 U7166 ( .A1(n5686), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7167 ( .A1(n5699), .A2(n5687), .ZN(n8890) );
  NAND2_X1 U7168 ( .A1(n8890), .A2(n4526), .ZN(n5692) );
  INV_X1 U7169 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U7170 ( .A1(n5733), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U7171 ( .A1(n5734), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5688) );
  OAI211_X1 U7172 ( .C1(n5738), .C2(n9055), .A(n5689), .B(n5688), .ZN(n5690)
         );
  INV_X1 U7173 ( .A(n5690), .ZN(n5691) );
  XNOR2_X1 U7174 ( .A(n5694), .B(n5693), .ZN(n6285) );
  NAND2_X1 U7175 ( .A1(n6285), .A2(n5730), .ZN(n5697) );
  OR2_X1 U7176 ( .A1(n4527), .A2(n5695), .ZN(n5696) );
  INV_X1 U7177 ( .A(n5699), .ZN(n5698) );
  INV_X1 U7178 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U7179 ( .A1(n5699), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7180 ( .A1(n5712), .A2(n5700), .ZN(n8875) );
  NAND2_X1 U7181 ( .A1(n8875), .A2(n4526), .ZN(n5705) );
  INV_X1 U7182 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U7183 ( .A1(n5734), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U7184 ( .A1(n5733), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5701) );
  OAI211_X1 U7185 ( .C1(n8530), .C2(n5738), .A(n5702), .B(n5701), .ZN(n5703)
         );
  INV_X1 U7186 ( .A(n5703), .ZN(n5704) );
  AND2_X2 U7187 ( .A1(n5705), .A2(n5704), .ZN(n8886) );
  INV_X2 U7188 ( .A(n8886), .ZN(n8728) );
  NAND2_X1 U7189 ( .A1(n8137), .A2(n5730), .ZN(n5711) );
  OR2_X1 U7190 ( .A1(n4527), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U7191 ( .A1(n5712), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7192 ( .A1(n8850), .A2(n5713), .ZN(n8869) );
  NAND2_X1 U7193 ( .A1(n8869), .A2(n4526), .ZN(n5718) );
  INV_X1 U7194 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U7195 ( .A1(n5734), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7196 ( .A1(n5733), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U7197 ( .C1(n5738), .C2(n9053), .A(n5715), .B(n5714), .ZN(n5716)
         );
  INV_X1 U7198 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7199 ( .A1(n9163), .A2(n5730), .ZN(n5721) );
  OR2_X1 U7200 ( .A1(n5319), .A2(n9166), .ZN(n5720) );
  INV_X1 U7201 ( .A(n8850), .ZN(n5722) );
  NAND2_X1 U7202 ( .A1(n5722), .A2(n4525), .ZN(n5745) );
  INV_X1 U7203 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U7204 ( .A1(n5734), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7205 ( .A1(n5733), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5723) );
  OAI211_X1 U7206 ( .C1(n6895), .C2(n5738), .A(n5724), .B(n5723), .ZN(n5725)
         );
  INV_X1 U7207 ( .A(n5725), .ZN(n5726) );
  INV_X1 U7208 ( .A(n5917), .ZN(n5727) );
  NAND2_X1 U7209 ( .A1(n8532), .A2(n5730), .ZN(n5732) );
  OR2_X1 U7210 ( .A1(n4527), .A2(n8578), .ZN(n5731) );
  INV_X1 U7211 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7212 ( .A1(n5733), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7213 ( .A1(n5734), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5735) );
  OAI211_X1 U7214 ( .C1(n5738), .C2(n5737), .A(n5736), .B(n5735), .ZN(n5739)
         );
  INV_X1 U7215 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U7216 ( .A1(n5745), .A2(n5740), .ZN(n8726) );
  INV_X1 U7217 ( .A(n8726), .ZN(n5746) );
  NAND2_X1 U7218 ( .A1(n9048), .A2(n5746), .ZN(n5933) );
  NAND2_X1 U7219 ( .A1(n5933), .A2(n5916), .ZN(n5929) );
  NAND2_X1 U7220 ( .A1(n5733), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7221 ( .A1(n4522), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7222 ( .A1(n5734), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5741) );
  AND3_X1 U7223 ( .A1(n5743), .A2(n5742), .A3(n5741), .ZN(n5744) );
  AND2_X1 U7224 ( .A1(n5745), .A2(n5744), .ZN(n5927) );
  OAI211_X1 U7225 ( .C1(n5747), .C2(n5929), .A(n8849), .B(n5932), .ZN(n5750)
         );
  NAND2_X1 U7226 ( .A1(n6804), .A2(n5916), .ZN(n5748) );
  AOI211_X1 U7227 ( .C1(n5748), .C2(n5917), .A(n8849), .B(n9048), .ZN(n5749)
         );
  AOI21_X1 U7228 ( .B1(n5926), .B2(n5750), .A(n5749), .ZN(n5940) );
  INV_X1 U7229 ( .A(n5751), .ZN(n5754) );
  INV_X1 U7230 ( .A(n5755), .ZN(n5781) );
  INV_X1 U7231 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7232 ( .A1(n6900), .A2(n7660), .ZN(n5776) );
  NOR3_X1 U7233 ( .A1(n5940), .A2(n7805), .A3(n5776), .ZN(n5779) );
  XNOR2_X1 U7234 ( .A(n9096), .B(n8849), .ZN(n5775) );
  NAND2_X1 U7235 ( .A1(n5932), .A2(n5917), .ZN(n5920) );
  NAND2_X1 U7236 ( .A1(n5910), .A2(n5911), .ZN(n8915) );
  INV_X1 U7237 ( .A(n8913), .ZN(n5759) );
  NAND2_X1 U7238 ( .A1(n5898), .A2(n5899), .ZN(n8938) );
  NAND2_X1 U7239 ( .A1(n8936), .A2(n5794), .ZN(n8948) );
  NAND2_X1 U7240 ( .A1(n5895), .A2(n8946), .ZN(n8961) );
  INV_X1 U7241 ( .A(n5880), .ZN(n5760) );
  AND2_X1 U7242 ( .A1(n5760), .A2(n5865), .ZN(n8006) );
  INV_X1 U7243 ( .A(n8006), .ZN(n8005) );
  AND2_X1 U7244 ( .A1(n5861), .A2(n5862), .ZN(n8071) );
  INV_X1 U7245 ( .A(n8071), .ZN(n8067) );
  NOR2_X1 U7246 ( .A1(n7930), .A2(n8731), .ZN(n5859) );
  OR2_X1 U7247 ( .A1(n5147), .A2(n5859), .ZN(n7971) );
  NAND2_X1 U7248 ( .A1(n5853), .A2(n5851), .ZN(n7817) );
  INV_X1 U7249 ( .A(n7817), .ZN(n5767) );
  NAND4_X1 U7250 ( .A1(n5761), .A2(n5325), .A3(n9042), .A4(n7374), .ZN(n5762)
         );
  INV_X1 U7251 ( .A(n7643), .ZN(n7649) );
  INV_X1 U7252 ( .A(n8583), .ZN(n7208) );
  NAND2_X1 U7253 ( .A1(n7208), .A2(n8739), .ZN(n5795) );
  NAND2_X1 U7254 ( .A1(n7114), .A2(n5795), .ZN(n8584) );
  NOR3_X1 U7255 ( .A1(n5762), .A2(n7649), .A3(n8584), .ZN(n5763) );
  XNOR2_X1 U7256 ( .A(n7394), .B(n6821), .ZN(n7426) );
  NAND3_X1 U7257 ( .A1(n5763), .A2(n10431), .A3(n7426), .ZN(n5765) );
  INV_X1 U7258 ( .A(n5846), .ZN(n5764) );
  OR2_X1 U7259 ( .A1(n5839), .A2(n5764), .ZN(n7778) );
  NAND2_X1 U7260 ( .A1(n5841), .A2(n5832), .ZN(n7700) );
  NOR4_X1 U7261 ( .A1(n5765), .A2(n7778), .A3(n7711), .A4(n7700), .ZN(n5766)
         );
  NAND4_X1 U7262 ( .A1(n7971), .A2(n7922), .A3(n5767), .A4(n5766), .ZN(n5768)
         );
  NOR4_X1 U7263 ( .A1(n9015), .A2(n8005), .A3(n8067), .A4(n5768), .ZN(n5769)
         );
  NAND4_X1 U7264 ( .A1(n8973), .A2(n6844), .A3(n5868), .A4(n5769), .ZN(n5770)
         );
  OR4_X1 U7265 ( .A1(n8938), .A2(n8948), .A3(n8961), .A4(n5770), .ZN(n5771) );
  NOR4_X1 U7266 ( .A1(n8901), .A2(n8915), .A3(n8922), .A4(n5771), .ZN(n5773)
         );
  INV_X1 U7267 ( .A(n5772), .ZN(n5787) );
  NAND4_X1 U7268 ( .A1(n5773), .A2(n8883), .A3(n5116), .A4(n8523), .ZN(n5774)
         );
  NOR4_X1 U7269 ( .A1(n5775), .A2(n5929), .A3(n5920), .A4(n5774), .ZN(n5942)
         );
  NOR3_X1 U7270 ( .A1(n5942), .A2(n5021), .A3(n5776), .ZN(n5778) );
  NAND2_X1 U7271 ( .A1(n5777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5948) );
  INV_X1 U7272 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5947) );
  XNOR2_X1 U7273 ( .A(n5948), .B(n5947), .ZN(n6693) );
  OR2_X1 U7274 ( .A1(n6693), .A2(P2_U3151), .ZN(n7894) );
  NOR3_X1 U7275 ( .A1(n5779), .A2(n5778), .A3(n7894), .ZN(n5946) );
  INV_X1 U7276 ( .A(n5905), .ZN(n5780) );
  AOI211_X1 U7277 ( .C1(n5787), .C2(n5912), .A(n5780), .B(n5123), .ZN(n5786)
         );
  NAND2_X1 U7278 ( .A1(n5706), .A2(n8886), .ZN(n5784) );
  NAND2_X1 U7279 ( .A1(n5781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5783) );
  XNOR2_X1 U7280 ( .A(n5783), .B(n5782), .ZN(n7878) );
  NOR2_X4 U7281 ( .A1(n7805), .A2(n7878), .ZN(n6884) );
  AOI21_X1 U7282 ( .B1(n5905), .B2(n5904), .A(n5914), .ZN(n5789) );
  NOR3_X1 U7283 ( .A1(n5789), .A2(n6884), .A3(n5788), .ZN(n5790) );
  OAI21_X1 U7284 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5915) );
  INV_X1 U7285 ( .A(n5794), .ZN(n5897) );
  NAND2_X1 U7286 ( .A1(n5795), .A2(n5021), .ZN(n5799) );
  NOR2_X1 U7287 ( .A1(n5799), .A2(n7878), .ZN(n5797) );
  INV_X1 U7288 ( .A(n5798), .ZN(n5803) );
  NAND3_X1 U7289 ( .A1(n5799), .A2(n7114), .A3(n5800), .ZN(n5801) );
  MUX2_X1 U7290 ( .A(n5801), .B(n5800), .S(n6884), .Z(n5802) );
  NAND3_X1 U7291 ( .A1(n5803), .A2(n5761), .A3(n5802), .ZN(n5810) );
  INV_X1 U7292 ( .A(n7168), .ZN(n10485) );
  NAND2_X1 U7293 ( .A1(n10485), .A2(n8738), .ZN(n5812) );
  NAND2_X1 U7294 ( .A1(n5812), .A2(n5804), .ZN(n5805) );
  NAND2_X1 U7295 ( .A1(n5805), .A2(n6884), .ZN(n5809) );
  NAND2_X1 U7296 ( .A1(n5806), .A2(n5819), .ZN(n5807) );
  NAND3_X1 U7297 ( .A1(n5810), .A2(n5809), .A3(n5808), .ZN(n5811) );
  NAND2_X1 U7298 ( .A1(n5811), .A2(n7374), .ZN(n5823) );
  INV_X1 U7299 ( .A(n5812), .ZN(n5815) );
  INV_X1 U7300 ( .A(n5813), .ZN(n5824) );
  OAI211_X1 U7301 ( .C1(n5823), .C2(n5815), .A(n5824), .B(n5814), .ZN(n5818)
         );
  AND2_X1 U7302 ( .A1(n5826), .A2(n5821), .ZN(n5817) );
  INV_X1 U7303 ( .A(n5828), .ZN(n5816) );
  AOI21_X1 U7304 ( .B1(n5818), .B2(n5817), .A(n5816), .ZN(n5831) );
  INV_X1 U7305 ( .A(n5819), .ZN(n5822) );
  NAND2_X1 U7306 ( .A1(n10489), .A2(n10428), .ZN(n5820) );
  OAI211_X1 U7307 ( .C1(n5823), .C2(n5822), .A(n5821), .B(n5820), .ZN(n5825)
         );
  NAND2_X1 U7308 ( .A1(n5825), .A2(n5824), .ZN(n5827) );
  NAND2_X1 U7309 ( .A1(n5827), .A2(n5826), .ZN(n5829) );
  NAND2_X1 U7310 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  MUX2_X1 U7311 ( .A(n5831), .B(n5830), .S(n6884), .Z(n5835) );
  NAND2_X1 U7312 ( .A1(n5840), .A2(n5841), .ZN(n5833) );
  INV_X1 U7313 ( .A(n5838), .ZN(n5834) );
  NAND3_X1 U7314 ( .A1(n5835), .A2(n5834), .A3(n7643), .ZN(n5845) );
  AND2_X1 U7315 ( .A1(n5841), .A2(n5836), .ZN(n5837) );
  OAI211_X1 U7316 ( .C1(n5838), .C2(n5837), .A(n5846), .B(n5840), .ZN(n5844)
         );
  NAND3_X1 U7317 ( .A1(n4578), .A2(n5841), .A3(n5840), .ZN(n5842) );
  AND2_X1 U7318 ( .A1(n5851), .A2(n5846), .ZN(n5848) );
  INV_X1 U7319 ( .A(n5853), .ZN(n5847) );
  NAND2_X1 U7320 ( .A1(n5850), .A2(n5849), .ZN(n5852) );
  MUX2_X1 U7321 ( .A(n5856), .B(n5855), .S(n5873), .Z(n5857) );
  INV_X1 U7322 ( .A(n5859), .ZN(n6836) );
  INV_X1 U7323 ( .A(n7930), .ZN(n8000) );
  MUX2_X1 U7324 ( .A(n7931), .B(n8000), .S(n6884), .Z(n5860) );
  MUX2_X1 U7325 ( .A(n5862), .B(n5861), .S(n6884), .Z(n5863) );
  NAND2_X1 U7326 ( .A1(n5864), .A2(n8006), .ZN(n5878) );
  AND2_X1 U7327 ( .A1(n5879), .A2(n5865), .ZN(n5866) );
  NAND2_X1 U7328 ( .A1(n5878), .A2(n5866), .ZN(n5867) );
  NAND2_X1 U7329 ( .A1(n5867), .A2(n5871), .ZN(n5869) );
  INV_X1 U7330 ( .A(n5871), .ZN(n5872) );
  NOR2_X1 U7331 ( .A1(n9001), .A2(n5872), .ZN(n5874) );
  INV_X1 U7332 ( .A(n5876), .ZN(n5877) );
  INV_X1 U7333 ( .A(n5878), .ZN(n5881) );
  OAI211_X1 U7334 ( .C1(n5881), .C2(n5880), .A(n5873), .B(n5879), .ZN(n5885)
         );
  INV_X1 U7335 ( .A(n5883), .ZN(n5884) );
  AOI211_X1 U7336 ( .C1(n5886), .C2(n5885), .A(n5080), .B(n5884), .ZN(n5888)
         );
  INV_X1 U7337 ( .A(n5891), .ZN(n5887) );
  INV_X1 U7338 ( .A(n8961), .ZN(n8958) );
  NAND2_X1 U7339 ( .A1(n8958), .A2(n5890), .ZN(n5893) );
  NAND2_X1 U7340 ( .A1(n8946), .A2(n5891), .ZN(n5892) );
  MUX2_X1 U7341 ( .A(n5893), .B(n5892), .S(n6884), .Z(n5894) );
  AOI21_X1 U7342 ( .B1(n8936), .B2(n5895), .A(n5873), .ZN(n5896) );
  INV_X1 U7343 ( .A(n5898), .ZN(n5901) );
  NAND2_X1 U7344 ( .A1(n8913), .A2(n5899), .ZN(n5900) );
  MUX2_X1 U7345 ( .A(n5901), .B(n5900), .S(n5873), .Z(n5902) );
  INV_X1 U7346 ( .A(n5903), .ZN(n5909) );
  NAND4_X1 U7347 ( .A1(n5905), .A2(n6884), .A3(n5904), .A4(n5910), .ZN(n5906)
         );
  INV_X1 U7348 ( .A(n5911), .ZN(n5913) );
  INV_X1 U7349 ( .A(n6862), .ZN(n5918) );
  INV_X1 U7350 ( .A(n8602), .ZN(n8727) );
  MUX2_X1 U7351 ( .A(n8727), .B(n8574), .S(n5873), .Z(n5922) );
  NAND2_X1 U7352 ( .A1(n5921), .A2(n5919), .ZN(n5928) );
  INV_X1 U7353 ( .A(n5928), .ZN(n5924) );
  NOR2_X1 U7354 ( .A1(n5920), .A2(n5873), .ZN(n5923) );
  OAI211_X1 U7355 ( .C1(n5924), .C2(n8574), .A(n5923), .B(n5931), .ZN(n5925)
         );
  OAI21_X1 U7356 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5937) );
  INV_X1 U7357 ( .A(n5932), .ZN(n5934) );
  OR2_X1 U7358 ( .A1(n6900), .A2(n7660), .ZN(n6906) );
  INV_X1 U7359 ( .A(n6906), .ZN(n5938) );
  NOR2_X1 U7360 ( .A1(n7660), .A2(n7722), .ZN(n5941) );
  NAND3_X1 U7361 ( .A1(n5940), .A2(n5021), .A3(n5941), .ZN(n5944) );
  NAND3_X1 U7362 ( .A1(n5942), .A2(n5941), .A3(n7805), .ZN(n5943) );
  INV_X1 U7363 ( .A(n7878), .ZN(n6887) );
  NAND2_X1 U7364 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  INV_X1 U7365 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5956) );
  INV_X1 U7366 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5950) );
  INV_X1 U7367 ( .A(n6885), .ZN(n5961) );
  NAND2_X1 U7368 ( .A1(n5952), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  MUX2_X1 U7369 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5953), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5955) );
  AND2_X1 U7370 ( .A1(n5955), .A2(n5954), .ZN(n6871) );
  NOR2_X1 U7371 ( .A1(n8099), .A2(n7996), .ZN(n5960) );
  NAND2_X1 U7372 ( .A1(n5961), .A2(n5960), .ZN(n7081) );
  AND2_X1 U7373 ( .A1(n6693), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6979) );
  AND2_X1 U7374 ( .A1(n7660), .A2(n6887), .ZN(n6805) );
  NAND2_X1 U7375 ( .A1(n7377), .A2(n6805), .ZN(n7093) );
  INV_X1 U7376 ( .A(n7093), .ZN(n7200) );
  AND2_X1 U7377 ( .A1(n7097), .A2(n7200), .ZN(n7088) );
  INV_X1 U7378 ( .A(n5962), .ZN(n6865) );
  NAND3_X1 U7379 ( .A1(n7088), .A2(n6865), .A3(n6773), .ZN(n5964) );
  OAI211_X1 U7380 ( .C1(n6887), .C2(n7894), .A(n5964), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5965) );
  INV_X1 U7381 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5969) );
  INV_X1 U7382 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5970) );
  INV_X1 U7383 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7384 ( .A1(n5970), .A2(n6405), .ZN(n5974) );
  AND2_X1 U7385 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5971) );
  NOR2_X1 U7386 ( .A1(n5991), .A2(n5971), .ZN(n5973) );
  OR2_X1 U7387 ( .A1(n5973), .A2(n5972), .ZN(n5981) );
  INV_X1 U7388 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5989) );
  INV_X1 U7389 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7390 ( .A1(n5989), .A2(n5975), .ZN(n5976) );
  INV_X1 U7391 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5982) );
  INV_X1 U7392 ( .A(n9756), .ZN(n5986) );
  NAND2_X1 U7393 ( .A1(n8163), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5987) );
  INV_X1 U7394 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7395 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5992) );
  NAND2_X1 U7396 ( .A1(n6008), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7397 ( .A1(n8163), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6333) );
  INV_X1 U7398 ( .A(SI_0_), .ZN(n5994) );
  NOR2_X1 U7399 ( .A1(n8151), .A2(n5994), .ZN(n5996) );
  INV_X1 U7400 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5995) );
  XNOR2_X1 U7401 ( .A(n5996), .B(n5995), .ZN(n9759) );
  MUX2_X1 U7402 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9759), .S(n6045), .Z(n6440) );
  NAND2_X1 U7403 ( .A1(n10265), .A2(n6440), .ZN(n10266) );
  NAND2_X1 U7404 ( .A1(n6171), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7405 ( .A1(n6008), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7406 ( .A1(n8163), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7407 ( .A1(n8162), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5998) );
  INV_X1 U7408 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6915) );
  OR2_X1 U7409 ( .A1(n6013), .A2(n6915), .ZN(n6006) );
  OR2_X1 U7410 ( .A1(n6071), .A2(n6948), .ZN(n6005) );
  INV_X1 U7411 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7412 ( .A1(n6029), .A2(n6003), .ZN(n6014) );
  OR2_X1 U7413 ( .A1(n6045), .A2(n7043), .ZN(n6004) );
  NAND2_X1 U7414 ( .A1(n9308), .A2(n10298), .ZN(n8445) );
  NAND2_X1 U7415 ( .A1(n6171), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6012) );
  INV_X1 U7416 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U7417 ( .A1(n6008), .A2(n7177), .ZN(n6011) );
  NAND2_X1 U7418 ( .A1(n8163), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7419 ( .A1(n8162), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6009) );
  NAND4_X1 U7420 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n9307)
         );
  OR2_X1 U7421 ( .A1(n6071), .A2(n6928), .ZN(n6018) );
  NAND2_X1 U7422 ( .A1(n6014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  INV_X1 U7423 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6015) );
  OR2_X1 U7424 ( .A1(n6045), .A2(n8224), .ZN(n6017) );
  INV_X1 U7425 ( .A(n8444), .ZN(n8231) );
  AND2_X1 U7426 ( .A1(n9307), .A2(n7609), .ZN(n8228) );
  INV_X1 U7427 ( .A(n8228), .ZN(n8250) );
  NAND2_X1 U7428 ( .A1(n8231), .A2(n8250), .ZN(n8360) );
  INV_X1 U7429 ( .A(n8360), .ZN(n7607) );
  NAND2_X1 U7430 ( .A1(n7606), .A2(n8231), .ZN(n10232) );
  INV_X2 U7431 ( .A(n6171), .ZN(n6193) );
  INV_X1 U7432 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6020) );
  INV_X1 U7433 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6019) );
  OAI22_X1 U7434 ( .A1(n6193), .A2(n6020), .B1(n6305), .B2(n6019), .ZN(n6026)
         );
  INV_X2 U7435 ( .A(n6008), .ZN(n6062) );
  INV_X1 U7436 ( .A(n6037), .ZN(n6023) );
  INV_X1 U7437 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7438 ( .A1(n7177), .A2(n6021), .ZN(n6022) );
  NAND2_X1 U7439 ( .A1(n6023), .A2(n6022), .ZN(n9242) );
  INV_X2 U7440 ( .A(n8162), .ZN(n6194) );
  INV_X1 U7441 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6024) );
  OAI22_X1 U7442 ( .A1(n6062), .A2(n9242), .B1(n6194), .B2(n6024), .ZN(n6025)
         );
  OR2_X1 U7443 ( .A1(n6013), .A2(n4668), .ZN(n6035) );
  OR2_X1 U7444 ( .A1(n6071), .A2(n6927), .ZN(n6034) );
  OR2_X1 U7445 ( .A1(n6027), .A2(n6103), .ZN(n6028) );
  AND2_X1 U7446 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  INV_X1 U7447 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U7448 ( .A1(n6030), .A2(n9858), .ZN(n6040) );
  INV_X1 U7449 ( .A(n6030), .ZN(n6031) );
  NAND2_X1 U7450 ( .A1(n6031), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6032) );
  INV_X1 U7451 ( .A(n7013), .ZN(n7055) );
  OR2_X1 U7452 ( .A1(n6045), .A2(n7055), .ZN(n6033) );
  NAND2_X1 U7453 ( .A1(n9306), .A2(n10311), .ZN(n8249) );
  NAND2_X1 U7454 ( .A1(n10232), .A2(n8249), .ZN(n7504) );
  INV_X1 U7455 ( .A(n10311), .ZN(n10236) );
  NAND2_X1 U7456 ( .A1(n6470), .A2(n10236), .ZN(n8230) );
  INV_X1 U7457 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7007) );
  INV_X1 U7458 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6036) );
  OAI22_X1 U7459 ( .A1(n6193), .A2(n7007), .B1(n6305), .B2(n6036), .ZN(n6039)
         );
  NAND2_X1 U7460 ( .A1(n6037), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6075) );
  OAI21_X1 U7461 ( .B1(n6037), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6075), .ZN(
        n7508) );
  INV_X1 U7462 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7509) );
  OAI22_X1 U7463 ( .A1(n6062), .A2(n7508), .B1(n6194), .B2(n7509), .ZN(n6038)
         );
  INV_X1 U7464 ( .A(n10323), .ZN(n8237) );
  NAND2_X1 U7465 ( .A1(n6040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6041) );
  XNOR2_X1 U7466 ( .A(n6041), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7006) );
  INV_X1 U7467 ( .A(n7006), .ZN(n9326) );
  INV_X1 U7468 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6917) );
  OR2_X1 U7469 ( .A1(n6013), .A2(n6917), .ZN(n6043) );
  OR2_X1 U7470 ( .A1(n6071), .A2(n6931), .ZN(n6042) );
  OAI211_X1 U7471 ( .C1(n6045), .C2(n9326), .A(n6043), .B(n6042), .ZN(n8236)
         );
  NAND2_X1 U7472 ( .A1(n8237), .A2(n8236), .ZN(n6343) );
  NAND2_X1 U7473 ( .A1(n7504), .A2(n4569), .ZN(n6044) );
  AND2_X1 U7474 ( .A1(n10323), .A2(n10318), .ZN(n8225) );
  INV_X1 U7475 ( .A(n8225), .ZN(n8450) );
  INV_X2 U7476 ( .A(n6071), .ZN(n8156) );
  NAND2_X1 U7477 ( .A1(n6950), .A2(n8156), .ZN(n6051) );
  OAI21_X1 U7478 ( .B1(n6047), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6048) );
  INV_X1 U7479 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7480 ( .A1(n6048), .A2(n6099), .ZN(n6082) );
  OR2_X1 U7481 ( .A1(n6048), .A2(n6099), .ZN(n6049) );
  AND2_X1 U7482 ( .A1(n6082), .A2(n6049), .ZN(n7216) );
  AOI22_X1 U7483 ( .A1(n6224), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6920), .B2(
        n7216), .ZN(n6050) );
  NAND2_X1 U7484 ( .A1(n6051), .A2(n6050), .ZN(n10223) );
  INV_X1 U7485 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7139) );
  INV_X1 U7486 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6052) );
  OAI22_X1 U7487 ( .A1(n6193), .A2(n7139), .B1(n6194), .B2(n6052), .ZN(n6057)
         );
  NAND2_X1 U7488 ( .A1(n6076), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6064) );
  INV_X1 U7489 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7490 ( .A1(n6064), .A2(n6053), .ZN(n6054) );
  NAND2_X1 U7491 ( .A1(n6088), .A2(n6054), .ZN(n10221) );
  INV_X1 U7492 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6055) );
  OAI22_X1 U7493 ( .A1(n6062), .A2(n10221), .B1(n6305), .B2(n6055), .ZN(n6056)
         );
  INV_X1 U7494 ( .A(n10341), .ZN(n7856) );
  NAND2_X1 U7495 ( .A1(n10223), .A2(n7856), .ZN(n8258) );
  OR2_X1 U7496 ( .A1(n6926), .A2(n6071), .ZN(n6060) );
  NAND2_X1 U7497 ( .A1(n6047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6058) );
  XNOR2_X1 U7498 ( .A(n6058), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7127) );
  AOI22_X1 U7499 ( .A1(n6224), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6920), .B2(
        n7127), .ZN(n6059) );
  INV_X1 U7500 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7137) );
  INV_X1 U7501 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6061) );
  OAI22_X1 U7502 ( .A1(n6193), .A2(n7137), .B1(n6194), .B2(n6061), .ZN(n6067)
         );
  OR2_X1 U7503 ( .A1(n6076), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7504 ( .A1(n6064), .A2(n6063), .ZN(n7496) );
  INV_X1 U7505 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6065) );
  OAI22_X1 U7506 ( .A1(n6062), .A2(n7496), .B1(n6305), .B2(n6065), .ZN(n6066)
         );
  INV_X1 U7507 ( .A(n10322), .ZN(n7755) );
  NAND2_X1 U7508 ( .A1(n7497), .A2(n7755), .ZN(n7633) );
  NAND2_X1 U7509 ( .A1(n8258), .A2(n7633), .ZN(n8369) );
  INV_X1 U7510 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7511 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U7512 ( .A(n6070), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9344) );
  AOI22_X1 U7513 ( .A1(n6224), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6920), .B2(
        n9344), .ZN(n6073) );
  OR2_X1 U7514 ( .A1(n6934), .A2(n6071), .ZN(n6072) );
  INV_X1 U7515 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7005) );
  INV_X1 U7516 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7523) );
  OAI22_X1 U7517 ( .A1(n6193), .A2(n7005), .B1(n6194), .B2(n7523), .ZN(n6080)
         );
  AND2_X1 U7518 ( .A1(n6075), .A2(n6074), .ZN(n6077) );
  OR2_X1 U7519 ( .A1(n6077), .A2(n6076), .ZN(n7522) );
  INV_X1 U7520 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6078) );
  OAI22_X1 U7521 ( .A1(n6062), .A2(n7522), .B1(n6305), .B2(n6078), .ZN(n6079)
         );
  NOR2_X1 U7522 ( .A1(n8369), .A2(n8449), .ZN(n6081) );
  NAND2_X1 U7523 ( .A1(n7517), .A2(n6081), .ZN(n6098) );
  NAND2_X1 U7524 ( .A1(n6955), .A2(n8156), .ZN(n6085) );
  NAND2_X1 U7525 ( .A1(n6082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7526 ( .A(n6083), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7339) );
  AOI22_X1 U7527 ( .A1(n6224), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6920), .B2(
        n7339), .ZN(n6084) );
  INV_X1 U7528 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6086) );
  INV_X1 U7529 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7629) );
  OAI22_X1 U7530 ( .A1(n6193), .A2(n6086), .B1(n6194), .B2(n7629), .ZN(n6092)
         );
  INV_X1 U7531 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6087) );
  AND2_X1 U7532 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  OR2_X1 U7533 ( .A1(n6089), .A2(n6111), .ZN(n7855) );
  INV_X1 U7534 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6090) );
  OAI22_X1 U7535 ( .A1(n6062), .A2(n7855), .B1(n6305), .B2(n6090), .ZN(n6091)
         );
  INV_X1 U7536 ( .A(n10349), .ZN(n7811) );
  OR2_X1 U7537 ( .A1(n10223), .A2(n7856), .ZN(n7637) );
  INV_X1 U7538 ( .A(n8257), .ZN(n6094) );
  INV_X1 U7539 ( .A(n8369), .ZN(n6093) );
  NAND2_X1 U7540 ( .A1(n10332), .A2(n10322), .ZN(n6347) );
  NAND2_X1 U7541 ( .A1(n7637), .A2(n6347), .ZN(n8256) );
  INV_X1 U7542 ( .A(n8256), .ZN(n6096) );
  AND2_X1 U7543 ( .A1(n10326), .A2(n9305), .ZN(n8226) );
  INV_X1 U7544 ( .A(n8226), .ZN(n6095) );
  AND3_X1 U7545 ( .A1(n8261), .A2(n6096), .A3(n6095), .ZN(n8372) );
  INV_X1 U7546 ( .A(n8372), .ZN(n8454) );
  NAND2_X1 U7547 ( .A1(n8452), .A2(n8454), .ZN(n6097) );
  NAND2_X1 U7548 ( .A1(n6098), .A2(n6097), .ZN(n7474) );
  NAND2_X1 U7549 ( .A1(n10342), .A2(n7811), .ZN(n8453) );
  NAND2_X1 U7550 ( .A1(n7474), .A2(n8453), .ZN(n6116) );
  OR2_X1 U7551 ( .A1(n6958), .A2(n6071), .ZN(n6109) );
  INV_X1 U7552 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6100) );
  INV_X1 U7553 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9966) );
  NAND3_X1 U7554 ( .A1(n6100), .A2(n9966), .A3(n6099), .ZN(n6101) );
  NOR2_X1 U7555 ( .A1(n6047), .A2(n6101), .ZN(n6105) );
  NOR2_X1 U7556 ( .A1(n6105), .A2(n6103), .ZN(n6102) );
  MUX2_X1 U7557 ( .A(n6103), .B(n6102), .S(P1_IR_REG_10__SCAN_IN), .Z(n6107)
         );
  INV_X1 U7558 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7559 ( .A1(n6105), .A2(n6104), .ZN(n6126) );
  INV_X1 U7560 ( .A(n6126), .ZN(n6106) );
  NOR2_X1 U7561 ( .A1(n6107), .A2(n6106), .ZN(n7433) );
  AOI22_X1 U7562 ( .A1(n6224), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6920), .B2(
        n7433), .ZN(n6108) );
  INV_X1 U7563 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7438) );
  INV_X1 U7564 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6110) );
  OAI22_X1 U7565 ( .A1(n6193), .A2(n7438), .B1(n6194), .B2(n6110), .ZN(n6115)
         );
  NOR2_X1 U7566 ( .A1(n6111), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6112) );
  OR2_X1 U7567 ( .A1(n6121), .A2(n6112), .ZN(n7810) );
  INV_X1 U7568 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6113) );
  OAI22_X1 U7569 ( .A1(n6062), .A2(n7810), .B1(n6305), .B2(n6113), .ZN(n6114)
         );
  AND2_X1 U7570 ( .A1(n10352), .A2(n9304), .ZN(n8271) );
  INV_X1 U7571 ( .A(n8271), .ZN(n8457) );
  INV_X1 U7572 ( .A(n9304), .ZN(n10359) );
  NAND2_X1 U7573 ( .A1(n7484), .A2(n10359), .ZN(n8273) );
  AND2_X1 U7574 ( .A1(n8457), .A2(n8273), .ZN(n6351) );
  NAND2_X1 U7575 ( .A1(n6963), .A2(n8156), .ZN(n6119) );
  NAND2_X1 U7576 ( .A1(n6126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6117) );
  XNOR2_X1 U7577 ( .A(n6117), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8187) );
  AOI22_X1 U7578 ( .A1(n6224), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6920), .B2(
        n8187), .ZN(n6118) );
  INV_X1 U7579 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7440) );
  INV_X1 U7580 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6120) );
  OAI22_X1 U7581 ( .A1(n6193), .A2(n7440), .B1(n6305), .B2(n6120), .ZN(n6124)
         );
  NAND2_X1 U7582 ( .A1(n6121), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7583 ( .A1(n6121), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7584 ( .A1(n6135), .A2(n6122), .ZN(n7882) );
  INV_X1 U7585 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7590) );
  OAI22_X1 U7586 ( .A1(n6062), .A2(n7882), .B1(n6194), .B2(n7590), .ZN(n6123)
         );
  AND2_X1 U7587 ( .A1(n7887), .A2(n10373), .ZN(n8275) );
  INV_X1 U7588 ( .A(n8275), .ZN(n8373) );
  INV_X1 U7589 ( .A(n7887), .ZN(n10362) );
  INV_X1 U7590 ( .A(n10373), .ZN(n7952) );
  NAND2_X1 U7591 ( .A1(n10362), .A2(n7952), .ZN(n8274) );
  NAND2_X1 U7592 ( .A1(n8373), .A2(n8274), .ZN(n7595) );
  INV_X1 U7593 ( .A(n8273), .ZN(n7596) );
  NOR2_X1 U7594 ( .A1(n7595), .A2(n7596), .ZN(n6125) );
  OR2_X1 U7595 ( .A1(n6126), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7596 ( .A1(n6127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  INV_X1 U7597 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7598 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7599 ( .A1(n6129), .A2(n6128), .ZN(n6140) );
  AND2_X1 U7600 ( .A1(n6130), .A2(n6140), .ZN(n8188) );
  AOI22_X1 U7601 ( .A1(n6224), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6920), .B2(
        n8188), .ZN(n6131) );
  INV_X1 U7602 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8175) );
  INV_X1 U7603 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6133) );
  OAI22_X1 U7604 ( .A1(n6193), .A2(n8175), .B1(n6305), .B2(n6133), .ZN(n6138)
         );
  INV_X1 U7605 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7606 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7607 ( .A1(n6144), .A2(n6136), .ZN(n7951) );
  INV_X1 U7608 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7688) );
  OAI22_X1 U7609 ( .A1(n6062), .A2(n7951), .B1(n6194), .B2(n7688), .ZN(n6137)
         );
  OR2_X1 U7610 ( .A1(n6138), .A2(n6137), .ZN(n9303) );
  INV_X1 U7611 ( .A(n9303), .ZN(n10357) );
  NOR2_X1 U7612 ( .A1(n7944), .A2(n10357), .ZN(n8276) );
  INV_X1 U7613 ( .A(n8276), .ZN(n6139) );
  NAND2_X1 U7614 ( .A1(n7944), .A2(n10357), .ZN(n8460) );
  NAND2_X1 U7615 ( .A1(n7684), .A2(n8460), .ZN(n7723) );
  INV_X1 U7616 ( .A(n7723), .ZN(n6150) );
  NAND2_X1 U7617 ( .A1(n6140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7618 ( .A(n6141), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8189) );
  AOI22_X1 U7619 ( .A1(n6224), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6920), .B2(
        n8189), .ZN(n6142) );
  INV_X1 U7620 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8172) );
  INV_X1 U7621 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7729) );
  OAI22_X1 U7622 ( .A1(n6193), .A2(n8172), .B1(n6194), .B2(n7729), .ZN(n6148)
         );
  INV_X1 U7623 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U7624 ( .A1(n6144), .A2(n9352), .ZN(n6145) );
  NAND2_X1 U7625 ( .A1(n6160), .A2(n6145), .ZN(n8041) );
  INV_X1 U7626 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6146) );
  OAI22_X1 U7627 ( .A1(n6062), .A2(n8041), .B1(n6305), .B2(n6146), .ZN(n6147)
         );
  OR2_X1 U7628 ( .A1(n6148), .A2(n6147), .ZN(n10372) );
  AND2_X1 U7629 ( .A1(n10383), .A2(n10372), .ZN(n8278) );
  INV_X1 U7630 ( .A(n10383), .ZN(n8048) );
  AND2_X1 U7631 ( .A1(n8048), .A2(n8104), .ZN(n8463) );
  INV_X1 U7632 ( .A(n8463), .ZN(n8267) );
  NAND2_X1 U7633 ( .A1(n7171), .A2(n8156), .ZN(n6157) );
  NOR2_X1 U7634 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6151) );
  NAND2_X1 U7635 ( .A1(n6068), .A2(n5144), .ZN(n6166) );
  NAND2_X1 U7636 ( .A1(n6166), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6155) );
  XNOR2_X1 U7637 ( .A(n6155), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9372) );
  AOI22_X1 U7638 ( .A1(n6224), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6920), .B2(
        n9372), .ZN(n6156) );
  INV_X1 U7639 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8177) );
  INV_X1 U7640 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6158) );
  OAI22_X1 U7641 ( .A1(n6193), .A2(n8177), .B1(n6194), .B2(n6158), .ZN(n6164)
         );
  INV_X1 U7642 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6159) );
  AND2_X1 U7643 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  OR2_X1 U7644 ( .A1(n6161), .A2(n6172), .ZN(n10208) );
  INV_X1 U7645 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6162) );
  OAI22_X1 U7646 ( .A1(n6062), .A2(n10208), .B1(n6305), .B2(n6162), .ZN(n6163)
         );
  OR2_X1 U7647 ( .A1(n6164), .A2(n6163), .ZN(n9302) );
  INV_X1 U7648 ( .A(n9302), .ZN(n6541) );
  OR2_X1 U7649 ( .A1(n10210), .A2(n6541), .ZN(n8281) );
  NAND2_X1 U7650 ( .A1(n10210), .A2(n6541), .ZN(n8466) );
  NAND2_X1 U7651 ( .A1(n8281), .A2(n8466), .ZN(n10202) );
  NAND2_X1 U7652 ( .A1(n10205), .A2(n8466), .ZN(n7900) );
  NAND2_X1 U7653 ( .A1(n7277), .A2(n8156), .ZN(n6170) );
  NAND2_X1 U7654 ( .A1(n6205), .A2(n6167), .ZN(n6178) );
  OR2_X1 U7655 ( .A1(n6205), .A2(n6167), .ZN(n6168) );
  AND2_X1 U7656 ( .A1(n6178), .A2(n6168), .ZN(n9382) );
  AOI22_X1 U7657 ( .A1(n6224), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6920), .B2(
        n9382), .ZN(n6169) );
  NAND2_X1 U7658 ( .A1(n6171), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6177) );
  OR2_X1 U7659 ( .A1(n6172), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7660 ( .A1(n6172), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6183) );
  AND2_X1 U7661 ( .A1(n6173), .A2(n6183), .ZN(n8089) );
  NAND2_X1 U7662 ( .A1(n6008), .A2(n8089), .ZN(n6176) );
  NAND2_X1 U7663 ( .A1(n8163), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7664 ( .A1(n8162), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6174) );
  NAND4_X1 U7665 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n9301)
         );
  INV_X1 U7666 ( .A(n9301), .ZN(n9207) );
  NOR2_X1 U7667 ( .A1(n8284), .A2(n9207), .ZN(n8282) );
  INV_X1 U7668 ( .A(n8282), .ZN(n8470) );
  NAND2_X1 U7669 ( .A1(n8284), .A2(n9207), .ZN(n8467) );
  NAND2_X1 U7670 ( .A1(n8470), .A2(n8467), .ZN(n8378) );
  INV_X1 U7671 ( .A(n8378), .ZN(n7899) );
  NAND2_X1 U7672 ( .A1(n7900), .A2(n7899), .ZN(n7898) );
  NAND2_X1 U7673 ( .A1(n7898), .A2(n8467), .ZN(n7956) );
  NAND2_X1 U7674 ( .A1(n7348), .A2(n8156), .ZN(n6181) );
  NAND2_X1 U7675 ( .A1(n6178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7676 ( .A(n6179), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9417) );
  AOI22_X1 U7677 ( .A1(n6224), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6920), .B2(
        n9417), .ZN(n6180) );
  INV_X1 U7678 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9390) );
  INV_X1 U7679 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9392) );
  OAI22_X1 U7680 ( .A1(n6193), .A2(n9390), .B1(n6194), .B2(n9392), .ZN(n6188)
         );
  INV_X1 U7681 ( .A(n6183), .ZN(n6182) );
  INV_X1 U7682 ( .A(n6195), .ZN(n6197) );
  INV_X1 U7683 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7684 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U7685 ( .A1(n6197), .A2(n6185), .ZN(n9206) );
  INV_X1 U7686 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6186) );
  OAI22_X1 U7687 ( .A1(n6062), .A2(n9206), .B1(n6305), .B2(n6186), .ZN(n6187)
         );
  OR2_X1 U7688 ( .A1(n6188), .A2(n6187), .ZN(n9300) );
  INV_X1 U7689 ( .A(n8474), .ZN(n8285) );
  INV_X1 U7690 ( .A(n10196), .ZN(n7961) );
  INV_X1 U7691 ( .A(n9300), .ZN(n8092) );
  NAND2_X1 U7692 ( .A1(n8285), .A2(n8476), .ZN(n8381) );
  NAND2_X1 U7693 ( .A1(n7956), .A2(n7963), .ZN(n6189) );
  NAND2_X1 U7694 ( .A1(n6189), .A2(n8476), .ZN(n8017) );
  INV_X1 U7695 ( .A(n8017), .ZN(n6202) );
  NAND2_X1 U7696 ( .A1(n7400), .A2(n8156), .ZN(n6192) );
  OAI21_X1 U7697 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7698 ( .A1(n6205), .A2(n6203), .ZN(n6190) );
  INV_X1 U7699 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10097) );
  XNOR2_X1 U7700 ( .A(n6190), .B(n10097), .ZN(n9427) );
  AOI22_X1 U7701 ( .A1(n6224), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6920), .B2(
        n9427), .ZN(n6191) );
  INV_X1 U7702 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9405) );
  INV_X1 U7703 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8025) );
  OAI22_X1 U7704 ( .A1(n6193), .A2(n9405), .B1(n6194), .B2(n8025), .ZN(n6201)
         );
  INV_X1 U7705 ( .A(n6213), .ZN(n6215) );
  INV_X1 U7706 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7707 ( .A1(n6197), .A2(n6196), .ZN(n6198) );
  NAND2_X1 U7708 ( .A1(n6215), .A2(n6198), .ZN(n9220) );
  INV_X1 U7709 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6199) );
  OAI22_X1 U7710 ( .A1(n6062), .A2(n9220), .B1(n6305), .B2(n6199), .ZN(n6200)
         );
  OR2_X1 U7711 ( .A1(n6201), .A2(n6200), .ZN(n9299) );
  INV_X1 U7712 ( .A(n9299), .ZN(n9272) );
  OR2_X1 U7713 ( .A1(n9222), .A2(n9272), .ZN(n8472) );
  NAND2_X1 U7714 ( .A1(n9222), .A2(n9272), .ZN(n8477) );
  INV_X1 U7715 ( .A(n8384), .ZN(n8018) );
  NAND2_X1 U7716 ( .A1(n6202), .A2(n8384), .ZN(n8015) );
  NAND2_X1 U7717 ( .A1(n8015), .A2(n8472), .ZN(n8054) );
  INV_X1 U7718 ( .A(n8054), .ZN(n6221) );
  NAND2_X1 U7719 ( .A1(n7567), .A2(n8156), .ZN(n6212) );
  AND2_X1 U7720 ( .A1(n6203), .A2(n10097), .ZN(n6204) );
  NAND2_X1 U7721 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  INV_X1 U7722 ( .A(n6209), .ZN(n6207) );
  NAND2_X1 U7723 ( .A1(n6207), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6210) );
  INV_X1 U7724 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7725 ( .A1(n6209), .A2(n6208), .ZN(n6222) );
  AND2_X1 U7726 ( .A1(n6210), .A2(n6222), .ZN(n9455) );
  AOI22_X1 U7727 ( .A1(n6224), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6920), .B2(
        n9455), .ZN(n6211) );
  INV_X1 U7728 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9432) );
  INV_X1 U7729 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9441) );
  OAI22_X1 U7730 ( .A1(n6193), .A2(n9432), .B1(n6194), .B2(n9441), .ZN(n6220)
         );
  INV_X1 U7731 ( .A(n6228), .ZN(n6217) );
  INV_X1 U7732 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7733 ( .A1(n6215), .A2(n6214), .ZN(n6216) );
  NAND2_X1 U7734 ( .A1(n6217), .A2(n6216), .ZN(n9271) );
  INV_X1 U7735 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6218) );
  OAI22_X1 U7736 ( .A1(n6062), .A2(n9271), .B1(n6305), .B2(n6218), .ZN(n6219)
         );
  OR2_X1 U7737 ( .A1(n6220), .A2(n6219), .ZN(n9298) );
  INV_X1 U7738 ( .A(n9298), .ZN(n9181) );
  OR2_X1 U7739 ( .A1(n9275), .A2(n9181), .ZN(n8295) );
  NAND2_X1 U7740 ( .A1(n9275), .A2(n9181), .ZN(n8294) );
  NAND2_X1 U7741 ( .A1(n6221), .A2(n8383), .ZN(n8056) );
  NAND2_X1 U7742 ( .A1(n7656), .A2(n8156), .ZN(n6226) );
  NAND2_X1 U7743 ( .A1(n6222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6223) );
  AOI22_X1 U7744 ( .A1(n6224), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8434), .B2(
        n6920), .ZN(n6225) );
  INV_X1 U7745 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6227) );
  INV_X1 U7746 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8130) );
  OAI22_X1 U7747 ( .A1(n6193), .A2(n6227), .B1(n6194), .B2(n8130), .ZN(n6231)
         );
  OAI21_X1 U7748 ( .B1(n6228), .B2(P1_REG3_REG_19__SCAN_IN), .A(n6235), .ZN(
        n9180) );
  INV_X1 U7749 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6229) );
  OAI22_X1 U7750 ( .A1(n6062), .A2(n9180), .B1(n6305), .B2(n6229), .ZN(n6230)
         );
  OR2_X1 U7751 ( .A1(n6231), .A2(n6230), .ZN(n9297) );
  INV_X1 U7752 ( .A(n9297), .ZN(n9623) );
  OR2_X1 U7753 ( .A1(n8129), .A2(n9623), .ZN(n8296) );
  NAND2_X1 U7754 ( .A1(n8129), .A2(n9623), .ZN(n8484) );
  INV_X1 U7755 ( .A(n8296), .ZN(n6232) );
  NAND2_X1 U7756 ( .A1(n7707), .A2(n8156), .ZN(n6234) );
  INV_X1 U7757 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9835) );
  OR2_X1 U7758 ( .A1(n6013), .A2(n9835), .ZN(n6233) );
  INV_X1 U7759 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9252) );
  AOI21_X1 U7760 ( .B1(n6235), .B2(n9252), .A(n6241), .ZN(n9628) );
  INV_X1 U7761 ( .A(n9628), .ZN(n9253) );
  INV_X1 U7762 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6236) );
  OAI22_X1 U7763 ( .A1(n6062), .A2(n9253), .B1(n6194), .B2(n6236), .ZN(n6238)
         );
  INV_X1 U7764 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9704) );
  INV_X1 U7765 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9742) );
  OAI22_X1 U7766 ( .A1(n6193), .A2(n9704), .B1(n6305), .B2(n9742), .ZN(n6237)
         );
  OR2_X1 U7767 ( .A1(n6238), .A2(n6237), .ZN(n9693) );
  INV_X1 U7768 ( .A(n9693), .ZN(n9188) );
  OR2_X1 U7769 ( .A1(n9627), .A2(n9188), .ZN(n8305) );
  NAND2_X1 U7770 ( .A1(n9627), .A2(n9188), .ZN(n8304) );
  NAND2_X1 U7771 ( .A1(n8305), .A2(n8304), .ZN(n9620) );
  NAND2_X1 U7772 ( .A1(n7760), .A2(n8156), .ZN(n6240) );
  OR2_X1 U7773 ( .A1(n6013), .A2(n7761), .ZN(n6239) );
  NAND2_X2 U7774 ( .A1(n6240), .A2(n6239), .ZN(n9615) );
  INV_X1 U7775 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9699) );
  INV_X1 U7776 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9605) );
  OAI22_X1 U7777 ( .A1(n6193), .A2(n9699), .B1(n6194), .B2(n9605), .ZN(n6245)
         );
  INV_X1 U7778 ( .A(n6248), .ZN(n6249) );
  INV_X1 U7779 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9187) );
  INV_X1 U7780 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U7781 ( .A1(n9187), .A2(n6242), .ZN(n6243) );
  NAND2_X1 U7782 ( .A1(n6249), .A2(n6243), .ZN(n9604) );
  INV_X1 U7783 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9738) );
  OAI22_X1 U7784 ( .A1(n6062), .A2(n9604), .B1(n6305), .B2(n9738), .ZN(n6244)
         );
  OR2_X1 U7785 ( .A1(n6245), .A2(n6244), .ZN(n9684) );
  XNOR2_X1 U7786 ( .A(n9615), .B(n9684), .ZN(n9602) );
  NAND2_X1 U7787 ( .A1(n9599), .A2(n9602), .ZN(n9598) );
  INV_X1 U7788 ( .A(n9684), .ZN(n9624) );
  NAND2_X1 U7789 ( .A1(n9615), .A2(n9624), .ZN(n8307) );
  NAND2_X1 U7790 ( .A1(n9598), .A2(n8307), .ZN(n9583) );
  NAND2_X1 U7791 ( .A1(n7876), .A2(n8156), .ZN(n6247) );
  OR2_X1 U7792 ( .A1(n6013), .A2(n10072), .ZN(n6246) );
  INV_X1 U7793 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9690) );
  INV_X1 U7794 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9587) );
  OAI22_X1 U7795 ( .A1(n6193), .A2(n9690), .B1(n6194), .B2(n9587), .ZN(n6253)
         );
  INV_X1 U7796 ( .A(n6258), .ZN(n6251) );
  INV_X1 U7797 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U7798 ( .A1(n6249), .A2(n9262), .ZN(n6250) );
  NAND2_X1 U7799 ( .A1(n6251), .A2(n6250), .ZN(n9586) );
  INV_X1 U7800 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9735) );
  OAI22_X1 U7801 ( .A1(n6062), .A2(n9586), .B1(n6305), .B2(n9735), .ZN(n6252)
         );
  OR2_X1 U7802 ( .A1(n6253), .A2(n6252), .ZN(n9692) );
  INV_X1 U7803 ( .A(n9692), .ZN(n9610) );
  XNOR2_X1 U7804 ( .A(n9595), .B(n9610), .ZN(n9582) );
  INV_X1 U7805 ( .A(n9582), .ZN(n9585) );
  NAND2_X1 U7806 ( .A1(n9583), .A2(n9585), .ZN(n6254) );
  NAND2_X1 U7807 ( .A1(n9595), .A2(n9610), .ZN(n8315) );
  NAND2_X1 U7808 ( .A1(n6254), .A2(n8315), .ZN(n9566) );
  NAND2_X1 U7809 ( .A1(n7893), .A2(n8156), .ZN(n6256) );
  OR2_X1 U7810 ( .A1(n6013), .A2(n7891), .ZN(n6255) );
  INV_X1 U7811 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9681) );
  INV_X1 U7812 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6257) );
  OAI22_X1 U7813 ( .A1(n6193), .A2(n9681), .B1(n6194), .B2(n6257), .ZN(n6260)
         );
  NAND2_X1 U7814 ( .A1(n6258), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6266) );
  OAI21_X1 U7815 ( .B1(n6258), .B2(P1_REG3_REG_23__SCAN_IN), .A(n6266), .ZN(
        n9571) );
  INV_X1 U7816 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9731) );
  OAI22_X1 U7817 ( .A1(n6062), .A2(n9571), .B1(n6305), .B2(n9731), .ZN(n6259)
         );
  OR2_X1 U7818 ( .A1(n6260), .A2(n6259), .ZN(n9683) );
  INV_X1 U7819 ( .A(n9683), .ZN(n9590) );
  NAND2_X1 U7820 ( .A1(n9576), .A2(n9590), .ZN(n8397) );
  NAND2_X1 U7821 ( .A1(n9566), .A2(n9574), .ZN(n6261) );
  NAND2_X1 U7822 ( .A1(n7991), .A2(n8156), .ZN(n6263) );
  OR2_X1 U7823 ( .A1(n6013), .A2(n7992), .ZN(n6262) );
  INV_X1 U7824 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6265) );
  INV_X1 U7825 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6264) );
  OAI22_X1 U7826 ( .A1(n6193), .A2(n6265), .B1(n6194), .B2(n6264), .ZN(n6271)
         );
  INV_X1 U7827 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U7828 ( .A1(n6266), .A2(n9230), .ZN(n6268) );
  INV_X1 U7829 ( .A(n6274), .ZN(n6267) );
  NAND2_X1 U7830 ( .A1(n6268), .A2(n6267), .ZN(n9553) );
  INV_X1 U7831 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6269) );
  OAI22_X1 U7832 ( .A1(n6062), .A2(n9553), .B1(n6305), .B2(n6269), .ZN(n6270)
         );
  NAND2_X1 U7833 ( .A1(n6378), .A2(n9197), .ZN(n8406) );
  NAND2_X1 U7834 ( .A1(n8399), .A2(n8406), .ZN(n9557) );
  NAND2_X1 U7835 ( .A1(n8035), .A2(n8156), .ZN(n6273) );
  OR2_X1 U7836 ( .A1(n6013), .A2(n8037), .ZN(n6272) );
  INV_X1 U7837 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9670) );
  INV_X1 U7838 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9543) );
  OAI22_X1 U7839 ( .A1(n6193), .A2(n9670), .B1(n6194), .B2(n9543), .ZN(n6276)
         );
  INV_X1 U7840 ( .A(n6279), .ZN(n6281) );
  OAI21_X1 U7841 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6274), .A(n6281), .ZN(
        n9542) );
  INV_X1 U7842 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9726) );
  OAI22_X1 U7843 ( .A1(n6062), .A2(n9542), .B1(n6305), .B2(n9726), .ZN(n6275)
         );
  INV_X1 U7844 ( .A(n9728), .ZN(n9541) );
  INV_X1 U7845 ( .A(n8320), .ZN(n8410) );
  NAND2_X1 U7846 ( .A1(n8081), .A2(n8156), .ZN(n6278) );
  OR2_X1 U7847 ( .A1(n6013), .A2(n8083), .ZN(n6277) );
  INV_X1 U7848 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9665) );
  INV_X1 U7849 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9525) );
  OAI22_X1 U7850 ( .A1(n6193), .A2(n9665), .B1(n6194), .B2(n9525), .ZN(n6284)
         );
  NAND2_X1 U7851 ( .A1(n6279), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6290) );
  INV_X1 U7852 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7853 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U7854 ( .A1(n6290), .A2(n6282), .ZN(n9524) );
  INV_X1 U7855 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9722) );
  OAI22_X1 U7856 ( .A1(n6062), .A2(n9524), .B1(n6305), .B2(n9722), .ZN(n6283)
         );
  XNOR2_X1 U7857 ( .A(n9532), .B(n9649), .ZN(n9523) );
  INV_X1 U7858 ( .A(n9649), .ZN(n9196) );
  NAND2_X1 U7859 ( .A1(n9519), .A2(n8488), .ZN(n9515) );
  NAND2_X1 U7860 ( .A1(n6285), .A2(n8156), .ZN(n6287) );
  OR2_X1 U7861 ( .A1(n6013), .A2(n10101), .ZN(n6286) );
  INV_X1 U7862 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9656) );
  INV_X1 U7863 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9718) );
  OAI22_X1 U7864 ( .A1(n6193), .A2(n9656), .B1(n6305), .B2(n9718), .ZN(n6294)
         );
  INV_X1 U7865 ( .A(n6290), .ZN(n6288) );
  NAND2_X1 U7866 ( .A1(n6288), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6306) );
  INV_X1 U7867 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7868 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NAND2_X1 U7869 ( .A1(n6306), .A2(n6291), .ZN(n6649) );
  INV_X1 U7870 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6292) );
  OAI22_X1 U7871 ( .A1(n6062), .A2(n6649), .B1(n6194), .B2(n6292), .ZN(n6293)
         );
  INV_X1 U7872 ( .A(n9659), .ZN(n9528) );
  NAND2_X1 U7873 ( .A1(n9513), .A2(n9528), .ZN(n8330) );
  NAND2_X1 U7874 ( .A1(n9515), .A2(n9514), .ZN(n6295) );
  NAND2_X1 U7875 ( .A1(n6295), .A2(n8330), .ZN(n9502) );
  NAND2_X1 U7876 ( .A1(n8137), .A2(n8156), .ZN(n6297) );
  OR2_X1 U7877 ( .A1(n6013), .A2(n8576), .ZN(n6296) );
  INV_X1 U7878 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6299) );
  INV_X1 U7879 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6298) );
  OAI22_X1 U7880 ( .A1(n6193), .A2(n6299), .B1(n6305), .B2(n6298), .ZN(n6301)
         );
  INV_X1 U7881 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6789) );
  XNOR2_X1 U7882 ( .A(n6306), .B(n6789), .ZN(n9492) );
  INV_X1 U7883 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9493) );
  OAI22_X1 U7884 ( .A1(n6062), .A2(n9492), .B1(n6194), .B2(n9493), .ZN(n6300)
         );
  INV_X1 U7885 ( .A(n9650), .ZN(n9509) );
  NOR2_X1 U7886 ( .A1(n6387), .A2(n9509), .ZN(n8332) );
  INV_X1 U7887 ( .A(n8332), .ZN(n8418) );
  NAND2_X1 U7888 ( .A1(n6387), .A2(n9509), .ZN(n8331) );
  NAND2_X1 U7889 ( .A1(n8418), .A2(n8331), .ZN(n9488) );
  NAND2_X1 U7890 ( .A1(n9502), .A2(n9501), .ZN(n6302) );
  NAND2_X1 U7891 ( .A1(n6302), .A2(n8331), .ZN(n6310) );
  NAND2_X1 U7892 ( .A1(n9163), .A2(n8156), .ZN(n6304) );
  OR2_X1 U7893 ( .A1(n6013), .A2(n9755), .ZN(n6303) );
  INV_X1 U7894 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6430) );
  INV_X1 U7895 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6658) );
  OAI22_X1 U7896 ( .A1(n6193), .A2(n6430), .B1(n6305), .B2(n6658), .ZN(n6309)
         );
  INV_X1 U7897 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7898 ( .A1(n6307), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9477) );
  INV_X1 U7899 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9478) );
  OAI22_X1 U7900 ( .A1(n6062), .A2(n9477), .B1(n6194), .B2(n9478), .ZN(n6308)
         );
  OR2_X1 U7901 ( .A1(n6309), .A2(n6308), .ZN(n9642) );
  INV_X1 U7902 ( .A(n9642), .ZN(n9496) );
  NAND2_X1 U7903 ( .A1(n9480), .A2(n9496), .ZN(n8421) );
  XNOR2_X1 U7904 ( .A(n6310), .B(n8393), .ZN(n6329) );
  NAND2_X1 U7905 ( .A1(n6311), .A2(n6312), .ZN(n6318) );
  NAND2_X1 U7906 ( .A1(n6317), .A2(n6316), .ZN(n6313) );
  NAND2_X1 U7907 ( .A1(n6314), .A2(n9899), .ZN(n6412) );
  NAND2_X1 U7908 ( .A1(n8434), .A2(n6393), .ZN(n6320) );
  NAND2_X1 U7909 ( .A1(n8439), .A2(n6390), .ZN(n8505) );
  NAND2_X1 U7910 ( .A1(n6320), .A2(n8505), .ZN(n10250) );
  INV_X1 U7911 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7912 ( .A1(n8162), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7913 ( .A1(n8163), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6321) );
  OAI211_X1 U7914 ( .C1(n6193), .C2(n6323), .A(n6322), .B(n6321), .ZN(n9296)
         );
  OR2_X1 U7915 ( .A1(n6391), .A2(n6325), .ZN(n8430) );
  INV_X1 U7916 ( .A(n8430), .ZN(n6921) );
  AND2_X1 U7917 ( .A1(n4524), .A2(n6921), .ZN(n10371) );
  INV_X1 U7918 ( .A(P1_B_REG_SCAN_IN), .ZN(n6400) );
  OR2_X1 U7919 ( .A1(n6326), .A2(n6400), .ZN(n6327) );
  AND2_X1 U7920 ( .A1(n10371), .A2(n6327), .ZN(n8166) );
  AND2_X1 U7921 ( .A1(n9296), .A2(n8166), .ZN(n6328) );
  AOI21_X1 U7922 ( .B1(n6329), .B2(n10250), .A(n6328), .ZN(n9487) );
  INV_X1 U7923 ( .A(n10298), .ZN(n10253) );
  XNOR2_X1 U7924 ( .A(n9308), .B(n10253), .ZN(n10248) );
  INV_X1 U7925 ( .A(n10248), .ZN(n10245) );
  NAND2_X1 U7926 ( .A1(n7032), .A2(n6440), .ZN(n10263) );
  NAND2_X1 U7927 ( .A1(n8361), .A2(n10263), .ZN(n6335) );
  NAND2_X1 U7928 ( .A1(n7068), .A2(n10290), .ZN(n6334) );
  NAND2_X1 U7929 ( .A1(n10245), .A2(n10246), .ZN(n6338) );
  INV_X1 U7930 ( .A(n9308), .ZN(n6336) );
  NAND2_X1 U7931 ( .A1(n6336), .A2(n10298), .ZN(n6337) );
  NAND2_X1 U7932 ( .A1(n6338), .A2(n6337), .ZN(n7605) );
  NAND2_X1 U7933 ( .A1(n7605), .A2(n8360), .ZN(n6340) );
  INV_X1 U7934 ( .A(n9307), .ZN(n7067) );
  NAND2_X1 U7935 ( .A1(n7067), .A2(n7609), .ZN(n6339) );
  NAND2_X1 U7936 ( .A1(n6340), .A2(n6339), .ZN(n10237) );
  NAND2_X1 U7937 ( .A1(n8230), .A2(n8249), .ZN(n10238) );
  NAND2_X1 U7938 ( .A1(n10237), .A2(n10238), .ZN(n6342) );
  NAND2_X1 U7939 ( .A1(n6470), .A2(n10311), .ZN(n6341) );
  NAND2_X1 U7940 ( .A1(n6342), .A2(n6341), .ZN(n7503) );
  NAND2_X1 U7941 ( .A1(n6343), .A2(n8450), .ZN(n8362) );
  NAND2_X1 U7942 ( .A1(n7503), .A2(n8362), .ZN(n6345) );
  NAND2_X1 U7943 ( .A1(n8237), .A2(n10318), .ZN(n6344) );
  OR2_X1 U7944 ( .A1(n8226), .A2(n8449), .ZN(n7516) );
  INV_X1 U7945 ( .A(n9305), .ZN(n8233) );
  NAND2_X1 U7946 ( .A1(n8233), .A2(n10326), .ZN(n6346) );
  AND2_X1 U7947 ( .A1(n6347), .A2(n7633), .ZN(n8245) );
  INV_X1 U7948 ( .A(n8245), .ZN(n7634) );
  NAND2_X1 U7949 ( .A1(n10332), .A2(n7755), .ZN(n6348) );
  NAND2_X1 U7950 ( .A1(n6349), .A2(n6348), .ZN(n10224) );
  NAND2_X1 U7951 ( .A1(n7637), .A2(n8258), .ZN(n10225) );
  OR2_X1 U7952 ( .A1(n10223), .A2(n10341), .ZN(n6350) );
  NAND2_X1 U7953 ( .A1(n8261), .A2(n8453), .ZN(n7639) );
  INV_X1 U7954 ( .A(n6351), .ZN(n7473) );
  NAND2_X1 U7955 ( .A1(n7463), .A2(n7473), .ZN(n6353) );
  NAND2_X1 U7956 ( .A1(n10352), .A2(n10359), .ZN(n6352) );
  NAND2_X1 U7957 ( .A1(n6353), .A2(n6352), .ZN(n7587) );
  NAND2_X1 U7958 ( .A1(n7587), .A2(n7595), .ZN(n6355) );
  NAND2_X1 U7959 ( .A1(n7887), .A2(n7952), .ZN(n6354) );
  NAND2_X1 U7960 ( .A1(n6355), .A2(n6354), .ZN(n7680) );
  NAND2_X1 U7961 ( .A1(n7680), .A2(n7681), .ZN(n6357) );
  OR2_X1 U7962 ( .A1(n7944), .A2(n9303), .ZN(n6356) );
  NAND2_X1 U7963 ( .A1(n6357), .A2(n6356), .ZN(n7728) );
  NAND2_X1 U7964 ( .A1(n10383), .A2(n8104), .ZN(n6358) );
  NAND2_X1 U7965 ( .A1(n10210), .A2(n9302), .ZN(n6359) );
  NAND2_X1 U7966 ( .A1(n6360), .A2(n6359), .ZN(n7897) );
  OR2_X1 U7967 ( .A1(n8284), .A2(n9301), .ZN(n6361) );
  OR2_X1 U7968 ( .A1(n10196), .A2(n8092), .ZN(n6362) );
  OR2_X1 U7969 ( .A1(n9222), .A2(n9299), .ZN(n6363) );
  NAND2_X1 U7970 ( .A1(n6364), .A2(n6363), .ZN(n8052) );
  NAND2_X1 U7971 ( .A1(n9275), .A2(n9298), .ZN(n6365) );
  NAND2_X1 U7972 ( .A1(n8052), .A2(n6365), .ZN(n6367) );
  OR2_X1 U7973 ( .A1(n9275), .A2(n9298), .ZN(n6366) );
  NAND2_X1 U7974 ( .A1(n6367), .A2(n6366), .ZN(n8133) );
  INV_X1 U7975 ( .A(n8133), .ZN(n6368) );
  OR2_X1 U7976 ( .A1(n8129), .A2(n9297), .ZN(n8300) );
  NAND2_X1 U7977 ( .A1(n8129), .A2(n9297), .ZN(n6369) );
  OR2_X1 U7978 ( .A1(n9627), .A2(n9693), .ZN(n6370) );
  NOR2_X1 U7979 ( .A1(n9615), .A2(n9684), .ZN(n6373) );
  NAND2_X1 U7980 ( .A1(n9615), .A2(n9684), .ZN(n6372) );
  OR2_X1 U7981 ( .A1(n9595), .A2(n9692), .ZN(n6374) );
  NAND2_X1 U7982 ( .A1(n9584), .A2(n6374), .ZN(n6376) );
  NAND2_X1 U7983 ( .A1(n9595), .A2(n9692), .ZN(n6375) );
  NAND2_X1 U7984 ( .A1(n6376), .A2(n6375), .ZN(n9575) );
  AND2_X1 U7985 ( .A1(n9576), .A2(n9683), .ZN(n6377) );
  NAND2_X1 U7986 ( .A1(n6379), .A2(n5142), .ZN(n6381) );
  NAND2_X1 U7987 ( .A1(n9728), .A2(n9559), .ZN(n6380) );
  AND2_X1 U7988 ( .A1(n9724), .A2(n9196), .ZN(n6382) );
  OR2_X1 U7989 ( .A1(n9724), .A2(n9196), .ZN(n6383) );
  INV_X1 U7990 ( .A(n6383), .ZN(n6384) );
  INV_X1 U7991 ( .A(n9514), .ZN(n6386) );
  NOR2_X1 U7992 ( .A1(n9513), .A2(n9659), .ZN(n6385) );
  NAND2_X1 U7993 ( .A1(n9489), .A2(n9488), .ZN(n9491) );
  NAND2_X1 U7994 ( .A1(n6387), .A2(n9650), .ZN(n6388) );
  NAND2_X1 U7995 ( .A1(n9491), .A2(n6388), .ZN(n6389) );
  XNOR2_X1 U7996 ( .A(n6389), .B(n8393), .ZN(n9485) );
  OR2_X1 U7997 ( .A1(n6434), .A2(n8430), .ZN(n6639) );
  AND2_X1 U7998 ( .A1(n6391), .A2(n6325), .ZN(n6428) );
  INV_X1 U7999 ( .A(n6428), .ZN(n6968) );
  AND2_X1 U8000 ( .A1(n6639), .A2(n6968), .ZN(n7570) );
  NAND2_X1 U8001 ( .A1(n6434), .A2(n6435), .ZN(n6394) );
  NAND2_X1 U8002 ( .A1(n7570), .A2(n6394), .ZN(n7471) );
  OR2_X1 U8003 ( .A1(n4524), .A2(n8430), .ZN(n10358) );
  INV_X1 U8004 ( .A(n9627), .ZN(n9744) );
  NAND2_X1 U8005 ( .A1(n10240), .A2(n10311), .ZN(n10239) );
  INV_X1 U8006 ( .A(n10326), .ZN(n8240) );
  INV_X1 U8007 ( .A(n10223), .ZN(n10338) );
  INV_X1 U8008 ( .A(n10342), .ZN(n7476) );
  NAND3_X1 U8009 ( .A1(n10228), .A2(n10352), .A3(n7476), .ZN(n7588) );
  AND2_X2 U8010 ( .A1(n9728), .A2(n9552), .ZN(n9539) );
  NAND2_X1 U8011 ( .A1(n6428), .A2(n8512), .ZN(n9626) );
  AOI21_X1 U8012 ( .B1(n9480), .B2(n9498), .A(n9626), .ZN(n6397) );
  NAND2_X1 U8013 ( .A1(n6397), .A2(n9471), .ZN(n9483) );
  OAI21_X1 U8014 ( .B1(n9509), .B2(n10358), .A(n9483), .ZN(n6398) );
  AOI21_X1 U8015 ( .B1(n9485), .B2(n10385), .A(n6398), .ZN(n6399) );
  AND2_X1 U8016 ( .A1(n9487), .A2(n6399), .ZN(n6663) );
  XNOR2_X1 U8017 ( .A(n6406), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8036) );
  OR2_X1 U8018 ( .A1(n8036), .A2(n6400), .ZN(n6404) );
  NAND2_X1 U8019 ( .A1(n4575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6401) );
  MUX2_X1 U8020 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6401), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6403) );
  NAND2_X1 U8021 ( .A1(n6403), .A2(n6402), .ZN(n7993) );
  INV_X1 U8022 ( .A(n7993), .ZN(n6410) );
  MUX2_X1 U8023 ( .A(n6404), .B(P1_B_REG_SCAN_IN), .S(n6410), .Z(n6409) );
  NAND2_X1 U8024 ( .A1(n6406), .A2(n6405), .ZN(n6407) );
  NAND2_X1 U8025 ( .A1(n6409), .A2(n8082), .ZN(n9750) );
  OR2_X1 U8026 ( .A1(n8082), .A2(n6410), .ZN(n9753) );
  OAI21_X1 U8027 ( .B1(n9750), .B2(P1_D_REG_0__SCAN_IN), .A(n9753), .ZN(n7465)
         );
  NAND2_X1 U8028 ( .A1(n6412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6413) );
  XNOR2_X1 U8029 ( .A(n6413), .B(n10083), .ZN(n6922) );
  AND2_X1 U8030 ( .A1(n6922), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8031 ( .A1(n6437), .A2(n6912), .ZN(n9749) );
  NAND2_X1 U8032 ( .A1(n6434), .A2(n6921), .ZN(n6646) );
  INV_X1 U8033 ( .A(n6646), .ZN(n6414) );
  OR2_X1 U8034 ( .A1(n9749), .A2(n6414), .ZN(n6655) );
  NOR2_X1 U8035 ( .A1(n7465), .A2(n6655), .ZN(n6427) );
  INV_X1 U8036 ( .A(n9750), .ZN(n6424) );
  NOR4_X1 U8037 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6423) );
  NOR4_X1 U8038 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6422) );
  INV_X1 U8039 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10284) );
  INV_X1 U8040 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10286) );
  INV_X1 U8041 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10287) );
  INV_X1 U8042 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10285) );
  NAND4_X1 U8043 ( .A1(n10284), .A2(n10286), .A3(n10287), .A4(n10285), .ZN(
        n6420) );
  NOR4_X1 U8044 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6418) );
  NOR4_X1 U8045 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6417) );
  NOR4_X1 U8046 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6416) );
  NOR4_X1 U8047 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6415) );
  NAND4_X1 U8048 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n6419)
         );
  NOR4_X1 U8049 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6420), .A4(n6419), .ZN(n6421) );
  NAND3_X1 U8050 ( .A1(n6423), .A2(n6422), .A3(n6421), .ZN(n6632) );
  NAND2_X1 U8051 ( .A1(n6424), .A2(n6632), .ZN(n6426) );
  OR2_X1 U8052 ( .A1(n8082), .A2(n8036), .ZN(n9752) );
  OAI21_X1 U8053 ( .B1(n9750), .B2(P1_D_REG_1__SCAN_IN), .A(n9752), .ZN(n6425)
         );
  AND3_X1 U8054 ( .A1(n6426), .A2(n6425), .A3(n6635), .ZN(n6657) );
  AND2_X2 U8055 ( .A1(n6427), .A2(n6657), .ZN(n10413) );
  NAND2_X1 U8056 ( .A1(n6434), .A2(n6428), .ZN(n10388) );
  INV_X1 U8057 ( .A(n10388), .ZN(n10363) );
  NAND2_X1 U8058 ( .A1(n10413), .A2(n10363), .ZN(n9710) );
  OAI21_X1 U8059 ( .B1(n6663), .B2(n10411), .A(n6432), .ZN(P1_U3551) );
  INV_X1 U8060 ( .A(n6437), .ZN(n6439) );
  INV_X1 U8061 ( .A(n6433), .ZN(n7469) );
  NAND2_X1 U8062 ( .A1(n6434), .A2(n6433), .ZN(n6436) );
  NAND2_X1 U8063 ( .A1(n6436), .A2(n6435), .ZN(n6438) );
  INV_X1 U8064 ( .A(n6440), .ZN(n10274) );
  OAI22_X1 U8065 ( .A1(n10265), .A2(n6451), .B1(n6461), .B2(n10274), .ZN(n6441) );
  AOI21_X1 U8066 ( .B1(n6439), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6441), .ZN(
        n6983) );
  AOI222_X1 U8067 ( .A1(n7032), .A2(n6786), .B1(n6440), .B2(n6446), .C1(n6439), 
        .C2(P1_IR_REG_0__SCAN_IN), .ZN(n6984) );
  NOR2_X1 U8068 ( .A1(n6983), .A2(n6984), .ZN(n6982) );
  INV_X1 U8069 ( .A(n6441), .ZN(n6442) );
  NOR2_X1 U8070 ( .A1(n6982), .A2(n5138), .ZN(n7029) );
  NAND2_X1 U8071 ( .A1(n9310), .A2(n6446), .ZN(n6443) );
  NAND2_X1 U8072 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  XNOR2_X1 U8073 ( .A(n6445), .B(n6546), .ZN(n6450) );
  INV_X1 U8074 ( .A(n6450), .ZN(n6448) );
  AOI22_X1 U8075 ( .A1(n9310), .A2(n6786), .B1(n6446), .B2(n10276), .ZN(n6449)
         );
  NAND2_X1 U8076 ( .A1(n6448), .A2(n6447), .ZN(n7026) );
  AOI21_X1 U8077 ( .B1(n7029), .B2(n7026), .A(n7025), .ZN(n7066) );
  NAND2_X1 U8078 ( .A1(n9308), .A2(n6786), .ZN(n6453) );
  OR2_X1 U8079 ( .A1(n10298), .A2(n6451), .ZN(n6452) );
  AND2_X1 U8080 ( .A1(n6453), .A2(n6452), .ZN(n6458) );
  NAND2_X1 U8081 ( .A1(n9308), .A2(n6446), .ZN(n6455) );
  NAND2_X1 U8082 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  NOR2_X1 U8083 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  INV_X1 U8084 ( .A(n6459), .ZN(n6460) );
  AOI22_X1 U8085 ( .A1(n6446), .A2(n10303), .B1(n9307), .B2(n6786), .ZN(n6471)
         );
  NAND2_X1 U8086 ( .A1(n9307), .A2(n6446), .ZN(n6463) );
  OR2_X1 U8087 ( .A1(n7609), .A2(n6461), .ZN(n6462) );
  NAND2_X1 U8088 ( .A1(n6463), .A2(n6462), .ZN(n6465) );
  XNOR2_X1 U8089 ( .A(n6465), .B(n6612), .ZN(n6473) );
  XOR2_X1 U8090 ( .A(n6471), .B(n6473), .Z(n7174) );
  NAND2_X1 U8091 ( .A1(n9306), .A2(n6446), .ZN(n6467) );
  OR2_X1 U8092 ( .A1(n10311), .A2(n6461), .ZN(n6466) );
  NAND2_X1 U8093 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  XNOR2_X1 U8094 ( .A(n6468), .B(n6784), .ZN(n6477) );
  OAI22_X1 U8095 ( .A1(n6470), .A2(n6469), .B1(n10311), .B2(n6451), .ZN(n6476)
         );
  XNOR2_X1 U8096 ( .A(n6477), .B(n6476), .ZN(n9235) );
  INV_X1 U8097 ( .A(n6471), .ZN(n6472) );
  NOR2_X1 U8098 ( .A1(n6473), .A2(n6472), .ZN(n9236) );
  INV_X1 U8099 ( .A(n6482), .ZN(n6480) );
  AOI22_X1 U8100 ( .A1(n10323), .A2(n6446), .B1(n8236), .B2(n6781), .ZN(n6478)
         );
  INV_X1 U8101 ( .A(n6546), .ZN(n6612) );
  XNOR2_X1 U8102 ( .A(n6478), .B(n6612), .ZN(n6481) );
  INV_X1 U8103 ( .A(n6481), .ZN(n6479) );
  NAND2_X1 U8104 ( .A1(n6480), .A2(n6479), .ZN(n6483) );
  NAND2_X1 U8105 ( .A1(n6482), .A2(n6481), .ZN(n6484) );
  AOI22_X1 U8106 ( .A1(n10323), .A2(n6786), .B1(n6446), .B2(n8236), .ZN(n7450)
         );
  NAND2_X1 U8107 ( .A1(n9305), .A2(n6446), .ZN(n6485) );
  OAI21_X1 U8108 ( .B1(n10326), .B2(n6461), .A(n6485), .ZN(n6486) );
  XNOR2_X1 U8109 ( .A(n6486), .B(n6784), .ZN(n6490) );
  OR2_X1 U8110 ( .A1(n10326), .A2(n6451), .ZN(n6488) );
  NAND2_X1 U8111 ( .A1(n9305), .A2(n6786), .ZN(n6487) );
  NAND2_X1 U8112 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  NAND2_X1 U8113 ( .A1(n6490), .A2(n6489), .ZN(n7456) );
  OR2_X1 U8114 ( .A1(n10332), .A2(n6451), .ZN(n6492) );
  NAND2_X1 U8115 ( .A1(n10322), .A2(n6786), .ZN(n6491) );
  NAND2_X1 U8116 ( .A1(n6492), .A2(n6491), .ZN(n6495) );
  AOI22_X1 U8117 ( .A1(n7497), .A2(n6781), .B1(n6446), .B2(n10322), .ZN(n6493)
         );
  XNOR2_X1 U8118 ( .A(n6493), .B(n6784), .ZN(n6494) );
  XOR2_X1 U8119 ( .A(n6495), .B(n6494), .Z(n7580) );
  INV_X1 U8120 ( .A(n6494), .ZN(n6496) );
  AOI22_X1 U8121 ( .A1(n10342), .A2(n6781), .B1(n6446), .B2(n10349), .ZN(n6497) );
  XNOR2_X1 U8122 ( .A(n6497), .B(n6612), .ZN(n7851) );
  INV_X1 U8123 ( .A(n7851), .ZN(n6505) );
  NAND2_X1 U8124 ( .A1(n10342), .A2(n6446), .ZN(n6499) );
  NAND2_X1 U8125 ( .A1(n10349), .A2(n6786), .ZN(n6498) );
  AND2_X1 U8126 ( .A1(n6499), .A2(n6498), .ZN(n6507) );
  INV_X1 U8127 ( .A(n6507), .ZN(n7850) );
  NAND2_X1 U8128 ( .A1(n10223), .A2(n6781), .ZN(n6501) );
  NAND2_X1 U8129 ( .A1(n10341), .A2(n6446), .ZN(n6500) );
  NAND2_X1 U8130 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  XNOR2_X1 U8131 ( .A(n6502), .B(n6612), .ZN(n7847) );
  NAND2_X1 U8132 ( .A1(n10223), .A2(n6446), .ZN(n6504) );
  NAND2_X1 U8133 ( .A1(n10341), .A2(n6786), .ZN(n6503) );
  NAND2_X1 U8134 ( .A1(n6504), .A2(n6503), .ZN(n7753) );
  OAI22_X1 U8135 ( .A1(n6505), .A2(n7850), .B1(n7847), .B2(n7753), .ZN(n6511)
         );
  NAND2_X1 U8136 ( .A1(n7847), .A2(n7753), .ZN(n6506) );
  INV_X1 U8137 ( .A(n6506), .ZN(n6509) );
  AOI21_X1 U8138 ( .B1(n6507), .B2(n6506), .A(n7851), .ZN(n6508) );
  AOI21_X1 U8139 ( .B1(n6509), .B2(n7850), .A(n6508), .ZN(n6510) );
  AOI22_X1 U8140 ( .A1(n7484), .A2(n6781), .B1(n6446), .B2(n9304), .ZN(n6512)
         );
  XOR2_X1 U8141 ( .A(n6784), .B(n6512), .Z(n6513) );
  NOR2_X1 U8142 ( .A1(n6515), .A2(n6516), .ZN(n7807) );
  AOI22_X1 U8143 ( .A1(n7484), .A2(n6446), .B1(n6786), .B2(n9304), .ZN(n7808)
         );
  OAI22_X1 U8144 ( .A1(n7887), .A2(n6461), .B1(n7952), .B2(n6451), .ZN(n6517)
         );
  XNOR2_X1 U8145 ( .A(n6517), .B(n6546), .ZN(n6520) );
  OR2_X1 U8146 ( .A1(n7887), .A2(n6451), .ZN(n6519) );
  NAND2_X1 U8147 ( .A1(n10373), .A2(n6786), .ZN(n6518) );
  AND2_X1 U8148 ( .A1(n6519), .A2(n6518), .ZN(n6521) );
  NAND2_X1 U8149 ( .A1(n6520), .A2(n6521), .ZN(n7945) );
  INV_X1 U8150 ( .A(n6520), .ZN(n6523) );
  INV_X1 U8151 ( .A(n6521), .ZN(n6522) );
  NAND2_X1 U8152 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  AND2_X1 U8153 ( .A1(n7945), .A2(n6524), .ZN(n7879) );
  NAND2_X1 U8154 ( .A1(n7944), .A2(n6781), .ZN(n6526) );
  NAND2_X1 U8155 ( .A1(n9303), .A2(n6446), .ZN(n6525) );
  NAND2_X1 U8156 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  XNOR2_X1 U8157 ( .A(n6527), .B(n6546), .ZN(n6529) );
  AND2_X1 U8158 ( .A1(n9303), .A2(n6786), .ZN(n6528) );
  AOI21_X1 U8159 ( .B1(n7944), .B2(n6446), .A(n6528), .ZN(n6530) );
  NAND2_X1 U8160 ( .A1(n6529), .A2(n6530), .ZN(n8043) );
  INV_X1 U8161 ( .A(n6529), .ZN(n6532) );
  INV_X1 U8162 ( .A(n6530), .ZN(n6531) );
  NAND2_X1 U8163 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  NAND2_X1 U8164 ( .A1(n6534), .A2(n7946), .ZN(n7948) );
  OAI22_X1 U8165 ( .A1(n10383), .A2(n6461), .B1(n8104), .B2(n6451), .ZN(n6535)
         );
  XNOR2_X1 U8166 ( .A(n6535), .B(n6612), .ZN(n6537) );
  OAI22_X1 U8167 ( .A1(n10383), .A2(n6451), .B1(n8104), .B2(n6469), .ZN(n6536)
         );
  OR2_X1 U8168 ( .A1(n6537), .A2(n6536), .ZN(n6539) );
  NAND2_X1 U8169 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  AND2_X1 U8170 ( .A1(n6539), .A2(n6538), .ZN(n8042) );
  AOI22_X1 U8171 ( .A1(n10210), .A2(n6781), .B1(n6446), .B2(n9302), .ZN(n6540)
         );
  INV_X1 U8172 ( .A(n10210), .ZN(n10389) );
  OAI22_X1 U8173 ( .A1(n10389), .A2(n6451), .B1(n6541), .B2(n6469), .ZN(n8103)
         );
  NAND2_X1 U8174 ( .A1(n8100), .A2(n8103), .ZN(n6544) );
  INV_X1 U8175 ( .A(n6542), .ZN(n6543) );
  NAND2_X1 U8176 ( .A1(n6543), .A2(n4541), .ZN(n8101) );
  OAI22_X1 U8177 ( .A1(n4714), .A2(n6451), .B1(n9207), .B2(n6469), .ZN(n8087)
         );
  AOI22_X1 U8178 ( .A1(n8284), .A2(n6781), .B1(n6446), .B2(n9301), .ZN(n6545)
         );
  XOR2_X1 U8179 ( .A(n6784), .B(n6545), .Z(n8086) );
  OAI22_X1 U8180 ( .A1(n10196), .A2(n6461), .B1(n8092), .B2(n6451), .ZN(n6547)
         );
  INV_X1 U8181 ( .A(n6546), .ZN(n6784) );
  XNOR2_X1 U8182 ( .A(n6547), .B(n6784), .ZN(n6551) );
  OR2_X1 U8183 ( .A1(n10196), .A2(n6451), .ZN(n6549) );
  NAND2_X1 U8184 ( .A1(n9300), .A2(n6786), .ZN(n6548) );
  NAND2_X1 U8185 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NOR2_X1 U8186 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  AOI21_X1 U8187 ( .B1(n6551), .B2(n6550), .A(n6552), .ZN(n9204) );
  NAND2_X1 U8188 ( .A1(n9222), .A2(n6781), .ZN(n6554) );
  NAND2_X1 U8189 ( .A1(n9299), .A2(n6446), .ZN(n6553) );
  NAND2_X1 U8190 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  XNOR2_X1 U8191 ( .A(n6555), .B(n6784), .ZN(n6558) );
  NAND2_X1 U8192 ( .A1(n9222), .A2(n6446), .ZN(n6557) );
  NAND2_X1 U8193 ( .A1(n9299), .A2(n6786), .ZN(n6556) );
  NAND2_X1 U8194 ( .A1(n6557), .A2(n6556), .ZN(n6559) );
  NAND2_X1 U8195 ( .A1(n6558), .A2(n6559), .ZN(n9214) );
  NAND2_X1 U8196 ( .A1(n9213), .A2(n9214), .ZN(n9212) );
  INV_X1 U8197 ( .A(n6558), .ZN(n6561) );
  INV_X1 U8198 ( .A(n6559), .ZN(n6560) );
  NAND2_X1 U8199 ( .A1(n6561), .A2(n6560), .ZN(n9216) );
  NAND2_X1 U8200 ( .A1(n9212), .A2(n9216), .ZN(n6563) );
  AOI22_X1 U8201 ( .A1(n9275), .A2(n6781), .B1(n6446), .B2(n9298), .ZN(n6562)
         );
  XNOR2_X1 U8202 ( .A(n6562), .B(n6784), .ZN(n6564) );
  NAND2_X1 U8203 ( .A1(n6563), .A2(n6564), .ZN(n9267) );
  NAND2_X1 U8204 ( .A1(n9267), .A2(n9270), .ZN(n6567) );
  INV_X1 U8205 ( .A(n6563), .ZN(n6566) );
  INV_X1 U8206 ( .A(n6564), .ZN(n6565) );
  NAND2_X1 U8207 ( .A1(n6566), .A2(n6565), .ZN(n9268) );
  AND2_X1 U8208 ( .A1(n9297), .A2(n6786), .ZN(n6568) );
  AOI21_X1 U8209 ( .B1(n8129), .B2(n6446), .A(n6568), .ZN(n6571) );
  AOI22_X1 U8210 ( .A1(n8129), .A2(n6781), .B1(n6446), .B2(n9297), .ZN(n6569)
         );
  XNOR2_X1 U8211 ( .A(n6569), .B(n6612), .ZN(n6570) );
  XOR2_X1 U8212 ( .A(n6571), .B(n6570), .Z(n9178) );
  INV_X1 U8213 ( .A(n6570), .ZN(n6573) );
  NAND2_X1 U8214 ( .A1(n9627), .A2(n6781), .ZN(n6576) );
  NAND2_X1 U8215 ( .A1(n9693), .A2(n6446), .ZN(n6575) );
  NAND2_X1 U8216 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  XNOR2_X1 U8217 ( .A(n6577), .B(n6612), .ZN(n9249) );
  NAND2_X1 U8218 ( .A1(n9627), .A2(n6446), .ZN(n6579) );
  NAND2_X1 U8219 ( .A1(n9693), .A2(n6786), .ZN(n6578) );
  NAND2_X1 U8220 ( .A1(n6579), .A2(n6578), .ZN(n9250) );
  AND2_X1 U8221 ( .A1(n9684), .A2(n6786), .ZN(n6581) );
  AOI21_X1 U8222 ( .B1(n9615), .B2(n6446), .A(n6581), .ZN(n6584) );
  AOI22_X1 U8223 ( .A1(n9615), .A2(n6781), .B1(n6446), .B2(n9684), .ZN(n6582)
         );
  XNOR2_X1 U8224 ( .A(n6582), .B(n6784), .ZN(n6583) );
  XOR2_X1 U8225 ( .A(n6584), .B(n6583), .Z(n9186) );
  INV_X1 U8226 ( .A(n6583), .ZN(n6586) );
  INV_X1 U8227 ( .A(n6584), .ZN(n6585) );
  NAND2_X1 U8228 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  NAND2_X1 U8229 ( .A1(n6588), .A2(n6587), .ZN(n6590) );
  AOI22_X1 U8230 ( .A1(n9595), .A2(n6781), .B1(n6446), .B2(n9692), .ZN(n6589)
         );
  XOR2_X1 U8231 ( .A(n6784), .B(n6589), .Z(n6591) );
  NAND2_X1 U8232 ( .A1(n6590), .A2(n6591), .ZN(n9258) );
  AOI22_X1 U8233 ( .A1(n9595), .A2(n6446), .B1(n6786), .B2(n9692), .ZN(n9260)
         );
  NAND2_X1 U8234 ( .A1(n9576), .A2(n6781), .ZN(n6595) );
  NAND2_X1 U8235 ( .A1(n9683), .A2(n6446), .ZN(n6594) );
  NAND2_X1 U8236 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  XNOR2_X1 U8237 ( .A(n6596), .B(n6784), .ZN(n6600) );
  NAND2_X1 U8238 ( .A1(n9576), .A2(n6446), .ZN(n6598) );
  NAND2_X1 U8239 ( .A1(n9683), .A2(n6786), .ZN(n6597) );
  NAND2_X1 U8240 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  AOI21_X1 U8241 ( .B1(n6600), .B2(n6599), .A(n9225), .ZN(n9171) );
  INV_X1 U8242 ( .A(n9225), .ZN(n6601) );
  NAND2_X1 U8243 ( .A1(n6378), .A2(n6781), .ZN(n6603) );
  NAND2_X1 U8244 ( .A1(n9568), .A2(n6446), .ZN(n6602) );
  NAND2_X1 U8245 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  XNOR2_X1 U8246 ( .A(n6604), .B(n6546), .ZN(n6606) );
  AND2_X1 U8247 ( .A1(n9568), .A2(n6786), .ZN(n6605) );
  NAND2_X1 U8248 ( .A1(n6606), .A2(n6607), .ZN(n6611) );
  INV_X1 U8249 ( .A(n6606), .ZN(n6609) );
  INV_X1 U8250 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8251 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  OAI22_X1 U8252 ( .A1(n9728), .A2(n6451), .B1(n9559), .B2(n6469), .ZN(n6617)
         );
  OAI22_X1 U8253 ( .A1(n9728), .A2(n6461), .B1(n9559), .B2(n6451), .ZN(n6613)
         );
  XNOR2_X1 U8254 ( .A(n6613), .B(n6612), .ZN(n6618) );
  XOR2_X1 U8255 ( .A(n6617), .B(n6618), .Z(n9194) );
  OAI22_X1 U8256 ( .A1(n9724), .A2(n6461), .B1(n9196), .B2(n6451), .ZN(n6614)
         );
  XNOR2_X1 U8257 ( .A(n6614), .B(n6784), .ZN(n6629) );
  NAND2_X1 U8258 ( .A1(n9649), .A2(n6786), .ZN(n6615) );
  NAND2_X1 U8259 ( .A1(n6616), .A2(n6615), .ZN(n6628) );
  XNOR2_X1 U8260 ( .A(n6629), .B(n6628), .ZN(n9282) );
  NOR2_X1 U8261 ( .A1(n6618), .A2(n6617), .ZN(n9279) );
  NOR2_X1 U8262 ( .A1(n9282), .A2(n9279), .ZN(n6619) );
  NAND2_X1 U8263 ( .A1(n9513), .A2(n6781), .ZN(n6621) );
  NAND2_X1 U8264 ( .A1(n9659), .A2(n6446), .ZN(n6620) );
  NAND2_X1 U8265 ( .A1(n6621), .A2(n6620), .ZN(n6622) );
  XNOR2_X1 U8266 ( .A(n6622), .B(n6546), .ZN(n6625) );
  INV_X1 U8267 ( .A(n6625), .ZN(n6627) );
  AND2_X1 U8268 ( .A1(n9659), .A2(n6786), .ZN(n6623) );
  AOI21_X1 U8269 ( .B1(n9513), .B2(n6446), .A(n6623), .ZN(n6624) );
  INV_X1 U8270 ( .A(n6624), .ZN(n6626) );
  AOI21_X1 U8271 ( .B1(n6627), .B2(n6626), .A(n6798), .ZN(n6631) );
  NOR2_X1 U8272 ( .A1(n4646), .A2(n4553), .ZN(n6630) );
  INV_X1 U8273 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U8274 ( .A1(n6632), .A2(n9883), .ZN(n6633) );
  OAI21_X1 U8275 ( .B1(n9750), .B2(n6633), .A(n9752), .ZN(n7464) );
  OR2_X1 U8276 ( .A1(n7465), .A2(n7464), .ZN(n6645) );
  NAND2_X1 U8277 ( .A1(n10388), .A2(n8430), .ZN(n6642) );
  OR2_X1 U8278 ( .A1(n9749), .A2(n6642), .ZN(n6634) );
  NOR2_X2 U8279 ( .A1(n6645), .A2(n6634), .ZN(n9285) );
  OR2_X1 U8280 ( .A1(n6968), .A2(n8512), .ZN(n6641) );
  OR2_X1 U8281 ( .A1(n9749), .A2(n6641), .ZN(n6636) );
  NOR2_X2 U8282 ( .A1(n9749), .A2(n6635), .ZN(n10271) );
  NAND2_X1 U8283 ( .A1(n9513), .A2(n6637), .ZN(n6653) );
  OR2_X1 U8284 ( .A1(n9749), .A2(n6434), .ZN(n6638) );
  NOR2_X1 U8285 ( .A1(n6645), .A2(n6638), .ZN(n7030) );
  INV_X1 U8286 ( .A(n10371), .ZN(n10356) );
  AND2_X1 U8287 ( .A1(n7030), .A2(n10371), .ZN(n9209) );
  AOI22_X1 U8288 ( .A1(n9209), .A2(n9650), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6651) );
  NOR2_X1 U8289 ( .A1(n9749), .A2(n6639), .ZN(n8517) );
  INV_X1 U8290 ( .A(n8517), .ZN(n6640) );
  NOR2_X1 U8291 ( .A1(n6645), .A2(n6640), .ZN(n9241) );
  INV_X1 U8292 ( .A(n4524), .ZN(n6997) );
  AND2_X1 U8293 ( .A1(n9241), .A2(n6997), .ZN(n8090) );
  INV_X1 U8294 ( .A(n6641), .ZN(n10252) );
  INV_X1 U8295 ( .A(n6642), .ZN(n6643) );
  OR3_X1 U8296 ( .A1(n8517), .A2(n10252), .A3(n6643), .ZN(n6644) );
  NAND2_X1 U8297 ( .A1(n6645), .A2(n6644), .ZN(n6985) );
  AND3_X1 U8298 ( .A1(n6437), .A2(n6922), .A3(n6646), .ZN(n6647) );
  NAND2_X1 U8299 ( .A1(n6985), .A2(n6647), .ZN(n6648) );
  AND2_X1 U8300 ( .A1(n6648), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9243) );
  INV_X1 U8301 ( .A(n6649), .ZN(n9506) );
  AOI22_X1 U8302 ( .A1(n8090), .A2(n9649), .B1(n9243), .B2(n9506), .ZN(n6650)
         );
  AND2_X1 U8303 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND2_X1 U8304 ( .A1(n6654), .A2(n5148), .ZN(P1_U3214) );
  INV_X1 U8305 ( .A(n6655), .ZN(n7466) );
  AND2_X1 U8306 ( .A1(n7465), .A2(n7466), .ZN(n6656) );
  AND2_X2 U8307 ( .A1(n6657), .A2(n6656), .ZN(n10395) );
  NAND2_X1 U8308 ( .A1(n10395), .A2(n10363), .ZN(n9747) );
  NOR2_X1 U8309 ( .A1(n10395), .A2(n6658), .ZN(n6659) );
  OAI21_X1 U8310 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(P1_U3519) );
  NAND2_X1 U8311 ( .A1(n5873), .A2(n7081), .ZN(n6664) );
  NAND2_X1 U8312 ( .A1(n6664), .A2(n6693), .ZN(n6728) );
  NAND2_X1 U8313 ( .A1(n6728), .A2(n6866), .ZN(n6665) );
  NAND2_X1 U8314 ( .A1(n6665), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8315 ( .A(n8767), .ZN(n7238) );
  INV_X1 U8316 ( .A(n6763), .ZN(n7841) );
  INV_X1 U8317 ( .A(n7676), .ZN(n6959) );
  NOR2_X1 U8318 ( .A1(n7206), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8319 ( .A1(n5339), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U8320 ( .B1(n7263), .B2(n6666), .A(n6667), .ZN(n7269) );
  INV_X1 U8321 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10470) );
  NOR2_X1 U8322 ( .A1(n7269), .A2(n10470), .ZN(n7268) );
  INV_X1 U8323 ( .A(n6667), .ZN(n6668) );
  NOR2_X1 U8324 ( .A1(n7268), .A2(n6668), .ZN(n7282) );
  AOI21_X1 U8325 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6949), .A(n7281), .ZN(
        n6669) );
  NOR2_X1 U8326 ( .A1(n6669), .A2(n4993), .ZN(n6670) );
  AOI21_X1 U8327 ( .B1(n6669), .B2(n4993), .A(n6670), .ZN(n7186) );
  INV_X1 U8328 ( .A(n6670), .ZN(n7253) );
  INV_X1 U8329 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6671) );
  MUX2_X1 U8330 ( .A(n6671), .B(P2_REG2_REG_4__SCAN_IN), .S(n7261), .Z(n7254)
         );
  INV_X1 U8331 ( .A(n6932), .ZN(n7233) );
  NAND2_X1 U8332 ( .A1(n7228), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7227) );
  INV_X1 U8333 ( .A(n6672), .ZN(n7298) );
  XNOR2_X1 U8334 ( .A(n6935), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7299) );
  INV_X1 U8335 ( .A(n7363), .ZN(n6745) );
  INV_X1 U8336 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7652) );
  INV_X1 U8337 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U8338 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7416), .B1(n6952), .B2(
        n6675), .ZN(n7411) );
  NOR2_X1 U8339 ( .A1(n7563), .A2(n6676), .ZN(n6677) );
  INV_X1 U8340 ( .A(n7563), .ZN(n6962) );
  INV_X1 U8341 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7716) );
  NOR2_X2 U8342 ( .A1(n6677), .A2(n7558), .ZN(n7672) );
  INV_X1 U8343 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7786) );
  AOI22_X1 U8344 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7676), .B1(n6959), .B2(
        n7786), .ZN(n7671) );
  NOR2_X1 U8345 ( .A1(n7745), .A2(n6678), .ZN(n6679) );
  INV_X1 U8346 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7824) );
  INV_X1 U8347 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6680) );
  AOI22_X1 U8348 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6763), .B1(n7841), .B2(
        n6680), .ZN(n7829) );
  NOR2_X1 U8349 ( .A1(n8754), .A2(n6681), .ZN(n6682) );
  INV_X1 U8350 ( .A(n8754), .ZN(n7075) );
  INV_X1 U8351 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8742) );
  INV_X1 U8352 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U8353 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8767), .B1(n7238), .B2(
        n6683), .ZN(n8759) );
  AOI21_X2 U8354 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7238), .A(n8758), .ZN(
        n6684) );
  NOR2_X1 U8355 ( .A1(n8785), .A2(n6684), .ZN(n6685) );
  INV_X1 U8356 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8777) );
  XNOR2_X1 U8357 ( .A(n6684), .B(n8785), .ZN(n8776) );
  NOR2_X1 U8358 ( .A1(n8777), .A2(n8776), .ZN(n8775) );
  NOR2_X1 U8359 ( .A1(n6685), .A2(n8775), .ZN(n8801) );
  NAND2_X1 U8360 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7385), .ZN(n6686) );
  OAI21_X1 U8361 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n7385), .A(n6686), .ZN(
        n8800) );
  NOR2_X1 U8362 ( .A1(n8801), .A2(n8800), .ZN(n8799) );
  NOR2_X1 U8363 ( .A1(n8822), .A2(n6687), .ZN(n6688) );
  INV_X1 U8364 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8810) );
  INV_X1 U8365 ( .A(n8844), .ZN(n7568) );
  NAND2_X1 U8366 ( .A1(n7568), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6689) );
  OAI21_X1 U8367 ( .B1(n7568), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6689), .ZN(
        n8826) );
  INV_X1 U8368 ( .A(n6689), .ZN(n6690) );
  NOR2_X1 U8369 ( .A1(n8825), .A2(n6690), .ZN(n6691) );
  XNOR2_X1 U8370 ( .A(n7660), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6733) );
  XNOR2_X1 U8371 ( .A(n6691), .B(n6733), .ZN(n6692) );
  NOR2_X1 U8372 ( .A1(n5962), .A2(P2_U3151), .ZN(n8138) );
  AND2_X1 U8373 ( .A1(n6728), .A2(n8138), .ZN(n10420) );
  AND2_X1 U8374 ( .A1(n10420), .A2(n6864), .ZN(n7255) );
  NAND2_X1 U8375 ( .A1(n6692), .A2(n7255), .ZN(n6780) );
  INV_X1 U8376 ( .A(n6693), .ZN(n6694) );
  NOR2_X1 U8377 ( .A1(n7081), .A2(n6694), .ZN(n6695) );
  OR2_X1 U8378 ( .A1(P2_U3150), .A2(n6695), .ZN(n8816) );
  INV_X1 U8379 ( .A(n8816), .ZN(n10414) );
  INV_X1 U8380 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10550) );
  INV_X1 U8381 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6696) );
  AND2_X1 U8382 ( .A1(n6696), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8383 ( .A1(n5339), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6698) );
  OAI21_X1 U8384 ( .B1(n7263), .B2(n6697), .A(n6698), .ZN(n7266) );
  INV_X1 U8385 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10548) );
  NAND2_X1 U8386 ( .A1(n7286), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8387 ( .A1(n6949), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6699) );
  INV_X1 U8388 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U8389 ( .A1(n7250), .A2(n7245), .ZN(n6700) );
  INV_X1 U8390 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U8391 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10554), .S(n7261), .Z(n7246)
         );
  NAND2_X1 U8392 ( .A1(n6700), .A2(n7246), .ZN(n7248) );
  NAND2_X1 U8393 ( .A1(n7261), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U8394 ( .A1(n7248), .A2(n6701), .ZN(n6703) );
  INV_X1 U8395 ( .A(n6703), .ZN(n6702) );
  INV_X1 U8396 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8397 ( .A1(n6935), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8398 ( .A1(n7305), .A2(n6705), .ZN(n6706) );
  NOR2_X1 U8399 ( .A1(n6706), .A2(n7363), .ZN(n6707) );
  INV_X1 U8400 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10558) );
  INV_X1 U8401 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U8402 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7416), .B1(n6952), .B2(
        n10560), .ZN(n7402) );
  INV_X1 U8403 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U8404 ( .A1(n7563), .A2(n6709), .ZN(n6710) );
  INV_X1 U8405 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U8406 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7676), .B1(n6959), .B2(
        n10564), .ZN(n7662) );
  NOR2_X1 U8407 ( .A1(n7745), .A2(n6711), .ZN(n6712) );
  INV_X1 U8408 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10566) );
  INV_X1 U8409 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6713) );
  MUX2_X1 U8410 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6713), .S(n6763), .Z(n7837)
         );
  NOR2_X1 U8411 ( .A1(n8754), .A2(n6714), .ZN(n6715) );
  INV_X1 U8412 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8748) );
  XNOR2_X1 U8413 ( .A(n8754), .B(n6714), .ZN(n8749) );
  NOR2_X1 U8414 ( .A1(n8748), .A2(n8749), .ZN(n8747) );
  XNOR2_X1 U8415 ( .A(n7238), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8764) );
  NOR2_X1 U8416 ( .A1(n8765), .A2(n8764), .ZN(n8763) );
  NOR2_X1 U8417 ( .A1(n8785), .A2(n6716), .ZN(n6717) );
  INV_X1 U8418 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8781) );
  XNOR2_X1 U8419 ( .A(n7385), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8793) );
  INV_X1 U8420 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U8421 ( .A1(n7568), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6721) );
  OAI21_X1 U8422 ( .B1(n7568), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6721), .ZN(
        n8834) );
  INV_X1 U8423 ( .A(n6721), .ZN(n6722) );
  NOR2_X1 U8424 ( .A1(n8833), .A2(n6722), .ZN(n6723) );
  XNOR2_X1 U8425 ( .A(n7660), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6732) );
  XNOR2_X1 U8426 ( .A(n6723), .B(n6732), .ZN(n6726) );
  INV_X1 U8427 ( .A(n10420), .ZN(n6724) );
  OR2_X1 U8428 ( .A1(n6724), .A2(n6864), .ZN(n8837) );
  NAND2_X1 U8429 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  NAND2_X1 U8430 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U8431 ( .A1(n6727), .A2(n8615), .ZN(n6731) );
  INV_X1 U8432 ( .A(n6979), .ZN(n7092) );
  NOR2_X1 U8433 ( .A1(n6773), .A2(P2_U3151), .ZN(n8124) );
  NAND2_X1 U8434 ( .A1(n6728), .A2(n8124), .ZN(n6729) );
  MUX2_X1 U8435 ( .A(n8831), .B(n6729), .S(n5962), .Z(n8830) );
  NOR2_X1 U8436 ( .A1(n8830), .A2(n7660), .ZN(n6730) );
  MUX2_X1 U8437 ( .A(n6733), .B(n6732), .S(n6773), .Z(n6777) );
  MUX2_X1 U8438 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6773), .Z(n6767) );
  MUX2_X1 U8439 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6773), .Z(n6766) );
  MUX2_X1 U8440 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6773), .Z(n6761) );
  INV_X1 U8441 ( .A(n6761), .ZN(n6762) );
  MUX2_X1 U8442 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6773), .Z(n6739) );
  MUX2_X1 U8443 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6773), .Z(n6735) );
  XOR2_X1 U8444 ( .A(n7263), .B(n6735), .Z(n7262) );
  INV_X1 U8445 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6734) );
  MUX2_X1 U8446 ( .A(n7206), .B(n6734), .S(n6773), .Z(n10417) );
  NAND2_X1 U8447 ( .A1(n10417), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U8448 ( .A1(n7262), .A2(n10416), .B1(n6735), .B2(n7263), .ZN(n7280)
         );
  MUX2_X1 U8449 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6773), .Z(n6736) );
  XNOR2_X1 U8450 ( .A(n6736), .B(n6949), .ZN(n7279) );
  INV_X1 U8451 ( .A(n6949), .ZN(n7292) );
  INV_X1 U8452 ( .A(n6736), .ZN(n6737) );
  OAI22_X1 U8453 ( .A1(n7280), .A2(n7279), .B1(n7292), .B2(n6737), .ZN(n7181)
         );
  MUX2_X1 U8454 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6773), .Z(n6738) );
  XNOR2_X1 U8455 ( .A(n6738), .B(n6929), .ZN(n7182) );
  NOR2_X1 U8456 ( .A1(n7181), .A2(n7182), .ZN(n7242) );
  NOR2_X1 U8457 ( .A1(n6738), .A2(n6929), .ZN(n7241) );
  XNOR2_X1 U8458 ( .A(n6739), .B(n7261), .ZN(n7240) );
  NOR3_X1 U8459 ( .A1(n7242), .A2(n7241), .A3(n7240), .ZN(n7239) );
  AOI21_X1 U8460 ( .B1(n6739), .B2(n7261), .A(n7239), .ZN(n7225) );
  MUX2_X1 U8461 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6773), .Z(n6740) );
  XNOR2_X1 U8462 ( .A(n6740), .B(n6932), .ZN(n7224) );
  INV_X1 U8463 ( .A(n6740), .ZN(n6741) );
  OAI22_X1 U8464 ( .A1(n7225), .A2(n7224), .B1(n7233), .B2(n6741), .ZN(n7296)
         );
  INV_X1 U8465 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9038) );
  MUX2_X1 U8466 ( .A(n9038), .B(n6742), .S(n6773), .Z(n6743) );
  INV_X1 U8467 ( .A(n6935), .ZN(n7311) );
  NAND2_X1 U8468 ( .A1(n6743), .A2(n7311), .ZN(n6744) );
  OAI21_X1 U8469 ( .B1(n6743), .B2(n7311), .A(n6744), .ZN(n7295) );
  NOR2_X1 U8470 ( .A1(n7296), .A2(n7295), .ZN(n7354) );
  INV_X1 U8471 ( .A(n6744), .ZN(n7353) );
  MUX2_X1 U8472 ( .A(n7652), .B(n10558), .S(n6773), .Z(n6746) );
  NAND2_X1 U8473 ( .A1(n6746), .A2(n6745), .ZN(n7405) );
  INV_X1 U8474 ( .A(n6746), .ZN(n6747) );
  NAND2_X1 U8475 ( .A1(n6747), .A2(n7363), .ZN(n6748) );
  AND2_X1 U8476 ( .A1(n7405), .A2(n6748), .ZN(n7352) );
  OAI21_X1 U8477 ( .B1(n7354), .B2(n7353), .A(n7352), .ZN(n7406) );
  MUX2_X1 U8478 ( .A(n6675), .B(n10560), .S(n6773), .Z(n6749) );
  NAND2_X1 U8479 ( .A1(n6749), .A2(n7416), .ZN(n6752) );
  INV_X1 U8480 ( .A(n6749), .ZN(n6750) );
  NAND2_X1 U8481 ( .A1(n6750), .A2(n6952), .ZN(n6751) );
  NAND2_X1 U8482 ( .A1(n6752), .A2(n6751), .ZN(n7404) );
  AOI21_X1 U8483 ( .B1(n7406), .B2(n7405), .A(n7404), .ZN(n7554) );
  INV_X1 U8484 ( .A(n6752), .ZN(n7553) );
  MUX2_X1 U8485 ( .A(n7716), .B(n10562), .S(n6773), .Z(n6753) );
  NAND2_X1 U8486 ( .A1(n6753), .A2(n7563), .ZN(n7665) );
  INV_X1 U8487 ( .A(n6753), .ZN(n6754) );
  NAND2_X1 U8488 ( .A1(n6754), .A2(n6962), .ZN(n6755) );
  AND2_X1 U8489 ( .A1(n7665), .A2(n6755), .ZN(n7552) );
  OAI21_X1 U8490 ( .B1(n7554), .B2(n7553), .A(n7552), .ZN(n7666) );
  MUX2_X1 U8491 ( .A(n7786), .B(n10564), .S(n6773), .Z(n6756) );
  NAND2_X1 U8492 ( .A1(n6756), .A2(n7676), .ZN(n6759) );
  INV_X1 U8493 ( .A(n6756), .ZN(n6757) );
  NAND2_X1 U8494 ( .A1(n6757), .A2(n6959), .ZN(n6758) );
  NAND2_X1 U8495 ( .A1(n6759), .A2(n6758), .ZN(n7664) );
  AOI21_X1 U8496 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7668) );
  INV_X1 U8497 ( .A(n6759), .ZN(n6760) );
  NOR2_X1 U8498 ( .A1(n7668), .A2(n6760), .ZN(n7741) );
  XNOR2_X1 U8499 ( .A(n6761), .B(n4893), .ZN(n7740) );
  NOR2_X1 U8500 ( .A1(n7741), .A2(n7740), .ZN(n7739) );
  AOI21_X1 U8501 ( .B1(n7745), .B2(n6762), .A(n7739), .ZN(n7835) );
  MUX2_X1 U8502 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6773), .Z(n6765) );
  INV_X1 U8503 ( .A(n6765), .ZN(n6764) );
  NAND2_X1 U8504 ( .A1(n6764), .A2(n6763), .ZN(n7832) );
  AND2_X1 U8505 ( .A1(n6765), .A2(n7841), .ZN(n7831) );
  AOI21_X1 U8506 ( .B1(n7835), .B2(n7832), .A(n7831), .ZN(n8745) );
  XNOR2_X1 U8507 ( .A(n6766), .B(n8754), .ZN(n8744) );
  NAND2_X1 U8508 ( .A1(n8745), .A2(n8744), .ZN(n8743) );
  OAI21_X1 U8509 ( .B1(n6766), .B2(n7075), .A(n8743), .ZN(n8762) );
  XNOR2_X1 U8510 ( .A(n6767), .B(n8767), .ZN(n8761) );
  NAND2_X1 U8511 ( .A1(n8762), .A2(n8761), .ZN(n8760) );
  OAI21_X1 U8512 ( .B1(n6767), .B2(n7238), .A(n8760), .ZN(n8779) );
  MUX2_X1 U8513 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6773), .Z(n6768) );
  XNOR2_X1 U8514 ( .A(n8785), .B(n6768), .ZN(n8778) );
  INV_X1 U8515 ( .A(n6768), .ZN(n6769) );
  AOI22_X1 U8516 ( .A1(n8779), .A2(n8778), .B1(n8785), .B2(n6769), .ZN(n8795)
         );
  MUX2_X1 U8517 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6773), .Z(n6770) );
  XNOR2_X1 U8518 ( .A(n6770), .B(n7385), .ZN(n8794) );
  OAI22_X1 U8519 ( .A1(n8795), .A2(n8794), .B1(n6770), .B2(n7385), .ZN(n8817)
         );
  MUX2_X1 U8520 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n6773), .Z(n6771) );
  XNOR2_X1 U8521 ( .A(n6771), .B(n8822), .ZN(n8818) );
  INV_X1 U8522 ( .A(n6771), .ZN(n6772) );
  AOI22_X1 U8523 ( .A1(n8817), .A2(n8818), .B1(n8822), .B2(n6772), .ZN(n6775)
         );
  MUX2_X1 U8524 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6773), .Z(n6774) );
  NAND2_X1 U8525 ( .A1(n6775), .A2(n6774), .ZN(n8827) );
  NOR2_X1 U8526 ( .A1(n6775), .A2(n6774), .ZN(n8829) );
  AOI21_X1 U8527 ( .B1(n8844), .B2(n8827), .A(n8829), .ZN(n6776) );
  XOR2_X1 U8528 ( .A(n6777), .B(n6776), .Z(n6778) );
  OR2_X1 U8529 ( .A1(n8831), .A2(n6865), .ZN(n8839) );
  NAND3_X1 U8530 ( .A1(n6780), .A2(n6779), .A3(n5145), .ZN(P2_U3201) );
  NAND2_X1 U8531 ( .A1(n6387), .A2(n6781), .ZN(n6783) );
  NAND2_X1 U8532 ( .A1(n9650), .A2(n6446), .ZN(n6782) );
  NAND2_X1 U8533 ( .A1(n6783), .A2(n6782), .ZN(n6785) );
  XNOR2_X1 U8534 ( .A(n6785), .B(n6784), .ZN(n6788) );
  AOI22_X1 U8535 ( .A1(n6387), .A2(n6446), .B1(n6786), .B2(n9650), .ZN(n6787)
         );
  XNOR2_X1 U8536 ( .A(n6788), .B(n6787), .ZN(n6797) );
  NAND3_X1 U8537 ( .A1(n6797), .A2(n9285), .A3(n6798), .ZN(n6793) );
  INV_X1 U8538 ( .A(n9209), .ZN(n9287) );
  OAI22_X1 U8539 ( .A1(n9287), .A2(n9496), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6789), .ZN(n6791) );
  INV_X1 U8540 ( .A(n8090), .ZN(n9289) );
  OAI22_X1 U8541 ( .A1(n9289), .A2(n9528), .B1(n9288), .B2(n9492), .ZN(n6790)
         );
  AOI211_X1 U8542 ( .C1(n6387), .C2(n6637), .A(n6791), .B(n6790), .ZN(n6792)
         );
  AOI21_X1 U8543 ( .B1(n6796), .B2(n6795), .A(n6794), .ZN(n6803) );
  INV_X1 U8544 ( .A(n6797), .ZN(n6800) );
  INV_X1 U8545 ( .A(n6798), .ZN(n6799) );
  NAND2_X1 U8546 ( .A1(n6801), .A2(n5149), .ZN(n6802) );
  NAND2_X1 U8547 ( .A1(n6803), .A2(n6802), .ZN(P1_U3220) );
  XNOR2_X1 U8548 ( .A(n6804), .B(n6862), .ZN(n6868) );
  INV_X1 U8549 ( .A(n6868), .ZN(n8854) );
  INV_X1 U8550 ( .A(n6805), .ZN(n6806) );
  NAND2_X1 U8551 ( .A1(n7102), .A2(n6806), .ZN(n6807) );
  NAND2_X1 U8552 ( .A1(n7805), .A2(n7878), .ZN(n10539) );
  AND2_X1 U8553 ( .A1(n6807), .A2(n10539), .ZN(n6808) );
  NAND2_X1 U8554 ( .A1(n7093), .A2(n6808), .ZN(n10451) );
  NAND2_X1 U8555 ( .A1(n8739), .A2(n8583), .ZN(n10458) );
  NAND2_X1 U8556 ( .A1(n6809), .A2(n10458), .ZN(n6813) );
  NAND2_X1 U8557 ( .A1(n6810), .A2(n6811), .ZN(n6812) );
  NAND2_X1 U8558 ( .A1(n6813), .A2(n6812), .ZN(n10439) );
  NAND2_X1 U8559 ( .A1(n10439), .A2(n10440), .ZN(n6815) );
  NAND2_X1 U8560 ( .A1(n10455), .A2(n10479), .ZN(n6814) );
  NOR2_X1 U8561 ( .A1(n8738), .A2(n7168), .ZN(n6817) );
  NAND2_X1 U8562 ( .A1(n8738), .A2(n7168), .ZN(n6816) );
  OAI21_X1 U8563 ( .B1(n7369), .B2(n6820), .A(n6818), .ZN(n7421) );
  AND2_X1 U8564 ( .A1(n6818), .A2(n10495), .ZN(n6819) );
  OR2_X1 U8565 ( .A1(n6821), .A2(n7394), .ZN(n6822) );
  AND2_X1 U8566 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  AND2_X1 U8567 ( .A1(n8737), .A2(n10505), .ZN(n6826) );
  NOR2_X1 U8568 ( .A1(n9036), .A2(n8592), .ZN(n6828) );
  NAND2_X1 U8569 ( .A1(n9036), .A2(n8592), .ZN(n6827) );
  NAND2_X1 U8570 ( .A1(n10513), .A2(n8736), .ZN(n6829) );
  NAND2_X1 U8571 ( .A1(n6830), .A2(n6829), .ZN(n7712) );
  AND2_X1 U8572 ( .A1(n10518), .A2(n8735), .ZN(n6831) );
  OAI22_X1 U8573 ( .A1(n7712), .A2(n6831), .B1(n8735), .B2(n10518), .ZN(n7779)
         );
  NOR2_X1 U8574 ( .A1(n7788), .A2(n8734), .ZN(n6833) );
  NAND2_X1 U8575 ( .A1(n7788), .A2(n8734), .ZN(n6832) );
  OAI21_X1 U8576 ( .B1(n7779), .B2(n6833), .A(n6832), .ZN(n7818) );
  NAND2_X1 U8577 ( .A1(n7818), .A2(n7817), .ZN(n6835) );
  INV_X1 U8578 ( .A(n7921), .ZN(n8733) );
  NAND2_X1 U8579 ( .A1(n10536), .A2(n8733), .ZN(n6834) );
  NAND2_X1 U8580 ( .A1(n6835), .A2(n6834), .ZN(n7919) );
  AND2_X1 U8581 ( .A1(n7863), .A2(n8732), .ZN(n7967) );
  OR2_X1 U8582 ( .A1(n7967), .A2(n5147), .ZN(n8068) );
  AND2_X1 U8583 ( .A1(n8078), .A2(n8730), .ZN(n6839) );
  OR2_X1 U8584 ( .A1(n8078), .A2(n8730), .ZN(n6837) );
  OR2_X1 U8585 ( .A1(n7863), .A2(n8732), .ZN(n7969) );
  AND2_X1 U8586 ( .A1(n6836), .A2(n7969), .ZN(n7968) );
  OR2_X1 U8587 ( .A1(n5147), .A2(n7968), .ZN(n8069) );
  AND2_X1 U8588 ( .A1(n6837), .A2(n8069), .ZN(n6838) );
  AND2_X1 U8589 ( .A1(n9012), .A2(n9017), .ZN(n9013) );
  INV_X1 U8590 ( .A(n8718), .ZN(n9004) );
  NAND2_X1 U8591 ( .A1(n9158), .A2(n9004), .ZN(n6842) );
  NAND2_X1 U8592 ( .A1(n9002), .A2(n9001), .ZN(n9000) );
  INV_X1 U8593 ( .A(n8638), .ZN(n9018) );
  NAND2_X1 U8594 ( .A1(n9151), .A2(n9018), .ZN(n6843) );
  NAND2_X1 U8595 ( .A1(n4543), .A2(n8996), .ZN(n8987) );
  INV_X1 U8596 ( .A(n8977), .ZN(n9003) );
  OR2_X1 U8597 ( .A1(n8994), .A2(n9003), .ZN(n8972) );
  AND2_X1 U8598 ( .A1(n6845), .A2(n8972), .ZN(n6846) );
  NAND2_X1 U8599 ( .A1(n8987), .A2(n6846), .ZN(n8975) );
  INV_X1 U8600 ( .A(n8697), .ZN(n8988) );
  NAND2_X1 U8601 ( .A1(n8984), .A2(n8988), .ZN(n6847) );
  INV_X1 U8602 ( .A(n9138), .ZN(n8681) );
  NAND2_X1 U8603 ( .A1(n8681), .A2(n8978), .ZN(n6848) );
  INV_X1 U8604 ( .A(n8932), .ZN(n8963) );
  OR2_X1 U8605 ( .A1(n9072), .A2(n8963), .ZN(n6849) );
  NAND2_X1 U8606 ( .A1(n6850), .A2(n6849), .ZN(n8930) );
  NAND2_X1 U8607 ( .A1(n8930), .A2(n8938), .ZN(n6852) );
  INV_X1 U8608 ( .A(n8951), .ZN(n8924) );
  OR2_X1 U8609 ( .A1(n8940), .A2(n8924), .ZN(n6851) );
  NAND2_X1 U8610 ( .A1(n6852), .A2(n6851), .ZN(n8921) );
  NOR2_X1 U8611 ( .A1(n9124), .A2(n8908), .ZN(n6854) );
  NAND2_X1 U8612 ( .A1(n9124), .A2(n8908), .ZN(n6853) );
  AND2_X1 U8613 ( .A1(n9118), .A2(n8923), .ZN(n6856) );
  OR2_X1 U8614 ( .A1(n9118), .A2(n8923), .ZN(n6855) );
  NAND2_X1 U8615 ( .A1(n8566), .A2(n8526), .ZN(n6857) );
  AOI21_X1 U8616 ( .B1(n8602), .B2(n9103), .A(n8861), .ZN(n6861) );
  NOR2_X1 U8617 ( .A1(n6861), .A2(n6860), .ZN(n6863) );
  NAND2_X1 U8618 ( .A1(n7376), .A2(n6887), .ZN(n6901) );
  XNOR2_X1 U8619 ( .A(n6865), .B(n6864), .ZN(n7099) );
  INV_X1 U8620 ( .A(n7099), .ZN(n7095) );
  NAND2_X1 U8621 ( .A1(n7099), .A2(n6884), .ZN(n10454) );
  AOI21_X1 U8622 ( .B1(P2_B_REG_SCAN_IN), .B2(n6866), .A(n10454), .ZN(n8848)
         );
  AOI22_X1 U8623 ( .A1(n10425), .A2(n8727), .B1(n8726), .B2(n8848), .ZN(n6867)
         );
  AND3_X1 U8624 ( .A1(n7376), .A2(n7878), .A3(n7722), .ZN(n10474) );
  XNOR2_X1 U8625 ( .A(n7996), .B(P2_B_REG_SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8626 ( .A1(n6885), .A2(n6870), .ZN(n6872) );
  NOR2_X1 U8627 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6876) );
  NOR4_X1 U8628 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6875) );
  NOR4_X1 U8629 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6874) );
  NOR4_X1 U8630 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6873) );
  NAND4_X1 U8631 ( .A1(n6876), .A2(n6875), .A3(n6874), .A4(n6873), .ZN(n6882)
         );
  NOR4_X1 U8632 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6880) );
  NOR4_X1 U8633 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6879) );
  NOR4_X1 U8634 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6878) );
  NOR4_X1 U8635 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6877) );
  NAND4_X1 U8636 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6881)
         );
  NOR2_X1 U8637 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  OR2_X1 U8638 ( .A1(n6889), .A2(n6883), .ZN(n6904) );
  NAND2_X1 U8639 ( .A1(n6884), .A2(n7102), .ZN(n7082) );
  NAND3_X1 U8640 ( .A1(n6904), .A2(n7097), .A3(n7082), .ZN(n7196) );
  AND2_X1 U8641 ( .A1(n10474), .A2(n7805), .ZN(n7096) );
  NOR2_X1 U8642 ( .A1(n7196), .A2(n7096), .ZN(n6894) );
  OR2_X1 U8643 ( .A1(n6889), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8644 ( .A1(n6885), .A2(n8099), .ZN(n6974) );
  NAND2_X1 U8645 ( .A1(n6886), .A2(n6974), .ZN(n7195) );
  NAND3_X1 U8646 ( .A1(n7660), .A2(n6887), .A3(n6900), .ZN(n6888) );
  AND2_X1 U8647 ( .A1(n5873), .A2(n6888), .ZN(n6890) );
  OR2_X1 U8648 ( .A1(n7195), .A2(n6890), .ZN(n6893) );
  NAND2_X1 U8649 ( .A1(n8099), .A2(n7996), .ZN(n6977) );
  OAI21_X1 U8650 ( .B1(n6889), .B2(P2_D_REG_0__SCAN_IN), .A(n6977), .ZN(n7104)
         );
  INV_X1 U8651 ( .A(n6890), .ZN(n6891) );
  OR2_X1 U8652 ( .A1(n7104), .A2(n6891), .ZN(n6892) );
  NAND2_X1 U8653 ( .A1(n6893), .A2(n6892), .ZN(n7194) );
  OR2_X1 U8654 ( .A1(n7195), .A2(n7104), .ZN(n6899) );
  AND3_X2 U8655 ( .A1(n6894), .A2(n7194), .A3(n6899), .ZN(n10570) );
  INV_X1 U8656 ( .A(n10539), .ZN(n10537) );
  NAND2_X1 U8657 ( .A1(n10570), .A2(n10537), .ZN(n9078) );
  NAND2_X1 U8658 ( .A1(n6897), .A2(n5136), .ZN(P2_U3488) );
  INV_X1 U8659 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6910) );
  INV_X1 U8660 ( .A(n6904), .ZN(n6898) );
  NOR2_X1 U8661 ( .A1(n6899), .A2(n6898), .ZN(n7086) );
  NAND2_X1 U8662 ( .A1(n7086), .A2(n7097), .ZN(n7118) );
  INV_X1 U8663 ( .A(n6901), .ZN(n6902) );
  NAND2_X1 U8664 ( .A1(n7105), .A2(n6902), .ZN(n7080) );
  AND2_X1 U8665 ( .A1(n7093), .A2(n7080), .ZN(n6903) );
  OR2_X1 U8666 ( .A1(n7118), .A2(n6903), .ZN(n6908) );
  NAND3_X1 U8667 ( .A1(n7195), .A2(n7104), .A3(n6904), .ZN(n7089) );
  INV_X1 U8668 ( .A(n7097), .ZN(n6905) );
  OR2_X1 U8669 ( .A1(n7089), .A2(n6905), .ZN(n7094) );
  INV_X1 U8670 ( .A(n7094), .ZN(n7120) );
  NAND3_X1 U8671 ( .A1(n5873), .A2(n7080), .A3(n10539), .ZN(n7117) );
  NAND2_X1 U8672 ( .A1(n10537), .A2(n6906), .ZN(n10438) );
  NAND2_X1 U8673 ( .A1(n7117), .A2(n10438), .ZN(n7079) );
  NAND2_X1 U8674 ( .A1(n7120), .A2(n7079), .ZN(n6907) );
  INV_X2 U8675 ( .A(n10547), .ZN(n10545) );
  NAND2_X1 U8676 ( .A1(n10545), .A2(n10537), .ZN(n9143) );
  NAND2_X1 U8677 ( .A1(n6911), .A2(n5140), .ZN(P2_U3456) );
  INV_X1 U8678 ( .A(n8831), .ZN(P2_U3893) );
  INV_X1 U8679 ( .A(n6912), .ZN(n6913) );
  OR2_X2 U8680 ( .A1(n6437), .A2(n6913), .ZN(n9309) );
  INV_X1 U8681 ( .A(n9309), .ZN(P1_U3973) );
  XNOR2_X1 U8682 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8683 ( .A1(n8151), .A2(P1_U3086), .ZN(n8143) );
  AND2_X1 U8684 ( .A1(n6914), .A2(P1_U3086), .ZN(n7888) );
  INV_X2 U8685 ( .A(n7888), .ZN(n9758) );
  OAI222_X1 U8686 ( .A1(n9754), .A2(n4668), .B1(n7055), .B2(P1_U3086), .C1(
        n9758), .C2(n6927), .ZN(P1_U3351) );
  OAI222_X1 U8687 ( .A1(n9754), .A2(n6915), .B1(n7043), .B2(P1_U3086), .C1(
        n9758), .C2(n6948), .ZN(P1_U3353) );
  OAI222_X1 U8688 ( .A1(n9754), .A2(n4709), .B1(n8224), .B2(P1_U3086), .C1(
        n9758), .C2(n6928), .ZN(P1_U3352) );
  OAI222_X1 U8689 ( .A1(n9754), .A2(n6916), .B1(n9315), .B2(P1_U3086), .C1(
        n9758), .C2(n6936), .ZN(P1_U3354) );
  OAI222_X1 U8690 ( .A1(n9754), .A2(n6917), .B1(n9326), .B2(P1_U3086), .C1(
        n9758), .C2(n6931), .ZN(P1_U3350) );
  AOI22_X1 U8691 ( .A1(n9344), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n8143), .ZN(n6918) );
  OAI21_X1 U8692 ( .B1(n6934), .B2(n9758), .A(n6918), .ZN(P1_U3349) );
  INV_X1 U8693 ( .A(n6922), .ZN(n7889) );
  OR2_X1 U8694 ( .A1(n6437), .A2(n7889), .ZN(n6919) );
  NAND2_X1 U8695 ( .A1(n6919), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6941) );
  INV_X1 U8696 ( .A(n6941), .ZN(n6924) );
  NAND2_X1 U8697 ( .A1(n6922), .A2(n6921), .ZN(n6923) );
  NAND2_X1 U8698 ( .A1(n6045), .A2(n6923), .ZN(n6940) );
  AND2_X1 U8699 ( .A1(n6924), .A2(n6940), .ZN(n9467) );
  NOR2_X1 U8700 ( .A1(n9467), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8701 ( .A(n7127), .ZN(n7138) );
  INV_X1 U8702 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9921) );
  OAI222_X1 U8703 ( .A1(n9758), .A2(n6926), .B1(n7138), .B2(P1_U3086), .C1(
        n9921), .C2(n9754), .ZN(P1_U3348) );
  NAND2_X1 U8704 ( .A1(n8151), .A2(P2_U3151), .ZN(n8098) );
  NOR2_X1 U8705 ( .A1(n8151), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8149) );
  OAI222_X1 U8706 ( .A1(P2_U3151), .A2(n7363), .B1(n8098), .B2(n6926), .C1(
        n6925), .C2(n9167), .ZN(P2_U3288) );
  INV_X1 U8707 ( .A(n8098), .ZN(n7892) );
  INV_X1 U8708 ( .A(n7892), .ZN(n9164) );
  OAI222_X1 U8709 ( .A1(P2_U3151), .A2(n7261), .B1(n9164), .B2(n6927), .C1(
        n5173), .C2(n9167), .ZN(P2_U3291) );
  OAI222_X1 U8710 ( .A1(P2_U3151), .A2(n6929), .B1(n9164), .B2(n6928), .C1(
        n5169), .C2(n9167), .ZN(P2_U3292) );
  OAI222_X1 U8711 ( .A1(P2_U3151), .A2(n6932), .B1(n9164), .B2(n6931), .C1(
        n6930), .C2(n9167), .ZN(P2_U3290) );
  OAI222_X1 U8712 ( .A1(P2_U3151), .A2(n6935), .B1(n9164), .B2(n6934), .C1(
        n6933), .C2(n9167), .ZN(P2_U3289) );
  OAI222_X1 U8713 ( .A1(n7263), .A2(P2_U3151), .B1(n9167), .B2(n6937), .C1(
        n9164), .C2(n6936), .ZN(P2_U3294) );
  INV_X1 U8714 ( .A(n6326), .ZN(n7036) );
  INV_X1 U8715 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9318) );
  NOR2_X1 U8716 ( .A1(n6326), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8717 ( .B1(n7036), .B2(P1_REG1_REG_0__SCAN_IN), .A(n5141), .ZN(
        n6939) );
  MUX2_X1 U8718 ( .A(n6939), .B(n5141), .S(P1_IR_REG_0__SCAN_IN), .Z(n6945) );
  NOR2_X1 U8719 ( .A1(n6941), .A2(n6940), .ZN(n7000) );
  INV_X1 U8720 ( .A(n7000), .ZN(n6944) );
  AND2_X1 U8721 ( .A1(n7000), .A2(n6326), .ZN(n9435) );
  NAND3_X1 U8722 ( .A1(n9435), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9318), .ZN(
        n6943) );
  AOI22_X1 U8723 ( .A1(n9467), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6942) );
  OAI211_X1 U8724 ( .C1(n6945), .C2(n6944), .A(n6943), .B(n6942), .ZN(P1_U3243) );
  INV_X1 U8725 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8726 ( .A1(n7032), .A2(P1_U3973), .ZN(n6946) );
  OAI21_X1 U8727 ( .B1(P1_U3973), .B2(n6947), .A(n6946), .ZN(P1_U3554) );
  OAI222_X1 U8728 ( .A1(P2_U3151), .A2(n6949), .B1(n9164), .B2(n6948), .C1(
        n5156), .C2(n9167), .ZN(P2_U3293) );
  INV_X1 U8729 ( .A(n6950), .ZN(n6953) );
  OAI222_X1 U8730 ( .A1(n6952), .A2(P2_U3151), .B1(n9164), .B2(n6953), .C1(
        n6951), .C2(n9167), .ZN(P2_U3287) );
  INV_X1 U8731 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6954) );
  INV_X1 U8732 ( .A(n7216), .ZN(n7133) );
  OAI222_X1 U8733 ( .A1(n9754), .A2(n6954), .B1(n9758), .B2(n6953), .C1(
        P1_U3086), .C2(n7133), .ZN(P1_U3347) );
  NAND2_X1 U8734 ( .A1(n7097), .A2(n6889), .ZN(n6973) );
  AND2_X1 U8735 ( .A1(n6973), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8736 ( .A1(n6973), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8737 ( .A1(n6973), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8738 ( .A1(n6973), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8739 ( .A1(n6973), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8740 ( .A1(n6973), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8741 ( .A1(n6973), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8742 ( .A1(n6973), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8743 ( .A1(n6973), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8744 ( .A1(n6973), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8745 ( .A1(n6973), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8746 ( .A1(n6973), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8747 ( .A1(n6973), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  INV_X1 U8748 ( .A(n7433), .ZN(n7439) );
  INV_X1 U8749 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9938) );
  OAI222_X1 U8750 ( .A1(n9758), .A2(n6958), .B1(n7439), .B2(P1_U3086), .C1(
        n9938), .C2(n9754), .ZN(P1_U3345) );
  INV_X1 U8751 ( .A(n6955), .ZN(n6961) );
  INV_X1 U8752 ( .A(n7339), .ZN(n7209) );
  INV_X1 U8753 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6956) );
  OAI222_X1 U8754 ( .A1(n9758), .A2(n6961), .B1(n7209), .B2(P1_U3086), .C1(
        n6956), .C2(n9754), .ZN(P1_U3346) );
  INV_X1 U8755 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6957) );
  OAI222_X1 U8756 ( .A1(P2_U3151), .A2(n6959), .B1(n8098), .B2(n6958), .C1(
        n6957), .C2(n9167), .ZN(P2_U3285) );
  INV_X1 U8757 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6960) );
  OAI222_X1 U8758 ( .A1(P2_U3151), .A2(n6962), .B1(n8098), .B2(n6961), .C1(
        n6960), .C2(n9167), .ZN(P2_U3286) );
  INV_X1 U8759 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6964) );
  INV_X1 U8760 ( .A(n6963), .ZN(n6966) );
  INV_X1 U8761 ( .A(n8187), .ZN(n8174) );
  OAI222_X1 U8762 ( .A1(n9754), .A2(n6964), .B1(n9758), .B2(n6966), .C1(
        P1_U3086), .C2(n8174), .ZN(P1_U3344) );
  INV_X1 U8763 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6965) );
  OAI222_X1 U8764 ( .A1(n4893), .A2(P2_U3151), .B1(n8098), .B2(n6966), .C1(
        n6965), .C2(n9167), .ZN(P2_U3284) );
  NAND2_X1 U8765 ( .A1(n7032), .A2(n10274), .ZN(n8440) );
  NAND2_X1 U8766 ( .A1(n10266), .A2(n8440), .ZN(n8365) );
  INV_X1 U8767 ( .A(n8365), .ZN(n7573) );
  NOR2_X1 U8768 ( .A1(n10385), .A2(n10250), .ZN(n6967) );
  OAI222_X1 U8769 ( .A1(n10274), .A2(n6968), .B1(n7573), .B2(n6967), .C1(
        n10356), .C2(n7068), .ZN(n6970) );
  NAND2_X1 U8770 ( .A1(n6970), .A2(n10413), .ZN(n6969) );
  OAI21_X1 U8771 ( .B1(n10413), .B2(n9318), .A(n6969), .ZN(P1_U3522) );
  INV_X1 U8772 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8773 ( .A1(n6970), .A2(n10395), .ZN(n6971) );
  OAI21_X1 U8774 ( .B1(n10395), .B2(n6972), .A(n6971), .ZN(P1_U3453) );
  INV_X1 U8775 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6976) );
  INV_X1 U8776 ( .A(n6974), .ZN(n6975) );
  AOI22_X1 U8777 ( .A1(n6973), .A2(n6976), .B1(n6979), .B2(n6975), .ZN(
        P2_U3377) );
  INV_X1 U8778 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6980) );
  INV_X1 U8779 ( .A(n6977), .ZN(n6978) );
  AOI22_X1 U8780 ( .A1(n6973), .A2(n6980), .B1(n6979), .B2(n6978), .ZN(
        P2_U3376) );
  AND2_X1 U8781 ( .A1(n6973), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8782 ( .A1(n6973), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8783 ( .A1(n6973), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8784 ( .A1(n6973), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8785 ( .A1(n6973), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8786 ( .A1(n6973), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8787 ( .A1(n6973), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8788 ( .A1(n6973), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8789 ( .A1(n6973), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8790 ( .A1(n6973), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8791 ( .A1(n6973), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8792 ( .A1(n6973), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8793 ( .A1(n6973), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8794 ( .A1(n6973), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8795 ( .A1(n6973), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8796 ( .A1(n6973), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8797 ( .A1(n6973), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AOI22_X1 U8798 ( .A1(n8188), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n8143), .ZN(n6981) );
  OAI21_X1 U8799 ( .B1(n7024), .B2(n9758), .A(n6981), .ZN(P1_U3343) );
  AOI21_X1 U8800 ( .B1(n6984), .B2(n6983), .A(n6982), .ZN(n7037) );
  NAND2_X1 U8801 ( .A1(n7037), .A2(n9285), .ZN(n6987) );
  NAND2_X1 U8802 ( .A1(n6985), .A2(n7466), .ZN(n7069) );
  AOI22_X1 U8803 ( .A1(n6637), .A2(n6440), .B1(n7069), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6986) );
  OAI211_X1 U8804 ( .C1(n7068), .C2(n9287), .A(n6987), .B(n6986), .ZN(P1_U3232) );
  INV_X1 U8805 ( .A(n8224), .ZN(n6993) );
  INV_X1 U8806 ( .A(n7043), .ZN(n6990) );
  INV_X1 U8807 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10260) );
  MUX2_X1 U8808 ( .A(n10260), .B(P1_REG2_REG_2__SCAN_IN), .S(n7043), .Z(n7045)
         );
  INV_X1 U8809 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6988) );
  MUX2_X1 U8810 ( .A(n6988), .B(P1_REG2_REG_1__SCAN_IN), .S(n9315), .Z(n9313)
         );
  AND2_X1 U8811 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9312) );
  NAND2_X1 U8812 ( .A1(n9313), .A2(n9312), .ZN(n9311) );
  INV_X1 U8813 ( .A(n9315), .ZN(n9314) );
  NAND2_X1 U8814 ( .A1(n9314), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U8815 ( .A1(n9311), .A2(n6989), .ZN(n7044) );
  INV_X1 U8816 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6991) );
  MUX2_X1 U8817 ( .A(n6991), .B(P1_REG2_REG_3__SCAN_IN), .S(n8224), .Z(n6992)
         );
  INV_X1 U8818 ( .A(n6992), .ZN(n8217) );
  NAND2_X1 U8819 ( .A1(n7013), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6994) );
  OAI21_X1 U8820 ( .B1(n7013), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6994), .ZN(
        n7057) );
  NOR2_X1 U8821 ( .A1(n7058), .A2(n7057), .ZN(n7056) );
  AOI21_X1 U8822 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n7013), .A(n7056), .ZN(
        n9331) );
  NAND2_X1 U8823 ( .A1(n7006), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U8824 ( .B1(n7006), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6995), .ZN(
        n9330) );
  NAND2_X1 U8825 ( .A1(n9344), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6996) );
  OAI21_X1 U8826 ( .B1(n9344), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6996), .ZN(
        n9340) );
  XNOR2_X1 U8827 ( .A(n7127), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8828 ( .A1(n6998), .A2(n6999), .ZN(n7126) );
  AND2_X1 U8829 ( .A1(n6997), .A2(n7036), .ZN(n8516) );
  NAND2_X1 U8830 ( .A1(n7000), .A2(n8516), .ZN(n9458) );
  AOI211_X1 U8831 ( .C1(n6999), .C2(n6998), .A(n7126), .B(n9458), .ZN(n7004)
         );
  NAND2_X1 U8832 ( .A1(n7000), .A2(n4524), .ZN(n9447) );
  NAND2_X1 U8833 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7581) );
  INV_X1 U8834 ( .A(n7581), .ZN(n7001) );
  AOI21_X1 U8835 ( .B1(n9467), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7001), .ZN(
        n7002) );
  OAI21_X1 U8836 ( .B1(n9447), .B2(n7138), .A(n7002), .ZN(n7003) );
  NOR2_X1 U8837 ( .A1(n7004), .A2(n7003), .ZN(n7022) );
  NAND2_X1 U8838 ( .A1(n9344), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7018) );
  MUX2_X1 U8839 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7005), .S(n9344), .Z(n9346)
         );
  NAND2_X1 U8840 ( .A1(n7006), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U8841 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7007), .S(n7006), .Z(n9334)
         );
  NAND2_X1 U8842 ( .A1(n7013), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7016) );
  INV_X1 U8843 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10399) );
  INV_X1 U8844 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10397) );
  MUX2_X1 U8845 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10397), .S(n7043), .Z(n7040)
         );
  INV_X1 U8846 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7008) );
  MUX2_X1 U8847 ( .A(n7008), .B(P1_REG1_REG_1__SCAN_IN), .S(n9315), .Z(n7010)
         );
  AND2_X1 U8848 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7009) );
  NAND2_X1 U8849 ( .A1(n7010), .A2(n7009), .ZN(n9320) );
  OR2_X1 U8850 ( .A1(n9315), .A2(n7008), .ZN(n7011) );
  AND2_X1 U8851 ( .A1(n9320), .A2(n7011), .ZN(n7041) );
  OAI22_X1 U8852 ( .A1(n7040), .A2(n7041), .B1(n10397), .B2(n7043), .ZN(n8211)
         );
  MUX2_X1 U8853 ( .A(n10399), .B(P1_REG1_REG_3__SCAN_IN), .S(n8224), .Z(n7012)
         );
  NAND2_X1 U8854 ( .A1(n8211), .A2(n7012), .ZN(n8212) );
  OAI21_X1 U8855 ( .B1(n10399), .B2(n8224), .A(n8212), .ZN(n7053) );
  MUX2_X1 U8856 ( .A(n6020), .B(P1_REG1_REG_4__SCAN_IN), .S(n7013), .Z(n7052)
         );
  INV_X1 U8857 ( .A(n7052), .ZN(n7014) );
  NAND2_X1 U8858 ( .A1(n7053), .A2(n7014), .ZN(n7015) );
  NAND2_X1 U8859 ( .A1(n7016), .A2(n7015), .ZN(n9335) );
  NAND2_X1 U8860 ( .A1(n9334), .A2(n9335), .ZN(n9333) );
  NAND2_X1 U8861 ( .A1(n7017), .A2(n9333), .ZN(n9347) );
  NAND2_X1 U8862 ( .A1(n9346), .A2(n9347), .ZN(n9345) );
  NAND2_X1 U8863 ( .A1(n7018), .A2(n9345), .ZN(n7020) );
  MUX2_X1 U8864 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7137), .S(n7127), .Z(n7019)
         );
  NAND2_X1 U8865 ( .A1(n7020), .A2(n7019), .ZN(n7136) );
  OAI211_X1 U8866 ( .C1(n7020), .C2(n7019), .A(n7136), .B(n9435), .ZN(n7021)
         );
  NAND2_X1 U8867 ( .A1(n7022), .A2(n7021), .ZN(P1_U3250) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7023) );
  OAI222_X1 U8869 ( .A1(P2_U3151), .A2(n7841), .B1(n8098), .B2(n7024), .C1(
        n7023), .C2(n9167), .ZN(P2_U3283) );
  INV_X1 U8870 ( .A(n7025), .ZN(n7027) );
  NAND2_X1 U8871 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  XNOR2_X1 U8872 ( .A(n7029), .B(n7028), .ZN(n7035) );
  INV_X1 U8873 ( .A(n9285), .ZN(n9277) );
  NAND2_X1 U8874 ( .A1(n9308), .A2(n10371), .ZN(n10264) );
  INV_X1 U8875 ( .A(n10264), .ZN(n7031) );
  AOI22_X1 U8876 ( .A1(n7031), .A2(n7030), .B1(n6637), .B2(n10276), .ZN(n7034)
         );
  AOI22_X1 U8877 ( .A1(n8090), .A2(n7032), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7069), .ZN(n7033) );
  OAI211_X1 U8878 ( .C1(n7035), .C2(n9277), .A(n7034), .B(n7033), .ZN(P1_U3222) );
  OR3_X1 U8879 ( .A1(n7037), .A2(n4524), .A3(n7036), .ZN(n7039) );
  AOI21_X1 U8880 ( .B1(n8516), .B2(n9312), .A(n9309), .ZN(n7038) );
  OAI211_X1 U8881 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n5141), .A(n7039), .B(n7038), .ZN(n7063) );
  XOR2_X1 U8882 ( .A(n7041), .B(n7040), .Z(n7050) );
  AOI22_X1 U8883 ( .A1(n9467), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7042) );
  OAI21_X1 U8884 ( .B1(n7043), .B2(n9447), .A(n7042), .ZN(n7049) );
  NOR2_X1 U8885 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  NOR3_X1 U8886 ( .A1(n9458), .A2(n7047), .A3(n7046), .ZN(n7048) );
  AOI211_X1 U8887 ( .C1(n9435), .C2(n7050), .A(n7049), .B(n7048), .ZN(n7051)
         );
  NAND2_X1 U8888 ( .A1(n7063), .A2(n7051), .ZN(P1_U3245) );
  XNOR2_X1 U8889 ( .A(n7053), .B(n7052), .ZN(n7061) );
  AND2_X1 U8890 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9240) );
  AOI21_X1 U8891 ( .B1(n9467), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9240), .ZN(
        n7054) );
  OAI21_X1 U8892 ( .B1(n9447), .B2(n7055), .A(n7054), .ZN(n7060) );
  AOI211_X1 U8893 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n9458), .ZN(n7059)
         );
  AOI211_X1 U8894 ( .C1(n9435), .C2(n7061), .A(n7060), .B(n7059), .ZN(n7062)
         );
  NAND2_X1 U8895 ( .A1(n7063), .A2(n7062), .ZN(P1_U3247) );
  AOI21_X1 U8896 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7072) );
  OAI22_X1 U8897 ( .A1(n7068), .A2(n10358), .B1(n7067), .B2(n10356), .ZN(
        n10249) );
  AOI22_X1 U8898 ( .A1(n10249), .A2(n9241), .B1(n10253), .B2(n6637), .ZN(n7071) );
  NAND2_X1 U8899 ( .A1(n7069), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7070) );
  OAI211_X1 U8900 ( .C1(n7072), .C2(n9277), .A(n7071), .B(n7070), .ZN(P1_U3237) );
  INV_X1 U8901 ( .A(n8189), .ZN(n9353) );
  INV_X1 U8902 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10089) );
  OAI222_X1 U8903 ( .A1(n9758), .A2(n7074), .B1(n9353), .B2(P1_U3086), .C1(
        n10089), .C2(n9754), .ZN(P1_U3342) );
  INV_X1 U8904 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7073) );
  OAI222_X1 U8905 ( .A1(P2_U3151), .A2(n7075), .B1(n8098), .B2(n7074), .C1(
        n7073), .C2(n9167), .ZN(P2_U3282) );
  INV_X1 U8906 ( .A(n10474), .ZN(n10527) );
  NAND2_X1 U8907 ( .A1(n10451), .A2(n10527), .ZN(n10544) );
  OAI21_X1 U8908 ( .B1(n10544), .B2(n10443), .A(n8584), .ZN(n7077) );
  NOR2_X1 U8909 ( .A1(n6810), .A2(n10454), .ZN(n7203) );
  INV_X1 U8910 ( .A(n7203), .ZN(n7076) );
  OAI211_X1 U8911 ( .C1(n7208), .C2(n10539), .A(n7077), .B(n7076), .ZN(n7153)
         );
  NAND2_X1 U8912 ( .A1(n7153), .A2(n10570), .ZN(n7078) );
  OAI21_X1 U8913 ( .B1(n10570), .B2(n6734), .A(n7078), .ZN(P2_U3459) );
  INV_X1 U8914 ( .A(n7079), .ZN(n7085) );
  INV_X1 U8915 ( .A(n7080), .ZN(n7119) );
  NAND2_X1 U8916 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  AOI21_X1 U8917 ( .B1(n7089), .B2(n7119), .A(n7083), .ZN(n7084) );
  OAI21_X1 U8918 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7087) );
  NAND2_X1 U8919 ( .A1(n7087), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7091) );
  NAND2_X1 U8920 ( .A1(n7089), .A2(n7088), .ZN(n7090) );
  NAND2_X1 U8921 ( .A1(n7091), .A2(n7090), .ZN(n7157) );
  NOR2_X1 U8922 ( .A1(n7157), .A2(n7092), .ZN(n8581) );
  INV_X1 U8923 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10465) );
  NOR2_X1 U8924 ( .A1(n7094), .A2(n7093), .ZN(n7100) );
  OR2_X1 U8925 ( .A1(n7118), .A2(n10539), .ZN(n7098) );
  NAND2_X1 U8926 ( .A1(n7097), .A2(n7096), .ZN(n10464) );
  NAND2_X1 U8927 ( .A1(n7098), .A2(n10464), .ZN(n8707) );
  INV_X1 U8928 ( .A(n8707), .ZN(n8724) );
  NAND2_X1 U8929 ( .A1(n7100), .A2(n7099), .ZN(n8717) );
  OAI22_X1 U8930 ( .A1(n8724), .A2(n6811), .B1(n10455), .B2(n8717), .ZN(n7101)
         );
  AOI21_X1 U8931 ( .B1(n8715), .B2(n8739), .A(n7101), .ZN(n7125) );
  INV_X1 U8932 ( .A(n7102), .ZN(n7103) );
  INV_X1 U8933 ( .A(n7104), .ZN(n7106) );
  NAND2_X4 U8934 ( .A1(n7108), .A2(n7107), .ZN(n8569) );
  XNOR2_X1 U8935 ( .A(n8569), .B(n10473), .ZN(n7111) );
  INV_X1 U8936 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U8937 ( .A1(n7110), .A2(n7109), .ZN(n7112) );
  NAND2_X1 U8938 ( .A1(n7111), .A2(n6810), .ZN(n7145) );
  NAND2_X1 U8939 ( .A1(n7208), .A2(n8556), .ZN(n7113) );
  NAND2_X1 U8940 ( .A1(n7114), .A2(n7113), .ZN(n7115) );
  NAND2_X1 U8941 ( .A1(n7116), .A2(n7115), .ZN(n7146) );
  OAI21_X1 U8942 ( .B1(n7116), .B2(n7115), .A(n7146), .ZN(n7123) );
  OR2_X1 U8943 ( .A1(n7118), .A2(n7117), .ZN(n7122) );
  NAND2_X1 U8944 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  NAND2_X1 U8945 ( .A1(n7123), .A2(n8693), .ZN(n7124) );
  OAI211_X1 U8946 ( .C1(n8581), .C2(n10465), .A(n7125), .B(n7124), .ZN(
        P2_U3162) );
  NAND2_X1 U8947 ( .A1(n7216), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7128) );
  OAI21_X1 U8948 ( .B1(n7216), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7128), .ZN(
        n7129) );
  AOI211_X1 U8949 ( .C1(n7130), .C2(n7129), .A(n7215), .B(n9458), .ZN(n7135)
         );
  AND2_X1 U8950 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7131) );
  AOI21_X1 U8951 ( .B1(n9467), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7131), .ZN(
        n7132) );
  OAI21_X1 U8952 ( .B1(n9447), .B2(n7133), .A(n7132), .ZN(n7134) );
  NOR2_X1 U8953 ( .A1(n7135), .A2(n7134), .ZN(n7143) );
  OAI21_X1 U8954 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7141) );
  MUX2_X1 U8955 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7139), .S(n7216), .Z(n7140)
         );
  NAND2_X1 U8956 ( .A1(n7140), .A2(n7141), .ZN(n7210) );
  OAI211_X1 U8957 ( .C1(n7141), .C2(n7140), .A(n9435), .B(n7210), .ZN(n7142)
         );
  NAND2_X1 U8958 ( .A1(n7143), .A2(n7142), .ZN(P1_U3251) );
  INV_X1 U8959 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10437) );
  XNOR2_X1 U8960 ( .A(n8569), .B(n7144), .ZN(n7158) );
  XNOR2_X1 U8961 ( .A(n7158), .B(n10426), .ZN(n7148) );
  NAND2_X1 U8962 ( .A1(n7146), .A2(n7145), .ZN(n7147) );
  NAND2_X1 U8963 ( .A1(n7147), .A2(n7148), .ZN(n7163) );
  OAI21_X1 U8964 ( .B1(n7148), .B2(n7147), .A(n7163), .ZN(n7149) );
  NAND2_X1 U8965 ( .A1(n7149), .A2(n8693), .ZN(n7152) );
  OAI22_X1 U8966 ( .A1(n8724), .A2(n10479), .B1(n10441), .B2(n8717), .ZN(n7150) );
  AOI21_X1 U8967 ( .B1(n8715), .B2(n7109), .A(n7150), .ZN(n7151) );
  OAI211_X1 U8968 ( .C1(n8581), .C2(n10437), .A(n7152), .B(n7151), .ZN(
        P2_U3177) );
  INV_X1 U8969 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8970 ( .A1(n10545), .A2(n7153), .ZN(n7154) );
  OAI21_X1 U8971 ( .B1(n10545), .B2(n7155), .A(n7154), .ZN(P2_U3390) );
  INV_X1 U8972 ( .A(n7894), .ZN(n7156) );
  INV_X1 U8973 ( .A(n8720), .ZN(n7775) );
  NAND2_X1 U8974 ( .A1(n7158), .A2(n10455), .ZN(n7160) );
  NAND2_X1 U8975 ( .A1(n7163), .A2(n7160), .ZN(n7159) );
  XNOR2_X1 U8976 ( .A(n7315), .B(n10441), .ZN(n7162) );
  AOI21_X1 U8977 ( .B1(n7159), .B2(n7162), .A(n8711), .ZN(n7165) );
  INV_X1 U8978 ( .A(n7160), .ZN(n7161) );
  NOR2_X1 U8979 ( .A1(n7162), .A2(n7161), .ZN(n7164) );
  NAND2_X1 U8980 ( .A1(n7164), .A2(n7163), .ZN(n7318) );
  NAND2_X1 U8981 ( .A1(n7165), .A2(n7318), .ZN(n7170) );
  NAND2_X1 U8982 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7188) );
  INV_X1 U8983 ( .A(n7188), .ZN(n7167) );
  INV_X1 U8984 ( .A(n8715), .ZN(n8677) );
  OAI22_X1 U8985 ( .A1(n8677), .A2(n10455), .B1(n7330), .B2(n8717), .ZN(n7166)
         );
  AOI211_X1 U8986 ( .C1(n7168), .C2(n8707), .A(n7167), .B(n7166), .ZN(n7169)
         );
  OAI211_X1 U8987 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7775), .A(n7170), .B(
        n7169), .ZN(P2_U3158) );
  INV_X1 U8988 ( .A(n7171), .ZN(n7237) );
  AOI22_X1 U8989 ( .A1(n9372), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n8143), .ZN(n7172) );
  OAI21_X1 U8990 ( .B1(n7237), .B2(n9758), .A(n7172), .ZN(P1_U3341) );
  AOI21_X1 U8991 ( .B1(n7175), .B2(n7174), .A(n7173), .ZN(n7180) );
  AOI22_X1 U8992 ( .A1(n8090), .A2(n9308), .B1(n9209), .B2(n9306), .ZN(n7179)
         );
  AND2_X1 U8993 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8221) );
  NOR2_X1 U8994 ( .A1(n9294), .A2(n7609), .ZN(n7176) );
  AOI211_X1 U8995 ( .C1(n9243), .C2(n7177), .A(n8221), .B(n7176), .ZN(n7178)
         );
  OAI211_X1 U8996 ( .C1(n7180), .C2(n9277), .A(n7179), .B(n7178), .ZN(P1_U3218) );
  AOI21_X1 U8997 ( .B1(n7182), .B2(n7181), .A(n7242), .ZN(n7193) );
  INV_X1 U8998 ( .A(n8830), .ZN(n10415) );
  INV_X1 U8999 ( .A(n7250), .ZN(n7183) );
  AOI21_X1 U9000 ( .B1(n10552), .B2(n7184), .A(n7183), .ZN(n7190) );
  OAI21_X1 U9001 ( .B1(n7186), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7185), .ZN(
        n7187) );
  AOI22_X1 U9002 ( .A1(n10414), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n7255), .B2(
        n7187), .ZN(n7189) );
  OAI211_X1 U9003 ( .C1(n7190), .C2(n8837), .A(n7189), .B(n7188), .ZN(n7191)
         );
  AOI21_X1 U9004 ( .B1(n4993), .B2(n10415), .A(n7191), .ZN(n7192) );
  OAI21_X1 U9005 ( .B1(n7193), .B2(n8839), .A(n7192), .ZN(P2_U3185) );
  INV_X1 U9006 ( .A(n7194), .ZN(n7199) );
  AND2_X1 U9007 ( .A1(n7195), .A2(n7104), .ZN(n7197) );
  NOR2_X1 U9008 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  NAND2_X1 U9009 ( .A1(n7199), .A2(n7198), .ZN(n7204) );
  OR2_X1 U9010 ( .A1(n7204), .A2(n10438), .ZN(n10466) );
  INV_X1 U9011 ( .A(n10464), .ZN(n9040) );
  INV_X1 U9012 ( .A(n8584), .ZN(n7201) );
  NOR3_X1 U9013 ( .A1(n7201), .A2(n10537), .A3(n7200), .ZN(n7202) );
  AOI211_X1 U9014 ( .C1(n9040), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7203), .B(
        n7202), .ZN(n7205) );
  NAND2_X2 U9015 ( .A1(n7204), .A2(n10464), .ZN(n10471) );
  MUX2_X1 U9016 ( .A(n7206), .B(n7205), .S(n10471), .Z(n7207) );
  OAI21_X1 U9017 ( .B1(n10466), .B2(n7208), .A(n7207), .ZN(P2_U3233) );
  AOI22_X1 U9018 ( .A1(n7339), .A2(n6086), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7209), .ZN(n7213) );
  NAND2_X1 U9019 ( .A1(n7216), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U9020 ( .A1(n7211), .A2(n7210), .ZN(n7212) );
  NOR2_X1 U9021 ( .A1(n7213), .A2(n7212), .ZN(n7340) );
  AOI21_X1 U9022 ( .B1(n7213), .B2(n7212), .A(n7340), .ZN(n7223) );
  INV_X1 U9023 ( .A(n9435), .ZN(n9464) );
  NOR2_X1 U9024 ( .A1(n7339), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7214) );
  AOI21_X1 U9025 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7339), .A(n7214), .ZN(
        n7218) );
  OAI21_X1 U9026 ( .B1(n7218), .B2(n7217), .A(n7336), .ZN(n7219) );
  INV_X1 U9027 ( .A(n9458), .ZN(n9462) );
  NAND2_X1 U9028 ( .A1(n7219), .A2(n9462), .ZN(n7222) );
  INV_X1 U9029 ( .A(n9447), .ZN(n9460) );
  INV_X1 U9030 ( .A(n9467), .ZN(n9370) );
  INV_X1 U9031 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U9032 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7854) );
  OAI21_X1 U9033 ( .B1(n9370), .B2(n10152), .A(n7854), .ZN(n7220) );
  AOI21_X1 U9034 ( .B1(n7339), .B2(n9460), .A(n7220), .ZN(n7221) );
  OAI211_X1 U9035 ( .C1(n7223), .C2(n9464), .A(n7222), .B(n7221), .ZN(P1_U3252) );
  XNOR2_X1 U9036 ( .A(n7225), .B(n7224), .ZN(n7235) );
  INV_X1 U9037 ( .A(n7303), .ZN(n7226) );
  AOI21_X1 U9038 ( .B1(n4995), .B2(n4618), .A(n7226), .ZN(n7231) );
  OAI21_X1 U9039 ( .B1(n7228), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7227), .ZN(
        n7229) );
  AOI22_X1 U9040 ( .A1(n7229), .A2(n7255), .B1(n10414), .B2(
        P2_ADDR_REG_5__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U9041 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7329) );
  OAI211_X1 U9042 ( .C1(n7231), .C2(n8837), .A(n7230), .B(n7329), .ZN(n7232)
         );
  AOI21_X1 U9043 ( .B1(n7233), .B2(n10415), .A(n7232), .ZN(n7234) );
  OAI21_X1 U9044 ( .B1(n7235), .B2(n8839), .A(n7234), .ZN(P2_U3187) );
  INV_X1 U9045 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7236) );
  OAI222_X1 U9046 ( .A1(n7238), .A2(P2_U3151), .B1(n9164), .B2(n7237), .C1(
        n7236), .C2(n9167), .ZN(P2_U3281) );
  INV_X1 U9047 ( .A(n7239), .ZN(n7244) );
  INV_X1 U9048 ( .A(n8839), .ZN(n10419) );
  OAI21_X1 U9049 ( .B1(n7242), .B2(n7241), .A(n7240), .ZN(n7243) );
  NAND3_X1 U9050 ( .A1(n7244), .A2(n10419), .A3(n7243), .ZN(n7260) );
  INV_X1 U9051 ( .A(n7245), .ZN(n7247) );
  NOR2_X1 U9052 ( .A1(n7247), .A2(n7246), .ZN(n7251) );
  INV_X1 U9053 ( .A(n7248), .ZN(n7249) );
  AOI21_X1 U9054 ( .B1(n7251), .B2(n7250), .A(n7249), .ZN(n7252) );
  NAND2_X1 U9055 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8661) );
  OAI21_X1 U9056 ( .B1(n8837), .B2(n7252), .A(n8661), .ZN(n7258) );
  NAND3_X1 U9057 ( .A1(n7185), .A2(n7254), .A3(n7253), .ZN(n7256) );
  INV_X1 U9058 ( .A(n7255), .ZN(n8846) );
  AOI21_X1 U9059 ( .B1(n4619), .B2(n7256), .A(n8846), .ZN(n7257) );
  AOI211_X1 U9060 ( .C1(n10414), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7258), .B(
        n7257), .ZN(n7259) );
  OAI211_X1 U9061 ( .C1(n8830), .C2(n7261), .A(n7260), .B(n7259), .ZN(P2_U3186) );
  XNOR2_X1 U9062 ( .A(n7262), .B(n10416), .ZN(n7276) );
  INV_X1 U9063 ( .A(n7263), .ZN(n7274) );
  INV_X1 U9064 ( .A(n7264), .ZN(n7265) );
  AOI21_X1 U9065 ( .B1(n10548), .B2(n7266), .A(n7265), .ZN(n7267) );
  OAI22_X1 U9066 ( .A1(n8837), .A2(n7267), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10465), .ZN(n7273) );
  AOI21_X1 U9067 ( .B1(n10470), .B2(n7269), .A(n7268), .ZN(n7271) );
  INV_X1 U9068 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7270) );
  OAI22_X1 U9069 ( .A1(n8846), .A2(n7271), .B1(n8816), .B2(n7270), .ZN(n7272)
         );
  AOI211_X1 U9070 ( .C1(n7274), .C2(n10415), .A(n7273), .B(n7272), .ZN(n7275)
         );
  OAI21_X1 U9071 ( .B1(n8839), .B2(n7276), .A(n7275), .ZN(P2_U3183) );
  INV_X1 U9072 ( .A(n7277), .ZN(n7314) );
  AOI22_X1 U9073 ( .A1(n8785), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8149), .ZN(n7278) );
  OAI21_X1 U9074 ( .B1(n7314), .B2(n9164), .A(n7278), .ZN(P2_U3280) );
  XNOR2_X1 U9075 ( .A(n7280), .B(n7279), .ZN(n7294) );
  AOI21_X1 U9076 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n7290) );
  OAI21_X1 U9077 ( .B1(n7286), .B2(n7285), .A(n7284), .ZN(n7287) );
  AOI22_X1 U9078 ( .A1(n6725), .A2(n7287), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7289) );
  NAND2_X1 U9079 ( .A1(n10414), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7288) );
  OAI211_X1 U9080 ( .C1(n8846), .C2(n7290), .A(n7289), .B(n7288), .ZN(n7291)
         );
  AOI21_X1 U9081 ( .B1(n7292), .B2(n10415), .A(n7291), .ZN(n7293) );
  OAI21_X1 U9082 ( .B1(n8839), .B2(n7294), .A(n7293), .ZN(P2_U3184) );
  AOI21_X1 U9083 ( .B1(n7296), .B2(n7295), .A(n7354), .ZN(n7313) );
  INV_X1 U9084 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7309) );
  INV_X1 U9085 ( .A(n7297), .ZN(n7301) );
  NAND3_X1 U9086 ( .A1(n7227), .A2(n7299), .A3(n7298), .ZN(n7300) );
  AOI21_X1 U9087 ( .B1(n7301), .B2(n7300), .A(n8846), .ZN(n7307) );
  NAND3_X1 U9088 ( .A1(n7303), .A2(n4623), .A3(n7302), .ZN(n7304) );
  AOI21_X1 U9089 ( .B1(n7305), .B2(n7304), .A(n8837), .ZN(n7306) );
  NOR2_X1 U9090 ( .A1(n7307), .A2(n7306), .ZN(n7308) );
  NAND2_X1 U9091 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7393) );
  OAI211_X1 U9092 ( .C1(n8816), .C2(n7309), .A(n7308), .B(n7393), .ZN(n7310)
         );
  AOI21_X1 U9093 ( .B1(n7311), .B2(n10415), .A(n7310), .ZN(n7312) );
  OAI21_X1 U9094 ( .B1(n7313), .B2(n8839), .A(n7312), .ZN(P2_U3188) );
  INV_X1 U9095 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9955) );
  INV_X1 U9096 ( .A(n9382), .ZN(n9373) );
  OAI222_X1 U9097 ( .A1(n9754), .A2(n9955), .B1(n9758), .B2(n7314), .C1(
        P1_U3086), .C2(n9373), .ZN(P1_U3340) );
  INV_X1 U9098 ( .A(n7427), .ZN(n7335) );
  INV_X1 U9099 ( .A(n7315), .ZN(n7316) );
  NAND2_X1 U9100 ( .A1(n7316), .A2(n8738), .ZN(n7317) );
  NAND2_X1 U9101 ( .A1(n7319), .A2(n7330), .ZN(n7324) );
  INV_X1 U9102 ( .A(n7319), .ZN(n7320) );
  NAND2_X1 U9103 ( .A1(n7320), .A2(n10428), .ZN(n7321) );
  INV_X1 U9104 ( .A(n7325), .ZN(n7323) );
  INV_X1 U9105 ( .A(n7324), .ZN(n7322) );
  XNOR2_X1 U9106 ( .A(n8569), .B(n10495), .ZN(n7386) );
  XNOR2_X1 U9107 ( .A(n7386), .B(n9035), .ZN(n7326) );
  NOR3_X1 U9108 ( .A1(n7323), .A2(n7322), .A3(n7326), .ZN(n7328) );
  INV_X1 U9109 ( .A(n7388), .ZN(n7327) );
  OAI21_X1 U9110 ( .B1(n7328), .B2(n7327), .A(n8693), .ZN(n7334) );
  INV_X1 U9111 ( .A(n7329), .ZN(n7332) );
  OAI22_X1 U9112 ( .A1(n8677), .A2(n7330), .B1(n7646), .B2(n8717), .ZN(n7331)
         );
  AOI211_X1 U9113 ( .C1(n10495), .C2(n8707), .A(n7332), .B(n7331), .ZN(n7333)
         );
  OAI211_X1 U9114 ( .C1(n7335), .C2(n7775), .A(n7334), .B(n7333), .ZN(P2_U3167) );
  OAI21_X1 U9115 ( .B1(n7339), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7336), .ZN(
        n7338) );
  XNOR2_X1 U9116 ( .A(n7433), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7337) );
  NOR2_X1 U9117 ( .A1(n7338), .A2(n7337), .ZN(n7432) );
  AOI211_X1 U9118 ( .C1(n7338), .C2(n7337), .A(n9458), .B(n7432), .ZN(n7347)
         );
  NOR2_X1 U9119 ( .A1(n7339), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7341) );
  NOR2_X1 U9120 ( .A1(n7341), .A2(n7340), .ZN(n7343) );
  MUX2_X1 U9121 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7438), .S(n7433), .Z(n7342)
         );
  NAND2_X1 U9122 ( .A1(n7343), .A2(n7342), .ZN(n7437) );
  OAI211_X1 U9123 ( .C1(n7343), .C2(n7342), .A(n7437), .B(n9435), .ZN(n7345)
         );
  AND2_X1 U9124 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7813) );
  AOI21_X1 U9125 ( .B1(n9467), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7813), .ZN(
        n7344) );
  OAI211_X1 U9126 ( .C1(n9447), .C2(n7439), .A(n7345), .B(n7344), .ZN(n7346)
         );
  OR2_X1 U9127 ( .A1(n7347), .A2(n7346), .ZN(P1_U3253) );
  INV_X1 U9128 ( .A(n7348), .ZN(n7384) );
  AOI22_X1 U9129 ( .A1(n9417), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n8143), .ZN(n7349) );
  OAI21_X1 U9130 ( .B1(n7384), .B2(n9758), .A(n7349), .ZN(P1_U3339) );
  AOI21_X1 U9131 ( .B1(n7351), .B2(n7652), .A(n7350), .ZN(n7368) );
  INV_X1 U9132 ( .A(n7406), .ZN(n7356) );
  NOR3_X1 U9133 ( .A1(n7354), .A2(n7353), .A3(n7352), .ZN(n7355) );
  OAI21_X1 U9134 ( .B1(n7356), .B2(n7355), .A(n10419), .ZN(n7367) );
  NAND2_X1 U9135 ( .A1(n7357), .A2(n10558), .ZN(n7360) );
  INV_X1 U9136 ( .A(n7358), .ZN(n7359) );
  AOI21_X1 U9137 ( .B1(n7360), .B2(n7359), .A(n8837), .ZN(n7365) );
  INV_X1 U9138 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10144) );
  OR2_X1 U9139 ( .A1(n8816), .A2(n10144), .ZN(n7362) );
  AND2_X1 U9140 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8591) );
  INV_X1 U9141 ( .A(n8591), .ZN(n7361) );
  OAI211_X1 U9142 ( .C1(n8830), .C2(n7363), .A(n7362), .B(n7361), .ZN(n7364)
         );
  NOR2_X1 U9143 ( .A1(n7365), .A2(n7364), .ZN(n7366) );
  OAI211_X1 U9144 ( .C1(n7368), .C2(n8846), .A(n7367), .B(n7366), .ZN(P2_U3189) );
  XNOR2_X1 U9145 ( .A(n7369), .B(n7374), .ZN(n7370) );
  NAND2_X1 U9146 ( .A1(n7370), .A2(n10443), .ZN(n7372) );
  AOI22_X1 U9147 ( .A1(n9035), .A2(n10427), .B1(n10425), .B2(n8738), .ZN(n7371) );
  NAND2_X1 U9148 ( .A1(n7372), .A2(n7371), .ZN(n10490) );
  INV_X1 U9149 ( .A(n10490), .ZN(n7382) );
  INV_X2 U9150 ( .A(n10471), .ZN(n10472) );
  OAI21_X1 U9151 ( .B1(n7375), .B2(n7374), .A(n7373), .ZN(n10492) );
  NAND2_X1 U9152 ( .A1(n7377), .A2(n7376), .ZN(n10463) );
  NAND2_X1 U9153 ( .A1(n10451), .A2(n10463), .ZN(n7378) );
  AOI22_X1 U9154 ( .A1(n9041), .A2(n8663), .B1(n9040), .B2(n8664), .ZN(n7379)
         );
  OAI21_X1 U9155 ( .B1(n6671), .B2(n10471), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9156 ( .B1(n10492), .B2(n10433), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9157 ( .B1(n7382), .B2(n10472), .A(n7381), .ZN(P2_U3229) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7383) );
  OAI222_X1 U9159 ( .A1(P2_U3151), .A2(n7385), .B1(n9164), .B2(n7384), .C1(
        n7383), .C2(n9167), .ZN(P2_U3279) );
  INV_X1 U9160 ( .A(n9039), .ZN(n7399) );
  NAND2_X1 U9161 ( .A1(n7386), .A2(n7394), .ZN(n7387) );
  NAND2_X1 U9162 ( .A1(n7388), .A2(n7387), .ZN(n7389) );
  XNOR2_X1 U9163 ( .A(n8569), .B(n10505), .ZN(n7533) );
  XNOR2_X1 U9164 ( .A(n7533), .B(n7646), .ZN(n7390) );
  AOI21_X1 U9165 ( .B1(n7389), .B2(n7390), .A(n8711), .ZN(n7392) );
  INV_X1 U9166 ( .A(n7390), .ZN(n7391) );
  NAND2_X1 U9167 ( .A1(n7392), .A2(n7536), .ZN(n7398) );
  INV_X1 U9168 ( .A(n7393), .ZN(n7396) );
  OAI22_X1 U9169 ( .A1(n8677), .A2(n7394), .B1(n7544), .B2(n8717), .ZN(n7395)
         );
  AOI211_X1 U9170 ( .C1(n10505), .C2(n8707), .A(n7396), .B(n7395), .ZN(n7397)
         );
  OAI211_X1 U9171 ( .C1(n7399), .C2(n7775), .A(n7398), .B(n7397), .ZN(P2_U3179) );
  INV_X1 U9172 ( .A(n7400), .ZN(n7448) );
  AOI22_X1 U9173 ( .A1(n8822), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8149), .ZN(n7401) );
  OAI21_X1 U9174 ( .B1(n7448), .B2(n9164), .A(n7401), .ZN(P2_U3278) );
  AOI21_X1 U9175 ( .B1(n7403), .B2(n7402), .A(n4621), .ZN(n7419) );
  AND3_X1 U9176 ( .A1(n7406), .A2(n7405), .A3(n7404), .ZN(n7407) );
  OAI21_X1 U9177 ( .B1(n7554), .B2(n7407), .A(n10419), .ZN(n7418) );
  INV_X1 U9178 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10147) );
  INV_X1 U9179 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7408) );
  NOR2_X1 U9180 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7408), .ZN(n7546) );
  INV_X1 U9181 ( .A(n7546), .ZN(n7409) );
  OAI21_X1 U9182 ( .B1(n8816), .B2(n10147), .A(n7409), .ZN(n7415) );
  AOI21_X1 U9183 ( .B1(n7412), .B2(n7411), .A(n7410), .ZN(n7413) );
  NOR2_X1 U9184 ( .A1(n7413), .A2(n8846), .ZN(n7414) );
  AOI211_X1 U9185 ( .C1(n10415), .C2(n7416), .A(n7415), .B(n7414), .ZN(n7417)
         );
  OAI211_X1 U9186 ( .C1(n7419), .C2(n8837), .A(n7418), .B(n7417), .ZN(P2_U3190) );
  INV_X1 U9187 ( .A(n7426), .ZN(n7420) );
  XNOR2_X1 U9188 ( .A(n7421), .B(n7420), .ZN(n7422) );
  NAND2_X1 U9189 ( .A1(n7422), .A2(n10443), .ZN(n7424) );
  AOI22_X1 U9190 ( .A1(n10427), .A2(n8737), .B1(n10428), .B2(n10425), .ZN(
        n7423) );
  AND2_X1 U9191 ( .A1(n7424), .A2(n7423), .ZN(n10498) );
  XNOR2_X1 U9192 ( .A(n7425), .B(n7426), .ZN(n10494) );
  INV_X1 U9193 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7429) );
  AOI22_X1 U9194 ( .A1(n9041), .A2(n10495), .B1(n9040), .B2(n7427), .ZN(n7428)
         );
  OAI21_X1 U9195 ( .B1(n7429), .B2(n10471), .A(n7428), .ZN(n7430) );
  AOI21_X1 U9196 ( .B1(n10494), .B2(n10433), .A(n7430), .ZN(n7431) );
  OAI21_X1 U9197 ( .B1(n10498), .B2(n10472), .A(n7431), .ZN(P2_U3228) );
  NAND2_X1 U9198 ( .A1(n8187), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7434) );
  OAI21_X1 U9199 ( .B1(n8187), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7434), .ZN(
        n7435) );
  AOI211_X1 U9200 ( .C1(n7436), .C2(n7435), .A(n8186), .B(n9458), .ZN(n7447)
         );
  OAI21_X1 U9201 ( .B1(n7439), .B2(n7438), .A(n7437), .ZN(n7442) );
  MUX2_X1 U9202 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7440), .S(n8187), .Z(n7441)
         );
  NAND2_X1 U9203 ( .A1(n7441), .A2(n7442), .ZN(n8173) );
  OAI211_X1 U9204 ( .C1(n7442), .C2(n7441), .A(n9435), .B(n8173), .ZN(n7445)
         );
  INV_X1 U9205 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7443) );
  NOR2_X1 U9206 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7443), .ZN(n7884) );
  AOI21_X1 U9207 ( .B1(n9467), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7884), .ZN(
        n7444) );
  OAI211_X1 U9208 ( .C1(n9447), .C2(n8174), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OR2_X1 U9209 ( .A1(n7447), .A2(n7446), .ZN(P1_U3254) );
  INV_X1 U9210 ( .A(n9427), .ZN(n9416) );
  OAI222_X1 U9211 ( .A1(n9754), .A2(n9970), .B1(P1_U3086), .B2(n9416), .C1(
        n9758), .C2(n7448), .ZN(P1_U3338) );
  NAND2_X1 U9212 ( .A1(n7451), .A2(n9285), .ZN(n7455) );
  INV_X1 U9213 ( .A(n10358), .ZN(n10374) );
  AOI22_X1 U9214 ( .A1(n10371), .A2(n9305), .B1(n9306), .B2(n10374), .ZN(n7506) );
  INV_X1 U9215 ( .A(n9241), .ZN(n7452) );
  INV_X1 U9216 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9325) );
  OAI22_X1 U9217 ( .A1(n7506), .A2(n7452), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9325), .ZN(n7453) );
  AOI21_X1 U9218 ( .B1(n8236), .B2(n6637), .A(n7453), .ZN(n7454) );
  OAI211_X1 U9219 ( .C1(n9288), .C2(n7508), .A(n7455), .B(n7454), .ZN(P1_U3227) );
  NAND2_X1 U9220 ( .A1(n4936), .A2(n7456), .ZN(n7457) );
  XNOR2_X1 U9221 ( .A(n7458), .B(n7457), .ZN(n7462) );
  AOI22_X1 U9222 ( .A1(n8090), .A2(n10323), .B1(n9209), .B2(n10322), .ZN(n7461) );
  AND2_X1 U9223 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9343) );
  NOR2_X1 U9224 ( .A1(n9288), .A2(n7522), .ZN(n7459) );
  AOI211_X1 U9225 ( .C1(n8240), .C2(n6637), .A(n9343), .B(n7459), .ZN(n7460)
         );
  OAI211_X1 U9226 ( .C1(n7462), .C2(n9277), .A(n7461), .B(n7460), .ZN(P1_U3239) );
  XNOR2_X1 U9227 ( .A(n7463), .B(n7473), .ZN(n10355) );
  INV_X1 U9228 ( .A(n10355), .ZN(n7488) );
  INV_X1 U9229 ( .A(n7464), .ZN(n7467) );
  NAND3_X1 U9230 ( .A1(n7467), .A2(n7466), .A3(n7465), .ZN(n7468) );
  AND2_X2 U9231 ( .A1(n7468), .A2(n9603), .ZN(n10282) );
  AND2_X1 U9232 ( .A1(n7469), .A2(n8434), .ZN(n7470) );
  NAND2_X1 U9233 ( .A1(n10261), .A2(n7470), .ZN(n10211) );
  INV_X1 U9234 ( .A(n7471), .ZN(n10370) );
  NAND2_X1 U9235 ( .A1(n10261), .A2(n10370), .ZN(n7472) );
  NAND2_X1 U9236 ( .A1(n10211), .A2(n7472), .ZN(n10242) );
  NAND3_X1 U9237 ( .A1(n7474), .A2(n8453), .A3(n7473), .ZN(n7475) );
  INV_X1 U9238 ( .A(n10250), .ZN(n10345) );
  AOI21_X1 U9239 ( .B1(n7594), .B2(n7475), .A(n10345), .ZN(n10354) );
  NAND2_X1 U9240 ( .A1(n10228), .A2(n7476), .ZN(n7477) );
  NAND2_X1 U9241 ( .A1(n7477), .A2(n7484), .ZN(n7478) );
  INV_X1 U9242 ( .A(n9626), .ZN(n10273) );
  NAND3_X1 U9243 ( .A1(n7588), .A2(n7478), .A3(n10273), .ZN(n10351) );
  NAND2_X1 U9244 ( .A1(n10261), .A2(n7479), .ZN(n9612) );
  AND2_X2 U9245 ( .A1(n10261), .A2(n10252), .ZN(n10275) );
  NAND2_X1 U9246 ( .A1(n10261), .A2(n10371), .ZN(n9609) );
  INV_X1 U9247 ( .A(n7810), .ZN(n7480) );
  AOI22_X1 U9248 ( .A1(n10282), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7480), .B2(
        n10271), .ZN(n7482) );
  AND2_X1 U9249 ( .A1(n10261), .A2(n10374), .ZN(n9607) );
  NAND2_X1 U9250 ( .A1(n9607), .A2(n10349), .ZN(n7481) );
  OAI211_X1 U9251 ( .C1(n7952), .C2(n9609), .A(n7482), .B(n7481), .ZN(n7483)
         );
  AOI21_X1 U9252 ( .B1(n7484), .B2(n10275), .A(n7483), .ZN(n7485) );
  OAI21_X1 U9253 ( .B1(n10351), .B2(n9612), .A(n7485), .ZN(n7486) );
  AOI21_X1 U9254 ( .B1(n10354), .B2(n10261), .A(n7486), .ZN(n7487) );
  OAI21_X1 U9255 ( .B1(n7488), .B2(n9635), .A(n7487), .ZN(P1_U3283) );
  OR2_X1 U9256 ( .A1(n7517), .A2(n8226), .ZN(n7489) );
  INV_X1 U9257 ( .A(n8449), .ZN(n8363) );
  AND2_X1 U9258 ( .A1(n7489), .A2(n8363), .ZN(n7635) );
  XNOR2_X1 U9259 ( .A(n7635), .B(n7634), .ZN(n7490) );
  NAND2_X1 U9260 ( .A1(n7490), .A2(n10250), .ZN(n7492) );
  AOI22_X1 U9261 ( .A1(n10374), .A2(n9305), .B1(n10341), .B2(n10371), .ZN(
        n7491) );
  NAND2_X1 U9262 ( .A1(n7492), .A2(n7491), .ZN(n10335) );
  INV_X1 U9263 ( .A(n10335), .ZN(n7502) );
  XNOR2_X1 U9264 ( .A(n7493), .B(n7634), .ZN(n10330) );
  INV_X1 U9265 ( .A(n10226), .ZN(n7495) );
  AOI21_X1 U9266 ( .B1(n7520), .B2(n7497), .A(n9626), .ZN(n7494) );
  NAND2_X1 U9267 ( .A1(n7495), .A2(n7494), .ZN(n10331) );
  INV_X1 U9268 ( .A(n7496), .ZN(n7584) );
  AOI22_X1 U9269 ( .A1(n10282), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7584), .B2(
        n10271), .ZN(n7499) );
  NAND2_X1 U9270 ( .A1(n7497), .A2(n10275), .ZN(n7498) );
  OAI211_X1 U9271 ( .C1(n10331), .C2(n9612), .A(n7499), .B(n7498), .ZN(n7500)
         );
  AOI21_X1 U9272 ( .B1(n10330), .B2(n10242), .A(n7500), .ZN(n7501) );
  OAI21_X1 U9273 ( .B1(n7502), .B2(n10282), .A(n7501), .ZN(P1_U3286) );
  XOR2_X1 U9274 ( .A(n8362), .B(n7503), .Z(n10316) );
  NAND2_X1 U9275 ( .A1(n7504), .A2(n8230), .ZN(n7505) );
  XNOR2_X1 U9276 ( .A(n8362), .B(n7505), .ZN(n7507) );
  OAI21_X1 U9277 ( .B1(n7507), .B2(n10345), .A(n7506), .ZN(n10319) );
  NAND2_X1 U9278 ( .A1(n10319), .A2(n10261), .ZN(n7514) );
  OAI22_X1 U9279 ( .A1(n10261), .A2(n7509), .B1(n7508), .B2(n9603), .ZN(n7512)
         );
  INV_X1 U9280 ( .A(n10239), .ZN(n7510) );
  OAI211_X1 U9281 ( .C1(n7510), .C2(n10318), .A(n10273), .B(n7519), .ZN(n10317) );
  NOR2_X1 U9282 ( .A1(n10317), .A2(n9612), .ZN(n7511) );
  AOI211_X1 U9283 ( .C1(n10275), .C2(n8236), .A(n7512), .B(n7511), .ZN(n7513)
         );
  OAI211_X1 U9284 ( .C1(n9635), .C2(n10316), .A(n7514), .B(n7513), .ZN(
        P1_U3288) );
  XNOR2_X1 U9285 ( .A(n7515), .B(n7516), .ZN(n10329) );
  INV_X1 U9286 ( .A(n10329), .ZN(n7529) );
  XOR2_X1 U9287 ( .A(n7517), .B(n7516), .Z(n7518) );
  NOR2_X1 U9288 ( .A1(n7518), .A2(n10345), .ZN(n10327) );
  AOI21_X1 U9289 ( .B1(n7519), .B2(n8240), .A(n9626), .ZN(n7521) );
  NAND2_X1 U9290 ( .A1(n7521), .A2(n7520), .ZN(n10325) );
  OAI22_X1 U9291 ( .A1(n10261), .A2(n7523), .B1(n7522), .B2(n9603), .ZN(n7524)
         );
  AOI21_X1 U9292 ( .B1(n10275), .B2(n8240), .A(n7524), .ZN(n7526) );
  INV_X1 U9293 ( .A(n9609), .ZN(n7576) );
  AOI22_X1 U9294 ( .A1(n7576), .A2(n10322), .B1(n9607), .B2(n10323), .ZN(n7525) );
  OAI211_X1 U9295 ( .C1(n10325), .C2(n9612), .A(n7526), .B(n7525), .ZN(n7527)
         );
  AOI21_X1 U9296 ( .B1(n10327), .B2(n10261), .A(n7527), .ZN(n7528) );
  OAI21_X1 U9297 ( .B1(n9635), .B2(n7529), .A(n7528), .ZN(P1_U3287) );
  INV_X1 U9298 ( .A(n7702), .ZN(n7549) );
  XNOR2_X1 U9299 ( .A(n8569), .B(n8592), .ZN(n7530) );
  NAND2_X1 U9300 ( .A1(n7530), .A2(n7544), .ZN(n7538) );
  INV_X1 U9301 ( .A(n7530), .ZN(n7531) );
  NAND2_X1 U9302 ( .A1(n7531), .A2(n9036), .ZN(n7532) );
  AND2_X1 U9303 ( .A1(n7538), .A2(n7532), .ZN(n8588) );
  INV_X1 U9304 ( .A(n7533), .ZN(n7534) );
  NAND2_X1 U9305 ( .A1(n7534), .A2(n8737), .ZN(n8587) );
  AND2_X1 U9306 ( .A1(n8588), .A2(n8587), .ZN(n7535) );
  INV_X1 U9307 ( .A(n7539), .ZN(n7537) );
  XNOR2_X1 U9308 ( .A(n10513), .B(n8569), .ZN(n7614) );
  XNOR2_X1 U9309 ( .A(n7614), .B(n8736), .ZN(n7540) );
  NOR3_X1 U9310 ( .A1(n7537), .A2(n5027), .A3(n7540), .ZN(n7543) );
  NAND2_X1 U9311 ( .A1(n7541), .A2(n7540), .ZN(n7616) );
  INV_X1 U9312 ( .A(n7616), .ZN(n7542) );
  OAI21_X1 U9313 ( .B1(n7543), .B2(n7542), .A(n8693), .ZN(n7548) );
  INV_X1 U9314 ( .A(n8717), .ZN(n8675) );
  OAI22_X1 U9315 ( .A1(n7544), .A2(n8677), .B1(n8724), .B2(n7704), .ZN(n7545)
         );
  AOI211_X1 U9316 ( .C1(n8675), .C2(n8735), .A(n7546), .B(n7545), .ZN(n7547)
         );
  OAI211_X1 U9317 ( .C1(n7549), .C2(n7775), .A(n7548), .B(n7547), .ZN(P2_U3161) );
  AOI21_X1 U9318 ( .B1(n10562), .B2(n7551), .A(n7550), .ZN(n7566) );
  INV_X1 U9319 ( .A(n7666), .ZN(n7556) );
  NOR3_X1 U9320 ( .A1(n7554), .A2(n7553), .A3(n7552), .ZN(n7555) );
  OAI21_X1 U9321 ( .B1(n7556), .B2(n7555), .A(n10419), .ZN(n7565) );
  INV_X1 U9322 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U9323 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5444), .ZN(n7621) );
  INV_X1 U9324 ( .A(n7621), .ZN(n7557) );
  OAI21_X1 U9325 ( .B1(n8816), .B2(n10151), .A(n7557), .ZN(n7562) );
  AOI21_X1 U9326 ( .B1(n7716), .B2(n7559), .A(n7558), .ZN(n7560) );
  NOR2_X1 U9327 ( .A1(n7560), .A2(n8846), .ZN(n7561) );
  AOI211_X1 U9328 ( .C1(n10415), .C2(n7563), .A(n7562), .B(n7561), .ZN(n7564)
         );
  OAI211_X1 U9329 ( .C1(n7566), .C2(n8837), .A(n7565), .B(n7564), .ZN(P2_U3191) );
  INV_X1 U9330 ( .A(n7567), .ZN(n7603) );
  OAI222_X1 U9331 ( .A1(n9167), .A2(n7569), .B1(n9164), .B2(n7603), .C1(
        P2_U3151), .C2(n7568), .ZN(P2_U3277) );
  AOI21_X1 U9332 ( .B1(n10278), .B2(n10273), .A(n10275), .ZN(n7578) );
  INV_X1 U9333 ( .A(n7570), .ZN(n7572) );
  INV_X1 U9334 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7571) );
  OAI22_X1 U9335 ( .A1(n7573), .A2(n7572), .B1(n7571), .B2(n9603), .ZN(n7574)
         );
  MUX2_X1 U9336 ( .A(P1_REG2_REG_0__SCAN_IN), .B(n7574), .S(n10261), .Z(n7575)
         );
  AOI21_X1 U9337 ( .B1(n7576), .B2(n9310), .A(n7575), .ZN(n7577) );
  OAI21_X1 U9338 ( .B1(n7578), .B2(n10274), .A(n7577), .ZN(P1_U3293) );
  XOR2_X1 U9339 ( .A(n7579), .B(n7580), .Z(n7586) );
  OAI21_X1 U9340 ( .B1(n9294), .B2(n10332), .A(n7581), .ZN(n7583) );
  OAI22_X1 U9341 ( .A1(n8233), .A2(n9289), .B1(n9287), .B2(n7856), .ZN(n7582)
         );
  AOI211_X1 U9342 ( .C1(n7584), .C2(n9243), .A(n7583), .B(n7582), .ZN(n7585)
         );
  OAI21_X1 U9343 ( .B1(n7586), .B2(n9277), .A(n7585), .ZN(P1_U3213) );
  XOR2_X1 U9344 ( .A(n7595), .B(n7587), .Z(n10367) );
  AOI21_X1 U9345 ( .B1(n7588), .B2(n10362), .A(n9626), .ZN(n7589) );
  AND2_X1 U9346 ( .A1(n7589), .A2(n7685), .ZN(n10360) );
  INV_X1 U9347 ( .A(n10275), .ZN(n9631) );
  OAI22_X1 U9348 ( .A1(n10261), .A2(n7590), .B1(n7882), .B2(n9603), .ZN(n7592)
         );
  NOR2_X1 U9349 ( .A1(n9609), .A2(n10357), .ZN(n7591) );
  AOI211_X1 U9350 ( .C1(n9607), .C2(n9304), .A(n7592), .B(n7591), .ZN(n7593)
         );
  OAI21_X1 U9351 ( .B1(n7887), .B2(n9631), .A(n7593), .ZN(n7601) );
  INV_X1 U9352 ( .A(n7594), .ZN(n7597) );
  OAI21_X1 U9353 ( .B1(n7597), .B2(n7596), .A(n7595), .ZN(n7599) );
  NAND3_X1 U9354 ( .A1(n7599), .A2(n7598), .A3(n10250), .ZN(n10364) );
  NOR2_X1 U9355 ( .A1(n10364), .A2(n10282), .ZN(n7600) );
  AOI211_X1 U9356 ( .C1(n10360), .C2(n10278), .A(n7601), .B(n7600), .ZN(n7602)
         );
  OAI21_X1 U9357 ( .B1(n10367), .B2(n9635), .A(n7602), .ZN(P1_U3282) );
  INV_X1 U9358 ( .A(n9455), .ZN(n9446) );
  OAI222_X1 U9359 ( .A1(n9754), .A2(n9837), .B1(n9446), .B2(P1_U3086), .C1(
        n9758), .C2(n7603), .ZN(P1_U3337) );
  NAND2_X1 U9360 ( .A1(n8831), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7604) );
  OAI21_X1 U9361 ( .B1(n8862), .B2(n8831), .A(n7604), .ZN(P2_U3520) );
  XNOR2_X1 U9362 ( .A(n7605), .B(n7607), .ZN(n10306) );
  OAI21_X1 U9363 ( .B1(n8229), .B2(n7607), .A(n7606), .ZN(n7608) );
  AOI222_X1 U9364 ( .A1(n10250), .A2(n7608), .B1(n9308), .B2(n10374), .C1(
        n9306), .C2(n10371), .ZN(n10305) );
  MUX2_X1 U9365 ( .A(n6991), .B(n10305), .S(n10261), .Z(n7612) );
  AOI211_X1 U9366 ( .C1(n10303), .C2(n10256), .A(n9626), .B(n10240), .ZN(
        n10302) );
  OAI22_X1 U9367 ( .A1(n9631), .A2(n7609), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9603), .ZN(n7610) );
  AOI21_X1 U9368 ( .B1(n10302), .B2(n10278), .A(n7610), .ZN(n7611) );
  OAI211_X1 U9369 ( .C1(n9635), .C2(n10306), .A(n7612), .B(n7611), .ZN(
        P1_U3290) );
  INV_X1 U9370 ( .A(n7613), .ZN(n7715) );
  NAND2_X1 U9371 ( .A1(n7614), .A2(n7714), .ZN(n7615) );
  XNOR2_X1 U9372 ( .A(n10518), .B(n8569), .ZN(n7763) );
  XNOR2_X1 U9373 ( .A(n7763), .B(n7780), .ZN(n7618) );
  AOI21_X1 U9374 ( .B1(n7617), .B2(n7618), .A(n8711), .ZN(n7620) );
  INV_X1 U9375 ( .A(n7618), .ZN(n7619) );
  NAND2_X1 U9376 ( .A1(n7620), .A2(n7766), .ZN(n7625) );
  AOI21_X1 U9377 ( .B1(n8675), .B2(n8734), .A(n7621), .ZN(n7622) );
  OAI21_X1 U9378 ( .B1(n7714), .B2(n8677), .A(n7622), .ZN(n7623) );
  AOI21_X1 U9379 ( .B1(n10518), .B2(n8707), .A(n7623), .ZN(n7624) );
  OAI211_X1 U9380 ( .C1(n7715), .C2(n7775), .A(n7625), .B(n7624), .ZN(P2_U3171) );
  XNOR2_X1 U9381 ( .A(n7626), .B(n7639), .ZN(n10348) );
  XNOR2_X1 U9382 ( .A(n10228), .B(n10342), .ZN(n7628) );
  AND2_X1 U9383 ( .A1(n9304), .A2(n10371), .ZN(n7627) );
  AOI21_X1 U9384 ( .B1(n7628), .B2(n10273), .A(n7627), .ZN(n10344) );
  OAI22_X1 U9385 ( .A1(n10261), .A2(n7629), .B1(n7855), .B2(n9603), .ZN(n7630)
         );
  AOI21_X1 U9386 ( .B1(n9607), .B2(n10341), .A(n7630), .ZN(n7632) );
  NAND2_X1 U9387 ( .A1(n10342), .A2(n10275), .ZN(n7631) );
  OAI211_X1 U9388 ( .C1(n10344), .C2(n9612), .A(n7632), .B(n7631), .ZN(n7641)
         );
  OAI21_X1 U9389 ( .B1(n7635), .B2(n7634), .A(n7633), .ZN(n10218) );
  INV_X1 U9390 ( .A(n8258), .ZN(n7636) );
  AOI21_X1 U9391 ( .B1(n10218), .B2(n7637), .A(n7636), .ZN(n7638) );
  XOR2_X1 U9392 ( .A(n7639), .B(n7638), .Z(n10346) );
  AND2_X1 U9393 ( .A1(n10261), .A2(n10250), .ZN(n9516) );
  INV_X1 U9394 ( .A(n9516), .ZN(n9618) );
  NOR2_X1 U9395 ( .A1(n10346), .A2(n9618), .ZN(n7640) );
  AOI211_X1 U9396 ( .C1(n10242), .C2(n10348), .A(n7641), .B(n7640), .ZN(n7642)
         );
  INV_X1 U9397 ( .A(n7642), .ZN(P1_U3284) );
  INV_X1 U9398 ( .A(n10425), .ZN(n10456) );
  INV_X1 U9399 ( .A(n10443), .ZN(n10459) );
  XNOR2_X1 U9400 ( .A(n7644), .B(n7643), .ZN(n7645) );
  OAI222_X1 U9401 ( .A1(n10454), .A2(n7714), .B1(n10456), .B2(n7646), .C1(
        n10459), .C2(n7645), .ZN(n10509) );
  INV_X1 U9402 ( .A(n10509), .ZN(n7655) );
  INV_X1 U9403 ( .A(n7647), .ZN(n7650) );
  INV_X1 U9404 ( .A(n7699), .ZN(n7648) );
  AOI21_X1 U9405 ( .B1(n7650), .B2(n7649), .A(n7648), .ZN(n10511) );
  AOI22_X1 U9406 ( .A1(n9041), .A2(n8592), .B1(n9040), .B2(n8593), .ZN(n7651)
         );
  OAI21_X1 U9407 ( .B1(n7652), .B2(n10471), .A(n7651), .ZN(n7653) );
  AOI21_X1 U9408 ( .B1(n10511), .B2(n10433), .A(n7653), .ZN(n7654) );
  OAI21_X1 U9409 ( .B1(n7655), .B2(n10472), .A(n7654), .ZN(P2_U3226) );
  INV_X1 U9410 ( .A(n7656), .ZN(n7659) );
  OAI222_X1 U9411 ( .A1(n9754), .A2(n7657), .B1(n9758), .B2(n7659), .C1(
        P1_U3086), .C2(n7479), .ZN(P1_U3336) );
  OAI222_X1 U9412 ( .A1(P2_U3151), .A2(n7660), .B1(n9164), .B2(n7659), .C1(
        n7658), .C2(n9167), .ZN(P2_U3276) );
  AOI21_X1 U9413 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7679) );
  AND3_X1 U9414 ( .A1(n7666), .A2(n7665), .A3(n7664), .ZN(n7667) );
  OAI21_X1 U9415 ( .B1(n7668), .B2(n7667), .A(n10419), .ZN(n7678) );
  INV_X1 U9416 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10155) );
  INV_X1 U9417 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U9418 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10103), .ZN(n7770) );
  INV_X1 U9419 ( .A(n7770), .ZN(n7669) );
  OAI21_X1 U9420 ( .B1(n8816), .B2(n10155), .A(n7669), .ZN(n7675) );
  AOI21_X1 U9421 ( .B1(n7672), .B2(n7671), .A(n7670), .ZN(n7673) );
  NOR2_X1 U9422 ( .A1(n7673), .A2(n8846), .ZN(n7674) );
  AOI211_X1 U9423 ( .C1(n10415), .C2(n7676), .A(n7675), .B(n7674), .ZN(n7677)
         );
  OAI211_X1 U9424 ( .C1(n7679), .C2(n8837), .A(n7678), .B(n7677), .ZN(P2_U3192) );
  XNOR2_X1 U9425 ( .A(n7680), .B(n7681), .ZN(n10380) );
  INV_X1 U9426 ( .A(n10380), .ZN(n7695) );
  NAND2_X1 U9427 ( .A1(n7682), .A2(n7681), .ZN(n7683) );
  AOI21_X1 U9428 ( .B1(n7684), .B2(n7683), .A(n10345), .ZN(n10379) );
  NAND2_X1 U9429 ( .A1(n7685), .A2(n7944), .ZN(n7686) );
  NAND2_X1 U9430 ( .A1(n7686), .A2(n10273), .ZN(n7687) );
  OR2_X1 U9431 ( .A1(n7687), .A2(n7730), .ZN(n10376) );
  OAI22_X1 U9432 ( .A1(n10261), .A2(n7688), .B1(n7951), .B2(n9603), .ZN(n7690)
         );
  NOR2_X1 U9433 ( .A1(n9609), .A2(n8104), .ZN(n7689) );
  AOI211_X1 U9434 ( .C1(n9607), .C2(n10373), .A(n7690), .B(n7689), .ZN(n7692)
         );
  NAND2_X1 U9435 ( .A1(n7944), .A2(n10275), .ZN(n7691) );
  OAI211_X1 U9436 ( .C1(n10376), .C2(n9612), .A(n7692), .B(n7691), .ZN(n7693)
         );
  AOI21_X1 U9437 ( .B1(n10379), .B2(n10261), .A(n7693), .ZN(n7694) );
  OAI21_X1 U9438 ( .B1(n7695), .B2(n9635), .A(n7694), .ZN(P1_U3281) );
  XOR2_X1 U9439 ( .A(n7696), .B(n7700), .Z(n7697) );
  AOI222_X1 U9440 ( .A1(n10443), .A2(n7697), .B1(n8735), .B2(n10427), .C1(
        n9036), .C2(n10425), .ZN(n10516) );
  NAND2_X1 U9441 ( .A1(n7699), .A2(n7698), .ZN(n7701) );
  XNOR2_X1 U9442 ( .A(n7701), .B(n7700), .ZN(n10514) );
  AOI22_X1 U9443 ( .A1(n10472), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9040), .B2(
        n7702), .ZN(n7703) );
  OAI21_X1 U9444 ( .B1(n7704), .B2(n10466), .A(n7703), .ZN(n7705) );
  AOI21_X1 U9445 ( .B1(n10514), .B2(n10433), .A(n7705), .ZN(n7706) );
  OAI21_X1 U9446 ( .B1(n10516), .B2(n10472), .A(n7706), .ZN(P2_U3225) );
  INV_X1 U9447 ( .A(n7707), .ZN(n7721) );
  OAI222_X1 U9448 ( .A1(n9758), .A2(n7721), .B1(n8512), .B2(P1_U3086), .C1(
        n9835), .C2(n9754), .ZN(P1_U3335) );
  INV_X1 U9449 ( .A(n7709), .ZN(n7710) );
  AOI21_X1 U9450 ( .B1(n7708), .B2(n7711), .A(n7710), .ZN(n10523) );
  INV_X1 U9451 ( .A(n10523), .ZN(n10520) );
  XNOR2_X1 U9452 ( .A(n7712), .B(n7711), .ZN(n7713) );
  OAI222_X1 U9453 ( .A1(n10454), .A2(n7820), .B1(n10456), .B2(n7714), .C1(
        n7713), .C2(n10459), .ZN(n10521) );
  NAND2_X1 U9454 ( .A1(n10521), .A2(n10471), .ZN(n7719) );
  OAI22_X1 U9455 ( .A1(n10471), .A2(n7716), .B1(n7715), .B2(n10464), .ZN(n7717) );
  AOI21_X1 U9456 ( .B1(n9041), .B2(n10518), .A(n7717), .ZN(n7718) );
  OAI211_X1 U9457 ( .C1(n9024), .C2(n10520), .A(n7719), .B(n7718), .ZN(
        P2_U3224) );
  OAI222_X1 U9458 ( .A1(n7722), .A2(P2_U3151), .B1(n9164), .B2(n7721), .C1(
        n7720), .C2(n9167), .ZN(P2_U3275) );
  AOI21_X1 U9459 ( .B1(n7723), .B2(n8379), .A(n10345), .ZN(n7727) );
  NAND2_X1 U9460 ( .A1(n9302), .A2(n10371), .ZN(n7725) );
  NAND2_X1 U9461 ( .A1(n9303), .A2(n10374), .ZN(n7724) );
  NAND2_X1 U9462 ( .A1(n7725), .A2(n7724), .ZN(n8039) );
  AOI21_X1 U9463 ( .B1(n7727), .B2(n7726), .A(n8039), .ZN(n10382) );
  XNOR2_X1 U9464 ( .A(n7728), .B(n8379), .ZN(n10386) );
  NAND2_X1 U9465 ( .A1(n10386), .A2(n10242), .ZN(n7734) );
  OAI22_X1 U9466 ( .A1(n10261), .A2(n7729), .B1(n8041), .B2(n9603), .ZN(n7732)
         );
  OAI211_X1 U9467 ( .C1(n7730), .C2(n10383), .A(n10212), .B(n10273), .ZN(
        n10381) );
  NOR2_X1 U9468 ( .A1(n10381), .A2(n9612), .ZN(n7731) );
  AOI211_X1 U9469 ( .C1(n10275), .C2(n8048), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI211_X1 U9470 ( .C1(n10282), .C2(n10382), .A(n7734), .B(n7733), .ZN(
        P1_U3280) );
  AOI21_X1 U9471 ( .B1(n7824), .B2(n7736), .A(n7735), .ZN(n7751) );
  INV_X1 U9472 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10159) );
  INV_X1 U9473 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7737) );
  NOR2_X1 U9474 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7737), .ZN(n7796) );
  INV_X1 U9475 ( .A(n7796), .ZN(n7738) );
  OAI21_X1 U9476 ( .B1(n8816), .B2(n10159), .A(n7738), .ZN(n7744) );
  AOI21_X1 U9477 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7742) );
  NOR2_X1 U9478 ( .A1(n7742), .A2(n8839), .ZN(n7743) );
  AOI211_X1 U9479 ( .C1(n10415), .C2(n7745), .A(n7744), .B(n7743), .ZN(n7750)
         );
  AOI21_X1 U9480 ( .B1(n10566), .B2(n7747), .A(n7746), .ZN(n7748) );
  OR2_X1 U9481 ( .A1(n7748), .A2(n8837), .ZN(n7749) );
  OAI211_X1 U9482 ( .C1(n7751), .C2(n8846), .A(n7750), .B(n7749), .ZN(P2_U3193) );
  XOR2_X1 U9483 ( .A(n7752), .B(n7847), .Z(n7754) );
  NOR2_X1 U9484 ( .A1(n7754), .A2(n7753), .ZN(n7848) );
  AOI21_X1 U9485 ( .B1(n7754), .B2(n7753), .A(n7848), .ZN(n7759) );
  OAI22_X1 U9486 ( .A1(n7755), .A2(n10358), .B1(n7811), .B2(n10356), .ZN(
        n10219) );
  AOI22_X1 U9487 ( .A1(n10219), .A2(n9241), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7756) );
  OAI21_X1 U9488 ( .B1(n10221), .B2(n9288), .A(n7756), .ZN(n7757) );
  AOI21_X1 U9489 ( .B1(n10223), .B2(n6637), .A(n7757), .ZN(n7758) );
  OAI21_X1 U9490 ( .B1(n7759), .B2(n9277), .A(n7758), .ZN(P1_U3221) );
  INV_X1 U9491 ( .A(n7760), .ZN(n7804) );
  OAI222_X1 U9492 ( .A1(n9758), .A2(n7804), .B1(n6325), .B2(P1_U3086), .C1(
        n7761), .C2(n9754), .ZN(P1_U3334) );
  INV_X1 U9493 ( .A(n7762), .ZN(n7785) );
  INV_X1 U9494 ( .A(n7763), .ZN(n7764) );
  NAND2_X1 U9495 ( .A1(n7764), .A2(n8735), .ZN(n7765) );
  XNOR2_X1 U9496 ( .A(n7788), .B(n8569), .ZN(n7767) );
  NAND2_X1 U9497 ( .A1(n7768), .A2(n7767), .ZN(n7794) );
  OAI21_X1 U9498 ( .B1(n7768), .B2(n7767), .A(n7794), .ZN(n7769) );
  NAND2_X1 U9499 ( .A1(n7769), .A2(n8693), .ZN(n7774) );
  AOI21_X1 U9500 ( .B1(n8675), .B2(n8733), .A(n7770), .ZN(n7771) );
  OAI21_X1 U9501 ( .B1(n7780), .B2(n8677), .A(n7771), .ZN(n7772) );
  AOI21_X1 U9502 ( .B1(n7788), .B2(n8707), .A(n7772), .ZN(n7773) );
  OAI211_X1 U9503 ( .C1(n7775), .C2(n7785), .A(n7774), .B(n7773), .ZN(P2_U3157) );
  INV_X1 U9504 ( .A(n10463), .ZN(n10448) );
  INV_X1 U9505 ( .A(n7778), .ZN(n7776) );
  XNOR2_X1 U9506 ( .A(n7777), .B(n7776), .ZN(n10528) );
  INV_X1 U9507 ( .A(n10528), .ZN(n7784) );
  XNOR2_X1 U9508 ( .A(n7779), .B(n7778), .ZN(n7782) );
  OAI22_X1 U9509 ( .A1(n7780), .A2(n10456), .B1(n7921), .B2(n10454), .ZN(n7781) );
  AOI21_X1 U9510 ( .B1(n7782), .B2(n10443), .A(n7781), .ZN(n7783) );
  OAI21_X1 U9511 ( .B1(n10528), .B2(n10451), .A(n7783), .ZN(n10530) );
  AOI21_X1 U9512 ( .B1(n10448), .B2(n7784), .A(n10530), .ZN(n7790) );
  OAI22_X1 U9513 ( .A1(n10471), .A2(n7786), .B1(n7785), .B2(n10464), .ZN(n7787) );
  AOI21_X1 U9514 ( .B1(n9041), .B2(n7788), .A(n7787), .ZN(n7789) );
  OAI21_X1 U9515 ( .B1(n7790), .B2(n10472), .A(n7789), .ZN(P2_U3223) );
  INV_X1 U9516 ( .A(n7791), .ZN(n7792) );
  NAND2_X1 U9517 ( .A1(n7792), .A2(n7820), .ZN(n7795) );
  XNOR2_X1 U9518 ( .A(n7817), .B(n8556), .ZN(n7861) );
  NAND2_X1 U9519 ( .A1(n7866), .A2(n8693), .ZN(n7802) );
  AOI21_X1 U9520 ( .B1(n7794), .B2(n7795), .A(n7861), .ZN(n7801) );
  NAND2_X1 U9521 ( .A1(n8720), .A2(n7822), .ZN(n7798) );
  AOI21_X1 U9522 ( .B1(n8675), .B2(n8732), .A(n7796), .ZN(n7797) );
  OAI211_X1 U9523 ( .C1(n7820), .C2(n8677), .A(n7798), .B(n7797), .ZN(n7799)
         );
  AOI21_X1 U9524 ( .B1(n10536), .B2(n8707), .A(n7799), .ZN(n7800) );
  OAI21_X1 U9525 ( .B1(n7802), .B2(n7801), .A(n7800), .ZN(P2_U3176) );
  OAI222_X1 U9526 ( .A1(n7805), .A2(P2_U3151), .B1(n9164), .B2(n7804), .C1(
        n7803), .C2(n9167), .ZN(P2_U3274) );
  OAI21_X1 U9527 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7809) );
  NAND2_X1 U9528 ( .A1(n7809), .A2(n9285), .ZN(n7815) );
  OAI22_X1 U9529 ( .A1(n9289), .A2(n7811), .B1(n9288), .B2(n7810), .ZN(n7812)
         );
  AOI211_X1 U9530 ( .C1(n9209), .C2(n10373), .A(n7813), .B(n7812), .ZN(n7814)
         );
  OAI211_X1 U9531 ( .C1(n10352), .C2(n9294), .A(n7815), .B(n7814), .ZN(
        P1_U3217) );
  XNOR2_X1 U9532 ( .A(n7816), .B(n7817), .ZN(n10533) );
  XNOR2_X1 U9533 ( .A(n7818), .B(n7817), .ZN(n7819) );
  OAI222_X1 U9534 ( .A1(n10454), .A2(n7821), .B1(n10456), .B2(n7820), .C1(
        n7819), .C2(n10459), .ZN(n10534) );
  NAND2_X1 U9535 ( .A1(n10534), .A2(n10471), .ZN(n7827) );
  INV_X1 U9536 ( .A(n7822), .ZN(n7823) );
  OAI22_X1 U9537 ( .A1(n10471), .A2(n7824), .B1(n7823), .B2(n10464), .ZN(n7825) );
  AOI21_X1 U9538 ( .B1(n10536), .B2(n9041), .A(n7825), .ZN(n7826) );
  OAI211_X1 U9539 ( .C1(n9024), .C2(n10533), .A(n7827), .B(n7826), .ZN(
        P2_U3222) );
  AOI21_X1 U9540 ( .B1(n7830), .B2(n7829), .A(n7828), .ZN(n7846) );
  INV_X1 U9541 ( .A(n7831), .ZN(n7833) );
  NAND2_X1 U9542 ( .A1(n7833), .A2(n7832), .ZN(n7834) );
  XNOR2_X1 U9543 ( .A(n7835), .B(n7834), .ZN(n7844) );
  AOI21_X1 U9544 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7839) );
  NOR2_X1 U9545 ( .A1(n7839), .A2(n8837), .ZN(n7843) );
  AND2_X1 U9546 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7871) );
  AOI21_X1 U9547 ( .B1(n10414), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7871), .ZN(
        n7840) );
  OAI21_X1 U9548 ( .B1(n7841), .B2(n8830), .A(n7840), .ZN(n7842) );
  AOI211_X1 U9549 ( .C1(n7844), .C2(n10419), .A(n7843), .B(n7842), .ZN(n7845)
         );
  OAI21_X1 U9550 ( .B1(n7846), .B2(n8846), .A(n7845), .ZN(P2_U3194) );
  INV_X1 U9551 ( .A(n7847), .ZN(n7849) );
  AOI21_X1 U9552 ( .B1(n7849), .B2(n7752), .A(n7848), .ZN(n7853) );
  XNOR2_X1 U9553 ( .A(n7851), .B(n7850), .ZN(n7852) );
  XNOR2_X1 U9554 ( .A(n7853), .B(n7852), .ZN(n7860) );
  OAI21_X1 U9555 ( .B1(n9287), .B2(n10359), .A(n7854), .ZN(n7858) );
  OAI22_X1 U9556 ( .A1(n9289), .A2(n7856), .B1(n9288), .B2(n7855), .ZN(n7857)
         );
  OAI21_X1 U9557 ( .B1(n7860), .B2(n9277), .A(n7859), .ZN(P1_U3231) );
  INV_X1 U9558 ( .A(n7863), .ZN(n10540) );
  INV_X1 U9559 ( .A(n7861), .ZN(n7862) );
  NAND2_X1 U9560 ( .A1(n7862), .A2(n8733), .ZN(n7868) );
  XNOR2_X1 U9561 ( .A(n7863), .B(n8556), .ZN(n7864) );
  NOR2_X1 U9562 ( .A1(n7864), .A2(n8732), .ZN(n7929) );
  AOI21_X1 U9563 ( .B1(n7864), .B2(n8732), .A(n7929), .ZN(n7867) );
  INV_X1 U9564 ( .A(n7935), .ZN(n7870) );
  AOI21_X1 U9565 ( .B1(n7866), .B2(n7868), .A(n7867), .ZN(n7869) );
  OAI21_X1 U9566 ( .B1(n7870), .B2(n7869), .A(n8693), .ZN(n7875) );
  AOI21_X1 U9567 ( .B1(n8675), .B2(n8731), .A(n7871), .ZN(n7872) );
  OAI21_X1 U9568 ( .B1(n7921), .B2(n8677), .A(n7872), .ZN(n7873) );
  AOI21_X1 U9569 ( .B1(n7924), .B2(n8720), .A(n7873), .ZN(n7874) );
  OAI211_X1 U9570 ( .C1(n10540), .C2(n8724), .A(n7875), .B(n7874), .ZN(
        P2_U3164) );
  INV_X1 U9571 ( .A(n7876), .ZN(n8140) );
  OAI222_X1 U9572 ( .A1(P2_U3151), .A2(n7878), .B1(n9164), .B2(n8140), .C1(
        n7877), .C2(n9167), .ZN(P2_U3273) );
  INV_X1 U9573 ( .A(n7806), .ZN(n7880) );
  NOR3_X1 U9574 ( .A1(n7880), .A2(n6516), .A3(n7879), .ZN(n7881) );
  OAI21_X1 U9575 ( .B1(n7881), .B2(n4602), .A(n9285), .ZN(n7886) );
  OAI22_X1 U9576 ( .A1(n9289), .A2(n10359), .B1(n9288), .B2(n7882), .ZN(n7883)
         );
  AOI211_X1 U9577 ( .C1(n9209), .C2(n9303), .A(n7884), .B(n7883), .ZN(n7885)
         );
  OAI211_X1 U9578 ( .C1(n7887), .C2(n9294), .A(n7886), .B(n7885), .ZN(P1_U3236) );
  NAND2_X1 U9579 ( .A1(n7893), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U9580 ( .A1(n7889), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8520) );
  OAI211_X1 U9581 ( .C1(n7891), .C2(n9754), .A(n7890), .B(n8520), .ZN(P1_U3332) );
  NAND2_X1 U9582 ( .A1(n7893), .A2(n7892), .ZN(n7895) );
  OAI211_X1 U9583 ( .C1(n7896), .C2(n9167), .A(n7895), .B(n7894), .ZN(P2_U3272) );
  INV_X1 U9584 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7905) );
  XNOR2_X1 U9585 ( .A(n7897), .B(n7899), .ZN(n7910) );
  OAI21_X1 U9586 ( .B1(n7900), .B2(n7899), .A(n7898), .ZN(n7901) );
  INV_X1 U9587 ( .A(n7901), .ZN(n7918) );
  AOI22_X1 U9588 ( .A1(n10374), .A2(n9302), .B1(n9300), .B2(n10371), .ZN(n7903) );
  INV_X1 U9589 ( .A(n10213), .ZN(n7902) );
  OAI211_X1 U9590 ( .C1(n4714), .C2(n7902), .A(n4716), .B(n10273), .ZN(n7913)
         );
  OAI211_X1 U9591 ( .C1(n7918), .C2(n10345), .A(n7903), .B(n7913), .ZN(n7904)
         );
  AOI21_X1 U9592 ( .B1(n7910), .B2(n10385), .A(n7904), .ZN(n7907) );
  MUX2_X1 U9593 ( .A(n7905), .B(n7907), .S(n10395), .Z(n7906) );
  OAI21_X1 U9594 ( .B1(n4714), .B2(n9747), .A(n7906), .ZN(P1_U3498) );
  INV_X1 U9595 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7908) );
  MUX2_X1 U9596 ( .A(n7908), .B(n7907), .S(n10413), .Z(n7909) );
  OAI21_X1 U9597 ( .B1(n4714), .B2(n9710), .A(n7909), .ZN(P1_U3537) );
  NAND2_X1 U9598 ( .A1(n7910), .A2(n10242), .ZN(n7917) );
  AOI22_X1 U9599 ( .A1(n10282), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8089), .B2(
        n10271), .ZN(n7912) );
  NAND2_X1 U9600 ( .A1(n9607), .A2(n9302), .ZN(n7911) );
  OAI211_X1 U9601 ( .C1(n8092), .C2(n9609), .A(n7912), .B(n7911), .ZN(n7915)
         );
  NOR2_X1 U9602 ( .A1(n7913), .A2(n9612), .ZN(n7914) );
  AOI211_X1 U9603 ( .C1(n10275), .C2(n8284), .A(n7915), .B(n7914), .ZN(n7916)
         );
  OAI211_X1 U9604 ( .C1(n7918), .C2(n9618), .A(n7917), .B(n7916), .ZN(P1_U3278) );
  XOR2_X1 U9605 ( .A(n7919), .B(n7922), .Z(n7920) );
  OAI222_X1 U9606 ( .A1(n10454), .A2(n7931), .B1(n10456), .B2(n7921), .C1(
        n7920), .C2(n10459), .ZN(n10541) );
  INV_X1 U9607 ( .A(n10541), .ZN(n7928) );
  XOR2_X1 U9608 ( .A(n7923), .B(n7922), .Z(n10543) );
  AOI22_X1 U9609 ( .A1(n10472), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9040), .B2(
        n7924), .ZN(n7925) );
  OAI21_X1 U9610 ( .B1(n10540), .B2(n10466), .A(n7925), .ZN(n7926) );
  AOI21_X1 U9611 ( .B1(n10543), .B2(n10433), .A(n7926), .ZN(n7927) );
  OAI21_X1 U9612 ( .B1(n7928), .B2(n10472), .A(n7927), .ZN(P2_U3221) );
  INV_X1 U9613 ( .A(n7929), .ZN(n7937) );
  XNOR2_X1 U9614 ( .A(n7930), .B(n8569), .ZN(n7932) );
  NAND2_X1 U9615 ( .A1(n7932), .A2(n7931), .ZN(n7981) );
  INV_X1 U9616 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U9617 ( .A1(n7933), .A2(n8731), .ZN(n7934) );
  NAND2_X1 U9618 ( .A1(n7981), .A2(n7934), .ZN(n7936) );
  AND3_X1 U9619 ( .A1(n7935), .A2(n7937), .A3(n7936), .ZN(n7938) );
  OAI21_X1 U9620 ( .B1(n7984), .B2(n7938), .A(n8693), .ZN(n7943) );
  NAND2_X1 U9621 ( .A1(n8715), .A2(n8732), .ZN(n7939) );
  NAND2_X1 U9622 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8750) );
  OAI211_X1 U9623 ( .C1(n7940), .C2(n8717), .A(n7939), .B(n8750), .ZN(n7941)
         );
  AOI21_X1 U9624 ( .B1(n7978), .B2(n8720), .A(n7941), .ZN(n7942) );
  OAI211_X1 U9625 ( .C1(n8000), .C2(n8724), .A(n7943), .B(n7942), .ZN(P2_U3174) );
  INV_X1 U9626 ( .A(n7944), .ZN(n10377) );
  INV_X1 U9627 ( .A(n7945), .ZN(n7947) );
  NOR3_X1 U9628 ( .A1(n4602), .A2(n7947), .A3(n7946), .ZN(n7950) );
  INV_X1 U9629 ( .A(n7948), .ZN(n7949) );
  OAI21_X1 U9630 ( .B1(n7950), .B2(n7949), .A(n9285), .ZN(n7955) );
  AND2_X1 U9631 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8207) );
  OAI22_X1 U9632 ( .A1(n9289), .A2(n7952), .B1(n9288), .B2(n7951), .ZN(n7953)
         );
  AOI211_X1 U9633 ( .C1(n9209), .C2(n10372), .A(n8207), .B(n7953), .ZN(n7954)
         );
  OAI211_X1 U9634 ( .C1(n10377), .C2(n9294), .A(n7955), .B(n7954), .ZN(
        P1_U3224) );
  XNOR2_X1 U9635 ( .A(n7956), .B(n7963), .ZN(n7957) );
  AOI222_X1 U9636 ( .A1(n10250), .A2(n7957), .B1(n9299), .B2(n10371), .C1(
        n9301), .C2(n10374), .ZN(n10195) );
  OAI22_X1 U9637 ( .A1(n10261), .A2(n9392), .B1(n9206), .B2(n9603), .ZN(n7960)
         );
  OAI211_X1 U9638 ( .C1(n10196), .C2(n7958), .A(n10273), .B(n8024), .ZN(n10194) );
  NOR2_X1 U9639 ( .A1(n10194), .A2(n9612), .ZN(n7959) );
  AOI211_X1 U9640 ( .C1(n10275), .C2(n7961), .A(n7960), .B(n7959), .ZN(n7965)
         );
  XNOR2_X1 U9641 ( .A(n7962), .B(n7963), .ZN(n10198) );
  NAND2_X1 U9642 ( .A1(n10198), .A2(n10242), .ZN(n7964) );
  OAI211_X1 U9643 ( .C1(n10195), .C2(n10282), .A(n7965), .B(n7964), .ZN(
        P1_U3277) );
  XNOR2_X1 U9644 ( .A(n7966), .B(n7971), .ZN(n8001) );
  OR2_X1 U9645 ( .A1(n7919), .A2(n7967), .ZN(n7970) );
  NAND2_X1 U9646 ( .A1(n7970), .A2(n7968), .ZN(n7974) );
  NAND2_X1 U9647 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  AOI21_X1 U9648 ( .B1(n7972), .B2(n7971), .A(n10459), .ZN(n7973) );
  OAI21_X1 U9649 ( .B1(n7974), .B2(n5147), .A(n7973), .ZN(n7976) );
  AOI22_X1 U9650 ( .A1(n10427), .A2(n8730), .B1(n8732), .B2(n10425), .ZN(n7975) );
  NAND2_X1 U9651 ( .A1(n7976), .A2(n7975), .ZN(n7999) );
  NOR2_X1 U9652 ( .A1(n8000), .A2(n10438), .ZN(n7977) );
  OAI21_X1 U9653 ( .B1(n7999), .B2(n7977), .A(n10471), .ZN(n7980) );
  AOI22_X1 U9654 ( .A1(n10472), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n9040), .B2(
        n7978), .ZN(n7979) );
  OAI211_X1 U9655 ( .C1(n8001), .C2(n9024), .A(n7980), .B(n7979), .ZN(P2_U3220) );
  INV_X1 U9656 ( .A(n8078), .ZN(n9025) );
  INV_X1 U9657 ( .A(n7981), .ZN(n7983) );
  XNOR2_X1 U9658 ( .A(n8078), .B(n8569), .ZN(n8533) );
  XNOR2_X1 U9659 ( .A(n8533), .B(n8730), .ZN(n7982) );
  INV_X1 U9660 ( .A(n8535), .ZN(n7986) );
  NOR3_X1 U9661 ( .A1(n7984), .A2(n7983), .A3(n7982), .ZN(n7985) );
  OAI21_X1 U9662 ( .B1(n7986), .B2(n7985), .A(n8693), .ZN(n7990) );
  NAND2_X1 U9663 ( .A1(n8715), .A2(n8731), .ZN(n7987) );
  NAND2_X1 U9664 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8768) );
  OAI211_X1 U9665 ( .C1(n8536), .C2(n8717), .A(n7987), .B(n8768), .ZN(n7988)
         );
  AOI21_X1 U9666 ( .B1(n9029), .B2(n8720), .A(n7988), .ZN(n7989) );
  OAI211_X1 U9667 ( .C1(n9025), .C2(n8724), .A(n7990), .B(n7989), .ZN(P2_U3155) );
  INV_X1 U9668 ( .A(n7991), .ZN(n7995) );
  OAI222_X1 U9669 ( .A1(n9758), .A2(n7995), .B1(P1_U3086), .B2(n7993), .C1(
        n7992), .C2(n9754), .ZN(P1_U3331) );
  OAI222_X1 U9670 ( .A1(n7996), .A2(P2_U3151), .B1(n8098), .B2(n7995), .C1(
        n7994), .C2(n9167), .ZN(P2_U3271) );
  MUX2_X1 U9671 ( .A(n7999), .B(P2_REG1_REG_13__SCAN_IN), .S(n10568), .Z(n7998) );
  NAND2_X1 U9672 ( .A1(n10570), .A2(n10544), .ZN(n9093) );
  OAI22_X1 U9673 ( .A1(n8001), .A2(n9093), .B1(n8000), .B2(n9078), .ZN(n7997)
         );
  OR2_X1 U9674 ( .A1(n7998), .A2(n7997), .ZN(P2_U3472) );
  MUX2_X1 U9675 ( .A(n7999), .B(P2_REG0_REG_13__SCAN_IN), .S(n10547), .Z(n8003) );
  NAND2_X1 U9676 ( .A1(n10545), .A2(n10544), .ZN(n9161) );
  OAI22_X1 U9677 ( .A1(n8001), .A2(n9161), .B1(n8000), .B2(n9143), .ZN(n8002)
         );
  OR2_X1 U9678 ( .A1(n8003), .A2(n8002), .ZN(P2_U3429) );
  XNOR2_X1 U9679 ( .A(n8004), .B(n8005), .ZN(n8034) );
  XNOR2_X1 U9680 ( .A(n9014), .B(n8006), .ZN(n8009) );
  NAND2_X1 U9681 ( .A1(n8730), .A2(n10425), .ZN(n8007) );
  OAI21_X1 U9682 ( .B1(n8718), .B2(n10454), .A(n8007), .ZN(n8008) );
  AOI21_X1 U9683 ( .B1(n8009), .B2(n10443), .A(n8008), .ZN(n8031) );
  MUX2_X1 U9684 ( .A(n8777), .B(n8031), .S(n10471), .Z(n8011) );
  AOI22_X1 U9685 ( .A1(n9012), .A2(n9041), .B1(n9040), .B2(n8721), .ZN(n8010)
         );
  OAI211_X1 U9686 ( .C1(n8034), .C2(n9024), .A(n8011), .B(n8010), .ZN(P2_U3218) );
  INV_X1 U9687 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8012) );
  MUX2_X1 U9688 ( .A(n8012), .B(n8031), .S(n10545), .Z(n8014) );
  INV_X1 U9689 ( .A(n9143), .ZN(n9157) );
  NAND2_X1 U9690 ( .A1(n9012), .A2(n9157), .ZN(n8013) );
  OAI211_X1 U9691 ( .C1(n8034), .C2(n9161), .A(n8014), .B(n8013), .ZN(P2_U3435) );
  INV_X1 U9692 ( .A(n9220), .ZN(n8022) );
  INV_X1 U9693 ( .A(n8015), .ZN(n8016) );
  AOI211_X1 U9694 ( .C1(n8018), .C2(n8017), .A(n10345), .B(n8016), .ZN(n8021)
         );
  NAND2_X1 U9695 ( .A1(n9298), .A2(n10371), .ZN(n8020) );
  NAND2_X1 U9696 ( .A1(n9300), .A2(n10374), .ZN(n8019) );
  NAND2_X1 U9697 ( .A1(n8020), .A2(n8019), .ZN(n9218) );
  OR2_X1 U9698 ( .A1(n8021), .A2(n9218), .ZN(n8109) );
  AOI21_X1 U9699 ( .B1(n8022), .B2(n10271), .A(n8109), .ZN(n8030) );
  INV_X1 U9700 ( .A(n8023), .ZN(n8057) );
  AOI211_X1 U9701 ( .C1(n9222), .C2(n8024), .A(n9626), .B(n8023), .ZN(n8110)
         );
  INV_X1 U9702 ( .A(n9222), .ZN(n8115) );
  OAI22_X1 U9703 ( .A1(n8115), .A2(n9631), .B1(n10261), .B2(n8025), .ZN(n8026)
         );
  AOI21_X1 U9704 ( .B1(n8110), .B2(n10278), .A(n8026), .ZN(n8029) );
  XNOR2_X1 U9705 ( .A(n8027), .B(n8384), .ZN(n8111) );
  NAND2_X1 U9706 ( .A1(n8111), .A2(n10242), .ZN(n8028) );
  OAI211_X1 U9707 ( .C1(n8030), .C2(n10282), .A(n8029), .B(n8028), .ZN(
        P1_U3276) );
  MUX2_X1 U9708 ( .A(n8781), .B(n8031), .S(n10570), .Z(n8033) );
  INV_X1 U9709 ( .A(n9078), .ZN(n9090) );
  NAND2_X1 U9710 ( .A1(n9012), .A2(n9090), .ZN(n8032) );
  OAI211_X1 U9711 ( .C1(n9093), .C2(n8034), .A(n8033), .B(n8032), .ZN(P2_U3474) );
  INV_X1 U9712 ( .A(n8035), .ZN(n8051) );
  INV_X1 U9713 ( .A(n8036), .ZN(n8038) );
  OAI222_X1 U9714 ( .A1(n9758), .A2(n8051), .B1(P1_U3086), .B2(n8038), .C1(
        n8037), .C2(n9754), .ZN(P1_U3330) );
  AOI22_X1 U9715 ( .A1(n8039), .A2(n9241), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8040) );
  OAI21_X1 U9716 ( .B1(n9288), .B2(n8041), .A(n8040), .ZN(n8047) );
  NAND3_X1 U9717 ( .A1(n7948), .A2(n8043), .A3(n4910), .ZN(n8044) );
  AOI21_X1 U9718 ( .B1(n8045), .B2(n8044), .A(n9277), .ZN(n8046) );
  AOI211_X1 U9719 ( .C1(n8048), .C2(n6637), .A(n8047), .B(n8046), .ZN(n8049)
         );
  INV_X1 U9720 ( .A(n8049), .ZN(P1_U3234) );
  OAI222_X1 U9721 ( .A1(n6885), .A2(P2_U3151), .B1(n8098), .B2(n8051), .C1(
        n8050), .C2(n9167), .ZN(P2_U3270) );
  XNOR2_X1 U9722 ( .A(n8052), .B(n8053), .ZN(n8120) );
  INV_X1 U9723 ( .A(n8120), .ZN(n8065) );
  NAND2_X1 U9724 ( .A1(n8054), .A2(n8053), .ZN(n8055) );
  AOI21_X1 U9725 ( .B1(n8056), .B2(n8055), .A(n10345), .ZN(n8118) );
  AOI21_X1 U9726 ( .B1(n9275), .B2(n8057), .A(n9626), .ZN(n8058) );
  NAND2_X1 U9727 ( .A1(n8058), .A2(n8128), .ZN(n8117) );
  OAI22_X1 U9728 ( .A1(n10261), .A2(n9441), .B1(n9271), .B2(n9603), .ZN(n8060)
         );
  NOR2_X1 U9729 ( .A1(n9609), .A2(n9623), .ZN(n8059) );
  AOI211_X1 U9730 ( .C1(n9607), .C2(n9299), .A(n8060), .B(n8059), .ZN(n8062)
         );
  NAND2_X1 U9731 ( .A1(n9275), .A2(n10275), .ZN(n8061) );
  OAI211_X1 U9732 ( .C1(n8117), .C2(n9612), .A(n8062), .B(n8061), .ZN(n8063)
         );
  AOI21_X1 U9733 ( .B1(n8118), .B2(n10261), .A(n8063), .ZN(n8064) );
  OAI21_X1 U9734 ( .B1(n8065), .B2(n9635), .A(n8064), .ZN(P1_U3275) );
  XNOR2_X1 U9735 ( .A(n8066), .B(n8067), .ZN(n9030) );
  INV_X1 U9736 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8074) );
  OR2_X1 U9737 ( .A1(n7919), .A2(n8068), .ZN(n8070) );
  AND2_X1 U9738 ( .A1(n8070), .A2(n8069), .ZN(n8072) );
  XNOR2_X1 U9739 ( .A(n8072), .B(n8071), .ZN(n8073) );
  AOI222_X1 U9740 ( .A1(n10443), .A2(n8073), .B1(n9017), .B2(n10427), .C1(
        n8731), .C2(n10425), .ZN(n9026) );
  MUX2_X1 U9741 ( .A(n8074), .B(n9026), .S(n10570), .Z(n8076) );
  NAND2_X1 U9742 ( .A1(n8078), .A2(n9090), .ZN(n8075) );
  OAI211_X1 U9743 ( .C1(n9093), .C2(n9030), .A(n8076), .B(n8075), .ZN(P2_U3473) );
  INV_X1 U9744 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8077) );
  MUX2_X1 U9745 ( .A(n8077), .B(n9026), .S(n10545), .Z(n8080) );
  NAND2_X1 U9746 ( .A1(n8078), .A2(n9157), .ZN(n8079) );
  OAI211_X1 U9747 ( .C1(n9030), .C2(n9161), .A(n8080), .B(n8079), .ZN(P2_U3432) );
  INV_X1 U9748 ( .A(n8081), .ZN(n8097) );
  INV_X1 U9749 ( .A(n8082), .ZN(n8084) );
  OAI222_X1 U9750 ( .A1(n9758), .A2(n8097), .B1(P1_U3086), .B2(n8084), .C1(
        n8083), .C2(n9754), .ZN(P1_U3329) );
  XOR2_X1 U9751 ( .A(n8087), .B(n8086), .Z(n8088) );
  XNOR2_X1 U9752 ( .A(n8085), .B(n8088), .ZN(n8095) );
  AOI22_X1 U9753 ( .A1(n8090), .A2(n9302), .B1(n9243), .B2(n8089), .ZN(n8091)
         );
  NAND2_X1 U9754 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9368) );
  OAI211_X1 U9755 ( .C1(n8092), .C2(n9287), .A(n8091), .B(n9368), .ZN(n8093)
         );
  AOI21_X1 U9756 ( .B1(n8284), .B2(n6637), .A(n8093), .ZN(n8094) );
  OAI21_X1 U9757 ( .B1(n8095), .B2(n9277), .A(n8094), .ZN(P1_U3241) );
  OAI222_X1 U9758 ( .A1(n8099), .A2(P2_U3151), .B1(n8098), .B2(n8097), .C1(
        n8096), .C2(n9167), .ZN(P2_U3269) );
  NAND2_X1 U9759 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  XOR2_X1 U9760 ( .A(n8103), .B(n8102), .Z(n8108) );
  OAI22_X1 U9761 ( .A1(n9207), .A2(n10356), .B1(n8104), .B2(n10358), .ZN(
        n10206) );
  AOI22_X1 U9762 ( .A1(n10206), .A2(n9241), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8105) );
  OAI21_X1 U9763 ( .B1(n10208), .B2(n9288), .A(n8105), .ZN(n8106) );
  AOI21_X1 U9764 ( .B1(n10210), .B2(n6637), .A(n8106), .ZN(n8107) );
  OAI21_X1 U9765 ( .B1(n8108), .B2(n9277), .A(n8107), .ZN(P1_U3215) );
  AOI211_X1 U9766 ( .C1(n8111), .C2(n10385), .A(n8110), .B(n8109), .ZN(n8113)
         );
  MUX2_X1 U9767 ( .A(n6199), .B(n8113), .S(n10395), .Z(n8112) );
  OAI21_X1 U9768 ( .B1(n8115), .B2(n9747), .A(n8112), .ZN(P1_U3504) );
  MUX2_X1 U9769 ( .A(n9405), .B(n8113), .S(n10413), .Z(n8114) );
  OAI21_X1 U9770 ( .B1(n8115), .B2(n9710), .A(n8114), .ZN(P1_U3539) );
  AOI22_X1 U9771 ( .A1(n10374), .A2(n9299), .B1(n9297), .B2(n10371), .ZN(n8116) );
  NAND2_X1 U9772 ( .A1(n8117), .A2(n8116), .ZN(n8119) );
  AOI211_X1 U9773 ( .C1(n8120), .C2(n10385), .A(n8119), .B(n8118), .ZN(n8122)
         );
  MUX2_X1 U9774 ( .A(n6218), .B(n8122), .S(n10395), .Z(n8121) );
  OAI21_X1 U9775 ( .B1(n6395), .B2(n9747), .A(n8121), .ZN(P1_U3507) );
  MUX2_X1 U9776 ( .A(n9432), .B(n8122), .S(n10413), .Z(n8123) );
  OAI21_X1 U9777 ( .B1(n6395), .B2(n9710), .A(n8123), .ZN(P1_U3540) );
  INV_X1 U9778 ( .A(n6285), .ZN(n8126) );
  AOI21_X1 U9779 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8149), .A(n8124), .ZN(
        n8125) );
  OAI21_X1 U9780 ( .B1(n8126), .B2(n9164), .A(n8125), .ZN(P2_U3268) );
  OAI222_X1 U9781 ( .A1(n9758), .A2(n8126), .B1(n6326), .B2(P1_U3086), .C1(
        n10101), .C2(n9754), .ZN(P1_U3328) );
  XNOR2_X1 U9782 ( .A(n4586), .B(n8385), .ZN(n8127) );
  OAI222_X1 U9783 ( .A1(n10356), .A2(n9188), .B1(n10358), .B2(n9181), .C1(
        n8127), .C2(n10345), .ZN(n9706) );
  INV_X1 U9784 ( .A(n9706), .ZN(n8136) );
  AOI211_X1 U9785 ( .C1(n8129), .C2(n8128), .A(n9626), .B(n9625), .ZN(n9707)
         );
  INV_X1 U9786 ( .A(n8129), .ZN(n9748) );
  NOR2_X1 U9787 ( .A1(n9748), .A2(n9631), .ZN(n8132) );
  OAI22_X1 U9788 ( .A1(n10261), .A2(n8130), .B1(n9180), .B2(n9603), .ZN(n8131)
         );
  AOI211_X1 U9789 ( .C1(n9707), .C2(n10278), .A(n8132), .B(n8131), .ZN(n8135)
         );
  XOR2_X1 U9790 ( .A(n8133), .B(n8385), .Z(n9708) );
  NAND2_X1 U9791 ( .A1(n9708), .A2(n10242), .ZN(n8134) );
  OAI211_X1 U9792 ( .C1(n8136), .C2(n10282), .A(n8135), .B(n8134), .ZN(
        P1_U3274) );
  INV_X1 U9793 ( .A(n8137), .ZN(n8577) );
  AOI21_X1 U9794 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8149), .A(n8138), .ZN(
        n8139) );
  OAI21_X1 U9795 ( .B1(n8577), .B2(n9164), .A(n8139), .ZN(P2_U3267) );
  OAI222_X1 U9796 ( .A1(n9754), .A2(n10072), .B1(n9758), .B2(n8140), .C1(
        P1_U3086), .C2(n6391), .ZN(P1_U3333) );
  NOR4_X1 U9797 ( .A1(n8141), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n6103), .ZN(n8142) );
  AOI21_X1 U9798 ( .B1(n8143), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n8142), .ZN(
        n8144) );
  OAI21_X1 U9799 ( .B1(n8153), .B2(n9758), .A(n8144), .ZN(P1_U3324) );
  INV_X1 U9800 ( .A(n8145), .ZN(n8147) );
  NOR4_X1 U9801 ( .A1(n8147), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8146), .ZN(n8148) );
  AOI21_X1 U9802 ( .B1(n8149), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8148), .ZN(
        n8150) );
  OAI21_X1 U9803 ( .B1(n8153), .B2(n9164), .A(n8150), .ZN(P2_U3264) );
  INV_X1 U9804 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8152) );
  MUX2_X1 U9805 ( .A(n8153), .B(n8152), .S(n8151), .Z(n8154) );
  INV_X1 U9806 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8167) );
  OR2_X1 U9807 ( .A1(n6013), .A2(n9951), .ZN(n8157) );
  INV_X1 U9808 ( .A(n9713), .ZN(n8160) );
  INV_X1 U9809 ( .A(n9471), .ZN(n8159) );
  XNOR2_X1 U9810 ( .A(n8359), .B(n9472), .ZN(n8161) );
  NAND2_X1 U9811 ( .A1(n8161), .A2(n10273), .ZN(n9470) );
  INV_X1 U9812 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U9813 ( .A1(n8162), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U9814 ( .A1(n8163), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8164) );
  OAI211_X1 U9815 ( .C1(n6193), .C2(n8170), .A(n8165), .B(n8164), .ZN(n9295)
         );
  NAND2_X1 U9816 ( .A1(n9295), .A2(n8166), .ZN(n9636) );
  MUX2_X1 U9817 ( .A(n8167), .B(n8169), .S(n10395), .Z(n8168) );
  OAI21_X1 U9818 ( .B1(n8359), .B2(n9747), .A(n8168), .ZN(P1_U3521) );
  MUX2_X1 U9819 ( .A(n8170), .B(n8169), .S(n10413), .Z(n8171) );
  OAI21_X1 U9820 ( .B1(n8359), .B2(n9710), .A(n8171), .ZN(P1_U3553) );
  INV_X1 U9821 ( .A(n9372), .ZN(n8197) );
  MUX2_X1 U9822 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n8172), .S(n8189), .Z(n9357)
         );
  INV_X1 U9823 ( .A(n8188), .ZN(n8210) );
  OAI21_X1 U9824 ( .B1(n8174), .B2(n7440), .A(n8173), .ZN(n8202) );
  MUX2_X1 U9825 ( .A(n8175), .B(P1_REG1_REG_12__SCAN_IN), .S(n8188), .Z(n8203)
         );
  NOR2_X1 U9826 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  AOI21_X1 U9827 ( .B1(n8210), .B2(n8175), .A(n8201), .ZN(n9358) );
  NAND2_X1 U9828 ( .A1(n9357), .A2(n9358), .ZN(n9356) );
  OAI21_X1 U9829 ( .B1(n9372), .B2(n8177), .A(n9356), .ZN(n8176) );
  AOI21_X1 U9830 ( .B1(n9372), .B2(n8177), .A(n8176), .ZN(n8183) );
  NAND2_X1 U9831 ( .A1(n8189), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9832 ( .A1(n8182), .A2(n9356), .ZN(n8180) );
  NAND2_X1 U9833 ( .A1(n9372), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9366) );
  OAI21_X1 U9834 ( .B1(n9372), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9366), .ZN(
        n8178) );
  INV_X1 U9835 ( .A(n8178), .ZN(n8179) );
  NAND2_X1 U9836 ( .A1(n8180), .A2(n8179), .ZN(n9367) );
  INV_X1 U9837 ( .A(n9367), .ZN(n8181) );
  AOI211_X1 U9838 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n9464), .ZN(n8193)
         );
  NAND2_X1 U9839 ( .A1(n8189), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8184) );
  OAI21_X1 U9840 ( .B1(n8189), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8184), .ZN(
        n9360) );
  NOR2_X1 U9841 ( .A1(n8188), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8185) );
  AOI21_X1 U9842 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8188), .A(n8185), .ZN(
        n8200) );
  OAI21_X1 U9843 ( .B1(n8188), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8198), .ZN(
        n9361) );
  NOR2_X1 U9844 ( .A1(n9360), .A2(n9361), .ZN(n9359) );
  XNOR2_X1 U9845 ( .A(n9372), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n8190) );
  AOI211_X1 U9846 ( .C1(n8191), .C2(n8190), .A(n9371), .B(n9458), .ZN(n8192)
         );
  NOR2_X1 U9847 ( .A1(n8193), .A2(n8192), .ZN(n8196) );
  AND2_X1 U9848 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8194) );
  AOI21_X1 U9849 ( .B1(n9467), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n8194), .ZN(
        n8195) );
  OAI211_X1 U9850 ( .C1(n8197), .C2(n9447), .A(n8196), .B(n8195), .ZN(P1_U3257) );
  OAI21_X1 U9851 ( .B1(n8200), .B2(n8199), .A(n8198), .ZN(n8206) );
  AOI21_X1 U9852 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8204) );
  NOR2_X1 U9853 ( .A1(n9464), .A2(n8204), .ZN(n8205) );
  AOI21_X1 U9854 ( .B1(n9462), .B2(n8206), .A(n8205), .ZN(n8209) );
  AOI21_X1 U9855 ( .B1(n9467), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8207), .ZN(
        n8208) );
  OAI211_X1 U9856 ( .C1(n8210), .C2(n9447), .A(n8209), .B(n8208), .ZN(P1_U3255) );
  INV_X1 U9857 ( .A(n8211), .ZN(n8215) );
  MUX2_X1 U9858 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10399), .S(n8224), .Z(n8214)
         );
  INV_X1 U9859 ( .A(n8212), .ZN(n8213) );
  AOI211_X1 U9860 ( .C1(n8215), .C2(n8214), .A(n8213), .B(n9464), .ZN(n8220)
         );
  AOI211_X1 U9861 ( .C1(n8218), .C2(n8217), .A(n8216), .B(n9458), .ZN(n8219)
         );
  NOR2_X1 U9862 ( .A1(n8220), .A2(n8219), .ZN(n8223) );
  AOI21_X1 U9863 ( .B1(n9467), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n8221), .ZN(
        n8222) );
  OAI211_X1 U9864 ( .C1(n8224), .C2(n9447), .A(n8223), .B(n8222), .ZN(P1_U3246) );
  AND2_X1 U9865 ( .A1(n9724), .A2(n9649), .ZN(n8490) );
  INV_X1 U9866 ( .A(n8490), .ZN(n8413) );
  INV_X1 U9867 ( .A(n8313), .ZN(n8316) );
  INV_X1 U9868 ( .A(n8249), .ZN(n8227) );
  NOR4_X1 U9869 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8508), .ZN(n8255)
         );
  INV_X1 U9870 ( .A(n8251), .ZN(n8232) );
  NAND3_X1 U9871 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(n8254) );
  NAND2_X1 U9872 ( .A1(n8233), .A2(n8351), .ZN(n8239) );
  INV_X1 U9873 ( .A(n8239), .ZN(n8234) );
  AOI21_X1 U9874 ( .B1(n8234), .B2(n8237), .A(n10318), .ZN(n8248) );
  NAND2_X1 U9875 ( .A1(n9305), .A2(n8508), .ZN(n8242) );
  INV_X1 U9876 ( .A(n8242), .ZN(n8235) );
  AOI21_X1 U9877 ( .B1(n8235), .B2(n10323), .A(n8236), .ZN(n8247) );
  NAND3_X1 U9878 ( .A1(n8237), .A2(n8351), .A3(n8236), .ZN(n8238) );
  AOI21_X1 U9879 ( .B1(n8239), .B2(n8238), .A(n10326), .ZN(n8244) );
  NAND3_X1 U9880 ( .A1(n10323), .A2(n10318), .A3(n8508), .ZN(n8241) );
  AOI21_X1 U9881 ( .B1(n8242), .B2(n8241), .A(n8240), .ZN(n8243) );
  NOR2_X1 U9882 ( .A1(n8244), .A2(n8243), .ZN(n8246) );
  OAI211_X1 U9883 ( .C1(n8248), .C2(n8247), .A(n8246), .B(n8245), .ZN(n8253)
         );
  NAND2_X1 U9884 ( .A1(n8250), .A2(n8249), .ZN(n8447) );
  NOR2_X1 U9885 ( .A1(n8251), .A2(n8447), .ZN(n8252) );
  MUX2_X1 U9886 ( .A(n8256), .B(n8369), .S(n8508), .Z(n8260) );
  MUX2_X1 U9887 ( .A(n8258), .B(n8257), .S(n8508), .Z(n8259) );
  INV_X1 U9888 ( .A(n8453), .ZN(n8262) );
  OAI21_X1 U9889 ( .B1(n8272), .B2(n8262), .A(n8261), .ZN(n8263) );
  AOI211_X1 U9890 ( .C1(n8263), .C2(n8273), .A(n8271), .B(n8275), .ZN(n8266)
         );
  INV_X1 U9891 ( .A(n8460), .ZN(n8265) );
  INV_X1 U9892 ( .A(n8274), .ZN(n8264) );
  NOR3_X1 U9893 ( .A1(n8266), .A2(n8265), .A3(n8264), .ZN(n8268) );
  OAI21_X1 U9894 ( .B1(n8268), .B2(n8276), .A(n8267), .ZN(n8269) );
  NAND3_X1 U9895 ( .A1(n8269), .A2(n6165), .A3(n8464), .ZN(n8270) );
  NAND4_X1 U9896 ( .A1(n8270), .A2(n8351), .A3(n8466), .A4(n8467), .ZN(n8288)
         );
  NAND2_X1 U9897 ( .A1(n8274), .A2(n8273), .ZN(n8456) );
  NOR2_X1 U9898 ( .A1(n8276), .A2(n8275), .ZN(n8459) );
  OAI21_X1 U9899 ( .B1(n8277), .B2(n8456), .A(n8459), .ZN(n8279) );
  AOI21_X1 U9900 ( .B1(n8279), .B2(n8460), .A(n8278), .ZN(n8280) );
  NOR3_X1 U9901 ( .A1(n8280), .A2(n8463), .A3(n10202), .ZN(n8283) );
  INV_X1 U9902 ( .A(n8281), .ZN(n8468) );
  OAI22_X1 U9903 ( .A1(n8474), .A2(n8467), .B1(n8508), .B2(n8284), .ZN(n8286)
         );
  NAND3_X1 U9904 ( .A1(n8286), .A2(n9301), .A3(n8476), .ZN(n8287) );
  NAND2_X1 U9905 ( .A1(n8295), .A2(n8472), .ZN(n8291) );
  NAND2_X1 U9906 ( .A1(n8294), .A2(n8477), .ZN(n8290) );
  MUX2_X1 U9907 ( .A(n8291), .B(n8290), .S(n8508), .Z(n8292) );
  AOI21_X1 U9908 ( .B1(n8293), .B2(n8384), .A(n8292), .ZN(n8303) );
  NAND2_X1 U9909 ( .A1(n8484), .A2(n8294), .ZN(n8479) );
  NAND2_X1 U9910 ( .A1(n8296), .A2(n8295), .ZN(n8485) );
  MUX2_X1 U9911 ( .A(n8479), .B(n8485), .S(n8508), .Z(n8302) );
  NAND2_X1 U9912 ( .A1(n8305), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U9913 ( .A1(n8304), .A2(n9297), .ZN(n8297) );
  MUX2_X1 U9914 ( .A(n8298), .B(n8297), .S(n8508), .Z(n8299) );
  OAI21_X1 U9915 ( .B1(n9620), .B2(n8300), .A(n8299), .ZN(n8301) );
  OAI21_X1 U9916 ( .B1(n8303), .B2(n8302), .A(n8301), .ZN(n8311) );
  AND2_X1 U9917 ( .A1(n8307), .A2(n8304), .ZN(n8407) );
  OR2_X1 U9918 ( .A1(n9615), .A2(n9624), .ZN(n8306) );
  AND2_X1 U9919 ( .A1(n8306), .A2(n8305), .ZN(n8481) );
  MUX2_X1 U9920 ( .A(n8407), .B(n8481), .S(n8508), .Z(n8310) );
  INV_X1 U9921 ( .A(n8306), .ZN(n8408) );
  INV_X1 U9922 ( .A(n8307), .ZN(n8308) );
  MUX2_X1 U9923 ( .A(n8408), .B(n8308), .S(n8508), .Z(n8309) );
  AOI21_X1 U9924 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8314) );
  OR2_X1 U9925 ( .A1(n9595), .A2(n9610), .ZN(n8312) );
  AND2_X1 U9926 ( .A1(n8313), .A2(n8312), .ZN(n8396) );
  NAND2_X1 U9927 ( .A1(n8397), .A2(n8315), .ZN(n8404) );
  INV_X1 U9928 ( .A(n8399), .ZN(n8318) );
  INV_X1 U9929 ( .A(n8406), .ZN(n8317) );
  MUX2_X1 U9930 ( .A(n8318), .B(n8317), .S(n8508), .Z(n8319) );
  NOR2_X1 U9931 ( .A1(n8321), .A2(n8320), .ZN(n8326) );
  INV_X1 U9932 ( .A(n8326), .ZN(n8327) );
  NAND3_X1 U9933 ( .A1(n8327), .A2(n8351), .A3(n8413), .ZN(n8328) );
  OAI211_X1 U9934 ( .C1(n8351), .C2(n8413), .A(n8329), .B(n8328), .ZN(n8337)
         );
  INV_X1 U9935 ( .A(n8496), .ZN(n8416) );
  OAI21_X1 U9936 ( .B1(n8337), .B2(n8416), .A(n8335), .ZN(n8334) );
  OAI21_X1 U9937 ( .B1(n8334), .B2(n8338), .A(n8421), .ZN(n8344) );
  NOR2_X1 U9938 ( .A1(n8344), .A2(n9713), .ZN(n8350) );
  INV_X1 U9939 ( .A(n8335), .ZN(n8336) );
  AOI21_X1 U9940 ( .B1(n9713), .B2(n8508), .A(n9295), .ZN(n8340) );
  OAI21_X1 U9941 ( .B1(n8342), .B2(n8351), .A(n8340), .ZN(n8341) );
  INV_X1 U9942 ( .A(n8342), .ZN(n8352) );
  NAND2_X1 U9943 ( .A1(n9296), .A2(n8508), .ZN(n8346) );
  NOR2_X1 U9944 ( .A1(n8352), .A2(n8346), .ZN(n8348) );
  NAND2_X1 U9945 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  OAI211_X1 U9946 ( .C1(n8346), .C2(n9713), .A(n8345), .B(n9295), .ZN(n8347)
         );
  OAI22_X1 U9947 ( .A1(n8349), .A2(n8358), .B1(n8348), .B2(n8347), .ZN(n8356)
         );
  NOR2_X1 U9948 ( .A1(n8350), .A2(n8508), .ZN(n8354) );
  INV_X1 U9949 ( .A(n9296), .ZN(n8391) );
  OAI211_X1 U9950 ( .C1(n8354), .C2(n8353), .A(n8391), .B(n8358), .ZN(n8355)
         );
  NAND2_X1 U9951 ( .A1(n8356), .A2(n8355), .ZN(n8507) );
  NAND2_X1 U9952 ( .A1(n8507), .A2(n6393), .ZN(n8395) );
  OR2_X1 U9953 ( .A1(n9713), .A2(n8391), .ZN(n8425) );
  NAND2_X1 U9954 ( .A1(n8509), .A2(n8425), .ZN(n8502) );
  NAND2_X1 U9955 ( .A1(n8359), .A2(n9295), .ZN(n8504) );
  INV_X1 U9956 ( .A(n8456), .ZN(n8375) );
  NOR2_X1 U9957 ( .A1(n8360), .A2(n10238), .ZN(n8368) );
  NOR2_X1 U9958 ( .A1(n8361), .A2(n8362), .ZN(n8367) );
  NAND2_X1 U9959 ( .A1(n8363), .A2(n6325), .ZN(n8364) );
  NOR2_X1 U9960 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  NAND4_X1 U9961 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n10248), .ZN(n8370)
         );
  NOR2_X1 U9962 ( .A1(n8370), .A2(n8369), .ZN(n8371) );
  AND4_X1 U9963 ( .A1(n8372), .A2(n8457), .A3(n8371), .A4(n8453), .ZN(n8374)
         );
  NAND4_X1 U9964 ( .A1(n8376), .A2(n8375), .A3(n8374), .A4(n8373), .ZN(n8377)
         );
  OR4_X1 U9965 ( .A1(n8379), .A2(n8378), .A3(n10202), .A4(n8377), .ZN(n8380)
         );
  NOR2_X1 U9966 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  NAND4_X1 U9967 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), .ZN(n8386)
         );
  NOR2_X1 U9968 ( .A1(n9620), .A2(n8386), .ZN(n8387) );
  NAND4_X1 U9969 ( .A1(n9574), .A2(n8387), .A3(n9585), .A4(n9602), .ZN(n8388)
         );
  NOR2_X1 U9970 ( .A1(n9557), .A2(n8388), .ZN(n8389) );
  NAND4_X1 U9971 ( .A1(n9514), .A2(n9546), .A3(n8389), .A4(n9523), .ZN(n8390)
         );
  NOR2_X1 U9972 ( .A1(n9488), .A2(n8390), .ZN(n8392) );
  NAND2_X1 U9973 ( .A1(n9713), .A2(n8391), .ZN(n8420) );
  NAND4_X1 U9974 ( .A1(n8504), .A2(n8393), .A3(n8392), .A4(n8420), .ZN(n8394)
         );
  NOR2_X1 U9975 ( .A1(n8502), .A2(n8394), .ZN(n8432) );
  AOI21_X1 U9976 ( .B1(n8395), .B2(n8439), .A(n8432), .ZN(n8437) );
  INV_X1 U9977 ( .A(n8396), .ZN(n8398) );
  NAND2_X1 U9978 ( .A1(n8398), .A2(n8397), .ZN(n8400) );
  NAND2_X1 U9979 ( .A1(n8400), .A2(n8399), .ZN(n8401) );
  NAND2_X1 U9980 ( .A1(n8401), .A2(n8406), .ZN(n8402) );
  NAND2_X1 U9981 ( .A1(n8403), .A2(n8402), .ZN(n8412) );
  INV_X1 U9982 ( .A(n8412), .ZN(n8487) );
  NAND3_X1 U9983 ( .A1(n8487), .A2(n8481), .A3(n9621), .ZN(n8415) );
  INV_X1 U9984 ( .A(n8404), .ZN(n8405) );
  OAI211_X1 U9985 ( .C1(n8408), .C2(n8407), .A(n8406), .B(n8405), .ZN(n8409)
         );
  INV_X1 U9986 ( .A(n8409), .ZN(n8411) );
  OAI21_X1 U9987 ( .B1(n8412), .B2(n8411), .A(n8410), .ZN(n8414) );
  NAND2_X1 U9988 ( .A1(n8414), .A2(n8413), .ZN(n8491) );
  OAI211_X1 U9989 ( .C1(n8490), .C2(n8415), .A(n8491), .B(n8488), .ZN(n8417)
         );
  AOI21_X1 U9990 ( .B1(n8492), .B2(n8417), .A(n8416), .ZN(n8424) );
  NAND2_X1 U9991 ( .A1(n8419), .A2(n8418), .ZN(n8438) );
  INV_X1 U9992 ( .A(n8420), .ZN(n8423) );
  INV_X1 U9993 ( .A(n8421), .ZN(n8422) );
  OAI21_X1 U9994 ( .B1(n8424), .B2(n8438), .A(n8497), .ZN(n8428) );
  INV_X1 U9995 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U9996 ( .A1(n8426), .A2(n9295), .ZN(n8427) );
  AOI22_X1 U9997 ( .A1(n8428), .A2(n8427), .B1(n8357), .B2(n9713), .ZN(n8431)
         );
  INV_X1 U9998 ( .A(n8509), .ZN(n8429) );
  AOI211_X1 U9999 ( .C1(n8431), .C2(n8504), .A(n8430), .B(n8429), .ZN(n8433)
         );
  OR2_X1 U10000 ( .A1(n8433), .A2(n8432), .ZN(n8435) );
  OAI211_X1 U10001 ( .C1(n8437), .C2(n7479), .A(n8436), .B(n6390), .ZN(n8515)
         );
  INV_X1 U10002 ( .A(n8438), .ZN(n8500) );
  INV_X1 U10003 ( .A(n10247), .ZN(n8443) );
  NAND3_X1 U10004 ( .A1(n8441), .A2(n8440), .A3(n8439), .ZN(n8442) );
  NAND3_X1 U10005 ( .A1(n8443), .A2(n5135), .A3(n8442), .ZN(n8446) );
  AOI21_X1 U10006 ( .B1(n8446), .B2(n8445), .A(n8444), .ZN(n8448) );
  OAI21_X1 U10007 ( .B1(n8448), .B2(n8447), .A(n4569), .ZN(n8451) );
  AOI21_X1 U10008 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8455) );
  OAI211_X1 U10009 ( .C1(n8455), .C2(n8454), .A(n8453), .B(n8452), .ZN(n8458)
         );
  AOI21_X1 U10010 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8462) );
  INV_X1 U10011 ( .A(n8459), .ZN(n8461) );
  OAI21_X1 U10012 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n8465) );
  AOI21_X1 U10013 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n8469) );
  OAI211_X1 U10014 ( .C1(n8469), .C2(n8468), .A(n8467), .B(n8466), .ZN(n8471)
         );
  NAND2_X1 U10015 ( .A1(n8471), .A2(n8470), .ZN(n8475) );
  INV_X1 U10016 ( .A(n8472), .ZN(n8473) );
  AOI211_X1 U10017 ( .C1(n8476), .C2(n8475), .A(n8474), .B(n8473), .ZN(n8480)
         );
  INV_X1 U10018 ( .A(n8477), .ZN(n8478) );
  NOR3_X1 U10019 ( .A1(n8480), .A2(n8479), .A3(n8478), .ZN(n8483) );
  INV_X1 U10020 ( .A(n8481), .ZN(n8482) );
  AOI211_X1 U10021 ( .C1(n8485), .C2(n8484), .A(n8483), .B(n8482), .ZN(n8486)
         );
  NAND2_X1 U10022 ( .A1(n8487), .A2(n8486), .ZN(n8489) );
  OAI21_X1 U10023 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8494) );
  INV_X1 U10024 ( .A(n8491), .ZN(n8493) );
  OAI21_X1 U10025 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n8495) );
  NAND2_X1 U10026 ( .A1(n8496), .A2(n8495), .ZN(n8499) );
  INV_X1 U10027 ( .A(n8497), .ZN(n8498) );
  AOI21_X1 U10028 ( .B1(n8500), .B2(n8499), .A(n8498), .ZN(n8501) );
  OAI21_X1 U10029 ( .B1(n8502), .B2(n8501), .A(n8504), .ZN(n8503) );
  XOR2_X1 U10030 ( .A(n8434), .B(n8503), .Z(n8513) );
  INV_X1 U10031 ( .A(n8504), .ZN(n8506) );
  AOI211_X1 U10032 ( .C1(n8506), .C2(n8434), .A(n6393), .B(n8505), .ZN(n8511)
         );
  OAI21_X1 U10033 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8510) );
  NAND2_X1 U10034 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  OAI211_X1 U10035 ( .C1(n6393), .C2(n8520), .A(n8518), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8519) );
  OAI21_X1 U10036 ( .B1(n8521), .B2(n8520), .A(n8519), .ZN(P1_U3242) );
  INV_X1 U10037 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8527) );
  XOR2_X1 U10038 ( .A(n8522), .B(n8523), .Z(n8879) );
  XNOR2_X1 U10039 ( .A(n8524), .B(n8523), .ZN(n8525) );
  OAI222_X1 U10040 ( .A1(n10456), .A2(n8526), .B1(n10454), .B2(n8602), .C1(
        n10459), .C2(n8525), .ZN(n8874) );
  AOI21_X1 U10041 ( .B1(n10544), .B2(n8879), .A(n8874), .ZN(n8529) );
  MUX2_X1 U10042 ( .A(n8527), .B(n8529), .S(n10545), .Z(n8528) );
  OAI21_X1 U10043 ( .B1(n8877), .B2(n9143), .A(n8528), .ZN(P2_U3454) );
  MUX2_X1 U10044 ( .A(n8530), .B(n8529), .S(n10570), .Z(n8531) );
  OAI21_X1 U10045 ( .B1(n8877), .B2(n9078), .A(n8531), .ZN(P2_U3486) );
  INV_X1 U10046 ( .A(n8532), .ZN(n8579) );
  OAI222_X1 U10047 ( .A1(n9754), .A2(n9951), .B1(n9758), .B2(n8579), .C1(
        P1_U3086), .C2(n5985), .ZN(P1_U3325) );
  XNOR2_X1 U10048 ( .A(n9012), .B(n8569), .ZN(n8537) );
  INV_X1 U10049 ( .A(n8537), .ZN(n8538) );
  NAND2_X1 U10050 ( .A1(n8533), .A2(n7940), .ZN(n8534) );
  NAND2_X1 U10051 ( .A1(n8535), .A2(n8534), .ZN(n8712) );
  XNOR2_X1 U10052 ( .A(n8537), .B(n8536), .ZN(n8713) );
  NOR2_X1 U10053 ( .A1(n8712), .A2(n8713), .ZN(n8710) );
  XNOR2_X1 U10054 ( .A(n9158), .B(n8569), .ZN(n8539) );
  XNOR2_X1 U10055 ( .A(n8539), .B(n8718), .ZN(n8636) );
  XNOR2_X1 U10056 ( .A(n9151), .B(n8569), .ZN(n8540) );
  NAND2_X1 U10057 ( .A1(n8540), .A2(n8638), .ZN(n8541) );
  OAI21_X1 U10058 ( .B1(n8540), .B2(n8638), .A(n8541), .ZN(n8645) );
  INV_X1 U10059 ( .A(n8541), .ZN(n8692) );
  XNOR2_X1 U10060 ( .A(n8994), .B(n8569), .ZN(n8542) );
  NAND2_X1 U10061 ( .A1(n8542), .A2(n8977), .ZN(n8613) );
  INV_X1 U10062 ( .A(n8542), .ZN(n8543) );
  NAND2_X1 U10063 ( .A1(n8543), .A2(n9003), .ZN(n8544) );
  XNOR2_X1 U10064 ( .A(n8984), .B(n8569), .ZN(n8545) );
  NAND2_X1 U10065 ( .A1(n8545), .A2(n8697), .ZN(n8548) );
  INV_X1 U10066 ( .A(n8545), .ZN(n8546) );
  NAND2_X1 U10067 ( .A1(n8546), .A2(n8988), .ZN(n8547) );
  NAND2_X1 U10068 ( .A1(n8548), .A2(n8547), .ZN(n8612) );
  INV_X1 U10069 ( .A(n8548), .ZN(n8671) );
  XNOR2_X1 U10070 ( .A(n9138), .B(n8569), .ZN(n8549) );
  NAND2_X1 U10071 ( .A1(n8549), .A2(n8978), .ZN(n8620) );
  INV_X1 U10072 ( .A(n8549), .ZN(n8550) );
  INV_X1 U10073 ( .A(n8978), .ZN(n8729) );
  NAND2_X1 U10074 ( .A1(n8550), .A2(n8729), .ZN(n8551) );
  XNOR2_X1 U10075 ( .A(n9072), .B(n8569), .ZN(n8552) );
  XNOR2_X1 U10076 ( .A(n8552), .B(n8932), .ZN(n8621) );
  NAND2_X1 U10077 ( .A1(n8553), .A2(n8951), .ZN(n8682) );
  INV_X1 U10078 ( .A(n8553), .ZN(n8554) );
  NAND2_X1 U10079 ( .A1(n8554), .A2(n8924), .ZN(n8683) );
  NAND2_X1 U10080 ( .A1(n8555), .A2(n8683), .ZN(n8557) );
  XNOR2_X1 U10081 ( .A(n9124), .B(n8556), .ZN(n8558) );
  XNOR2_X1 U10082 ( .A(n8557), .B(n8558), .ZN(n8606) );
  OAI22_X1 U10083 ( .A1(n8606), .A2(n8908), .B1(n8558), .B2(n8557), .ZN(n8651)
         );
  XNOR2_X1 U10084 ( .A(n9118), .B(n8569), .ZN(n8559) );
  XNOR2_X1 U10085 ( .A(n8559), .B(n8923), .ZN(n8652) );
  NAND2_X1 U10086 ( .A1(n8651), .A2(n8652), .ZN(n8562) );
  NAND2_X1 U10087 ( .A1(n8562), .A2(n8561), .ZN(n8629) );
  XNOR2_X1 U10088 ( .A(n9112), .B(n8569), .ZN(n8563) );
  XNOR2_X1 U10089 ( .A(n8563), .B(n8907), .ZN(n8630) );
  NAND2_X1 U10090 ( .A1(n8629), .A2(n8630), .ZN(n8565) );
  NAND2_X1 U10091 ( .A1(n8563), .A2(n8885), .ZN(n8564) );
  XNOR2_X1 U10092 ( .A(n8566), .B(n8569), .ZN(n8567) );
  NAND2_X1 U10093 ( .A1(n8567), .A2(n8895), .ZN(n8702) );
  XNOR2_X1 U10094 ( .A(n8877), .B(n8569), .ZN(n8568) );
  XNOR2_X1 U10095 ( .A(n8568), .B(n8886), .ZN(n8598) );
  XNOR2_X1 U10096 ( .A(n8867), .B(n8569), .ZN(n8570) );
  AOI22_X1 U10097 ( .A1(n8728), .A2(n8715), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8572) );
  NAND2_X1 U10098 ( .A1(n8869), .A2(n8720), .ZN(n8571) );
  OAI211_X1 U10099 ( .C1(n8862), .C2(n8717), .A(n8572), .B(n8571), .ZN(n8573)
         );
  AOI21_X1 U10100 ( .B1(n8574), .B2(n8707), .A(n8573), .ZN(n8575) );
  OAI222_X1 U10101 ( .A1(n9758), .A2(n8577), .B1(P1_U3086), .B2(n4524), .C1(
        n8576), .C2(n9754), .ZN(P1_U3327) );
  OAI222_X1 U10102 ( .A1(n8580), .A2(P2_U3151), .B1(n9164), .B2(n8579), .C1(
        n8578), .C2(n9167), .ZN(P2_U3265) );
  INV_X1 U10103 ( .A(n8581), .ZN(n8582) );
  NAND2_X1 U10104 ( .A1(n8582), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8586) );
  AOI22_X1 U10105 ( .A1(n8693), .A2(n8584), .B1(n8583), .B2(n8707), .ZN(n8585)
         );
  OAI211_X1 U10106 ( .C1(n6810), .C2(n8717), .A(n8586), .B(n8585), .ZN(
        P2_U3172) );
  AND2_X1 U10107 ( .A1(n7536), .A2(n8587), .ZN(n8589) );
  OAI21_X1 U10108 ( .B1(n8589), .B2(n8588), .A(n7539), .ZN(n8590) );
  NAND2_X1 U10109 ( .A1(n8590), .A2(n8693), .ZN(n8597) );
  AOI21_X1 U10110 ( .B1(n8707), .B2(n8592), .A(n8591), .ZN(n8596) );
  AOI22_X1 U10111 ( .A1(n8675), .A2(n8736), .B1(n8715), .B2(n8737), .ZN(n8595)
         );
  NAND2_X1 U10112 ( .A1(n8720), .A2(n8593), .ZN(n8594) );
  NAND4_X1 U10113 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(
        P2_U3153) );
  XNOR2_X1 U10114 ( .A(n8599), .B(n8598), .ZN(n8605) );
  AOI22_X1 U10115 ( .A1(n8895), .A2(n8715), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8601) );
  NAND2_X1 U10116 ( .A1(n8875), .A2(n8720), .ZN(n8600) );
  OAI211_X1 U10117 ( .C1(n8602), .C2(n8717), .A(n8601), .B(n8600), .ZN(n8603)
         );
  AOI21_X1 U10118 ( .B1(n5706), .B2(n8707), .A(n8603), .ZN(n8604) );
  OAI21_X1 U10119 ( .B1(n8605), .B2(n8711), .A(n8604), .ZN(P2_U3154) );
  XNOR2_X1 U10120 ( .A(n8606), .B(n8933), .ZN(n8611) );
  AOI22_X1 U10121 ( .A1(n8924), .A2(n8715), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8608) );
  NAND2_X1 U10122 ( .A1(n8720), .A2(n8927), .ZN(n8607) );
  OAI211_X1 U10123 ( .C1(n8560), .C2(n8717), .A(n8608), .B(n8607), .ZN(n8609)
         );
  AOI21_X1 U10124 ( .B1(n9124), .B2(n8707), .A(n8609), .ZN(n8610) );
  OAI21_X1 U10125 ( .B1(n8611), .B2(n8711), .A(n8610), .ZN(P2_U3156) );
  INV_X1 U10126 ( .A(n8984), .ZN(n9144) );
  AND3_X1 U10127 ( .A1(n8690), .A2(n8613), .A3(n8612), .ZN(n8614) );
  OAI21_X1 U10128 ( .B1(n8672), .B2(n8614), .A(n8693), .ZN(n8619) );
  NAND2_X1 U10129 ( .A1(n8715), .A2(n9003), .ZN(n8616) );
  OAI211_X1 U10130 ( .C1(n8978), .C2(n8717), .A(n8616), .B(n8615), .ZN(n8617)
         );
  AOI21_X1 U10131 ( .B1(n8983), .B2(n8720), .A(n8617), .ZN(n8618) );
  OAI211_X1 U10132 ( .C1(n9144), .C2(n8724), .A(n8619), .B(n8618), .ZN(
        P2_U3159) );
  INV_X1 U10133 ( .A(n9072), .ZN(n8628) );
  AND3_X1 U10134 ( .A1(n8669), .A2(n8621), .A3(n8620), .ZN(n8622) );
  OAI21_X1 U10135 ( .B1(n8623), .B2(n8622), .A(n8693), .ZN(n8627) );
  AOI22_X1 U10136 ( .A1(n8715), .A2(n8729), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8624) );
  OAI21_X1 U10137 ( .B1(n8951), .B2(n8717), .A(n8624), .ZN(n8625) );
  AOI21_X1 U10138 ( .B1(n8952), .B2(n8720), .A(n8625), .ZN(n8626) );
  OAI211_X1 U10139 ( .C1(n8628), .C2(n8724), .A(n8627), .B(n8626), .ZN(
        P2_U3163) );
  XOR2_X1 U10140 ( .A(n8630), .B(n8629), .Z(n8635) );
  AOI22_X1 U10141 ( .A1(n8895), .A2(n8675), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8632) );
  NAND2_X1 U10142 ( .A1(n8720), .A2(n8899), .ZN(n8631) );
  OAI211_X1 U10143 ( .C1(n8560), .C2(n8677), .A(n8632), .B(n8631), .ZN(n8633)
         );
  AOI21_X1 U10144 ( .B1(n9112), .B2(n8707), .A(n8633), .ZN(n8634) );
  OAI21_X1 U10145 ( .B1(n8635), .B2(n8711), .A(n8634), .ZN(P2_U3165) );
  XNOR2_X1 U10146 ( .A(n4611), .B(n8636), .ZN(n8642) );
  NAND2_X1 U10147 ( .A1(n8715), .A2(n9017), .ZN(n8637) );
  NAND2_X1 U10148 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U10149 ( .C1(n8638), .C2(n8717), .A(n8637), .B(n8797), .ZN(n8639)
         );
  AOI21_X1 U10150 ( .B1(n9021), .B2(n8720), .A(n8639), .ZN(n8641) );
  NAND2_X1 U10151 ( .A1(n9158), .A2(n8707), .ZN(n8640) );
  OAI211_X1 U10152 ( .C1(n8642), .C2(n8711), .A(n8641), .B(n8640), .ZN(
        P2_U3166) );
  AOI21_X1 U10153 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8650) );
  NAND2_X1 U10154 ( .A1(n8715), .A2(n9004), .ZN(n8646) );
  NAND2_X1 U10155 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8814) );
  OAI211_X1 U10156 ( .C1(n8977), .C2(n8717), .A(n8646), .B(n8814), .ZN(n8647)
         );
  AOI21_X1 U10157 ( .B1(n9007), .B2(n8720), .A(n8647), .ZN(n8649) );
  NAND2_X1 U10158 ( .A1(n9151), .A2(n8707), .ZN(n8648) );
  OAI211_X1 U10159 ( .C1(n8650), .C2(n8711), .A(n8649), .B(n8648), .ZN(
        P2_U3168) );
  XOR2_X1 U10160 ( .A(n8652), .B(n8651), .Z(n8657) );
  AOI22_X1 U10161 ( .A1(n8907), .A2(n8675), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8654) );
  NAND2_X1 U10162 ( .A1(n8720), .A2(n8912), .ZN(n8653) );
  OAI211_X1 U10163 ( .C1(n8933), .C2(n8677), .A(n8654), .B(n8653), .ZN(n8655)
         );
  AOI21_X1 U10164 ( .B1(n9118), .B2(n8707), .A(n8655), .ZN(n8656) );
  OAI21_X1 U10165 ( .B1(n8657), .B2(n8711), .A(n8656), .ZN(P2_U3169) );
  OAI21_X1 U10166 ( .B1(n8659), .B2(n8658), .A(n7325), .ZN(n8660) );
  NAND2_X1 U10167 ( .A1(n8660), .A2(n8693), .ZN(n8668) );
  INV_X1 U10168 ( .A(n8661), .ZN(n8662) );
  AOI21_X1 U10169 ( .B1(n8707), .B2(n8663), .A(n8662), .ZN(n8667) );
  AOI22_X1 U10170 ( .A1(n8675), .A2(n9035), .B1(n8715), .B2(n8738), .ZN(n8666)
         );
  NAND2_X1 U10171 ( .A1(n8720), .A2(n8664), .ZN(n8665) );
  NAND4_X1 U10172 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(
        P2_U3170) );
  INV_X1 U10173 ( .A(n8669), .ZN(n8674) );
  NOR3_X1 U10174 ( .A1(n8672), .A2(n8671), .A3(n8670), .ZN(n8673) );
  OAI21_X1 U10175 ( .B1(n8674), .B2(n8673), .A(n8693), .ZN(n8680) );
  AOI22_X1 U10176 ( .A1(n8675), .A2(n8963), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8676) );
  OAI21_X1 U10177 ( .B1(n8697), .B2(n8677), .A(n8676), .ZN(n8678) );
  AOI21_X1 U10178 ( .B1(n8966), .B2(n8720), .A(n8678), .ZN(n8679) );
  OAI211_X1 U10179 ( .C1(n8681), .C2(n8724), .A(n8680), .B(n8679), .ZN(
        P2_U3173) );
  NAND2_X1 U10180 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  XOR2_X1 U10181 ( .A(n8684), .B(n4587), .Z(n8689) );
  NAND2_X1 U10182 ( .A1(n8720), .A2(n8941), .ZN(n8686) );
  AOI22_X1 U10183 ( .A1(n8715), .A2(n8963), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8685) );
  OAI211_X1 U10184 ( .C1(n8933), .C2(n8717), .A(n8686), .B(n8685), .ZN(n8687)
         );
  AOI21_X1 U10185 ( .B1(n8940), .B2(n8707), .A(n8687), .ZN(n8688) );
  OAI21_X1 U10186 ( .B1(n8689), .B2(n8711), .A(n8688), .ZN(P2_U3175) );
  INV_X1 U10187 ( .A(n8994), .ZN(n9085) );
  INV_X1 U10188 ( .A(n8690), .ZN(n8695) );
  NOR3_X1 U10189 ( .A1(n8643), .A2(n8692), .A3(n8691), .ZN(n8694) );
  OAI21_X1 U10190 ( .B1(n8695), .B2(n8694), .A(n8693), .ZN(n8700) );
  NAND2_X1 U10191 ( .A1(n8715), .A2(n9018), .ZN(n8696) );
  NAND2_X1 U10192 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8835) );
  OAI211_X1 U10193 ( .C1(n8697), .C2(n8717), .A(n8696), .B(n8835), .ZN(n8698)
         );
  AOI21_X1 U10194 ( .B1(n8990), .B2(n8720), .A(n8698), .ZN(n8699) );
  OAI211_X1 U10195 ( .C1(n9085), .C2(n8724), .A(n8700), .B(n8699), .ZN(
        P2_U3178) );
  NAND2_X1 U10196 ( .A1(n4605), .A2(n8702), .ZN(n8703) );
  XNOR2_X1 U10197 ( .A(n8701), .B(n8703), .ZN(n8709) );
  AOI22_X1 U10198 ( .A1(n8907), .A2(n8715), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8705) );
  NAND2_X1 U10199 ( .A1(n8890), .A2(n8720), .ZN(n8704) );
  OAI211_X1 U10200 ( .C1(n8886), .C2(n8717), .A(n8705), .B(n8704), .ZN(n8706)
         );
  AOI21_X1 U10201 ( .B1(n9106), .B2(n8707), .A(n8706), .ZN(n8708) );
  OAI21_X1 U10202 ( .B1(n8709), .B2(n8711), .A(n8708), .ZN(P2_U3180) );
  INV_X1 U10203 ( .A(n9012), .ZN(n8725) );
  AOI211_X1 U10204 ( .C1(n8713), .C2(n8712), .A(n8711), .B(n8710), .ZN(n8714)
         );
  INV_X1 U10205 ( .A(n8714), .ZN(n8723) );
  NAND2_X1 U10206 ( .A1(n8715), .A2(n8730), .ZN(n8716) );
  NAND2_X1 U10207 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8783) );
  OAI211_X1 U10208 ( .C1(n8718), .C2(n8717), .A(n8716), .B(n8783), .ZN(n8719)
         );
  AOI21_X1 U10209 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8722) );
  OAI211_X1 U10210 ( .C1(n8725), .C2(n8724), .A(n8723), .B(n8722), .ZN(
        P2_U3181) );
  MUX2_X1 U10211 ( .A(n8849), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8831), .Z(
        P2_U3522) );
  MUX2_X1 U10212 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8726), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10213 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8727), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10214 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8728), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10215 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8895), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10216 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8907), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10217 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8923), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10218 ( .A(n8908), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8831), .Z(
        P2_U3514) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8924), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10220 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8963), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8729), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10222 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8988), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10223 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9003), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9018), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10225 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9004), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10226 ( .A(n9017), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8831), .Z(
        P2_U3506) );
  MUX2_X1 U10227 ( .A(n8730), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8831), .Z(
        P2_U3505) );
  MUX2_X1 U10228 ( .A(n8731), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8831), .Z(
        P2_U3504) );
  MUX2_X1 U10229 ( .A(n8732), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8831), .Z(
        P2_U3503) );
  MUX2_X1 U10230 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8733), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10231 ( .A(n8734), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8831), .Z(
        P2_U3501) );
  MUX2_X1 U10232 ( .A(n8735), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8831), .Z(
        P2_U3500) );
  MUX2_X1 U10233 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8736), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10234 ( .A(n9036), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8831), .Z(
        P2_U3498) );
  MUX2_X1 U10235 ( .A(n8737), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8831), .Z(
        P2_U3497) );
  MUX2_X1 U10236 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9035), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10237 ( .A(n10428), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8831), .Z(
        P2_U3495) );
  MUX2_X1 U10238 ( .A(n8738), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8831), .Z(
        P2_U3494) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10426), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7109), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10241 ( .A(n8739), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8831), .Z(
        P2_U3491) );
  AOI21_X1 U10242 ( .B1(n8742), .B2(n8741), .A(n8740), .ZN(n8757) );
  OAI21_X1 U10243 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n8746) );
  NAND2_X1 U10244 ( .A1(n8746), .A2(n10419), .ZN(n8756) );
  AOI21_X1 U10245 ( .B1(n8749), .B2(n8748), .A(n8747), .ZN(n8751) );
  OAI21_X1 U10246 ( .B1(n8837), .B2(n8751), .A(n8750), .ZN(n8753) );
  INV_X1 U10247 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10167) );
  NOR2_X1 U10248 ( .A1(n8816), .A2(n10167), .ZN(n8752) );
  AOI211_X1 U10249 ( .C1(n10415), .C2(n8754), .A(n8753), .B(n8752), .ZN(n8755)
         );
  OAI211_X1 U10250 ( .C1(n8757), .C2(n8846), .A(n8756), .B(n8755), .ZN(
        P2_U3195) );
  AOI21_X1 U10251 ( .B1(n4603), .B2(n8759), .A(n8758), .ZN(n8774) );
  OAI21_X1 U10252 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8772) );
  AOI21_X1 U10253 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8766) );
  NOR2_X1 U10254 ( .A1(n8766), .A2(n8837), .ZN(n8771) );
  INV_X1 U10255 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U10256 ( .A1(n10415), .A2(n8767), .ZN(n8769) );
  OAI211_X1 U10257 ( .C1(n10171), .C2(n8816), .A(n8769), .B(n8768), .ZN(n8770)
         );
  AOI211_X1 U10258 ( .C1(n8772), .C2(n10419), .A(n8771), .B(n8770), .ZN(n8773)
         );
  OAI21_X1 U10259 ( .B1(n8774), .B2(n8846), .A(n8773), .ZN(P2_U3196) );
  AOI21_X1 U10260 ( .B1(n8777), .B2(n8776), .A(n8775), .ZN(n8791) );
  XNOR2_X1 U10261 ( .A(n8779), .B(n8778), .ZN(n8789) );
  AOI21_X1 U10262 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8787) );
  INV_X1 U10263 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10175) );
  OAI21_X1 U10264 ( .B1(n8816), .B2(n10175), .A(n8783), .ZN(n8784) );
  AOI21_X1 U10265 ( .B1(n8785), .B2(n10415), .A(n8784), .ZN(n8786) );
  OAI21_X1 U10266 ( .B1(n8787), .B2(n8837), .A(n8786), .ZN(n8788) );
  AOI21_X1 U10267 ( .B1(n8789), .B2(n10419), .A(n8788), .ZN(n8790) );
  OAI21_X1 U10268 ( .B1(n8791), .B2(n8846), .A(n8790), .ZN(P2_U3197) );
  AOI21_X1 U10269 ( .B1(n4607), .B2(n8793), .A(n8792), .ZN(n8807) );
  XNOR2_X1 U10270 ( .A(n8795), .B(n8794), .ZN(n8805) );
  INV_X1 U10271 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U10272 ( .A1(n10415), .A2(n8796), .ZN(n8798) );
  OAI211_X1 U10273 ( .C1(n10178), .C2(n8816), .A(n8798), .B(n8797), .ZN(n8804)
         );
  AOI21_X1 U10274 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8802) );
  NOR2_X1 U10275 ( .A1(n8802), .A2(n8846), .ZN(n8803) );
  AOI211_X1 U10276 ( .C1(n10419), .C2(n8805), .A(n8804), .B(n8803), .ZN(n8806)
         );
  OAI21_X1 U10277 ( .B1(n8807), .B2(n8837), .A(n8806), .ZN(P2_U3198) );
  AOI21_X1 U10278 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n8824) );
  INV_X1 U10279 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U10280 ( .A1(n8811), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8812) );
  OAI21_X1 U10281 ( .B1(n8813), .B2(n8812), .A(n6725), .ZN(n8815) );
  OAI211_X1 U10282 ( .C1(n10182), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8821)
         );
  XOR2_X1 U10283 ( .A(n8818), .B(n8817), .Z(n8819) );
  NOR2_X1 U10284 ( .A1(n8819), .A2(n8839), .ZN(n8820) );
  AOI211_X1 U10285 ( .C1(n10415), .C2(n8822), .A(n8821), .B(n8820), .ZN(n8823)
         );
  OAI21_X1 U10286 ( .B1(n8824), .B2(n8846), .A(n8823), .ZN(P2_U3199) );
  AOI21_X1 U10287 ( .B1(n4559), .B2(n8826), .A(n8825), .ZN(n8847) );
  INV_X1 U10288 ( .A(n8827), .ZN(n8828) );
  NOR2_X1 U10289 ( .A1(n8829), .A2(n8828), .ZN(n8840) );
  INV_X1 U10290 ( .A(n8840), .ZN(n8832) );
  OAI21_X1 U10291 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8843) );
  AOI21_X1 U10292 ( .B1(n4563), .B2(n8834), .A(n8833), .ZN(n8838) );
  NAND2_X1 U10293 ( .A1(n10414), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8836) );
  OAI211_X1 U10294 ( .C1(n8838), .C2(n8837), .A(n8836), .B(n8835), .ZN(n8842)
         );
  NOR3_X1 U10295 ( .A1(n8840), .A2(n8844), .A3(n8839), .ZN(n8841) );
  AOI211_X1 U10296 ( .C1(n8844), .C2(n8843), .A(n8842), .B(n8841), .ZN(n8845)
         );
  OAI21_X1 U10297 ( .B1(n8847), .B2(n8846), .A(n8845), .ZN(P2_U3200) );
  AND2_X1 U10298 ( .A1(n8849), .A2(n8848), .ZN(n9094) );
  NOR2_X1 U10299 ( .A1(n8850), .A2(n10464), .ZN(n8857) );
  AOI21_X1 U10300 ( .B1(n9094), .B2(n10471), .A(n8857), .ZN(n8853) );
  NAND2_X1 U10301 ( .A1(n10472), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8851) );
  OAI211_X1 U10302 ( .C1(n9096), .C2(n10466), .A(n8853), .B(n8851), .ZN(
        P2_U3202) );
  INV_X1 U10303 ( .A(n9048), .ZN(n9099) );
  NAND2_X1 U10304 ( .A1(n10472), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8852) );
  OAI211_X1 U10305 ( .C1(n9099), .C2(n10466), .A(n8853), .B(n8852), .ZN(
        P2_U3203) );
  NOR2_X1 U10306 ( .A1(n8854), .A2(n10463), .ZN(n8855) );
  OAI21_X1 U10307 ( .B1(n8856), .B2(n8855), .A(n10471), .ZN(n8859) );
  AOI21_X1 U10308 ( .B1(n10472), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8857), .ZN(
        n8858) );
  OAI211_X1 U10309 ( .C1(n8860), .C2(n10466), .A(n8859), .B(n8858), .ZN(
        P2_U3204) );
  INV_X1 U10310 ( .A(n9051), .ZN(n8873) );
  XOR2_X1 U10311 ( .A(n8868), .B(n8867), .Z(n9052) );
  AOI22_X1 U10312 ( .A1(n8869), .A2(n9040), .B1(n10472), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8870) );
  OAI21_X1 U10313 ( .B1(n9103), .B2(n10466), .A(n8870), .ZN(n8871) );
  AOI21_X1 U10314 ( .B1(n9052), .B2(n10433), .A(n8871), .ZN(n8872) );
  OAI21_X1 U10315 ( .B1(n8873), .B2(n10472), .A(n8872), .ZN(P2_U3205) );
  INV_X1 U10316 ( .A(n8874), .ZN(n8881) );
  AOI22_X1 U10317 ( .A1(n8875), .A2(n9040), .B1(n10472), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8876) );
  OAI21_X1 U10318 ( .B1(n8877), .B2(n10466), .A(n8876), .ZN(n8878) );
  AOI21_X1 U10319 ( .B1(n8879), .B2(n10433), .A(n8878), .ZN(n8880) );
  OAI21_X1 U10320 ( .B1(n8881), .B2(n10472), .A(n8880), .ZN(P2_U3206) );
  INV_X1 U10321 ( .A(n8883), .ZN(n8882) );
  XNOR2_X1 U10322 ( .A(n4549), .B(n8882), .ZN(n9109) );
  INV_X1 U10323 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8889) );
  XNOR2_X1 U10324 ( .A(n8884), .B(n8883), .ZN(n8888) );
  OAI22_X1 U10325 ( .A1(n8886), .A2(n10454), .B1(n8885), .B2(n10456), .ZN(
        n8887) );
  AOI21_X1 U10326 ( .B1(n8888), .B2(n10443), .A(n8887), .ZN(n9104) );
  MUX2_X1 U10327 ( .A(n8889), .B(n9104), .S(n10471), .Z(n8892) );
  AOI22_X1 U10328 ( .A1(n9106), .A2(n9041), .B1(n9040), .B2(n8890), .ZN(n8891)
         );
  OAI211_X1 U10329 ( .C1(n9109), .C2(n9024), .A(n8892), .B(n8891), .ZN(
        P2_U3207) );
  INV_X1 U10330 ( .A(n9112), .ZN(n8893) );
  NOR2_X1 U10331 ( .A1(n8893), .A2(n10438), .ZN(n8898) );
  XNOR2_X1 U10332 ( .A(n8894), .B(n8901), .ZN(n8896) );
  AOI222_X1 U10333 ( .A1(n10443), .A2(n8896), .B1(n8895), .B2(n10427), .C1(
        n8923), .C2(n10425), .ZN(n9110) );
  INV_X1 U10334 ( .A(n9110), .ZN(n8897) );
  AOI211_X1 U10335 ( .C1(n9040), .C2(n8899), .A(n8898), .B(n8897), .ZN(n8904)
         );
  XOR2_X1 U10336 ( .A(n8901), .B(n8900), .Z(n9115) );
  INV_X1 U10337 ( .A(n9115), .ZN(n8902) );
  AOI22_X1 U10338 ( .A1(n8902), .A2(n10433), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10472), .ZN(n8903) );
  OAI21_X1 U10339 ( .B1(n8904), .B2(n10472), .A(n8903), .ZN(P2_U3208) );
  INV_X1 U10340 ( .A(n9118), .ZN(n8905) );
  NOR2_X1 U10341 ( .A1(n8905), .A2(n10438), .ZN(n8911) );
  XOR2_X1 U10342 ( .A(n8915), .B(n8906), .Z(n8909) );
  AOI222_X1 U10343 ( .A1(n10443), .A2(n8909), .B1(n8908), .B2(n10425), .C1(
        n8907), .C2(n10427), .ZN(n9116) );
  INV_X1 U10344 ( .A(n9116), .ZN(n8910) );
  AOI211_X1 U10345 ( .C1(n9040), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8919)
         );
  NAND2_X1 U10346 ( .A1(n8914), .A2(n8913), .ZN(n8916) );
  XNOR2_X1 U10347 ( .A(n8916), .B(n8915), .ZN(n9121) );
  INV_X1 U10348 ( .A(n9121), .ZN(n8917) );
  AOI22_X1 U10349 ( .A1(n8917), .A2(n10433), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10472), .ZN(n8918) );
  OAI21_X1 U10350 ( .B1(n8919), .B2(n10472), .A(n8918), .ZN(P2_U3209) );
  XOR2_X1 U10351 ( .A(n8920), .B(n8922), .Z(n9127) );
  INV_X1 U10352 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8926) );
  XNOR2_X1 U10353 ( .A(n8921), .B(n8922), .ZN(n8925) );
  AOI222_X1 U10354 ( .A1(n10443), .A2(n8925), .B1(n8924), .B2(n10425), .C1(
        n8923), .C2(n10427), .ZN(n9122) );
  MUX2_X1 U10355 ( .A(n8926), .B(n9122), .S(n10471), .Z(n8929) );
  AOI22_X1 U10356 ( .A1(n9124), .A2(n9041), .B1(n9040), .B2(n8927), .ZN(n8928)
         );
  OAI211_X1 U10357 ( .C1(n9127), .C2(n9024), .A(n8929), .B(n8928), .ZN(
        P2_U3210) );
  XOR2_X1 U10358 ( .A(n8930), .B(n8938), .Z(n8931) );
  OAI222_X1 U10359 ( .A1(n10454), .A2(n8933), .B1(n10456), .B2(n8932), .C1(
        n10459), .C2(n8931), .ZN(n9067) );
  INV_X1 U10360 ( .A(n9067), .ZN(n8945) );
  NAND2_X1 U10361 ( .A1(n8934), .A2(n8935), .ZN(n8937) );
  NAND2_X1 U10362 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  XNOR2_X1 U10363 ( .A(n8939), .B(n8938), .ZN(n9068) );
  INV_X1 U10364 ( .A(n8940), .ZN(n9131) );
  AOI22_X1 U10365 ( .A1(n10472), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9040), 
        .B2(n8941), .ZN(n8942) );
  OAI21_X1 U10366 ( .B1(n9131), .B2(n10466), .A(n8942), .ZN(n8943) );
  AOI21_X1 U10367 ( .B1(n9068), .B2(n10433), .A(n8943), .ZN(n8944) );
  OAI21_X1 U10368 ( .B1(n8945), .B2(n10472), .A(n8944), .ZN(P2_U3211) );
  NAND2_X1 U10369 ( .A1(n8934), .A2(n8946), .ZN(n8947) );
  XNOR2_X1 U10370 ( .A(n8947), .B(n8948), .ZN(n9135) );
  XOR2_X1 U10371 ( .A(n8949), .B(n8948), .Z(n8950) );
  OAI222_X1 U10372 ( .A1(n10454), .A2(n8951), .B1(n10456), .B2(n8978), .C1(
        n10459), .C2(n8950), .ZN(n9071) );
  NAND2_X1 U10373 ( .A1(n9071), .A2(n10471), .ZN(n8957) );
  INV_X1 U10374 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8954) );
  INV_X1 U10375 ( .A(n8952), .ZN(n8953) );
  OAI22_X1 U10376 ( .A1(n10471), .A2(n8954), .B1(n8953), .B2(n10464), .ZN(
        n8955) );
  AOI21_X1 U10377 ( .B1(n9072), .B2(n9041), .A(n8955), .ZN(n8956) );
  OAI211_X1 U10378 ( .C1(n9135), .C2(n9024), .A(n8957), .B(n8956), .ZN(
        P2_U3212) );
  XNOR2_X1 U10379 ( .A(n8959), .B(n8958), .ZN(n9141) );
  INV_X1 U10380 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8965) );
  OAI21_X1 U10381 ( .B1(n8962), .B2(n8961), .A(n8960), .ZN(n8964) );
  AOI222_X1 U10382 ( .A1(n10443), .A2(n8964), .B1(n8988), .B2(n10425), .C1(
        n8963), .C2(n10427), .ZN(n9136) );
  MUX2_X1 U10383 ( .A(n8965), .B(n9136), .S(n10471), .Z(n8968) );
  AOI22_X1 U10384 ( .A1(n9138), .A2(n9041), .B1(n9040), .B2(n8966), .ZN(n8967)
         );
  OAI211_X1 U10385 ( .C1(n9141), .C2(n9024), .A(n8968), .B(n8967), .ZN(
        P2_U3213) );
  OR2_X1 U10386 ( .A1(n8969), .A2(n8973), .ZN(n8970) );
  NAND2_X1 U10387 ( .A1(n8971), .A2(n8970), .ZN(n9145) );
  NAND2_X1 U10388 ( .A1(n8987), .A2(n8972), .ZN(n8974) );
  NAND2_X1 U10389 ( .A1(n8974), .A2(n8973), .ZN(n8976) );
  NAND3_X1 U10390 ( .A1(n8976), .A2(n10443), .A3(n8975), .ZN(n8981) );
  OAI22_X1 U10391 ( .A1(n8978), .A2(n10454), .B1(n8977), .B2(n10456), .ZN(
        n8979) );
  INV_X1 U10392 ( .A(n8979), .ZN(n8980) );
  NAND2_X1 U10393 ( .A1(n8981), .A2(n8980), .ZN(n9142) );
  MUX2_X1 U10394 ( .A(n9142), .B(P2_REG2_REG_19__SCAN_IN), .S(n10472), .Z(
        n8982) );
  INV_X1 U10395 ( .A(n8982), .ZN(n8986) );
  AOI22_X1 U10396 ( .A1(n8984), .A2(n9041), .B1(n9040), .B2(n8983), .ZN(n8985)
         );
  OAI211_X1 U10397 ( .C1(n9145), .C2(n9024), .A(n8986), .B(n8985), .ZN(
        P2_U3214) );
  OAI21_X1 U10398 ( .B1(n4543), .B2(n8996), .A(n8987), .ZN(n8989) );
  AOI222_X1 U10399 ( .A1(n10443), .A2(n8989), .B1(n8988), .B2(n10427), .C1(
        n9018), .C2(n10425), .ZN(n9084) );
  INV_X1 U10400 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8992) );
  INV_X1 U10401 ( .A(n8990), .ZN(n8991) );
  OAI22_X1 U10402 ( .A1(n10471), .A2(n8992), .B1(n8991), .B2(n10464), .ZN(
        n8993) );
  AOI21_X1 U10403 ( .B1(n8994), .B2(n9041), .A(n8993), .ZN(n8998) );
  NAND2_X1 U10404 ( .A1(n8995), .A2(n8996), .ZN(n9081) );
  NAND3_X1 U10405 ( .A1(n9082), .A2(n9081), .A3(n10433), .ZN(n8997) );
  OAI211_X1 U10406 ( .C1(n9084), .C2(n10472), .A(n8998), .B(n8997), .ZN(
        P2_U3215) );
  XNOR2_X1 U10407 ( .A(n8999), .B(n9001), .ZN(n9154) );
  OAI211_X1 U10408 ( .C1(n9002), .C2(n9001), .A(n9000), .B(n10443), .ZN(n9006)
         );
  AOI22_X1 U10409 ( .A1(n10425), .A2(n9004), .B1(n9003), .B2(n10427), .ZN(
        n9005) );
  MUX2_X1 U10410 ( .A(n9150), .B(n8810), .S(n10472), .Z(n9009) );
  AOI22_X1 U10411 ( .A1(n9151), .A2(n9041), .B1(n9040), .B2(n9007), .ZN(n9008)
         );
  OAI211_X1 U10412 ( .C1(n9154), .C2(n9024), .A(n9009), .B(n9008), .ZN(
        P2_U3216) );
  XNOR2_X1 U10413 ( .A(n9011), .B(n9010), .ZN(n9162) );
  INV_X1 U10414 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9020) );
  OAI22_X1 U10415 ( .A1(n9014), .A2(n9013), .B1(n9017), .B2(n9012), .ZN(n9016)
         );
  XNOR2_X1 U10416 ( .A(n9016), .B(n9015), .ZN(n9019) );
  AOI222_X1 U10417 ( .A1(n10443), .A2(n9019), .B1(n9018), .B2(n10427), .C1(
        n9017), .C2(n10425), .ZN(n9155) );
  MUX2_X1 U10418 ( .A(n9020), .B(n9155), .S(n10471), .Z(n9023) );
  AOI22_X1 U10419 ( .A1(n9158), .A2(n9041), .B1(n9040), .B2(n9021), .ZN(n9022)
         );
  OAI211_X1 U10420 ( .C1(n9162), .C2(n9024), .A(n9023), .B(n9022), .ZN(
        P2_U3217) );
  NOR2_X1 U10421 ( .A1(n9025), .A2(n10438), .ZN(n9028) );
  INV_X1 U10422 ( .A(n9026), .ZN(n9027) );
  AOI211_X1 U10423 ( .C1(n9040), .C2(n9029), .A(n9028), .B(n9027), .ZN(n9033)
         );
  INV_X1 U10424 ( .A(n9030), .ZN(n9031) );
  AOI22_X1 U10425 ( .A1(n9031), .A2(n10433), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n10472), .ZN(n9032) );
  OAI21_X1 U10426 ( .B1(n9033), .B2(n10472), .A(n9032), .ZN(P2_U3219) );
  XNOR2_X1 U10427 ( .A(n9034), .B(n9042), .ZN(n9037) );
  AOI222_X1 U10428 ( .A1(n10443), .A2(n9037), .B1(n9036), .B2(n10427), .C1(
        n9035), .C2(n10425), .ZN(n10502) );
  MUX2_X1 U10429 ( .A(n9038), .B(n10502), .S(n10471), .Z(n9046) );
  AOI22_X1 U10430 ( .A1(n9041), .A2(n10505), .B1(n9040), .B2(n9039), .ZN(n9045) );
  OR2_X1 U10431 ( .A1(n9043), .A2(n9042), .ZN(n10501) );
  NAND3_X1 U10432 ( .A1(n10501), .A2(n10500), .A3(n10433), .ZN(n9044) );
  NAND3_X1 U10433 ( .A1(n9046), .A2(n9045), .A3(n9044), .ZN(P2_U3227) );
  NAND2_X1 U10434 ( .A1(n10568), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10435 ( .A1(n9094), .A2(n10570), .ZN(n9049) );
  OAI211_X1 U10436 ( .C1(n9096), .C2(n9078), .A(n9047), .B(n9049), .ZN(
        P2_U3490) );
  NAND2_X1 U10437 ( .A1(n9048), .A2(n9090), .ZN(n9050) );
  OAI211_X1 U10438 ( .C1(n10570), .C2(n5737), .A(n9050), .B(n9049), .ZN(
        P2_U3489) );
  AOI21_X1 U10439 ( .B1(n9052), .B2(n10544), .A(n9051), .ZN(n9100) );
  MUX2_X1 U10440 ( .A(n9053), .B(n9100), .S(n10570), .Z(n9054) );
  OAI21_X1 U10441 ( .B1(n9103), .B2(n9078), .A(n9054), .ZN(P2_U3487) );
  MUX2_X1 U10442 ( .A(n9055), .B(n9104), .S(n10570), .Z(n9057) );
  NAND2_X1 U10443 ( .A1(n9106), .A2(n9090), .ZN(n9056) );
  OAI211_X1 U10444 ( .C1(n9109), .C2(n9093), .A(n9057), .B(n9056), .ZN(
        P2_U3485) );
  MUX2_X1 U10445 ( .A(n9058), .B(n9110), .S(n10570), .Z(n9060) );
  NAND2_X1 U10446 ( .A1(n9112), .A2(n9090), .ZN(n9059) );
  OAI211_X1 U10447 ( .C1(n9115), .C2(n9093), .A(n9060), .B(n9059), .ZN(
        P2_U3484) );
  MUX2_X1 U10448 ( .A(n9061), .B(n9116), .S(n10570), .Z(n9063) );
  NAND2_X1 U10449 ( .A1(n9118), .A2(n9090), .ZN(n9062) );
  OAI211_X1 U10450 ( .C1(n9093), .C2(n9121), .A(n9063), .B(n9062), .ZN(
        P2_U3483) );
  MUX2_X1 U10451 ( .A(n9064), .B(n9122), .S(n10570), .Z(n9066) );
  NAND2_X1 U10452 ( .A1(n9124), .A2(n9090), .ZN(n9065) );
  OAI211_X1 U10453 ( .C1(n9127), .C2(n9093), .A(n9066), .B(n9065), .ZN(
        P2_U3482) );
  INV_X1 U10454 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9069) );
  AOI21_X1 U10455 ( .B1(n10544), .B2(n9068), .A(n9067), .ZN(n9128) );
  MUX2_X1 U10456 ( .A(n9069), .B(n9128), .S(n10570), .Z(n9070) );
  OAI21_X1 U10457 ( .B1(n9131), .B2(n9078), .A(n9070), .ZN(P2_U3481) );
  INV_X1 U10458 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9073) );
  AOI21_X1 U10459 ( .B1(n10537), .B2(n9072), .A(n9071), .ZN(n9132) );
  MUX2_X1 U10460 ( .A(n9073), .B(n9132), .S(n10570), .Z(n9074) );
  OAI21_X1 U10461 ( .B1(n9093), .B2(n9135), .A(n9074), .ZN(P2_U3480) );
  INV_X1 U10462 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9075) );
  MUX2_X1 U10463 ( .A(n9075), .B(n9136), .S(n10570), .Z(n9077) );
  NAND2_X1 U10464 ( .A1(n9138), .A2(n9090), .ZN(n9076) );
  OAI211_X1 U10465 ( .C1(n9141), .C2(n9093), .A(n9077), .B(n9076), .ZN(
        P2_U3479) );
  MUX2_X1 U10466 ( .A(n9142), .B(P2_REG1_REG_19__SCAN_IN), .S(n10568), .Z(
        n9080) );
  OAI22_X1 U10467 ( .A1(n9145), .A2(n9093), .B1(n9144), .B2(n9078), .ZN(n9079)
         );
  OR2_X1 U10468 ( .A1(n9080), .A2(n9079), .ZN(P2_U3478) );
  NAND3_X1 U10469 ( .A1(n9082), .A2(n9081), .A3(n10544), .ZN(n9083) );
  OAI211_X1 U10470 ( .C1(n9085), .C2(n10539), .A(n9084), .B(n9083), .ZN(n9148)
         );
  MUX2_X1 U10471 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9148), .S(n10570), .Z(
        P2_U3477) );
  MUX2_X1 U10472 ( .A(n9150), .B(n9086), .S(n10568), .Z(n9088) );
  NAND2_X1 U10473 ( .A1(n9151), .A2(n9090), .ZN(n9087) );
  OAI211_X1 U10474 ( .C1(n9093), .C2(n9154), .A(n9088), .B(n9087), .ZN(
        P2_U3476) );
  INV_X1 U10475 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9089) );
  MUX2_X1 U10476 ( .A(n9089), .B(n9155), .S(n10570), .Z(n9092) );
  NAND2_X1 U10477 ( .A1(n9158), .A2(n9090), .ZN(n9091) );
  OAI211_X1 U10478 ( .C1(n9162), .C2(n9093), .A(n9092), .B(n9091), .ZN(
        P2_U3475) );
  NAND2_X1 U10479 ( .A1(n10547), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U10480 ( .A1(n9094), .A2(n10545), .ZN(n9098) );
  OAI211_X1 U10481 ( .C1(n9096), .C2(n9143), .A(n9095), .B(n9098), .ZN(
        P2_U3458) );
  NAND2_X1 U10482 ( .A1(n10547), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9097) );
  OAI211_X1 U10483 ( .C1(n9099), .C2(n9143), .A(n9098), .B(n9097), .ZN(
        P2_U3457) );
  INV_X1 U10484 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9101) );
  MUX2_X1 U10485 ( .A(n9101), .B(n9100), .S(n10545), .Z(n9102) );
  OAI21_X1 U10486 ( .B1(n9103), .B2(n9143), .A(n9102), .ZN(P2_U3455) );
  INV_X1 U10487 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9105) );
  MUX2_X1 U10488 ( .A(n9105), .B(n9104), .S(n10545), .Z(n9108) );
  NAND2_X1 U10489 ( .A1(n9106), .A2(n9157), .ZN(n9107) );
  OAI211_X1 U10490 ( .C1(n9109), .C2(n9161), .A(n9108), .B(n9107), .ZN(
        P2_U3453) );
  INV_X1 U10491 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9111) );
  MUX2_X1 U10492 ( .A(n9111), .B(n9110), .S(n10545), .Z(n9114) );
  NAND2_X1 U10493 ( .A1(n9112), .A2(n9157), .ZN(n9113) );
  OAI211_X1 U10494 ( .C1(n9115), .C2(n9161), .A(n9114), .B(n9113), .ZN(
        P2_U3452) );
  INV_X1 U10495 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9117) );
  MUX2_X1 U10496 ( .A(n9117), .B(n9116), .S(n10545), .Z(n9120) );
  NAND2_X1 U10497 ( .A1(n9118), .A2(n9157), .ZN(n9119) );
  OAI211_X1 U10498 ( .C1(n9121), .C2(n9161), .A(n9120), .B(n9119), .ZN(
        P2_U3451) );
  INV_X1 U10499 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9123) );
  MUX2_X1 U10500 ( .A(n9123), .B(n9122), .S(n10545), .Z(n9126) );
  NAND2_X1 U10501 ( .A1(n9124), .A2(n9157), .ZN(n9125) );
  OAI211_X1 U10502 ( .C1(n9127), .C2(n9161), .A(n9126), .B(n9125), .ZN(
        P2_U3450) );
  INV_X1 U10503 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10504 ( .A(n9129), .B(n9128), .S(n10545), .Z(n9130) );
  OAI21_X1 U10505 ( .B1(n9131), .B2(n9143), .A(n9130), .ZN(P2_U3449) );
  INV_X1 U10506 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9133) );
  MUX2_X1 U10507 ( .A(n9133), .B(n9132), .S(n10545), .Z(n9134) );
  OAI21_X1 U10508 ( .B1(n9135), .B2(n9161), .A(n9134), .ZN(P2_U3448) );
  INV_X1 U10509 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9137) );
  MUX2_X1 U10510 ( .A(n9137), .B(n9136), .S(n10545), .Z(n9140) );
  NAND2_X1 U10511 ( .A1(n9138), .A2(n9157), .ZN(n9139) );
  OAI211_X1 U10512 ( .C1(n9141), .C2(n9161), .A(n9140), .B(n9139), .ZN(
        P2_U3447) );
  MUX2_X1 U10513 ( .A(n9142), .B(P2_REG0_REG_19__SCAN_IN), .S(n10547), .Z(
        n9147) );
  OAI22_X1 U10514 ( .A1(n9145), .A2(n9161), .B1(n9144), .B2(n9143), .ZN(n9146)
         );
  OR2_X1 U10515 ( .A1(n9147), .A2(n9146), .ZN(P2_U3446) );
  MUX2_X1 U10516 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9148), .S(n10545), .Z(
        P2_U3444) );
  INV_X1 U10517 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9149) );
  MUX2_X1 U10518 ( .A(n9150), .B(n9149), .S(n10547), .Z(n9153) );
  NAND2_X1 U10519 ( .A1(n9151), .A2(n9157), .ZN(n9152) );
  OAI211_X1 U10520 ( .C1(n9154), .C2(n9161), .A(n9153), .B(n9152), .ZN(
        P2_U3441) );
  INV_X1 U10521 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9156) );
  MUX2_X1 U10522 ( .A(n9156), .B(n9155), .S(n10545), .Z(n9160) );
  NAND2_X1 U10523 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  OAI211_X1 U10524 ( .C1(n9162), .C2(n9161), .A(n9160), .B(n9159), .ZN(
        P2_U3438) );
  INV_X1 U10525 ( .A(n9163), .ZN(n9757) );
  OAI222_X1 U10526 ( .A1(n9167), .A2(n9166), .B1(P2_U3151), .B2(n9165), .C1(
        n9757), .C2(n9164), .ZN(P2_U3266) );
  MUX2_X1 U10527 ( .A(n9168), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10528 ( .A(n9576), .ZN(n9733) );
  OAI21_X1 U10529 ( .B1(n9171), .B2(n9169), .A(n9170), .ZN(n9172) );
  NAND2_X1 U10530 ( .A1(n9172), .A2(n9285), .ZN(n9176) );
  NOR2_X1 U10531 ( .A1(n9287), .A2(n9197), .ZN(n9174) );
  OAI22_X1 U10532 ( .A1(n9289), .A2(n9610), .B1(n9288), .B2(n9571), .ZN(n9173)
         );
  AOI211_X1 U10533 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n9174), 
        .B(n9173), .ZN(n9175) );
  OAI211_X1 U10534 ( .C1(n9733), .C2(n9294), .A(n9176), .B(n9175), .ZN(
        P1_U3216) );
  OAI211_X1 U10535 ( .C1(n9179), .C2(n9178), .A(n9177), .B(n9285), .ZN(n9184)
         );
  AND2_X1 U10536 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9466) );
  OAI22_X1 U10537 ( .A1(n9289), .A2(n9181), .B1(n9288), .B2(n9180), .ZN(n9182)
         );
  AOI211_X1 U10538 ( .C1(n9209), .C2(n9693), .A(n9466), .B(n9182), .ZN(n9183)
         );
  OAI211_X1 U10539 ( .C1(n9748), .C2(n9294), .A(n9184), .B(n9183), .ZN(
        P1_U3219) );
  XNOR2_X1 U10540 ( .A(n9185), .B(n9186), .ZN(n9192) );
  OAI22_X1 U10541 ( .A1(n9287), .A2(n9610), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9187), .ZN(n9190) );
  OAI22_X1 U10542 ( .A1(n9289), .A2(n9188), .B1(n9288), .B2(n9604), .ZN(n9189)
         );
  AOI211_X1 U10543 ( .C1(n9615), .C2(n6637), .A(n9190), .B(n9189), .ZN(n9191)
         );
  OAI21_X1 U10544 ( .B1(n9192), .B2(n9277), .A(n9191), .ZN(P1_U3223) );
  OAI21_X1 U10545 ( .B1(n9194), .B2(n9193), .A(n9281), .ZN(n9195) );
  NAND2_X1 U10546 ( .A1(n9195), .A2(n9285), .ZN(n9201) );
  NOR2_X1 U10547 ( .A1(n9287), .A2(n9196), .ZN(n9199) );
  OAI22_X1 U10548 ( .A1(n9289), .A2(n9197), .B1(n9288), .B2(n9542), .ZN(n9198)
         );
  AOI211_X1 U10549 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n9199), 
        .B(n9198), .ZN(n9200) );
  OAI211_X1 U10550 ( .C1(n9728), .C2(n9294), .A(n9201), .B(n9200), .ZN(
        P1_U3225) );
  OAI21_X1 U10551 ( .B1(n9204), .B2(n9203), .A(n9202), .ZN(n9205) );
  NAND2_X1 U10552 ( .A1(n9205), .A2(n9285), .ZN(n9211) );
  AND2_X1 U10553 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9399) );
  OAI22_X1 U10554 ( .A1(n9289), .A2(n9207), .B1(n9288), .B2(n9206), .ZN(n9208)
         );
  AOI211_X1 U10555 ( .C1(n9209), .C2(n9299), .A(n9399), .B(n9208), .ZN(n9210)
         );
  OAI211_X1 U10556 ( .C1(n10196), .C2(n9294), .A(n9211), .B(n9210), .ZN(
        P1_U3226) );
  INV_X1 U10557 ( .A(n9212), .ZN(n9217) );
  AOI21_X1 U10558 ( .B1(n9216), .B2(n9214), .A(n9213), .ZN(n9215) );
  AOI21_X1 U10559 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9224) );
  NAND2_X1 U10560 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U10561 ( .A1(n9218), .A2(n9241), .ZN(n9219) );
  OAI211_X1 U10562 ( .C1(n9288), .C2(n9220), .A(n9414), .B(n9219), .ZN(n9221)
         );
  AOI21_X1 U10563 ( .B1(n9222), .B2(n6637), .A(n9221), .ZN(n9223) );
  OAI21_X1 U10564 ( .B1(n9224), .B2(n9277), .A(n9223), .ZN(P1_U3228) );
  NOR2_X1 U10565 ( .A1(n9226), .A2(n9225), .ZN(n9229) );
  INV_X1 U10566 ( .A(n9227), .ZN(n9228) );
  AOI21_X1 U10567 ( .B1(n9229), .B2(n9170), .A(n9228), .ZN(n9234) );
  OAI22_X1 U10568 ( .A1(n9287), .A2(n9559), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9230), .ZN(n9232) );
  OAI22_X1 U10569 ( .A1(n9288), .A2(n9553), .B1(n9590), .B2(n9289), .ZN(n9231)
         );
  AOI211_X1 U10570 ( .C1(n6378), .C2(n6637), .A(n9232), .B(n9231), .ZN(n9233)
         );
  OAI21_X1 U10571 ( .B1(n9234), .B2(n9277), .A(n9233), .ZN(P1_U3229) );
  OAI21_X1 U10572 ( .B1(n7173), .B2(n9236), .A(n9235), .ZN(n9237) );
  NAND3_X1 U10573 ( .A1(n4614), .A2(n9285), .A3(n9237), .ZN(n9247) );
  NAND2_X1 U10574 ( .A1(n9307), .A2(n10374), .ZN(n9239) );
  NAND2_X1 U10575 ( .A1(n10323), .A2(n10371), .ZN(n9238) );
  NAND2_X1 U10576 ( .A1(n9239), .A2(n9238), .ZN(n10233) );
  AOI21_X1 U10577 ( .B1(n10233), .B2(n9241), .A(n9240), .ZN(n9246) );
  INV_X1 U10578 ( .A(n9242), .ZN(n10235) );
  NAND2_X1 U10579 ( .A1(n9243), .A2(n10235), .ZN(n9245) );
  NAND2_X1 U10580 ( .A1(n6637), .A2(n10236), .ZN(n9244) );
  NAND4_X1 U10581 ( .A1(n9247), .A2(n9246), .A3(n9245), .A4(n9244), .ZN(
        P1_U3230) );
  XOR2_X1 U10582 ( .A(n9250), .B(n9249), .Z(n9251) );
  XNOR2_X1 U10583 ( .A(n9248), .B(n9251), .ZN(n9257) );
  OAI22_X1 U10584 ( .A1(n9287), .A2(n9624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9252), .ZN(n9255) );
  OAI22_X1 U10585 ( .A1(n9289), .A2(n9623), .B1(n9288), .B2(n9253), .ZN(n9254)
         );
  AOI211_X1 U10586 ( .C1(n9627), .C2(n6637), .A(n9255), .B(n9254), .ZN(n9256)
         );
  OAI21_X1 U10587 ( .B1(n9257), .B2(n9277), .A(n9256), .ZN(P1_U3233) );
  NAND2_X1 U10588 ( .A1(n9259), .A2(n9258), .ZN(n9261) );
  XNOR2_X1 U10589 ( .A(n9261), .B(n9260), .ZN(n9266) );
  OAI22_X1 U10590 ( .A1(n9287), .A2(n9590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9262), .ZN(n9264) );
  OAI22_X1 U10591 ( .A1(n9289), .A2(n9624), .B1(n9288), .B2(n9586), .ZN(n9263)
         );
  AOI211_X1 U10592 ( .C1(n9595), .C2(n6637), .A(n9264), .B(n9263), .ZN(n9265)
         );
  OAI21_X1 U10593 ( .B1(n9266), .B2(n9277), .A(n9265), .ZN(P1_U3235) );
  NAND2_X1 U10594 ( .A1(n9268), .A2(n9267), .ZN(n9269) );
  XOR2_X1 U10595 ( .A(n9270), .B(n9269), .Z(n9278) );
  NAND2_X1 U10596 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9437) );
  OAI21_X1 U10597 ( .B1(n9287), .B2(n9623), .A(n9437), .ZN(n9274) );
  OAI22_X1 U10598 ( .A1(n9289), .A2(n9272), .B1(n9288), .B2(n9271), .ZN(n9273)
         );
  AOI211_X1 U10599 ( .C1(n9275), .C2(n6637), .A(n9274), .B(n9273), .ZN(n9276)
         );
  OAI21_X1 U10600 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(P1_U3238) );
  INV_X1 U10601 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U10602 ( .A1(n9281), .A2(n9280), .ZN(n9283) );
  NAND2_X1 U10603 ( .A1(n9283), .A2(n9282), .ZN(n9286) );
  NAND3_X1 U10604 ( .A1(n9286), .A2(n9285), .A3(n9284), .ZN(n9293) );
  NOR2_X1 U10605 ( .A1(n9287), .A2(n9528), .ZN(n9291) );
  OAI22_X1 U10606 ( .A1(n9289), .A2(n9559), .B1(n9288), .B2(n9524), .ZN(n9290)
         );
  AOI211_X1 U10607 ( .C1(P1_REG3_REG_26__SCAN_IN), .C2(P1_U3086), .A(n9291), 
        .B(n9290), .ZN(n9292) );
  OAI211_X1 U10608 ( .C1(n9724), .C2(n9294), .A(n9293), .B(n9292), .ZN(
        P1_U3240) );
  MUX2_X1 U10609 ( .A(n9295), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9309), .Z(
        P1_U3585) );
  MUX2_X1 U10610 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9296), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10611 ( .A(n9642), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9309), .Z(
        P1_U3583) );
  MUX2_X1 U10612 ( .A(n9650), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9309), .Z(
        P1_U3582) );
  MUX2_X1 U10613 ( .A(n9659), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9309), .Z(
        P1_U3581) );
  MUX2_X1 U10614 ( .A(n9649), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9309), .Z(
        P1_U3580) );
  MUX2_X1 U10615 ( .A(n9658), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9309), .Z(
        P1_U3579) );
  MUX2_X1 U10616 ( .A(n9568), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9309), .Z(
        P1_U3578) );
  MUX2_X1 U10617 ( .A(n9683), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9309), .Z(
        P1_U3577) );
  MUX2_X1 U10618 ( .A(n9692), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9309), .Z(
        P1_U3576) );
  MUX2_X1 U10619 ( .A(n9684), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9309), .Z(
        P1_U3575) );
  MUX2_X1 U10620 ( .A(n9693), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9309), .Z(
        P1_U3574) );
  MUX2_X1 U10621 ( .A(n9297), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9309), .Z(
        P1_U3573) );
  MUX2_X1 U10622 ( .A(n9298), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9309), .Z(
        P1_U3572) );
  MUX2_X1 U10623 ( .A(n9299), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9309), .Z(
        P1_U3571) );
  MUX2_X1 U10624 ( .A(n9300), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9309), .Z(
        P1_U3570) );
  MUX2_X1 U10625 ( .A(n9301), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9309), .Z(
        P1_U3569) );
  MUX2_X1 U10626 ( .A(n9302), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9309), .Z(
        P1_U3568) );
  MUX2_X1 U10627 ( .A(n10372), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9309), .Z(
        P1_U3567) );
  MUX2_X1 U10628 ( .A(n9303), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9309), .Z(
        P1_U3566) );
  MUX2_X1 U10629 ( .A(n10373), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9309), .Z(
        P1_U3565) );
  MUX2_X1 U10630 ( .A(n9304), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9309), .Z(
        P1_U3564) );
  MUX2_X1 U10631 ( .A(n10349), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9309), .Z(
        P1_U3563) );
  MUX2_X1 U10632 ( .A(n10341), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9309), .Z(
        P1_U3562) );
  MUX2_X1 U10633 ( .A(n10322), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9309), .Z(
        P1_U3561) );
  MUX2_X1 U10634 ( .A(n9305), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9309), .Z(
        P1_U3560) );
  MUX2_X1 U10635 ( .A(n10323), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9309), .Z(
        P1_U3559) );
  MUX2_X1 U10636 ( .A(n9306), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9309), .Z(
        P1_U3558) );
  MUX2_X1 U10637 ( .A(n9307), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9309), .Z(
        P1_U3557) );
  MUX2_X1 U10638 ( .A(n9308), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9309), .Z(
        P1_U3556) );
  MUX2_X1 U10639 ( .A(n9310), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9309), .Z(
        P1_U3555) );
  OAI211_X1 U10640 ( .C1(n9313), .C2(n9312), .A(n9462), .B(n9311), .ZN(n9324)
         );
  AOI22_X1 U10641 ( .A1(n9467), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9323) );
  NAND2_X1 U10642 ( .A1(n9460), .A2(n9314), .ZN(n9322) );
  INV_X1 U10643 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9317) );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7008), .S(n9315), .Z(n9316)
         );
  OAI21_X1 U10645 ( .B1(n9318), .B2(n9317), .A(n9316), .ZN(n9319) );
  NAND3_X1 U10646 ( .A1(n9435), .A2(n9320), .A3(n9319), .ZN(n9321) );
  NAND4_X1 U10647 ( .A1(n9324), .A2(n9323), .A3(n9322), .A4(n9321), .ZN(
        P1_U3244) );
  NOR2_X1 U10648 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9325), .ZN(n9328) );
  NOR2_X1 U10649 ( .A1(n9447), .A2(n9326), .ZN(n9327) );
  AOI211_X1 U10650 ( .C1(n9467), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9328), .B(
        n9327), .ZN(n9338) );
  AOI211_X1 U10651 ( .C1(n9331), .C2(n9330), .A(n9329), .B(n9458), .ZN(n9332)
         );
  INV_X1 U10652 ( .A(n9332), .ZN(n9337) );
  OAI211_X1 U10653 ( .C1(n9335), .C2(n9334), .A(n9435), .B(n9333), .ZN(n9336)
         );
  NAND3_X1 U10654 ( .A1(n9338), .A2(n9337), .A3(n9336), .ZN(P1_U3248) );
  AOI211_X1 U10655 ( .C1(n9341), .C2(n9340), .A(n9339), .B(n9458), .ZN(n9342)
         );
  INV_X1 U10656 ( .A(n9342), .ZN(n9351) );
  AOI21_X1 U10657 ( .B1(n9467), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9343), .ZN(
        n9350) );
  NAND2_X1 U10658 ( .A1(n9460), .A2(n9344), .ZN(n9349) );
  OAI211_X1 U10659 ( .C1(n9347), .C2(n9346), .A(n9435), .B(n9345), .ZN(n9348)
         );
  NAND4_X1 U10660 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(
        P1_U3249) );
  NOR2_X1 U10661 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9352), .ZN(n9355) );
  NOR2_X1 U10662 ( .A1(n9447), .A2(n9353), .ZN(n9354) );
  AOI211_X1 U10663 ( .C1(n9467), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9355), .B(
        n9354), .ZN(n9365) );
  OAI211_X1 U10664 ( .C1(n9358), .C2(n9357), .A(n9435), .B(n9356), .ZN(n9364)
         );
  AOI211_X1 U10665 ( .C1(n9361), .C2(n9360), .A(n9359), .B(n9458), .ZN(n9362)
         );
  INV_X1 U10666 ( .A(n9362), .ZN(n9363) );
  NAND3_X1 U10667 ( .A1(n9365), .A2(n9364), .A3(n9363), .ZN(P1_U3256) );
  NAND2_X1 U10668 ( .A1(n9367), .A2(n9366), .ZN(n9383) );
  XNOR2_X1 U10669 ( .A(n9383), .B(n9373), .ZN(n9381) );
  XNOR2_X1 U10670 ( .A(n9381), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n9380) );
  INV_X1 U10671 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9369) );
  OAI21_X1 U10672 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9378) );
  INV_X1 U10673 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9376) );
  INV_X1 U10674 ( .A(n9374), .ZN(n9375) );
  NOR2_X1 U10675 ( .A1(n9376), .A2(n9375), .ZN(n9395) );
  AOI211_X1 U10676 ( .C1(n9376), .C2(n9375), .A(n9395), .B(n9458), .ZN(n9377)
         );
  AOI211_X1 U10677 ( .C1(n9460), .C2(n9382), .A(n9378), .B(n9377), .ZN(n9379)
         );
  OAI21_X1 U10678 ( .B1(n9380), .B2(n9464), .A(n9379), .ZN(P1_U3258) );
  NAND2_X1 U10679 ( .A1(n9381), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U10680 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  NAND2_X1 U10681 ( .A1(n9385), .A2(n9384), .ZN(n9389) );
  NOR2_X1 U10682 ( .A1(n9417), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9387) );
  AND2_X1 U10683 ( .A1(n9417), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U10684 ( .A1(n9417), .A2(n9390), .ZN(n9388) );
  OAI211_X1 U10685 ( .C1(n9417), .C2(n9390), .A(n9389), .B(n9388), .ZN(n9391)
         );
  AOI21_X1 U10686 ( .B1(n9412), .B2(n9391), .A(n9464), .ZN(n9404) );
  INV_X1 U10687 ( .A(n9417), .ZN(n9402) );
  OR2_X1 U10688 ( .A1(n9417), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U10689 ( .A1(n9417), .A2(n9392), .ZN(n9393) );
  NAND2_X1 U10690 ( .A1(n9394), .A2(n9393), .ZN(n9398) );
  OR2_X1 U10691 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U10692 ( .A1(n9398), .A2(n9397), .ZN(n9419) );
  OAI211_X1 U10693 ( .C1(n9398), .C2(n9397), .A(n9462), .B(n9419), .ZN(n9401)
         );
  AOI21_X1 U10694 ( .B1(n9467), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9399), .ZN(
        n9400) );
  OAI211_X1 U10695 ( .C1(n9447), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9403)
         );
  OR2_X1 U10696 ( .A1(n9404), .A2(n9403), .ZN(P1_U3259) );
  OR2_X1 U10697 ( .A1(n9417), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U10698 ( .A1(n9412), .A2(n9410), .ZN(n9408) );
  OR2_X1 U10699 ( .A1(n9427), .A2(n9405), .ZN(n9407) );
  NAND2_X1 U10700 ( .A1(n9427), .A2(n9405), .ZN(n9406) );
  NAND2_X1 U10701 ( .A1(n9407), .A2(n9406), .ZN(n9409) );
  NAND2_X1 U10702 ( .A1(n9408), .A2(n9409), .ZN(n9429) );
  INV_X1 U10703 ( .A(n9409), .ZN(n9411) );
  NAND3_X1 U10704 ( .A1(n9412), .A2(n9411), .A3(n9410), .ZN(n9413) );
  AOI21_X1 U10705 ( .B1(n9429), .B2(n9413), .A(n9464), .ZN(n9426) );
  NAND2_X1 U10706 ( .A1(n9467), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9415) );
  OAI211_X1 U10707 ( .C1(n9416), .C2(n9447), .A(n9415), .B(n9414), .ZN(n9425)
         );
  NAND2_X1 U10708 ( .A1(n9417), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U10709 ( .A1(n9419), .A2(n9418), .ZN(n9422) );
  OR2_X1 U10710 ( .A1(n9427), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U10711 ( .A1(n9427), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U10712 ( .A1(n9439), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U10713 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  AOI21_X1 U10714 ( .B1(n9440), .B2(n9423), .A(n9458), .ZN(n9424) );
  OR3_X1 U10715 ( .A1(n9426), .A2(n9425), .A3(n9424), .ZN(P1_U3260) );
  OR2_X1 U10716 ( .A1(n9427), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U10717 ( .A1(n9429), .A2(n9428), .ZN(n9434) );
  NOR2_X1 U10718 ( .A1(n9455), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9431) );
  AND2_X1 U10719 ( .A1(n9455), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9430) );
  OR3_X1 U10720 ( .A1(n9434), .A2(n9431), .A3(n9430), .ZN(n9453) );
  NAND2_X1 U10721 ( .A1(n9455), .A2(n9432), .ZN(n9433) );
  OAI211_X1 U10722 ( .C1(n9455), .C2(n9432), .A(n9434), .B(n9433), .ZN(n9436)
         );
  NAND3_X1 U10723 ( .A1(n9453), .A2(n9436), .A3(n9435), .ZN(n9451) );
  INV_X1 U10724 ( .A(n9437), .ZN(n9438) );
  AOI21_X1 U10725 ( .B1(n9467), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9438), .ZN(
        n9450) );
  OR2_X1 U10726 ( .A1(n9455), .A2(n9441), .ZN(n9443) );
  NAND2_X1 U10727 ( .A1(n9455), .A2(n9441), .ZN(n9442) );
  NAND2_X1 U10728 ( .A1(n9443), .A2(n9442), .ZN(n9444) );
  OAI211_X1 U10729 ( .C1(n9445), .C2(n9444), .A(n9462), .B(n9456), .ZN(n9449)
         );
  OR2_X1 U10730 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  NAND4_X1 U10731 ( .A1(n9451), .A2(n9450), .A3(n9449), .A4(n9448), .ZN(
        P1_U3261) );
  NAND2_X1 U10732 ( .A1(n9455), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U10733 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  XNOR2_X1 U10734 ( .A(n9454), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9459) );
  XNOR2_X1 U10735 ( .A(n9457), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9461) );
  INV_X1 U10736 ( .A(n9459), .ZN(n9465) );
  AOI21_X1 U10737 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9463) );
  NOR2_X1 U10738 ( .A1(n10282), .A2(n9636), .ZN(n9474) );
  AOI21_X1 U10739 ( .B1(n10282), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9474), .ZN(
        n9469) );
  NAND2_X1 U10740 ( .A1(n8358), .A2(n10275), .ZN(n9468) );
  OAI211_X1 U10741 ( .C1(n9470), .C2(n9612), .A(n9469), .B(n9468), .ZN(
        P1_U3263) );
  AOI21_X1 U10742 ( .B1(n9713), .B2(n9471), .A(n9626), .ZN(n9473) );
  NAND2_X1 U10743 ( .A1(n9473), .A2(n9472), .ZN(n9637) );
  AOI21_X1 U10744 ( .B1(n10282), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9474), .ZN(
        n9476) );
  NAND2_X1 U10745 ( .A1(n9713), .A2(n10275), .ZN(n9475) );
  OAI211_X1 U10746 ( .C1(n9637), .C2(n9612), .A(n9476), .B(n9475), .ZN(
        P1_U3264) );
  OAI22_X1 U10747 ( .A1(n10261), .A2(n9478), .B1(n9477), .B2(n9603), .ZN(n9479) );
  AOI21_X1 U10748 ( .B1(n9607), .B2(n9650), .A(n9479), .ZN(n9482) );
  NAND2_X1 U10749 ( .A1(n9480), .A2(n10275), .ZN(n9481) );
  OAI211_X1 U10750 ( .C1(n9483), .C2(n9612), .A(n9482), .B(n9481), .ZN(n9484)
         );
  AOI21_X1 U10751 ( .B1(n9485), .B2(n10242), .A(n9484), .ZN(n9486) );
  OAI21_X1 U10752 ( .B1(n9487), .B2(n10282), .A(n9486), .ZN(P1_U3356) );
  OR2_X1 U10753 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  OAI22_X1 U10754 ( .A1(n10261), .A2(n9493), .B1(n9492), .B2(n9603), .ZN(n9494) );
  AOI21_X1 U10755 ( .B1(n9607), .B2(n9659), .A(n9494), .ZN(n9495) );
  OAI21_X1 U10756 ( .B1(n9496), .B2(n9609), .A(n9495), .ZN(n9500) );
  AOI21_X1 U10757 ( .B1(n6387), .B2(n4544), .A(n9626), .ZN(n9497) );
  NAND2_X1 U10758 ( .A1(n9498), .A2(n9497), .ZN(n9644) );
  NOR2_X1 U10759 ( .A1(n9644), .A2(n9612), .ZN(n9499) );
  AOI211_X1 U10760 ( .C1(n10275), .C2(n6387), .A(n9500), .B(n9499), .ZN(n9504)
         );
  XNOR2_X1 U10761 ( .A(n9502), .B(n9501), .ZN(n9641) );
  NAND2_X1 U10762 ( .A1(n9641), .A2(n9516), .ZN(n9503) );
  OAI211_X1 U10763 ( .C1(n9646), .C2(n9635), .A(n9504), .B(n9503), .ZN(
        P1_U3265) );
  XNOR2_X1 U10764 ( .A(n9505), .B(n9514), .ZN(n9653) );
  AOI22_X1 U10765 ( .A1(n10282), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9506), 
        .B2(n10271), .ZN(n9508) );
  NAND2_X1 U10766 ( .A1(n9607), .A2(n9649), .ZN(n9507) );
  OAI211_X1 U10767 ( .C1(n9509), .C2(n9609), .A(n9508), .B(n9507), .ZN(n9512)
         );
  NAND2_X1 U10768 ( .A1(n9513), .A2(n9529), .ZN(n9510) );
  NAND3_X1 U10769 ( .A1(n4544), .A2(n10273), .A3(n9510), .ZN(n9651) );
  NOR2_X1 U10770 ( .A1(n9651), .A2(n9612), .ZN(n9511) );
  AOI211_X1 U10771 ( .C1(n10275), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9518)
         );
  XNOR2_X1 U10772 ( .A(n9515), .B(n9514), .ZN(n9655) );
  NAND2_X1 U10773 ( .A1(n9655), .A2(n9516), .ZN(n9517) );
  OAI211_X1 U10774 ( .C1(n9653), .C2(n9635), .A(n9518), .B(n9517), .ZN(
        P1_U3266) );
  OAI21_X1 U10775 ( .B1(n9520), .B2(n9523), .A(n9519), .ZN(n9521) );
  INV_X1 U10776 ( .A(n9521), .ZN(n9662) );
  XOR2_X1 U10777 ( .A(n9523), .B(n9522), .Z(n9664) );
  NAND2_X1 U10778 ( .A1(n9664), .A2(n10242), .ZN(n9534) );
  OAI22_X1 U10779 ( .A1(n10261), .A2(n9525), .B1(n9524), .B2(n9603), .ZN(n9526) );
  AOI21_X1 U10780 ( .B1(n9607), .B2(n9658), .A(n9526), .ZN(n9527) );
  OAI21_X1 U10781 ( .B1(n9528), .B2(n9609), .A(n9527), .ZN(n9531) );
  OAI211_X1 U10782 ( .C1(n9724), .C2(n9539), .A(n10273), .B(n9529), .ZN(n9660)
         );
  NOR2_X1 U10783 ( .A1(n9660), .A2(n9612), .ZN(n9530) );
  AOI211_X1 U10784 ( .C1(n10275), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  OAI211_X1 U10785 ( .C1(n9662), .C2(n9618), .A(n9534), .B(n9533), .ZN(
        P1_U3267) );
  OAI211_X1 U10786 ( .C1(n9536), .C2(n9546), .A(n9535), .B(n10250), .ZN(n9538)
         );
  AOI22_X1 U10787 ( .A1(n10374), .A2(n9568), .B1(n9649), .B2(n10371), .ZN(
        n9537) );
  NAND2_X1 U10788 ( .A1(n9538), .A2(n9537), .ZN(n9667) );
  INV_X1 U10789 ( .A(n9667), .ZN(n9550) );
  INV_X1 U10790 ( .A(n9552), .ZN(n9540) );
  AOI211_X1 U10791 ( .C1(n9541), .C2(n9540), .A(n9626), .B(n9539), .ZN(n9668)
         );
  NOR2_X1 U10792 ( .A1(n9728), .A2(n9631), .ZN(n9545) );
  OAI22_X1 U10793 ( .A1(n10261), .A2(n9543), .B1(n9542), .B2(n9603), .ZN(n9544) );
  AOI211_X1 U10794 ( .C1(n9668), .C2(n10278), .A(n9545), .B(n9544), .ZN(n9549)
         );
  XNOR2_X1 U10795 ( .A(n9547), .B(n9546), .ZN(n9669) );
  NAND2_X1 U10796 ( .A1(n9669), .A2(n10242), .ZN(n9548) );
  OAI211_X1 U10797 ( .C1(n9550), .C2(n10282), .A(n9549), .B(n9548), .ZN(
        P1_U3268) );
  XOR2_X1 U10798 ( .A(n9551), .B(n9557), .Z(n9675) );
  AOI211_X1 U10799 ( .C1(n6378), .C2(n9572), .A(n9626), .B(n9552), .ZN(n9672)
         );
  INV_X1 U10800 ( .A(n6378), .ZN(n9556) );
  INV_X1 U10801 ( .A(n9553), .ZN(n9554) );
  AOI22_X1 U10802 ( .A1(n10282), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9554), 
        .B2(n10271), .ZN(n9555) );
  OAI21_X1 U10803 ( .B1(n9556), .B2(n9631), .A(n9555), .ZN(n9564) );
  AOI21_X1 U10804 ( .B1(n9558), .B2(n9557), .A(n10345), .ZN(n9562) );
  OAI22_X1 U10805 ( .A1(n9590), .A2(n10358), .B1(n9559), .B2(n10356), .ZN(
        n9560) );
  AOI21_X1 U10806 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9674) );
  NOR2_X1 U10807 ( .A1(n9674), .A2(n10282), .ZN(n9563) );
  AOI211_X1 U10808 ( .C1(n9672), .C2(n10278), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OAI21_X1 U10809 ( .B1(n9635), .B2(n9675), .A(n9565), .ZN(P1_U3269) );
  XNOR2_X1 U10810 ( .A(n9566), .B(n9574), .ZN(n9567) );
  NAND2_X1 U10811 ( .A1(n9567), .A2(n10250), .ZN(n9678) );
  NAND2_X1 U10812 ( .A1(n9692), .A2(n10374), .ZN(n9570) );
  NAND2_X1 U10813 ( .A1(n9568), .A2(n10371), .ZN(n9569) );
  AND2_X1 U10814 ( .A1(n9570), .A2(n9569), .ZN(n9677) );
  OAI211_X1 U10815 ( .C1(n9603), .C2(n9571), .A(n9678), .B(n9677), .ZN(n9580)
         );
  AOI21_X1 U10816 ( .B1(n9576), .B2(n9592), .A(n9626), .ZN(n9573) );
  NAND2_X1 U10817 ( .A1(n9573), .A2(n9572), .ZN(n9676) );
  XNOR2_X1 U10818 ( .A(n9575), .B(n9574), .ZN(n9680) );
  NAND2_X1 U10819 ( .A1(n9680), .A2(n10242), .ZN(n9578) );
  AOI22_X1 U10820 ( .A1(n9576), .A2(n10275), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10282), .ZN(n9577) );
  OAI211_X1 U10821 ( .C1(n9676), .C2(n9612), .A(n9578), .B(n9577), .ZN(n9579)
         );
  AOI21_X1 U10822 ( .B1(n10261), .B2(n9580), .A(n9579), .ZN(n9581) );
  INV_X1 U10823 ( .A(n9581), .ZN(P1_U3270) );
  XNOR2_X1 U10824 ( .A(n9583), .B(n9582), .ZN(n9687) );
  XNOR2_X1 U10825 ( .A(n9584), .B(n9585), .ZN(n9689) );
  NAND2_X1 U10826 ( .A1(n9689), .A2(n10242), .ZN(n9597) );
  OAI22_X1 U10827 ( .A1(n10261), .A2(n9587), .B1(n9586), .B2(n9603), .ZN(n9588) );
  AOI21_X1 U10828 ( .B1(n9607), .B2(n9684), .A(n9588), .ZN(n9589) );
  OAI21_X1 U10829 ( .B1(n9590), .B2(n9609), .A(n9589), .ZN(n9594) );
  OAI211_X1 U10830 ( .C1(n6396), .C2(n9591), .A(n10273), .B(n9592), .ZN(n9685)
         );
  NOR2_X1 U10831 ( .A1(n9685), .A2(n9612), .ZN(n9593) );
  AOI211_X1 U10832 ( .C1(n10275), .C2(n9595), .A(n9594), .B(n9593), .ZN(n9596)
         );
  OAI211_X1 U10833 ( .C1(n9687), .C2(n9618), .A(n9597), .B(n9596), .ZN(
        P1_U3271) );
  OAI21_X1 U10834 ( .B1(n9599), .B2(n9602), .A(n9598), .ZN(n9600) );
  INV_X1 U10835 ( .A(n9600), .ZN(n9696) );
  XOR2_X1 U10836 ( .A(n9602), .B(n9601), .Z(n9698) );
  NAND2_X1 U10837 ( .A1(n9698), .A2(n10242), .ZN(n9617) );
  OAI22_X1 U10838 ( .A1(n10261), .A2(n9605), .B1(n9604), .B2(n9603), .ZN(n9606) );
  AOI21_X1 U10839 ( .B1(n9607), .B2(n9693), .A(n9606), .ZN(n9608) );
  OAI21_X1 U10840 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9614) );
  INV_X1 U10841 ( .A(n9615), .ZN(n9740) );
  OAI211_X1 U10842 ( .C1(n9740), .C2(n4540), .A(n10273), .B(n9611), .ZN(n9694)
         );
  NOR2_X1 U10843 ( .A1(n9694), .A2(n9612), .ZN(n9613) );
  AOI211_X1 U10844 ( .C1(n10275), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9616)
         );
  OAI211_X1 U10845 ( .C1(n9696), .C2(n9618), .A(n9617), .B(n9616), .ZN(
        P1_U3272) );
  XOR2_X1 U10846 ( .A(n9620), .B(n9619), .Z(n9703) );
  INV_X1 U10847 ( .A(n9703), .ZN(n9634) );
  XNOR2_X1 U10848 ( .A(n9621), .B(n9620), .ZN(n9622) );
  OAI222_X1 U10849 ( .A1(n10356), .A2(n9624), .B1(n10358), .B2(n9623), .C1(
        n10345), .C2(n9622), .ZN(n9701) );
  AOI211_X1 U10850 ( .C1(n9627), .C2(n4721), .A(n9626), .B(n4540), .ZN(n9702)
         );
  NAND2_X1 U10851 ( .A1(n9702), .A2(n10278), .ZN(n9630) );
  AOI22_X1 U10852 ( .A1(n10282), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9628), 
        .B2(n10271), .ZN(n9629) );
  OAI211_X1 U10853 ( .C1(n9744), .C2(n9631), .A(n9630), .B(n9629), .ZN(n9632)
         );
  AOI21_X1 U10854 ( .B1(n9701), .B2(n10261), .A(n9632), .ZN(n9633) );
  OAI21_X1 U10855 ( .B1(n9635), .B2(n9634), .A(n9633), .ZN(P1_U3273) );
  INV_X1 U10856 ( .A(n9710), .ZN(n9639) );
  NAND2_X1 U10857 ( .A1(n9637), .A2(n9636), .ZN(n9711) );
  MUX2_X1 U10858 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9711), .S(n10413), .Z(
        n9638) );
  AOI21_X1 U10859 ( .B1(n9639), .B2(n9713), .A(n9638), .ZN(n9640) );
  INV_X1 U10860 ( .A(n9640), .ZN(P1_U3552) );
  INV_X1 U10861 ( .A(n10385), .ZN(n10307) );
  NAND2_X1 U10862 ( .A1(n9641), .A2(n10250), .ZN(n9645) );
  AOI22_X1 U10863 ( .A1(n10374), .A2(n9659), .B1(n9642), .B2(n10371), .ZN(
        n9643) );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9715), .S(n10413), .Z(
        n9647) );
  INV_X1 U10865 ( .A(n9647), .ZN(n9648) );
  OAI21_X1 U10866 ( .B1(n9716), .B2(n9710), .A(n9648), .ZN(P1_U3550) );
  AOI22_X1 U10867 ( .A1(n10371), .A2(n9650), .B1(n9649), .B2(n10374), .ZN(
        n9652) );
  OAI211_X1 U10868 ( .C1(n9653), .C2(n10307), .A(n9652), .B(n9651), .ZN(n9654)
         );
  AOI21_X1 U10869 ( .B1(n9655), .B2(n10250), .A(n9654), .ZN(n9717) );
  MUX2_X1 U10870 ( .A(n9656), .B(n9717), .S(n10413), .Z(n9657) );
  OAI21_X1 U10871 ( .B1(n9720), .B2(n9710), .A(n9657), .ZN(P1_U3549) );
  AOI22_X1 U10872 ( .A1(n10371), .A2(n9659), .B1(n9658), .B2(n10374), .ZN(
        n9661) );
  OAI211_X1 U10873 ( .C1(n9662), .C2(n10345), .A(n9661), .B(n9660), .ZN(n9663)
         );
  AOI21_X1 U10874 ( .B1(n9664), .B2(n10385), .A(n9663), .ZN(n9721) );
  MUX2_X1 U10875 ( .A(n9665), .B(n9721), .S(n10413), .Z(n9666) );
  OAI21_X1 U10876 ( .B1(n9724), .B2(n9710), .A(n9666), .ZN(P1_U3548) );
  AOI211_X1 U10877 ( .C1(n9669), .C2(n10385), .A(n9668), .B(n9667), .ZN(n9725)
         );
  MUX2_X1 U10878 ( .A(n9670), .B(n9725), .S(n10413), .Z(n9671) );
  OAI21_X1 U10879 ( .B1(n9728), .B2(n9710), .A(n9671), .ZN(P1_U3547) );
  AOI21_X1 U10880 ( .B1(n10363), .B2(n6378), .A(n9672), .ZN(n9673) );
  OAI211_X1 U10881 ( .C1(n9675), .C2(n10307), .A(n9674), .B(n9673), .ZN(n9729)
         );
  MUX2_X1 U10882 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9729), .S(n10413), .Z(
        P1_U3546) );
  NAND3_X1 U10883 ( .A1(n9678), .A2(n9677), .A3(n9676), .ZN(n9679) );
  AOI21_X1 U10884 ( .B1(n9680), .B2(n10385), .A(n9679), .ZN(n9730) );
  MUX2_X1 U10885 ( .A(n9681), .B(n9730), .S(n10413), .Z(n9682) );
  OAI21_X1 U10886 ( .B1(n9733), .B2(n9710), .A(n9682), .ZN(P1_U3545) );
  AOI22_X1 U10887 ( .A1(n10374), .A2(n9684), .B1(n9683), .B2(n10371), .ZN(
        n9686) );
  OAI211_X1 U10888 ( .C1(n9687), .C2(n10345), .A(n9686), .B(n9685), .ZN(n9688)
         );
  AOI21_X1 U10889 ( .B1(n10385), .B2(n9689), .A(n9688), .ZN(n9734) );
  MUX2_X1 U10890 ( .A(n9690), .B(n9734), .S(n10413), .Z(n9691) );
  OAI21_X1 U10891 ( .B1(n6396), .B2(n9710), .A(n9691), .ZN(P1_U3544) );
  AOI22_X1 U10892 ( .A1(n10374), .A2(n9693), .B1(n9692), .B2(n10371), .ZN(
        n9695) );
  OAI211_X1 U10893 ( .C1(n9696), .C2(n10345), .A(n9695), .B(n9694), .ZN(n9697)
         );
  AOI21_X1 U10894 ( .B1(n9698), .B2(n10385), .A(n9697), .ZN(n9737) );
  MUX2_X1 U10895 ( .A(n9699), .B(n9737), .S(n10413), .Z(n9700) );
  OAI21_X1 U10896 ( .B1(n9740), .B2(n9710), .A(n9700), .ZN(P1_U3543) );
  AOI211_X1 U10897 ( .C1(n9703), .C2(n10385), .A(n9702), .B(n9701), .ZN(n9741)
         );
  MUX2_X1 U10898 ( .A(n9704), .B(n9741), .S(n10413), .Z(n9705) );
  OAI21_X1 U10899 ( .B1(n9744), .B2(n9710), .A(n9705), .ZN(P1_U3542) );
  AOI211_X1 U10900 ( .C1(n10385), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9745)
         );
  MUX2_X1 U10901 ( .A(n6227), .B(n9745), .S(n10413), .Z(n9709) );
  OAI21_X1 U10902 ( .B1(n9748), .B2(n9710), .A(n9709), .ZN(P1_U3541) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9711), .S(n10395), .Z(
        n9712) );
  AOI21_X1 U10904 ( .B1(n6660), .B2(n9713), .A(n9712), .ZN(n9714) );
  INV_X1 U10905 ( .A(n9714), .ZN(P1_U3520) );
  MUX2_X1 U10906 ( .A(n9718), .B(n9717), .S(n10395), .Z(n9719) );
  OAI21_X1 U10907 ( .B1(n9720), .B2(n9747), .A(n9719), .ZN(P1_U3517) );
  MUX2_X1 U10908 ( .A(n9722), .B(n9721), .S(n10395), .Z(n9723) );
  OAI21_X1 U10909 ( .B1(n9724), .B2(n9747), .A(n9723), .ZN(P1_U3516) );
  MUX2_X1 U10910 ( .A(n9726), .B(n9725), .S(n10395), .Z(n9727) );
  OAI21_X1 U10911 ( .B1(n9728), .B2(n9747), .A(n9727), .ZN(P1_U3515) );
  MUX2_X1 U10912 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9729), .S(n10395), .Z(
        P1_U3514) );
  MUX2_X1 U10913 ( .A(n9731), .B(n9730), .S(n10395), .Z(n9732) );
  OAI21_X1 U10914 ( .B1(n9733), .B2(n9747), .A(n9732), .ZN(P1_U3513) );
  MUX2_X1 U10915 ( .A(n9735), .B(n9734), .S(n10395), .Z(n9736) );
  OAI21_X1 U10916 ( .B1(n6396), .B2(n9747), .A(n9736), .ZN(P1_U3512) );
  MUX2_X1 U10917 ( .A(n9738), .B(n9737), .S(n10395), .Z(n9739) );
  OAI21_X1 U10918 ( .B1(n9740), .B2(n9747), .A(n9739), .ZN(P1_U3511) );
  MUX2_X1 U10919 ( .A(n9742), .B(n9741), .S(n10395), .Z(n9743) );
  OAI21_X1 U10920 ( .B1(n9744), .B2(n9747), .A(n9743), .ZN(P1_U3510) );
  MUX2_X1 U10921 ( .A(n6229), .B(n9745), .S(n10395), .Z(n9746) );
  OAI21_X1 U10922 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(P1_U3509) );
  INV_X1 U10923 ( .A(n9749), .ZN(n9751) );
  AND2_X1 U10924 ( .A1(n9751), .A2(n9750), .ZN(n10288) );
  MUX2_X1 U10925 ( .A(P1_D_REG_1__SCAN_IN), .B(n9752), .S(n10288), .Z(P1_U3440) );
  MUX2_X1 U10926 ( .A(P1_D_REG_0__SCAN_IN), .B(n9753), .S(n10288), .Z(P1_U3439) );
  OAI222_X1 U10927 ( .A1(n9758), .A2(n9757), .B1(n9756), .B2(P1_U3086), .C1(
        n9755), .C2(n9754), .ZN(P1_U3326) );
  MUX2_X1 U10928 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9759), .S(P1_U3086), .Z(
        P1_U3355) );
  OAI22_X1 U10929 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_g80), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .ZN(n9760) );
  AOI221_X1 U10930 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .C1(
        keyinput_g59), .C2(P2_REG3_REG_2__SCAN_IN), .A(n9760), .ZN(n9767) );
  OAI22_X1 U10931 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g107), .ZN(n9761) );
  AOI221_X1 U10932 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        keyinput_g107), .C2(P1_IR_REG_17__SCAN_IN), .A(n9761), .ZN(n9766) );
  OAI22_X1 U10933 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        keyinput_g117), .B2(P1_IR_REG_27__SCAN_IN), .ZN(n9762) );
  AOI221_X1 U10934 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_g117), .A(n9762), .ZN(n9765) );
  OAI22_X1 U10935 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g127), .B2(P1_D_REG_5__SCAN_IN), .ZN(n9763) );
  AOI221_X1 U10936 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput_g127), .A(n9763), .ZN(n9764) );
  NAND4_X1 U10937 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n9797)
         );
  OAI22_X1 U10938 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .ZN(n9768) );
  AOI221_X1 U10939 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        keyinput_g86), .C2(P2_DATAO_REG_10__SCAN_IN), .A(n9768), .ZN(n9775) );
  OAI22_X1 U10940 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        keyinput_g125), .B2(P1_D_REG_3__SCAN_IN), .ZN(n9769) );
  AOI221_X1 U10941 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput_g125), .A(n9769), .ZN(n9774) );
  OAI22_X1 U10942 ( .A1(SI_25_), .A2(keyinput_g7), .B1(SI_12_), .B2(
        keyinput_g20), .ZN(n9770) );
  AOI221_X1 U10943 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g20), .C2(
        SI_12_), .A(n9770), .ZN(n9773) );
  OAI22_X1 U10944 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g95), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput_g119), .ZN(n9771) );
  AOI221_X1 U10945 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g95), .C1(
        keyinput_g119), .C2(P1_IR_REG_29__SCAN_IN), .A(n9771), .ZN(n9772) );
  NAND4_X1 U10946 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(n9796)
         );
  OAI22_X1 U10947 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        keyinput_g104), .B2(P1_IR_REG_14__SCAN_IN), .ZN(n9776) );
  AOI221_X1 U10948 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g104), .A(n9776), .ZN(n9783) );
  OAI22_X1 U10949 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        keyinput_g98), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n9777) );
  AOI221_X1 U10950 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g98), .A(n9777), .ZN(n9782) );
  OAI22_X1 U10951 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        keyinput_g87), .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9778) );
  AOI221_X1 U10952 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_g87), .A(n9778), .ZN(n9781) );
  OAI22_X1 U10953 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_g71), .B1(
        keyinput_g81), .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9779) );
  AOI221_X1 U10954 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_g81), .A(n9779), .ZN(n9780) );
  NAND4_X1 U10955 ( .A1(n9783), .A2(n9782), .A3(n9781), .A4(n9780), .ZN(n9795)
         );
  INV_X1 U10956 ( .A(SI_14_), .ZN(n10086) );
  INV_X1 U10957 ( .A(SI_18_), .ZN(n10100) );
  AOI22_X1 U10958 ( .A1(n10086), .A2(keyinput_g18), .B1(n10100), .B2(
        keyinput_g14), .ZN(n9784) );
  OAI221_X1 U10959 ( .B1(n10086), .B2(keyinput_g18), .C1(n10100), .C2(
        keyinput_g14), .A(n9784), .ZN(n9793) );
  AOI22_X1 U10960 ( .A1(n5994), .A2(keyinput_g32), .B1(n9786), .B2(
        keyinput_g45), .ZN(n9785) );
  OAI221_X1 U10961 ( .B1(n5994), .B2(keyinput_g32), .C1(n9786), .C2(
        keyinput_g45), .A(n9785), .ZN(n9792) );
  XOR2_X1 U10962 ( .A(n8152), .B(keyinput_g65), .Z(n9790) );
  XNOR2_X1 U10963 ( .A(SI_6_), .B(keyinput_g26), .ZN(n9789) );
  XNOR2_X1 U10964 ( .A(SI_3_), .B(keyinput_g29), .ZN(n9788) );
  XNOR2_X1 U10965 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9787) );
  NAND4_X1 U10966 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n9791)
         );
  OR3_X1 U10967 ( .A1(n9793), .A2(n9792), .A3(n9791), .ZN(n9794) );
  NOR4_X1 U10968 ( .A1(n9797), .A2(n9796), .A3(n9795), .A4(n9794), .ZN(n10130)
         );
  OAI22_X1 U10969 ( .A1(SI_21_), .A2(keyinput_g11), .B1(keyinput_g16), .B2(
        SI_16_), .ZN(n9798) );
  AOI221_X1 U10970 ( .B1(SI_21_), .B2(keyinput_g11), .C1(SI_16_), .C2(
        keyinput_g16), .A(n9798), .ZN(n9805) );
  OAI22_X1 U10971 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .ZN(n9799) );
  AOI221_X1 U10972 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        keyinput_g66), .C2(P2_DATAO_REG_30__SCAN_IN), .A(n9799), .ZN(n9804) );
  OAI22_X1 U10973 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g99), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_g96), .ZN(n9800) );
  AOI221_X1 U10974 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g99), .C1(
        keyinput_g96), .C2(P1_IR_REG_6__SCAN_IN), .A(n9800), .ZN(n9803) );
  OAI22_X1 U10975 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g68), .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9801) );
  AOI221_X1 U10976 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_g68), .A(n9801), .ZN(n9802) );
  NAND4_X1 U10977 ( .A1(n9805), .A2(n9804), .A3(n9803), .A4(n9802), .ZN(n9935)
         );
  OAI22_X1 U10978 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n9806) );
  AOI221_X1 U10979 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g85), .C2(P2_DATAO_REG_11__SCAN_IN), .A(n9806), .ZN(n9831) );
  OAI22_X1 U10980 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(
        keyinput_g101), .B2(P1_IR_REG_11__SCAN_IN), .ZN(n9807) );
  AOI221_X1 U10981 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g101), .A(n9807), .ZN(n9810) );
  OAI22_X1 U10982 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput_g126), .ZN(n9808) );
  AOI221_X1 U10983 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        keyinput_g126), .C2(P1_D_REG_4__SCAN_IN), .A(n9808), .ZN(n9809) );
  OAI211_X1 U10984 ( .C1(n5444), .C2(keyinput_g53), .A(n9810), .B(n9809), .ZN(
        n9811) );
  AOI21_X1 U10985 ( .B1(n5444), .B2(keyinput_g53), .A(n9811), .ZN(n9830) );
  AOI22_X1 U10986 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_g102), .B1(SI_29_), .B2(keyinput_g3), .ZN(n9812) );
  OAI221_X1 U10987 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_g102), .C1(
        SI_29_), .C2(keyinput_g3), .A(n9812), .ZN(n9819) );
  AOI22_X1 U10988 ( .A1(SI_11_), .A2(keyinput_g21), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n9813) );
  OAI221_X1 U10989 ( .B1(SI_11_), .B2(keyinput_g21), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9813), .ZN(n9818) );
  AOI22_X1 U10990 ( .A1(SI_30_), .A2(keyinput_g2), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .ZN(n9814) );
  OAI221_X1 U10991 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_g70), .A(n9814), .ZN(n9817) );
  AOI22_X1 U10992 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9815) );
  OAI221_X1 U10993 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9815), .ZN(n9816) );
  NOR4_X1 U10994 ( .A1(n9819), .A2(n9818), .A3(n9817), .A4(n9816), .ZN(n9829)
         );
  AOI22_X1 U10995 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n9820) );
  OAI221_X1 U10996 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n9820), .ZN(n9827) );
  AOI22_X1 U10997 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g93), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n9821) );
  OAI221_X1 U10998 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n9821), .ZN(n9826) );
  AOI22_X1 U10999 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_g90), .B1(SI_10_), 
        .B2(keyinput_g22), .ZN(n9822) );
  OAI221_X1 U11000 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_g90), .C1(SI_10_), 
        .C2(keyinput_g22), .A(n9822), .ZN(n9825) );
  AOI22_X1 U11001 ( .A1(SI_17_), .A2(keyinput_g15), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n9823) );
  OAI221_X1 U11002 ( .B1(SI_17_), .B2(keyinput_g15), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_g69), .A(n9823), .ZN(n9824) );
  NOR4_X1 U11003 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9828)
         );
  NAND4_X1 U11004 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n9934)
         );
  AOI22_X1 U11005 ( .A1(n9950), .A2(keyinput_g56), .B1(keyinput_g40), .B2(
        n9833), .ZN(n9832) );
  OAI221_X1 U11006 ( .B1(n9950), .B2(keyinput_g56), .C1(n9833), .C2(
        keyinput_g40), .A(n9832), .ZN(n9843) );
  AOI22_X1 U11007 ( .A1(n9835), .A2(keyinput_g76), .B1(keyinput_g17), .B2(
        n5212), .ZN(n9834) );
  OAI221_X1 U11008 ( .B1(n9835), .B2(keyinput_g76), .C1(n5212), .C2(
        keyinput_g17), .A(n9834), .ZN(n9842) );
  AOI22_X1 U11009 ( .A1(n9940), .A2(keyinput_g25), .B1(n9837), .B2(
        keyinput_g78), .ZN(n9836) );
  OAI221_X1 U11010 ( .B1(n9940), .B2(keyinput_g25), .C1(n9837), .C2(
        keyinput_g78), .A(n9836), .ZN(n9841) );
  XNOR2_X1 U11011 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g118), .ZN(n9839)
         );
  XNOR2_X1 U11012 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n9838) );
  NAND2_X1 U11013 ( .A1(n9839), .A2(n9838), .ZN(n9840) );
  NOR4_X1 U11014 ( .A1(n9843), .A2(n9842), .A3(n9841), .A4(n9840), .ZN(n9881)
         );
  AOI22_X1 U11015 ( .A1(n9846), .A2(keyinput_g36), .B1(keyinput_g6), .B2(n9845), .ZN(n9844) );
  OAI221_X1 U11016 ( .B1(n9846), .B2(keyinput_g36), .C1(n9845), .C2(
        keyinput_g6), .A(n9844), .ZN(n9854) );
  XOR2_X1 U11017 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_g58), .Z(n9853) );
  XOR2_X1 U11018 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .Z(n9852) );
  XNOR2_X1 U11019 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_g83), .ZN(n9850)
         );
  XNOR2_X1 U11020 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9849) );
  XNOR2_X1 U11021 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g114), .ZN(n9848)
         );
  XNOR2_X1 U11022 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_g77), .ZN(n9847)
         );
  NAND4_X1 U11023 ( .A1(n9850), .A2(n9849), .A3(n9848), .A4(n9847), .ZN(n9851)
         );
  NOR4_X1 U11024 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n9851), .ZN(n9880)
         );
  INV_X1 U11025 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9954) );
  INV_X1 U11026 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U11027 ( .A1(n9954), .A2(keyinput_g55), .B1(keyinput_g122), .B2(
        n9856), .ZN(n9855) );
  OAI221_X1 U11028 ( .B1(n9954), .B2(keyinput_g55), .C1(n9856), .C2(
        keyinput_g122), .A(n9855), .ZN(n9861) );
  XNOR2_X1 U11029 ( .A(n9857), .B(keyinput_g19), .ZN(n9860) );
  XNOR2_X1 U11030 ( .A(n9858), .B(keyinput_g94), .ZN(n9859) );
  NOR3_X1 U11031 ( .A1(n9861), .A2(n9860), .A3(n9859), .ZN(n9865) );
  XNOR2_X1 U11032 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g120), .ZN(n9864)
         );
  XNOR2_X1 U11033 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g91), .ZN(n9863) );
  XNOR2_X1 U11034 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g100), .ZN(n9862)
         );
  NAND4_X1 U11035 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n9867)
         );
  INV_X1 U11036 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10200) );
  XNOR2_X1 U11037 ( .A(n10200), .B(keyinput_g0), .ZN(n9866) );
  NOR2_X1 U11038 ( .A1(n9867), .A2(n9866), .ZN(n9879) );
  XNOR2_X1 U11039 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g111), .ZN(n9871)
         );
  XNOR2_X1 U11040 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_g43), .ZN(n9870)
         );
  XNOR2_X1 U11041 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g109), .ZN(n9869)
         );
  XNOR2_X1 U11042 ( .A(SI_27_), .B(keyinput_g5), .ZN(n9868) );
  NAND4_X1 U11043 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n9877)
         );
  XNOR2_X1 U11044 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g121), .ZN(n9875)
         );
  XNOR2_X1 U11045 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n9874)
         );
  XNOR2_X1 U11046 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g92), .ZN(n9873) );
  XNOR2_X1 U11047 ( .A(SI_8_), .B(keyinput_g24), .ZN(n9872) );
  NAND4_X1 U11048 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n9876)
         );
  NOR2_X1 U11049 ( .A1(n9877), .A2(n9876), .ZN(n9878) );
  NAND4_X1 U11050 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n9933)
         );
  INV_X1 U11051 ( .A(SI_31_), .ZN(n9884) );
  AOI22_X1 U11052 ( .A1(n9884), .A2(keyinput_g1), .B1(n9883), .B2(
        keyinput_g123), .ZN(n9882) );
  OAI221_X1 U11053 ( .B1(n9884), .B2(keyinput_g1), .C1(n9883), .C2(
        keyinput_g123), .A(n9882), .ZN(n9893) );
  AOI22_X1 U11054 ( .A1(n5384), .A2(keyinput_g49), .B1(keyinput_g23), .B2(
        n9886), .ZN(n9885) );
  OAI221_X1 U11055 ( .B1(n5384), .B2(keyinput_g49), .C1(n9886), .C2(
        keyinput_g23), .A(n9885), .ZN(n9892) );
  XOR2_X1 U11056 ( .A(n5228), .B(keyinput_g13), .Z(n9890) );
  XNOR2_X1 U11057 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g103), .ZN(n9889)
         );
  XNOR2_X1 U11058 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g116), .ZN(n9888)
         );
  XNOR2_X1 U11059 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n9887)
         );
  NAND4_X1 U11060 ( .A1(n9890), .A2(n9889), .A3(n9888), .A4(n9887), .ZN(n9891)
         );
  NOR3_X1 U11061 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(n9931) );
  AOI22_X1 U11062 ( .A1(n9974), .A2(keyinput_g50), .B1(keyinput_g27), .B2(
        n9975), .ZN(n9894) );
  OAI221_X1 U11063 ( .B1(n9974), .B2(keyinput_g50), .C1(n9975), .C2(
        keyinput_g27), .A(n9894), .ZN(n9903) );
  XNOR2_X1 U11064 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g108), .ZN(n9898)
         );
  XNOR2_X1 U11065 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n9897) );
  XNOR2_X1 U11066 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g110), .ZN(n9896)
         );
  XNOR2_X1 U11067 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .ZN(n9895)
         );
  NAND4_X1 U11068 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n9902)
         );
  XNOR2_X1 U11069 ( .A(n9899), .B(keyinput_g112), .ZN(n9901) );
  INV_X1 U11070 ( .A(SI_24_), .ZN(n9937) );
  XNOR2_X1 U11071 ( .A(keyinput_g8), .B(n9937), .ZN(n9900) );
  NOR4_X1 U11072 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9930)
         );
  AOI22_X1 U11073 ( .A1(n9941), .A2(keyinput_g52), .B1(keyinput_g124), .B2(
        n10287), .ZN(n9904) );
  OAI221_X1 U11074 ( .B1(n9941), .B2(keyinput_g52), .C1(n10287), .C2(
        keyinput_g124), .A(n9904), .ZN(n9913) );
  AOI22_X1 U11075 ( .A1(n10070), .A2(keyinput_g4), .B1(keyinput_g10), .B2(
        n9906), .ZN(n9905) );
  OAI221_X1 U11076 ( .B1(n10070), .B2(keyinput_g4), .C1(n9906), .C2(
        keyinput_g10), .A(n9905), .ZN(n9912) );
  XNOR2_X1 U11077 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g105), .ZN(n9910)
         );
  XNOR2_X1 U11078 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_g113), .ZN(n9909)
         );
  XNOR2_X1 U11079 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g106), .ZN(n9908)
         );
  XNOR2_X1 U11080 ( .A(keyinput_g54), .B(P2_REG3_REG_0__SCAN_IN), .ZN(n9907)
         );
  NAND4_X1 U11081 ( .A1(n9910), .A2(n9909), .A3(n9908), .A4(n9907), .ZN(n9911)
         );
  NOR3_X1 U11082 ( .A1(n9913), .A2(n9912), .A3(n9911), .ZN(n9929) );
  INV_X1 U11083 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9916) );
  INV_X1 U11084 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U11085 ( .A1(n9916), .A2(keyinput_g60), .B1(n9915), .B2(
        keyinput_g42), .ZN(n9914) );
  OAI221_X1 U11086 ( .B1(n9916), .B2(keyinput_g60), .C1(n9915), .C2(
        keyinput_g42), .A(n9914), .ZN(n9927) );
  AOI22_X1 U11087 ( .A1(n9918), .A2(keyinput_g12), .B1(n5673), .B2(
        keyinput_g47), .ZN(n9917) );
  OAI221_X1 U11088 ( .B1(n9918), .B2(keyinput_g12), .C1(n5673), .C2(
        keyinput_g47), .A(n9917), .ZN(n9926) );
  AOI22_X1 U11089 ( .A1(n9921), .A2(keyinput_g89), .B1(n9920), .B2(
        keyinput_g51), .ZN(n9919) );
  OAI221_X1 U11090 ( .B1(n9921), .B2(keyinput_g89), .C1(n9920), .C2(
        keyinput_g51), .A(n9919), .ZN(n9925) );
  XNOR2_X1 U11091 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_g73), .ZN(n9923)
         );
  XNOR2_X1 U11092 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9922) );
  NAND2_X1 U11093 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  NOR4_X1 U11094 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9928)
         );
  NAND4_X1 U11095 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n9932)
         );
  NOR4_X1 U11096 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(n10129)
         );
  AOI22_X1 U11097 ( .A1(n9938), .A2(keyinput_f86), .B1(n9937), .B2(keyinput_f8), .ZN(n9936) );
  OAI221_X1 U11098 ( .B1(n9938), .B2(keyinput_f86), .C1(n9937), .C2(
        keyinput_f8), .A(n9936), .ZN(n9948) );
  AOI22_X1 U11099 ( .A1(n9941), .A2(keyinput_f52), .B1(keyinput_f25), .B2(
        n9940), .ZN(n9939) );
  OAI221_X1 U11100 ( .B1(n9941), .B2(keyinput_f52), .C1(n9940), .C2(
        keyinput_f25), .A(n9939), .ZN(n9947) );
  XNOR2_X1 U11101 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_f76), .ZN(n9945)
         );
  XNOR2_X1 U11102 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f104), .ZN(n9944)
         );
  XNOR2_X1 U11103 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f119), .ZN(n9943)
         );
  XNOR2_X1 U11104 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_f40), .ZN(n9942)
         );
  NAND4_X1 U11105 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9946)
         );
  NOR3_X1 U11106 ( .A1(n9948), .A2(n9947), .A3(n9946), .ZN(n10122) );
  AOI22_X1 U11107 ( .A1(n9951), .A2(keyinput_f66), .B1(n9950), .B2(
        keyinput_f56), .ZN(n9949) );
  OAI221_X1 U11108 ( .B1(n9951), .B2(keyinput_f66), .C1(n9950), .C2(
        keyinput_f56), .A(n9949), .ZN(n9952) );
  INV_X1 U11109 ( .A(n9952), .ZN(n9964) );
  AOI22_X1 U11110 ( .A1(n9955), .A2(keyinput_f81), .B1(n9954), .B2(
        keyinput_f55), .ZN(n9953) );
  OAI221_X1 U11111 ( .B1(n9955), .B2(keyinput_f81), .C1(n9954), .C2(
        keyinput_f55), .A(n9953), .ZN(n9956) );
  INV_X1 U11112 ( .A(n9956), .ZN(n9963) );
  XNOR2_X1 U11113 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f118), .ZN(n9959)
         );
  XNOR2_X1 U11114 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f93), .ZN(n9958) );
  XNOR2_X1 U11115 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_f36), .ZN(n9957)
         );
  AND3_X1 U11116 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n9962) );
  INV_X1 U11117 ( .A(keyinput_f124), .ZN(n9960) );
  XNOR2_X1 U11118 ( .A(n10287), .B(n9960), .ZN(n9961) );
  AND4_X1 U11119 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), .ZN(n10121)
         );
  OAI22_X1 U11120 ( .A1(n9966), .A2(keyinput_f99), .B1(n10285), .B2(
        keyinput_f126), .ZN(n9965) );
  AOI221_X1 U11121 ( .B1(n9966), .B2(keyinput_f99), .C1(keyinput_f126), .C2(
        n10285), .A(n9965), .ZN(n9990) );
  INV_X1 U11122 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10423) );
  INV_X1 U11123 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9968) );
  AOI22_X1 U11124 ( .A1(n10423), .A2(keyinput_f54), .B1(n9968), .B2(
        keyinput_f37), .ZN(n9967) );
  OAI221_X1 U11125 ( .B1(n10423), .B2(keyinput_f54), .C1(n9968), .C2(
        keyinput_f37), .A(n9967), .ZN(n9972) );
  AOI22_X1 U11126 ( .A1(n8152), .A2(keyinput_f65), .B1(n9970), .B2(
        keyinput_f79), .ZN(n9969) );
  OAI221_X1 U11127 ( .B1(n8152), .B2(keyinput_f65), .C1(n9970), .C2(
        keyinput_f79), .A(n9969), .ZN(n9971) );
  NOR2_X1 U11128 ( .A1(n9972), .A2(n9971), .ZN(n9989) );
  AOI22_X1 U11129 ( .A1(n9975), .A2(keyinput_f27), .B1(n9974), .B2(
        keyinput_f50), .ZN(n9973) );
  OAI221_X1 U11130 ( .B1(n9975), .B2(keyinput_f27), .C1(n9974), .C2(
        keyinput_f50), .A(n9973), .ZN(n9977) );
  XNOR2_X1 U11131 ( .A(keyinput_f0), .B(n10200), .ZN(n9976) );
  NOR2_X1 U11132 ( .A1(n9977), .A2(n9976), .ZN(n9988) );
  XNOR2_X1 U11133 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_f84), .ZN(n9981)
         );
  XNOR2_X1 U11134 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_f114), .ZN(n9980)
         );
  XNOR2_X1 U11135 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f110), .ZN(n9979)
         );
  XNOR2_X1 U11136 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_f89), .ZN(n9978)
         );
  NAND4_X1 U11137 ( .A1(n9981), .A2(n9980), .A3(n9979), .A4(n9978), .ZN(n9986)
         );
  XNOR2_X1 U11138 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_f117), .ZN(n9984)
         );
  XNOR2_X1 U11139 ( .A(SI_22_), .B(keyinput_f10), .ZN(n9983) );
  XNOR2_X1 U11140 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f100), .ZN(n9982)
         );
  NAND3_X1 U11141 ( .A1(n9984), .A2(n9983), .A3(n9982), .ZN(n9985) );
  NOR2_X1 U11142 ( .A1(n9986), .A2(n9985), .ZN(n9987) );
  AND4_X1 U11143 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n10120)
         );
  OAI22_X1 U11144 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P1_IR_REG_15__SCAN_IN), 
        .B2(keyinput_f105), .ZN(n9991) );
  AOI221_X1 U11145 ( .B1(SI_23_), .B2(keyinput_f9), .C1(keyinput_f105), .C2(
        P1_IR_REG_15__SCAN_IN), .A(n9991), .ZN(n9998) );
  OAI22_X1 U11146 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_f70), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n9992) );
  AOI221_X1 U11147 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .C1(
        keyinput_f13), .C2(SI_19_), .A(n9992), .ZN(n9997) );
  OAI22_X1 U11148 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .ZN(n9993) );
  AOI221_X1 U11149 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        keyinput_f103), .C2(P1_IR_REG_13__SCAN_IN), .A(n9993), .ZN(n9996) );
  OAI22_X1 U11150 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        keyinput_f71), .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9994) );
  AOI221_X1 U11151 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_f71), .A(n9994), .ZN(n9995) );
  NAND4_X1 U11152 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10118) );
  OAI22_X1 U11153 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f122), .B2(P1_D_REG_0__SCAN_IN), .ZN(n9999) );
  AOI221_X1 U11154 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_f122), .A(n9999), .ZN(n10024) );
  OAI22_X1 U11155 ( .A1(SI_13_), .A2(keyinput_f19), .B1(P1_IR_REG_5__SCAN_IN), 
        .B2(keyinput_f95), .ZN(n10000) );
  AOI221_X1 U11156 ( .B1(SI_13_), .B2(keyinput_f19), .C1(keyinput_f95), .C2(
        P1_IR_REG_5__SCAN_IN), .A(n10000), .ZN(n10003) );
  OAI22_X1 U11157 ( .A1(SI_25_), .A2(keyinput_f7), .B1(keyinput_f108), .B2(
        P1_IR_REG_18__SCAN_IN), .ZN(n10001) );
  AOI221_X1 U11158 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P1_IR_REG_18__SCAN_IN), 
        .C2(keyinput_f108), .A(n10001), .ZN(n10002) );
  OAI211_X1 U11159 ( .C1(n5444), .C2(keyinput_f53), .A(n10003), .B(n10002), 
        .ZN(n10004) );
  AOI21_X1 U11160 ( .B1(n5444), .B2(keyinput_f53), .A(n10004), .ZN(n10023) );
  AOI22_X1 U11161 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f91), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .ZN(n10005) );
  OAI221_X1 U11162 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f91), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n10005), .ZN(n10012)
         );
  AOI22_X1 U11163 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_f75), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10006) );
  OAI221_X1 U11164 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n10006), .ZN(n10011)
         );
  AOI22_X1 U11165 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n10007) );
  OAI221_X1 U11166 ( .B1(SI_29_), .B2(keyinput_f3), .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10007), .ZN(n10010) );
  AOI22_X1 U11167 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .ZN(n10008) );
  OAI221_X1 U11168 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_f68), .A(n10008), .ZN(n10009)
         );
  NOR4_X1 U11169 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10022) );
  AOI22_X1 U11170 ( .A1(SI_16_), .A2(keyinput_f16), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n10013) );
  OAI221_X1 U11171 ( .B1(SI_16_), .B2(keyinput_f16), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10013), .ZN(n10020)
         );
  AOI22_X1 U11172 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10014) );
  OAI221_X1 U11173 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n10014), .ZN(n10019) );
  AOI22_X1 U11174 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n10015) );
  OAI221_X1 U11175 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n10015), .ZN(n10018)
         );
  AOI22_X1 U11176 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f102), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n10016) );
  OAI221_X1 U11177 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n10016), .ZN(n10017)
         );
  NOR4_X1 U11178 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10021) );
  NAND4_X1 U11179 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10117) );
  AOI22_X1 U11180 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_f115), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_f112), .ZN(n10025) );
  OAI221_X1 U11181 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_f115), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_f112), .A(n10025), .ZN(n10032) );
  AOI22_X1 U11182 ( .A1(SI_0_), .A2(keyinput_f32), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n10026) );
  OAI221_X1 U11183 ( .B1(SI_0_), .B2(keyinput_f32), .C1(SI_20_), .C2(
        keyinput_f12), .A(n10026), .ZN(n10031) );
  AOI22_X1 U11184 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P1_IR_REG_7__SCAN_IN), 
        .B2(keyinput_f97), .ZN(n10027) );
  OAI221_X1 U11185 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P1_IR_REG_7__SCAN_IN), 
        .C2(keyinput_f97), .A(n10027), .ZN(n10030) );
  AOI22_X1 U11186 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_f121), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n10028) );
  OAI221_X1 U11187 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_f121), .C1(SI_2_), .C2(keyinput_f30), .A(n10028), .ZN(n10029) );
  NOR4_X1 U11188 ( .A1(n10032), .A2(n10031), .A3(n10030), .A4(n10029), .ZN(
        n10060) );
  AOI22_X1 U11189 ( .A1(SI_1_), .A2(keyinput_f31), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .ZN(n10033) );
  OAI221_X1 U11190 ( .B1(SI_1_), .B2(keyinput_f31), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_f82), .A(n10033), .ZN(n10040)
         );
  AOI22_X1 U11191 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f98), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .ZN(n10034) );
  OAI221_X1 U11192 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f98), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n10034), .ZN(n10039) );
  AOI22_X1 U11193 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f109), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n10035) );
  OAI221_X1 U11194 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n10035), .ZN(n10038) );
  AOI22_X1 U11195 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10036) );
  OAI221_X1 U11196 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10036), .ZN(n10037)
         );
  NOR4_X1 U11197 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10059) );
  AOI22_X1 U11198 ( .A1(SI_6_), .A2(keyinput_f26), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10041) );
  OAI221_X1 U11199 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10041), .ZN(n10048)
         );
  AOI22_X1 U11200 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f111), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .ZN(n10042) );
  OAI221_X1 U11201 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_f88), .A(n10042), .ZN(n10047)
         );
  AOI22_X1 U11202 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n10043) );
  OAI221_X1 U11203 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10043), .ZN(n10046) );
  AOI22_X1 U11204 ( .A1(SI_3_), .A2(keyinput_f29), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n10044) );
  OAI221_X1 U11205 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10044), .ZN(n10045)
         );
  NOR4_X1 U11206 ( .A1(n10048), .A2(n10047), .A3(n10046), .A4(n10045), .ZN(
        n10058) );
  AOI22_X1 U11207 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n10049) );
  OAI221_X1 U11208 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10049), .ZN(n10056)
         );
  AOI22_X1 U11209 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_f127), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .ZN(n10050) );
  OAI221_X1 U11210 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_f127), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n10050), .ZN(n10055)
         );
  AOI22_X1 U11211 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n10051) );
  OAI221_X1 U11212 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10051), .ZN(n10054)
         );
  AOI22_X1 U11213 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n10052) );
  OAI221_X1 U11214 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10052), .ZN(n10053) );
  NOR4_X1 U11215 ( .A1(n10056), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(
        n10057) );
  NAND4_X1 U11216 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10116) );
  AOI22_X1 U11217 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n10061) );
  OAI221_X1 U11218 ( .B1(SI_27_), .B2(keyinput_f5), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n10061), .ZN(n10068)
         );
  AOI22_X1 U11219 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f101), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n10062) );
  OAI221_X1 U11220 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n10062), .ZN(n10067)
         );
  AOI22_X1 U11221 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10063) );
  OAI221_X1 U11222 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n10063), .ZN(n10066)
         );
  AOI22_X1 U11223 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f116), .B1(SI_17_), .B2(keyinput_f15), .ZN(n10064) );
  OAI221_X1 U11224 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f116), .C1(
        SI_17_), .C2(keyinput_f15), .A(n10064), .ZN(n10065) );
  NOR4_X1 U11225 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        n10114) );
  AOI22_X1 U11226 ( .A1(n5212), .A2(keyinput_f17), .B1(n10070), .B2(
        keyinput_f4), .ZN(n10069) );
  OAI221_X1 U11227 ( .B1(n5212), .B2(keyinput_f17), .C1(n10070), .C2(
        keyinput_f4), .A(n10069), .ZN(n10081) );
  AOI22_X1 U11228 ( .A1(n10073), .A2(keyinput_f24), .B1(n10072), .B2(
        keyinput_f74), .ZN(n10071) );
  OAI221_X1 U11229 ( .B1(n10073), .B2(keyinput_f24), .C1(n10072), .C2(
        keyinput_f74), .A(n10071), .ZN(n10080) );
  AOI22_X1 U11230 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f96), .B1(SI_26_), 
        .B2(keyinput_f6), .ZN(n10074) );
  OAI221_X1 U11231 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f96), .C1(SI_26_), 
        .C2(keyinput_f6), .A(n10074), .ZN(n10079) );
  INV_X1 U11232 ( .A(SI_21_), .ZN(n10075) );
  XOR2_X1 U11233 ( .A(n10075), .B(keyinput_f11), .Z(n10077) );
  XNOR2_X1 U11234 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f90), .ZN(n10076) );
  NAND2_X1 U11235 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  NOR4_X1 U11236 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        n10113) );
  AOI22_X1 U11237 ( .A1(n10083), .A2(keyinput_f113), .B1(keyinput_f125), .B2(
        n10286), .ZN(n10082) );
  OAI221_X1 U11238 ( .B1(n10083), .B2(keyinput_f113), .C1(n10286), .C2(
        keyinput_f125), .A(n10082), .ZN(n10095) );
  AOI22_X1 U11239 ( .A1(n10086), .A2(keyinput_f18), .B1(keyinput_f22), .B2(
        n10085), .ZN(n10084) );
  OAI221_X1 U11240 ( .B1(n10086), .B2(keyinput_f18), .C1(n10085), .C2(
        keyinput_f22), .A(n10084), .ZN(n10094) );
  AOI22_X1 U11241 ( .A1(n10089), .A2(keyinput_f83), .B1(keyinput_f2), .B2(
        n10088), .ZN(n10087) );
  OAI221_X1 U11242 ( .B1(n10089), .B2(keyinput_f83), .C1(n10088), .C2(
        keyinput_f2), .A(n10087), .ZN(n10093) );
  XNOR2_X1 U11243 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f92), .ZN(n10091) );
  XNOR2_X1 U11244 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_f57), .ZN(n10090)
         );
  NAND2_X1 U11245 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  NOR4_X1 U11246 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n10112) );
  AOI22_X1 U11247 ( .A1(n10098), .A2(keyinput_f63), .B1(keyinput_f107), .B2(
        n10097), .ZN(n10096) );
  OAI221_X1 U11248 ( .B1(n10098), .B2(keyinput_f63), .C1(n10097), .C2(
        keyinput_f107), .A(n10096), .ZN(n10110) );
  AOI22_X1 U11249 ( .A1(n10101), .A2(keyinput_f69), .B1(keyinput_f14), .B2(
        n10100), .ZN(n10099) );
  OAI221_X1 U11250 ( .B1(n10101), .B2(keyinput_f69), .C1(n10100), .C2(
        keyinput_f14), .A(n10099), .ZN(n10109) );
  AOI22_X1 U11251 ( .A1(n10104), .A2(keyinput_f21), .B1(n10103), .B2(
        keyinput_f39), .ZN(n10102) );
  OAI221_X1 U11252 ( .B1(n10104), .B2(keyinput_f21), .C1(n10103), .C2(
        keyinput_f39), .A(n10102), .ZN(n10108) );
  XNOR2_X1 U11253 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f106), .ZN(n10106)
         );
  XNOR2_X1 U11254 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f94), .ZN(n10105) );
  NAND2_X1 U11255 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  NOR4_X1 U11256 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10111) );
  NAND4_X1 U11257 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10115) );
  NOR4_X1 U11258 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10119) );
  NAND4_X1 U11259 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10124) );
  AOI21_X1 U11260 ( .B1(keyinput_f28), .B2(n10124), .A(keyinput_g28), .ZN(
        n10126) );
  INV_X1 U11261 ( .A(keyinput_f28), .ZN(n10123) );
  AOI21_X1 U11262 ( .B1(n10124), .B2(n10123), .A(n10127), .ZN(n10125) );
  AOI22_X1 U11263 ( .A1(n10127), .A2(n10126), .B1(keyinput_g28), .B2(n10125), 
        .ZN(n10128) );
  AOI21_X1 U11264 ( .B1(n10130), .B2(n10129), .A(n10128), .ZN(n10189) );
  INV_X1 U11265 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10187) );
  NOR2_X1 U11266 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10185) );
  NOR2_X1 U11267 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10181) );
  NOR2_X1 U11268 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10177) );
  NOR2_X1 U11269 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10174) );
  NOR2_X1 U11270 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10170) );
  NOR2_X1 U11271 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10166) );
  NOR2_X1 U11272 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10162) );
  NOR2_X1 U11273 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10158) );
  NOR2_X1 U11274 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10154) );
  NOR2_X1 U11275 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10150) );
  NOR2_X1 U11276 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10146) );
  NOR2_X1 U11277 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10143) );
  NOR2_X1 U11278 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10141) );
  NOR2_X1 U11279 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10139) );
  NAND2_X1 U11280 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10137) );
  XOR2_X1 U11281 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10606) );
  NAND2_X1 U11282 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10135) );
  AOI21_X1 U11283 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10572) );
  INV_X1 U11284 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U11285 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10131) );
  NOR2_X1 U11286 ( .A1(n10132), .A2(n10131), .ZN(n10571) );
  NOR2_X1 U11287 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10571), .ZN(n10133) );
  NOR2_X1 U11288 ( .A1(n10572), .A2(n10133), .ZN(n10596) );
  XOR2_X1 U11289 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10595) );
  NAND2_X1 U11290 ( .A1(n10596), .A2(n10595), .ZN(n10134) );
  NAND2_X1 U11291 ( .A1(n10135), .A2(n10134), .ZN(n10605) );
  NAND2_X1 U11292 ( .A1(n10606), .A2(n10605), .ZN(n10136) );
  NAND2_X1 U11293 ( .A1(n10137), .A2(n10136), .ZN(n10608) );
  XNOR2_X1 U11294 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10607) );
  NOR2_X1 U11295 ( .A1(n10608), .A2(n10607), .ZN(n10138) );
  NOR2_X1 U11296 ( .A1(n10139), .A2(n10138), .ZN(n10598) );
  XNOR2_X1 U11297 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10597) );
  NOR2_X1 U11298 ( .A1(n10598), .A2(n10597), .ZN(n10140) );
  NOR2_X1 U11299 ( .A1(n10141), .A2(n10140), .ZN(n10604) );
  XNOR2_X1 U11300 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10603) );
  NOR2_X1 U11301 ( .A1(n10604), .A2(n10603), .ZN(n10142) );
  NOR2_X1 U11302 ( .A1(n10143), .A2(n10142), .ZN(n10600) );
  XOR2_X1 U11303 ( .A(n10144), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n10599) );
  NOR2_X1 U11304 ( .A1(n10600), .A2(n10599), .ZN(n10145) );
  NOR2_X1 U11305 ( .A1(n10146), .A2(n10145), .ZN(n10602) );
  INV_X1 U11306 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U11307 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10148), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10147), .ZN(n10601) );
  NOR2_X1 U11308 ( .A1(n10602), .A2(n10601), .ZN(n10149) );
  NOR2_X1 U11309 ( .A1(n10150), .A2(n10149), .ZN(n10594) );
  AOI22_X1 U11310 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10152), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10151), .ZN(n10593) );
  NOR2_X1 U11311 ( .A1(n10594), .A2(n10593), .ZN(n10153) );
  NOR2_X1 U11312 ( .A1(n10154), .A2(n10153), .ZN(n10592) );
  INV_X1 U11313 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U11314 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10156), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10155), .ZN(n10591) );
  NOR2_X1 U11315 ( .A1(n10592), .A2(n10591), .ZN(n10157) );
  NOR2_X1 U11316 ( .A1(n10158), .A2(n10157), .ZN(n10590) );
  INV_X1 U11317 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U11318 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10160), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10159), .ZN(n10589) );
  NOR2_X1 U11319 ( .A1(n10590), .A2(n10589), .ZN(n10161) );
  NOR2_X1 U11320 ( .A1(n10162), .A2(n10161), .ZN(n10588) );
  INV_X1 U11321 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10164) );
  INV_X1 U11322 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11323 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10164), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10163), .ZN(n10587) );
  NOR2_X1 U11324 ( .A1(n10588), .A2(n10587), .ZN(n10165) );
  NOR2_X1 U11325 ( .A1(n10166), .A2(n10165), .ZN(n10586) );
  INV_X1 U11326 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U11327 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10168), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10167), .ZN(n10585) );
  NOR2_X1 U11328 ( .A1(n10586), .A2(n10585), .ZN(n10169) );
  NOR2_X1 U11329 ( .A1(n10170), .A2(n10169), .ZN(n10584) );
  INV_X1 U11330 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11331 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10172), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10171), .ZN(n10583) );
  NOR2_X1 U11332 ( .A1(n10584), .A2(n10583), .ZN(n10173) );
  NOR2_X1 U11333 ( .A1(n10174), .A2(n10173), .ZN(n10582) );
  AOI22_X1 U11334 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9369), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10175), .ZN(n10581) );
  NOR2_X1 U11335 ( .A1(n10582), .A2(n10581), .ZN(n10176) );
  NOR2_X1 U11336 ( .A1(n10177), .A2(n10176), .ZN(n10580) );
  INV_X1 U11337 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U11338 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10179), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10178), .ZN(n10579) );
  NOR2_X1 U11339 ( .A1(n10580), .A2(n10579), .ZN(n10180) );
  NOR2_X1 U11340 ( .A1(n10181), .A2(n10180), .ZN(n10578) );
  INV_X1 U11341 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U11342 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10183), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10182), .ZN(n10577) );
  NOR2_X1 U11343 ( .A1(n10578), .A2(n10577), .ZN(n10184) );
  NOR2_X1 U11344 ( .A1(n10185), .A2(n10184), .ZN(n10575) );
  NAND2_X1 U11345 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10575), .ZN(n10186) );
  NOR2_X1 U11346 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10575), .ZN(n10574) );
  AOI21_X1 U11347 ( .B1(n10187), .B2(n10186), .A(n10574), .ZN(n10188) );
  XOR2_X1 U11348 ( .A(n10189), .B(n10188), .Z(n10193) );
  NOR2_X1 U11349 ( .A1(n10191), .A2(n10190), .ZN(n10192) );
  XOR2_X1 U11350 ( .A(n10193), .B(n10192), .Z(ADD_1068_U4) );
  OAI211_X1 U11351 ( .C1(n10196), .C2(n10388), .A(n10195), .B(n10194), .ZN(
        n10197) );
  AOI21_X1 U11352 ( .B1(n10198), .B2(n10385), .A(n10197), .ZN(n10199) );
  AOI22_X1 U11353 ( .A1(n10413), .A2(n10199), .B1(n9390), .B2(n10411), .ZN(
        P1_U3538) );
  AOI22_X1 U11354 ( .A1(n10395), .A2(n10199), .B1(n6186), .B2(n6662), .ZN(
        P1_U3501) );
  XOR2_X1 U11355 ( .A(n10200), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11356 ( .A(n10201), .B(n10202), .ZN(n10393) );
  NAND2_X1 U11357 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  AOI21_X1 U11358 ( .B1(n10205), .B2(n10204), .A(n10345), .ZN(n10207) );
  AOI211_X1 U11359 ( .C1(n10393), .C2(n10370), .A(n10207), .B(n10206), .ZN(
        n10390) );
  INV_X1 U11360 ( .A(n10208), .ZN(n10209) );
  AOI222_X1 U11361 ( .A1(n10210), .A2(n10275), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n10282), .C1(n10271), .C2(n10209), .ZN(n10217) );
  INV_X1 U11362 ( .A(n10211), .ZN(n10279) );
  INV_X1 U11363 ( .A(n10212), .ZN(n10214) );
  OAI211_X1 U11364 ( .C1(n10214), .C2(n10389), .A(n10273), .B(n10213), .ZN(
        n10387) );
  INV_X1 U11365 ( .A(n10387), .ZN(n10215) );
  AOI22_X1 U11366 ( .A1(n10393), .A2(n10279), .B1(n10278), .B2(n10215), .ZN(
        n10216) );
  OAI211_X1 U11367 ( .C1(n10282), .C2(n10390), .A(n10217), .B(n10216), .ZN(
        P1_U3279) );
  XOR2_X1 U11368 ( .A(n10225), .B(n10218), .Z(n10220) );
  AOI21_X1 U11369 ( .B1(n10220), .B2(n10250), .A(n10219), .ZN(n10337) );
  INV_X1 U11370 ( .A(n10221), .ZN(n10222) );
  AOI222_X1 U11371 ( .A1(n10223), .A2(n10275), .B1(n10222), .B2(n10271), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n10282), .ZN(n10231) );
  XNOR2_X1 U11372 ( .A(n10224), .B(n10225), .ZN(n10340) );
  OAI21_X1 U11373 ( .B1(n10226), .B2(n10338), .A(n10273), .ZN(n10227) );
  OR2_X1 U11374 ( .A1(n10228), .A2(n10227), .ZN(n10336) );
  INV_X1 U11375 ( .A(n10336), .ZN(n10229) );
  AOI22_X1 U11376 ( .A1(n10340), .A2(n10242), .B1(n10278), .B2(n10229), .ZN(
        n10230) );
  OAI211_X1 U11377 ( .C1(n10282), .C2(n10337), .A(n10231), .B(n10230), .ZN(
        P1_U3285) );
  XOR2_X1 U11378 ( .A(n10232), .B(n10238), .Z(n10234) );
  AOI21_X1 U11379 ( .B1(n10234), .B2(n10250), .A(n10233), .ZN(n10312) );
  AOI222_X1 U11380 ( .A1(n10236), .A2(n10275), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n10282), .C1(n10271), .C2(n10235), .ZN(n10244) );
  XNOR2_X1 U11381 ( .A(n10237), .B(n10238), .ZN(n10315) );
  OAI211_X1 U11382 ( .C1(n10240), .C2(n10311), .A(n10239), .B(n10273), .ZN(
        n10310) );
  INV_X1 U11383 ( .A(n10310), .ZN(n10241) );
  AOI22_X1 U11384 ( .A1(n10315), .A2(n10242), .B1(n10278), .B2(n10241), .ZN(
        n10243) );
  OAI211_X1 U11385 ( .C1(n10282), .C2(n10312), .A(n10244), .B(n10243), .ZN(
        P1_U3289) );
  XNOR2_X1 U11386 ( .A(n10246), .B(n10245), .ZN(n10300) );
  XNOR2_X1 U11387 ( .A(n10248), .B(n10247), .ZN(n10251) );
  AOI21_X1 U11388 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(n10297) );
  AOI22_X1 U11389 ( .A1(n10253), .A2(n10252), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10271), .ZN(n10254) );
  NAND2_X1 U11390 ( .A1(n10297), .A2(n10254), .ZN(n10255) );
  AOI21_X1 U11391 ( .B1(n10370), .B2(n10300), .A(n10255), .ZN(n10262) );
  OAI211_X1 U11392 ( .C1(n10257), .C2(n10298), .A(n10273), .B(n10256), .ZN(
        n10296) );
  INV_X1 U11393 ( .A(n10296), .ZN(n10258) );
  AOI22_X1 U11394 ( .A1(n10300), .A2(n10279), .B1(n10278), .B2(n10258), .ZN(
        n10259) );
  OAI221_X1 U11395 ( .B1(n10282), .B2(n10262), .C1(n10261), .C2(n10260), .A(
        n10259), .ZN(P1_U3291) );
  XNOR2_X1 U11396 ( .A(n8361), .B(n10263), .ZN(n10294) );
  OAI21_X1 U11397 ( .B1(n10265), .B2(n10358), .A(n10264), .ZN(n10270) );
  NAND2_X1 U11398 ( .A1(n8361), .A2(n10266), .ZN(n10267) );
  AOI21_X1 U11399 ( .B1(n10268), .B2(n10267), .A(n10345), .ZN(n10269) );
  AOI211_X1 U11400 ( .C1(n10370), .C2(n10294), .A(n10270), .B(n10269), .ZN(
        n10291) );
  AOI22_X1 U11401 ( .A1(n10271), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n10282), .ZN(n10281) );
  OAI211_X1 U11402 ( .C1(n10290), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10289) );
  INV_X1 U11403 ( .A(n10289), .ZN(n10277) );
  AOI222_X1 U11404 ( .A1(n10294), .A2(n10279), .B1(n10278), .B2(n10277), .C1(
        n10276), .C2(n10275), .ZN(n10280) );
  OAI211_X1 U11405 ( .C1(n10282), .C2(n10291), .A(n10281), .B(n10280), .ZN(
        P1_U3292) );
  INV_X1 U11406 ( .A(n10288), .ZN(n10283) );
  AND2_X1 U11407 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10283), .ZN(P1_U3294) );
  AND2_X1 U11408 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10283), .ZN(P1_U3295) );
  AND2_X1 U11409 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10283), .ZN(P1_U3296) );
  AND2_X1 U11410 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10283), .ZN(P1_U3297) );
  AND2_X1 U11411 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10283), .ZN(P1_U3298) );
  AND2_X1 U11412 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10283), .ZN(P1_U3299) );
  AND2_X1 U11413 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10283), .ZN(P1_U3300) );
  AND2_X1 U11414 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10283), .ZN(P1_U3301) );
  AND2_X1 U11415 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10283), .ZN(P1_U3302) );
  AND2_X1 U11416 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10283), .ZN(P1_U3303) );
  AND2_X1 U11417 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10283), .ZN(P1_U3304) );
  AND2_X1 U11418 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10283), .ZN(P1_U3305) );
  AND2_X1 U11419 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10283), .ZN(P1_U3306) );
  AND2_X1 U11420 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10283), .ZN(P1_U3307) );
  AND2_X1 U11421 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10283), .ZN(P1_U3308) );
  AND2_X1 U11422 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10283), .ZN(P1_U3309) );
  AND2_X1 U11423 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10283), .ZN(P1_U3310) );
  AND2_X1 U11424 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10283), .ZN(P1_U3311) );
  AND2_X1 U11425 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10283), .ZN(P1_U3312) );
  AND2_X1 U11426 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10283), .ZN(P1_U3313) );
  AND2_X1 U11427 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10283), .ZN(P1_U3314) );
  AND2_X1 U11428 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10283), .ZN(P1_U3315) );
  AND2_X1 U11429 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10283), .ZN(P1_U3316) );
  AND2_X1 U11430 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10283), .ZN(P1_U3317) );
  AND2_X1 U11431 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10283), .ZN(P1_U3318) );
  AND2_X1 U11432 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10283), .ZN(P1_U3319) );
  NOR2_X1 U11433 ( .A1(n10288), .A2(n10284), .ZN(P1_U3320) );
  NOR2_X1 U11434 ( .A1(n10288), .A2(n10285), .ZN(P1_U3321) );
  NOR2_X1 U11435 ( .A1(n10288), .A2(n10286), .ZN(P1_U3322) );
  NOR2_X1 U11436 ( .A1(n10288), .A2(n10287), .ZN(P1_U3323) );
  INV_X1 U11437 ( .A(n10366), .ZN(n10394) );
  OAI21_X1 U11438 ( .B1(n10290), .B2(n10388), .A(n10289), .ZN(n10293) );
  INV_X1 U11439 ( .A(n10291), .ZN(n10292) );
  AOI211_X1 U11440 ( .C1(n10394), .C2(n10294), .A(n10293), .B(n10292), .ZN(
        n10396) );
  INV_X1 U11441 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U11442 ( .A1(n10395), .A2(n10396), .B1(n10295), .B2(n6662), .ZN(
        P1_U3456) );
  OAI211_X1 U11443 ( .C1(n10298), .C2(n10388), .A(n10297), .B(n10296), .ZN(
        n10299) );
  AOI21_X1 U11444 ( .B1(n10300), .B2(n10385), .A(n10299), .ZN(n10398) );
  INV_X1 U11445 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U11446 ( .A1(n10395), .A2(n10398), .B1(n10301), .B2(n6662), .ZN(
        P1_U3459) );
  AOI21_X1 U11447 ( .B1(n10363), .B2(n10303), .A(n10302), .ZN(n10304) );
  OAI211_X1 U11448 ( .C1(n10307), .C2(n10306), .A(n10305), .B(n10304), .ZN(
        n10308) );
  INV_X1 U11449 ( .A(n10308), .ZN(n10400) );
  INV_X1 U11450 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U11451 ( .A1(n10395), .A2(n10400), .B1(n10309), .B2(n6662), .ZN(
        P1_U3462) );
  OAI21_X1 U11452 ( .B1(n10311), .B2(n10388), .A(n10310), .ZN(n10314) );
  INV_X1 U11453 ( .A(n10312), .ZN(n10313) );
  AOI211_X1 U11454 ( .C1(n10385), .C2(n10315), .A(n10314), .B(n10313), .ZN(
        n10401) );
  AOI22_X1 U11455 ( .A1(n10395), .A2(n10401), .B1(n6019), .B2(n6662), .ZN(
        P1_U3465) );
  INV_X1 U11456 ( .A(n10316), .ZN(n10321) );
  OAI21_X1 U11457 ( .B1(n10318), .B2(n10388), .A(n10317), .ZN(n10320) );
  AOI211_X1 U11458 ( .C1(n10385), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10402) );
  AOI22_X1 U11459 ( .A1(n10395), .A2(n10402), .B1(n6036), .B2(n6662), .ZN(
        P1_U3468) );
  AOI22_X1 U11460 ( .A1(n10374), .A2(n10323), .B1(n10322), .B2(n10371), .ZN(
        n10324) );
  OAI211_X1 U11461 ( .C1(n10326), .C2(n10388), .A(n10325), .B(n10324), .ZN(
        n10328) );
  AOI211_X1 U11462 ( .C1(n10385), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10403) );
  AOI22_X1 U11463 ( .A1(n10395), .A2(n10403), .B1(n6078), .B2(n6662), .ZN(
        P1_U3471) );
  AND2_X1 U11464 ( .A1(n10330), .A2(n10385), .ZN(n10334) );
  OAI21_X1 U11465 ( .B1(n10332), .B2(n10388), .A(n10331), .ZN(n10333) );
  NOR3_X1 U11466 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10404) );
  AOI22_X1 U11467 ( .A1(n10395), .A2(n10404), .B1(n6065), .B2(n6662), .ZN(
        P1_U3474) );
  OAI211_X1 U11468 ( .C1(n10338), .C2(n10388), .A(n10337), .B(n10336), .ZN(
        n10339) );
  AOI21_X1 U11469 ( .B1(n10385), .B2(n10340), .A(n10339), .ZN(n10405) );
  AOI22_X1 U11470 ( .A1(n10395), .A2(n10405), .B1(n6055), .B2(n6662), .ZN(
        P1_U3477) );
  AOI22_X1 U11471 ( .A1(n10342), .A2(n10363), .B1(n10374), .B2(n10341), .ZN(
        n10343) );
  OAI211_X1 U11472 ( .C1(n10346), .C2(n10345), .A(n10344), .B(n10343), .ZN(
        n10347) );
  AOI21_X1 U11473 ( .B1(n10385), .B2(n10348), .A(n10347), .ZN(n10406) );
  AOI22_X1 U11474 ( .A1(n10395), .A2(n10406), .B1(n6090), .B2(n6662), .ZN(
        P1_U3480) );
  AOI22_X1 U11475 ( .A1(n10371), .A2(n10373), .B1(n10349), .B2(n10374), .ZN(
        n10350) );
  OAI211_X1 U11476 ( .C1(n10352), .C2(n10388), .A(n10351), .B(n10350), .ZN(
        n10353) );
  AOI211_X1 U11477 ( .C1(n10355), .C2(n10385), .A(n10354), .B(n10353), .ZN(
        n10407) );
  AOI22_X1 U11478 ( .A1(n10395), .A2(n10407), .B1(n6113), .B2(n6662), .ZN(
        P1_U3483) );
  INV_X1 U11479 ( .A(n10367), .ZN(n10369) );
  OAI22_X1 U11480 ( .A1(n10359), .A2(n10358), .B1(n10357), .B2(n10356), .ZN(
        n10361) );
  AOI211_X1 U11481 ( .C1(n10363), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10365) );
  OAI211_X1 U11482 ( .C1(n10367), .C2(n10366), .A(n10365), .B(n10364), .ZN(
        n10368) );
  AOI21_X1 U11483 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(n10408) );
  AOI22_X1 U11484 ( .A1(n10395), .A2(n10408), .B1(n6120), .B2(n6662), .ZN(
        P1_U3486) );
  AOI22_X1 U11485 ( .A1(n10374), .A2(n10373), .B1(n10372), .B2(n10371), .ZN(
        n10375) );
  OAI211_X1 U11486 ( .C1(n10377), .C2(n10388), .A(n10376), .B(n10375), .ZN(
        n10378) );
  AOI211_X1 U11487 ( .C1(n10380), .C2(n10385), .A(n10379), .B(n10378), .ZN(
        n10409) );
  AOI22_X1 U11488 ( .A1(n10395), .A2(n10409), .B1(n6133), .B2(n6662), .ZN(
        P1_U3489) );
  OAI211_X1 U11489 ( .C1(n10383), .C2(n10388), .A(n10382), .B(n10381), .ZN(
        n10384) );
  AOI21_X1 U11490 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(n10410) );
  AOI22_X1 U11491 ( .A1(n10395), .A2(n10410), .B1(n6146), .B2(n6662), .ZN(
        P1_U3492) );
  OAI21_X1 U11492 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(n10392) );
  INV_X1 U11493 ( .A(n10390), .ZN(n10391) );
  AOI211_X1 U11494 ( .C1(n10394), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        n10412) );
  AOI22_X1 U11495 ( .A1(n10395), .A2(n10412), .B1(n6162), .B2(n6662), .ZN(
        P1_U3495) );
  AOI22_X1 U11496 ( .A1(n10413), .A2(n10396), .B1(n7008), .B2(n10411), .ZN(
        P1_U3523) );
  AOI22_X1 U11497 ( .A1(n10413), .A2(n10398), .B1(n10397), .B2(n10411), .ZN(
        P1_U3524) );
  AOI22_X1 U11498 ( .A1(n10413), .A2(n10400), .B1(n10399), .B2(n10411), .ZN(
        P1_U3525) );
  AOI22_X1 U11499 ( .A1(n10413), .A2(n10401), .B1(n6020), .B2(n10411), .ZN(
        P1_U3526) );
  AOI22_X1 U11500 ( .A1(n10413), .A2(n10402), .B1(n7007), .B2(n10411), .ZN(
        P1_U3527) );
  AOI22_X1 U11501 ( .A1(n10413), .A2(n10403), .B1(n7005), .B2(n10411), .ZN(
        P1_U3528) );
  AOI22_X1 U11502 ( .A1(n10413), .A2(n10404), .B1(n7137), .B2(n10411), .ZN(
        P1_U3529) );
  AOI22_X1 U11503 ( .A1(n10413), .A2(n10405), .B1(n7139), .B2(n10411), .ZN(
        P1_U3530) );
  AOI22_X1 U11504 ( .A1(n10413), .A2(n10406), .B1(n6086), .B2(n10411), .ZN(
        P1_U3531) );
  AOI22_X1 U11505 ( .A1(n10413), .A2(n10407), .B1(n7438), .B2(n10411), .ZN(
        P1_U3532) );
  AOI22_X1 U11506 ( .A1(n10413), .A2(n10408), .B1(n7440), .B2(n10411), .ZN(
        P1_U3533) );
  AOI22_X1 U11507 ( .A1(n10413), .A2(n10409), .B1(n8175), .B2(n10411), .ZN(
        P1_U3534) );
  AOI22_X1 U11508 ( .A1(n10413), .A2(n10410), .B1(n8172), .B2(n10411), .ZN(
        P1_U3535) );
  AOI22_X1 U11509 ( .A1(n10413), .A2(n10412), .B1(n8177), .B2(n10411), .ZN(
        P1_U3536) );
  AOI22_X1 U11510 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n10415), .B1(n10414), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10422) );
  OAI21_X1 U11511 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10417), .A(n10416), .ZN(
        n10418) );
  OAI21_X1 U11512 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(n10421) );
  OAI211_X1 U11513 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10423), .A(n10422), .B(
        n10421), .ZN(P2_U3182) );
  XOR2_X1 U11514 ( .A(n10424), .B(n10431), .Z(n10429) );
  AOI222_X1 U11515 ( .A1(n10443), .A2(n10429), .B1(n10428), .B2(n10427), .C1(
        n10426), .C2(n10425), .ZN(n10484) );
  INV_X1 U11516 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10435) );
  XNOR2_X1 U11517 ( .A(n10430), .B(n10431), .ZN(n10487) );
  OAI22_X1 U11518 ( .A1(n10466), .A2(n10485), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10464), .ZN(n10432) );
  AOI21_X1 U11519 ( .B1(n10487), .B2(n10433), .A(n10432), .ZN(n10434) );
  OAI221_X1 U11520 ( .B1(n10472), .B2(n10484), .C1(n10471), .C2(n10435), .A(
        n10434), .ZN(P2_U3230) );
  INV_X1 U11521 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10450) );
  XNOR2_X1 U11522 ( .A(n10436), .B(n10440), .ZN(n10480) );
  INV_X1 U11523 ( .A(n10480), .ZN(n10447) );
  OAI22_X1 U11524 ( .A1(n10479), .A2(n10438), .B1(n10437), .B2(n10464), .ZN(
        n10446) );
  XNOR2_X1 U11525 ( .A(n10440), .B(n10439), .ZN(n10444) );
  OAI22_X1 U11526 ( .A1(n10441), .A2(n10454), .B1(n6810), .B2(n10456), .ZN(
        n10442) );
  AOI21_X1 U11527 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(n10445) );
  OAI21_X1 U11528 ( .B1(n10480), .B2(n10451), .A(n10445), .ZN(n10482) );
  AOI211_X1 U11529 ( .C1(n10448), .C2(n10447), .A(n10446), .B(n10482), .ZN(
        n10449) );
  AOI22_X1 U11530 ( .A1(n10472), .A2(n10450), .B1(n10449), .B2(n10471), .ZN(
        P2_U3231) );
  INV_X1 U11531 ( .A(n10451), .ZN(n10524) );
  OAI21_X1 U11532 ( .B1(n5325), .B2(n10453), .A(n10452), .ZN(n10475) );
  OAI22_X1 U11533 ( .A1(n10457), .A2(n10456), .B1(n10455), .B2(n10454), .ZN(
        n10462) );
  XNOR2_X1 U11534 ( .A(n5325), .B(n10458), .ZN(n10460) );
  NOR2_X1 U11535 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  AOI211_X1 U11536 ( .C1(n10524), .C2(n10475), .A(n10462), .B(n10461), .ZN(
        n10477) );
  NOR2_X1 U11537 ( .A1(n10472), .A2(n10463), .ZN(n10468) );
  OAI22_X1 U11538 ( .A1(n10466), .A2(n6811), .B1(n10465), .B2(n10464), .ZN(
        n10467) );
  AOI21_X1 U11539 ( .B1(n10475), .B2(n10468), .A(n10467), .ZN(n10469) );
  OAI221_X1 U11540 ( .B1(n10472), .B2(n10477), .C1(n10471), .C2(n10470), .A(
        n10469), .ZN(P2_U3232) );
  INV_X1 U11541 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U11542 ( .A1(n10475), .A2(n10474), .B1(n10537), .B2(n10473), .ZN(
        n10476) );
  AND2_X1 U11543 ( .A1(n10477), .A2(n10476), .ZN(n10549) );
  AOI22_X1 U11544 ( .A1(n10547), .A2(n10478), .B1(n10549), .B2(n10545), .ZN(
        P2_U3393) );
  INV_X1 U11545 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10483) );
  OAI22_X1 U11546 ( .A1(n10480), .A2(n10527), .B1(n10479), .B2(n10539), .ZN(
        n10481) );
  NOR2_X1 U11547 ( .A1(n10482), .A2(n10481), .ZN(n10551) );
  AOI22_X1 U11548 ( .A1(n10547), .A2(n10483), .B1(n10551), .B2(n10545), .ZN(
        P2_U3396) );
  INV_X1 U11549 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10488) );
  OAI21_X1 U11550 ( .B1(n10485), .B2(n10539), .A(n10484), .ZN(n10486) );
  AOI21_X1 U11551 ( .B1(n10544), .B2(n10487), .A(n10486), .ZN(n10553) );
  AOI22_X1 U11552 ( .A1(n10547), .A2(n10488), .B1(n10553), .B2(n10545), .ZN(
        P2_U3399) );
  INV_X1 U11553 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10493) );
  NOR2_X1 U11554 ( .A1(n10489), .A2(n10539), .ZN(n10491) );
  AOI211_X1 U11555 ( .C1(n10544), .C2(n10492), .A(n10491), .B(n10490), .ZN(
        n10555) );
  AOI22_X1 U11556 ( .A1(n10547), .A2(n10493), .B1(n10555), .B2(n10545), .ZN(
        P2_U3402) );
  INV_X1 U11557 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U11558 ( .A1(n10494), .A2(n10544), .ZN(n10497) );
  NAND2_X1 U11559 ( .A1(n10495), .A2(n10537), .ZN(n10496) );
  AND3_X1 U11560 ( .A1(n10498), .A2(n10497), .A3(n10496), .ZN(n10556) );
  AOI22_X1 U11561 ( .A1(n10547), .A2(n10499), .B1(n10556), .B2(n10545), .ZN(
        P2_U3405) );
  INV_X1 U11562 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10506) );
  AND3_X1 U11563 ( .A1(n10501), .A2(n10500), .A3(n10544), .ZN(n10504) );
  INV_X1 U11564 ( .A(n10502), .ZN(n10503) );
  AOI211_X1 U11565 ( .C1(n10537), .C2(n10505), .A(n10504), .B(n10503), .ZN(
        n10557) );
  AOI22_X1 U11566 ( .A1(n10547), .A2(n10506), .B1(n10557), .B2(n10545), .ZN(
        P2_U3408) );
  INV_X1 U11567 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10512) );
  INV_X1 U11568 ( .A(n10511), .ZN(n10508) );
  OAI22_X1 U11569 ( .A1(n10508), .A2(n10527), .B1(n10507), .B2(n10539), .ZN(
        n10510) );
  AOI211_X1 U11570 ( .C1(n10524), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10559) );
  AOI22_X1 U11571 ( .A1(n10547), .A2(n10512), .B1(n10559), .B2(n10545), .ZN(
        P2_U3411) );
  INV_X1 U11572 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U11573 ( .A1(n10514), .A2(n10544), .B1(n10537), .B2(n10513), .ZN(
        n10515) );
  AND2_X1 U11574 ( .A1(n10516), .A2(n10515), .ZN(n10561) );
  AOI22_X1 U11575 ( .A1(n10547), .A2(n10517), .B1(n10561), .B2(n10545), .ZN(
        P2_U3414) );
  INV_X1 U11576 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10525) );
  INV_X1 U11577 ( .A(n10518), .ZN(n10519) );
  OAI22_X1 U11578 ( .A1(n10520), .A2(n10527), .B1(n10519), .B2(n10539), .ZN(
        n10522) );
  AOI211_X1 U11579 ( .C1(n10524), .C2(n10523), .A(n10522), .B(n10521), .ZN(
        n10563) );
  AOI22_X1 U11580 ( .A1(n10547), .A2(n10525), .B1(n10563), .B2(n10545), .ZN(
        P2_U3417) );
  INV_X1 U11581 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10531) );
  OAI22_X1 U11582 ( .A1(n10528), .A2(n10527), .B1(n10526), .B2(n10539), .ZN(
        n10529) );
  NOR2_X1 U11583 ( .A1(n10530), .A2(n10529), .ZN(n10565) );
  AOI22_X1 U11584 ( .A1(n10547), .A2(n10531), .B1(n10565), .B2(n10545), .ZN(
        P2_U3420) );
  INV_X1 U11585 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10538) );
  INV_X1 U11586 ( .A(n10544), .ZN(n10532) );
  NOR2_X1 U11587 ( .A1(n10533), .A2(n10532), .ZN(n10535) );
  AOI211_X1 U11588 ( .C1(n10537), .C2(n10536), .A(n10535), .B(n10534), .ZN(
        n10567) );
  AOI22_X1 U11589 ( .A1(n10547), .A2(n10538), .B1(n10567), .B2(n10545), .ZN(
        P2_U3423) );
  INV_X1 U11590 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10546) );
  NOR2_X1 U11591 ( .A1(n10540), .A2(n10539), .ZN(n10542) );
  AOI211_X1 U11592 ( .C1(n10544), .C2(n10543), .A(n10542), .B(n10541), .ZN(
        n10569) );
  AOI22_X1 U11593 ( .A1(n10547), .A2(n10546), .B1(n10569), .B2(n10545), .ZN(
        P2_U3426) );
  AOI22_X1 U11594 ( .A1(n10570), .A2(n10549), .B1(n10548), .B2(n10568), .ZN(
        P2_U3460) );
  AOI22_X1 U11595 ( .A1(n10570), .A2(n10551), .B1(n10550), .B2(n10568), .ZN(
        P2_U3461) );
  AOI22_X1 U11596 ( .A1(n10570), .A2(n10553), .B1(n10552), .B2(n10568), .ZN(
        P2_U3462) );
  AOI22_X1 U11597 ( .A1(n10570), .A2(n10555), .B1(n10554), .B2(n10568), .ZN(
        P2_U3463) );
  AOI22_X1 U11598 ( .A1(n10570), .A2(n10556), .B1(n4995), .B2(n10568), .ZN(
        P2_U3464) );
  AOI22_X1 U11599 ( .A1(n10570), .A2(n10557), .B1(n6742), .B2(n10568), .ZN(
        P2_U3465) );
  AOI22_X1 U11600 ( .A1(n10570), .A2(n10559), .B1(n10558), .B2(n10568), .ZN(
        P2_U3466) );
  AOI22_X1 U11601 ( .A1(n10570), .A2(n10561), .B1(n10560), .B2(n10568), .ZN(
        P2_U3467) );
  AOI22_X1 U11602 ( .A1(n10570), .A2(n10563), .B1(n10562), .B2(n10568), .ZN(
        P2_U3468) );
  AOI22_X1 U11603 ( .A1(n10570), .A2(n10565), .B1(n10564), .B2(n10568), .ZN(
        P2_U3469) );
  AOI22_X1 U11604 ( .A1(n10570), .A2(n10567), .B1(n10566), .B2(n10568), .ZN(
        P2_U3470) );
  AOI22_X1 U11605 ( .A1(n10570), .A2(n10569), .B1(n6713), .B2(n10568), .ZN(
        P2_U3471) );
  NOR2_X1 U11606 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  XOR2_X1 U11607 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10573), .Z(ADD_1068_U5) );
  XOR2_X1 U11608 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11609 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10575), .A(n10574), 
        .ZN(n10576) );
  XOR2_X1 U11610 ( .A(n10576), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11611 ( .A(n10578), .B(n10577), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11612 ( .A(n10580), .B(n10579), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11613 ( .A(n10582), .B(n10581), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11614 ( .A(n10584), .B(n10583), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11615 ( .A(n10586), .B(n10585), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11616 ( .A(n10588), .B(n10587), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11617 ( .A(n10590), .B(n10589), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11618 ( .A(n10592), .B(n10591), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11619 ( .A(n10594), .B(n10593), .ZN(ADD_1068_U47) );
  XOR2_X1 U11620 ( .A(n10596), .B(n10595), .Z(ADD_1068_U54) );
  XNOR2_X1 U11621 ( .A(n10598), .B(n10597), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11622 ( .A(n10600), .B(n10599), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11623 ( .A(n10602), .B(n10601), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11624 ( .A(n10604), .B(n10603), .ZN(ADD_1068_U50) );
  XOR2_X1 U11625 ( .A(n10606), .B(n10605), .Z(ADD_1068_U53) );
  XNOR2_X1 U11626 ( .A(n10608), .B(n10607), .ZN(ADD_1068_U52) );
  INV_X2 U5080 ( .A(n6884), .ZN(n5873) );
  CLKBUF_X3 U5127 ( .A(n8151), .Z(n4666) );
endmodule

