

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320;

  INV_X2 U11055 ( .A(n17810), .ZN(n17837) );
  INV_X2 U11056 ( .A(n17923), .ZN(n17908) );
  INV_X1 U11057 ( .A(n21191), .ZN(n17869) );
  NAND2_X2 U11058 ( .A1(n20931), .A2(n10951), .ZN(n21112) );
  XNOR2_X1 U11059 ( .A(n12785), .B(n12784), .ZN(n12786) );
  INV_X1 U11060 ( .A(n15212), .ZN(n11337) );
  NAND3_X1 U11061 ( .A1(n14838), .A2(n20028), .A3(n11622), .ZN(n20738) );
  XNOR2_X1 U11062 ( .A(n13172), .B(n13173), .ZN(n14191) );
  AND2_X2 U11063 ( .A1(n12440), .A2(n19183), .ZN(n12467) );
  CLKBUF_X2 U11064 ( .A(n14067), .Z(n10980) );
  AND2_X1 U11065 ( .A1(n12978), .A2(n14272), .ZN(n13684) );
  INV_X1 U11066 ( .A(n20625), .ZN(n20597) );
  AND2_X1 U11067 ( .A1(n11966), .A2(n11963), .ZN(n19027) );
  CLKBUF_X1 U11068 ( .A(n12946), .Z(n15139) );
  AND2_X1 U11069 ( .A1(n15897), .A2(n13958), .ZN(n15865) );
  INV_X1 U11070 ( .A(n14569), .ZN(n15883) );
  CLKBUF_X2 U11071 ( .A(n11988), .Z(n16036) );
  AND2_X1 U11072 ( .A1(n11260), .A2(n15891), .ZN(n15870) );
  AND2_X1 U11073 ( .A1(n11975), .A2(n15891), .ZN(n15871) );
  CLKBUF_X2 U11074 ( .A(n11482), .Z(n17262) );
  CLKBUF_X2 U11075 ( .A(n11433), .Z(n17497) );
  INV_X1 U11076 ( .A(n17261), .ZN(n17463) );
  CLKBUF_X1 U11077 ( .A(n11433), .Z(n17462) );
  CLKBUF_X2 U11078 ( .A(n11435), .Z(n10960) );
  CLKBUF_X2 U11079 ( .A(n14406), .Z(n15000) );
  CLKBUF_X2 U11080 ( .A(n12941), .Z(n10966) );
  NAND2_X1 U11081 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20712), .ZN(
        n11405) );
  INV_X2 U11082 ( .A(n19597), .ZN(n12379) );
  NAND2_X1 U11083 ( .A1(n11878), .A2(n11860), .ZN(n12420) );
  AND2_X1 U11084 ( .A1(n12826), .A2(n11213), .ZN(n12923) );
  AND2_X2 U11085 ( .A1(n14042), .A2(n14063), .ZN(n12941) );
  NOR2_X2 U11086 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12830) );
  INV_X1 U11087 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11352) );
  NOR2_X2 U11088 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13975) );
  CLKBUF_X2 U11090 ( .A(n12951), .Z(n15095) );
  CLKBUF_X2 U11091 ( .A(n12928), .Z(n15146) );
  AND2_X1 U11092 ( .A1(n15891), .A2(n13970), .ZN(n15876) );
  AND2_X1 U11093 ( .A1(n15891), .A2(n11980), .ZN(n15875) );
  OR2_X1 U11094 ( .A1(n15895), .A2(n13958), .ZN(n15874) );
  MUX2_X1 U11095 ( .A(n11875), .B(n11874), .S(n19410), .Z(n11876) );
  NOR2_X1 U11096 ( .A1(n11954), .A2(n11953), .ZN(n11972) );
  INV_X1 U11097 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13952) );
  CLKBUF_X2 U11098 ( .A(n12752), .Z(n15224) );
  BUF_X1 U11099 ( .A(n11885), .Z(n12374) );
  AND3_X2 U11100 ( .A1(n12168), .A2(n11752), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11979) );
  INV_X1 U11101 ( .A(n14571), .ZN(n15884) );
  AND2_X1 U11102 ( .A1(n15897), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14809) );
  INV_X1 U11103 ( .A(n11855), .ZN(n11084) );
  AND2_X1 U11104 ( .A1(n11986), .A2(n13958), .ZN(n15882) );
  INV_X1 U11105 ( .A(n13348), .ZN(n13390) );
  CLKBUF_X3 U11106 ( .A(n12855), .Z(n13315) );
  INV_X1 U11107 ( .A(n12970), .ZN(n13435) );
  NAND2_X1 U11108 ( .A1(n11083), .A2(n11927), .ZN(n12664) );
  AND2_X1 U11109 ( .A1(n11962), .A2(n11965), .ZN(n12087) );
  AND2_X1 U11110 ( .A1(n11966), .A2(n11960), .ZN(n12084) );
  NOR2_X1 U11111 ( .A1(n12978), .A2(n14272), .ZN(n12985) );
  NAND2_X1 U11112 ( .A1(n13315), .A2(n15511), .ZN(n12967) );
  AND2_X2 U11113 ( .A1(n14272), .A2(n21915), .ZN(n21195) );
  NOR2_X1 U11114 ( .A1(n14799), .A2(n13376), .ZN(n14791) );
  XNOR2_X1 U11115 ( .A(n13131), .B(n14070), .ZN(n21802) );
  INV_X1 U11116 ( .A(n12965), .ZN(n13056) );
  OR2_X1 U11117 ( .A1(n16167), .A2(n12655), .ZN(n16155) );
  NAND2_X1 U11118 ( .A1(n12438), .A2(n12437), .ZN(n15269) );
  INV_X1 U11119 ( .A(n12440), .ZN(n11871) );
  BUF_X1 U11120 ( .A(n11939), .Z(n11944) );
  NAND2_X1 U11121 ( .A1(n20028), .A2(n20721), .ZN(n14840) );
  NOR4_X1 U11122 ( .A1(n20597), .A2(n11686), .A3(n11619), .A4(n11618), .ZN(
        n11620) );
  AND2_X1 U11123 ( .A1(n14709), .A2(n14270), .ZN(n21586) );
  INV_X1 U11124 ( .A(n10970), .ZN(n14846) );
  INV_X1 U11125 ( .A(n20993), .ZN(n21063) );
  INV_X1 U11126 ( .A(n21586), .ZN(n21600) );
  NAND2_X1 U11127 ( .A1(n21164), .A2(n21163), .ZN(n21191) );
  NOR2_X2 U11128 ( .A1(n20527), .A2(n20708), .ZN(n20709) );
  INV_X1 U11129 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20761) );
  CLKBUF_X3 U11130 ( .A(n11440), .Z(n17499) );
  CLKBUF_X3 U11131 ( .A(n11440), .Z(n17435) );
  INV_X1 U11132 ( .A(n11758), .ZN(n11986) );
  INV_X1 U11133 ( .A(n13039), .ZN(n10959) );
  NAND2_X2 U11134 ( .A1(n11862), .A2(n14524), .ZN(n11854) );
  INV_X2 U11135 ( .A(n19410), .ZN(n11878) );
  INV_X2 U11136 ( .A(n16112), .ZN(n16046) );
  OAI21_X2 U11137 ( .B1(n12060), .B2(n12059), .A(n12058), .ZN(n12160) );
  OR2_X2 U11138 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  AND4_X4 U11139 ( .A1(n12897), .A2(n12896), .A3(n12895), .A4(n12894), .ZN(
        n12970) );
  AND4_X2 U11140 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        n12894) );
  NOR2_X2 U11141 ( .A1(n14127), .A2(n14128), .ZN(n14126) );
  OR2_X4 U11142 ( .A1(n16416), .A2(n16659), .ZN(n17007) );
  INV_X2 U11144 ( .A(n20739), .ZN(n10948) );
  INV_X1 U11145 ( .A(n15973), .ZN(n10949) );
  XNOR2_X2 U11146 ( .A(n13108), .B(n13107), .ZN(n14067) );
  OAI21_X2 U11147 ( .B1(n21850), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13091), 
        .ZN(n13108) );
  AND2_X4 U11148 ( .A1(n12830), .A2(n13698), .ZN(n13046) );
  AND3_X2 U11149 ( .A1(n12168), .A2(n11752), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10950) );
  XNOR2_X2 U11150 ( .A(n13104), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16953) );
  NAND2_X2 U11151 ( .A1(n13778), .A2(n13064), .ZN(n13104) );
  XNOR2_X2 U11152 ( .A(n15969), .B(n11375), .ZN(n16081) );
  NAND2_X2 U11153 ( .A1(n16085), .A2(n11376), .ZN(n15969) );
  AOI211_X2 U11154 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19958), .A(
        n19957), .B(n19956), .ZN(n19959) );
  XNOR2_X2 U11155 ( .A(n12222), .B(n12221), .ZN(n14610) );
  NAND2_X2 U11156 ( .A1(n12220), .A2(n18082), .ZN(n12222) );
  NOR2_X1 U11157 ( .A1(n11404), .A2(n20740), .ZN(n11440) );
  AOI22_X2 U11158 ( .A1(n17786), .A2(n17836), .B1(n17908), .B2(n20869), .ZN(
        n17821) );
  NOR2_X4 U11159 ( .A1(n11733), .A2(n17922), .ZN(n17836) );
  INV_X1 U11160 ( .A(n20946), .ZN(n10951) );
  CLKBUF_X3 U11161 ( .A(n11449), .Z(n10952) );
  CLKBUF_X3 U11162 ( .A(n11449), .Z(n10953) );
  INV_X1 U11163 ( .A(n11483), .ZN(n10954) );
  INV_X1 U11164 ( .A(n10954), .ZN(n10955) );
  INV_X1 U11165 ( .A(n10954), .ZN(n10956) );
  INV_X1 U11166 ( .A(n10954), .ZN(n10957) );
  NOR2_X1 U11167 ( .A1(n11405), .A2(n20740), .ZN(n11483) );
  NAND2_X1 U11168 ( .A1(n14387), .A2(n12789), .ZN(n12793) );
  BUF_X1 U11169 ( .A(n12791), .Z(n12795) );
  NAND2_X1 U11170 ( .A1(n11139), .A2(n12061), .ZN(n12785) );
  INV_X4 U11171 ( .A(n13221), .ZN(n13212) );
  AND2_X1 U11172 ( .A1(n11966), .A2(n11957), .ZN(n12190) );
  NOR2_X1 U11173 ( .A1(n17828), .A2(n17827), .ZN(n17826) );
  NAND2_X1 U11174 ( .A1(n20084), .A2(n20949), .ZN(n20995) );
  NAND2_X1 U11175 ( .A1(n20949), .A2(n20520), .ZN(n21132) );
  BUF_X1 U11176 ( .A(n13838), .Z(n18499) );
  NAND2_X1 U11177 ( .A1(n11218), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13065) );
  AND2_X1 U11178 ( .A1(n14030), .A2(n19597), .ZN(n12433) );
  AND2_X1 U11179 ( .A1(n12411), .A2(n11869), .ZN(n11877) );
  INV_X1 U11180 ( .A(n12420), .ZN(n12758) );
  NAND4_X2 U11182 ( .A1(n12957), .A2(n12958), .A3(n12959), .A4(n12956), .ZN(
        n14272) );
  NAND2_X1 U11183 ( .A1(n12853), .A2(n12852), .ZN(n12986) );
  AND4_X1 U11184 ( .A1(n12950), .A2(n12949), .A3(n12948), .A4(n12947), .ZN(
        n12957) );
  AND4_X1 U11185 ( .A1(n12945), .A2(n12944), .A3(n12943), .A4(n12942), .ZN(
        n12958) );
  INV_X2 U11186 ( .A(n21373), .ZN(n13790) );
  BUF_X2 U11187 ( .A(n13080), .Z(n10981) );
  CLKBUF_X2 U11188 ( .A(n14651), .Z(n15005) );
  BUF_X2 U11189 ( .A(n12923), .Z(n15145) );
  BUF_X2 U11190 ( .A(n12906), .Z(n15138) );
  INV_X2 U11191 ( .A(n21105), .ZN(n10958) );
  CLKBUF_X2 U11192 ( .A(n11461), .Z(n17220) );
  CLKBUF_X2 U11193 ( .A(n13045), .Z(n15147) );
  NAND2_X1 U11194 ( .A1(n11406), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11404) );
  AND2_X1 U11195 ( .A1(n11082), .A2(n12329), .ZN(n16245) );
  NAND2_X1 U11196 ( .A1(n16268), .A2(n10990), .ZN(n12329) );
  AND2_X1 U11197 ( .A1(n12817), .A2(n12816), .ZN(n12818) );
  NOR2_X1 U11198 ( .A1(n16327), .A2(n16326), .ZN(n16331) );
  OAI21_X1 U11199 ( .B1(n15593), .B2(n15592), .A(n15591), .ZN(n15721) );
  OAI21_X1 U11200 ( .B1(n16246), .B2(n11224), .A(n15216), .ZN(n11222) );
  NOR2_X1 U11201 ( .A1(n16246), .A2(n15271), .ZN(n16238) );
  OAI21_X1 U11202 ( .B1(n16351), .B2(n16323), .A(n16322), .ZN(n16325) );
  OAI21_X1 U11203 ( .B1(n16374), .B2(n16319), .A(n16320), .ZN(n16351) );
  NAND2_X1 U11204 ( .A1(n12810), .A2(n12809), .ZN(n16339) );
  AOI21_X1 U11205 ( .B1(n15257), .B2(n15317), .A(n15256), .ZN(n15304) );
  AND2_X1 U11206 ( .A1(n15317), .A2(n15316), .ZN(n15597) );
  XNOR2_X1 U11207 ( .A(n11244), .B(n11243), .ZN(n15295) );
  NAND2_X1 U11208 ( .A1(n12805), .A2(n12804), .ZN(n16977) );
  NAND2_X1 U11209 ( .A1(n12798), .A2(n12797), .ZN(n14723) );
  OAI211_X1 U11210 ( .C1(n12794), .C2(n12795), .A(n11369), .B(n11021), .ZN(
        n14608) );
  XNOR2_X1 U11211 ( .A(n16091), .B(n15949), .ZN(n16087) );
  NOR2_X2 U11212 ( .A1(n16103), .A2(n16095), .ZN(n16094) );
  NAND2_X1 U11213 ( .A1(n15175), .A2(n15174), .ZN(n15173) );
  NAND2_X1 U11214 ( .A1(n16100), .A2(n12742), .ZN(n16103) );
  NAND2_X1 U11215 ( .A1(n16093), .A2(n16092), .ZN(n16091) );
  AOI21_X1 U11216 ( .B1(n11109), .B2(n11055), .A(n13402), .ZN(n11107) );
  NOR2_X1 U11217 ( .A1(n14830), .A2(n16109), .ZN(n16100) );
  AND2_X1 U11218 ( .A1(n11309), .A2(n11308), .ZN(n11307) );
  NAND2_X1 U11219 ( .A1(n11254), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U11220 ( .A1(n12115), .A2(n12114), .ZN(n12799) );
  AND2_X2 U11221 ( .A1(n14239), .A2(n11051), .ZN(n14498) );
  NAND2_X1 U11222 ( .A1(n11163), .A2(n13212), .ZN(n11313) );
  AND2_X1 U11223 ( .A1(n12162), .A2(n12785), .ZN(n14353) );
  AND3_X1 U11224 ( .A1(n17665), .A2(n17597), .A3(n11246), .ZN(n17660) );
  NOR2_X2 U11225 ( .A1(n14240), .A2(n14241), .ZN(n14239) );
  NAND2_X1 U11226 ( .A1(n13220), .A2(n11164), .ZN(n11163) );
  NAND2_X1 U11227 ( .A1(n12160), .A2(n12161), .ZN(n12162) );
  OR2_X1 U11228 ( .A1(n14155), .A2(n14154), .ZN(n14240) );
  NAND2_X1 U11229 ( .A1(n17667), .A2(n17666), .ZN(n17665) );
  AND2_X1 U11230 ( .A1(n15680), .A2(n13223), .ZN(n15669) );
  AND2_X1 U11231 ( .A1(n15693), .A2(n15696), .ZN(n15680) );
  NOR2_X1 U11232 ( .A1(n14107), .A2(n14158), .ZN(n14237) );
  AND2_X1 U11233 ( .A1(n12216), .A2(n12215), .ZN(n12800) );
  AND2_X1 U11234 ( .A1(n12112), .A2(n12111), .ZN(n12114) );
  OR2_X1 U11235 ( .A1(n12197), .A2(n12196), .ZN(n12216) );
  NAND2_X1 U11236 ( .A1(n13204), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13205) );
  AND2_X1 U11237 ( .A1(n13221), .A2(n13217), .ZN(n19933) );
  OR2_X1 U11238 ( .A1(n16585), .A2(n16197), .ZN(n16560) );
  NAND2_X1 U11239 ( .A1(n20520), .A2(n17869), .ZN(n17922) );
  NAND2_X1 U11240 ( .A1(n20084), .A2(n17869), .ZN(n17923) );
  AOI22_X1 U11241 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19136), .B1(
        n12191), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12037) );
  OAI22_X1 U11242 ( .A1(n19038), .A2(n14568), .B1(n11946), .B2(n19161), .ZN(
        n11947) );
  OAI22_X1 U11243 ( .A1(n14565), .A2(n19053), .B1(n11950), .B2(n11949), .ZN(
        n11954) );
  NAND2_X1 U11244 ( .A1(n14087), .A2(n14086), .ZN(n14131) );
  INV_X1 U11245 ( .A(n19161), .ZN(n12191) );
  XNOR2_X1 U11246 ( .A(n13198), .B(n13197), .ZN(n14251) );
  INV_X1 U11247 ( .A(n12185), .ZN(n19080) );
  NAND2_X1 U11248 ( .A1(n13869), .A2(n13868), .ZN(n13943) );
  AOI22_X1 U11249 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n12190), .B1(
        n19116), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12039) );
  OAI21_X2 U11250 ( .B1(n20018), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21191), 
        .ZN(n17918) );
  INV_X1 U11251 ( .A(n12036), .ZN(n19184) );
  INV_X1 U11252 ( .A(n12190), .ZN(n19038) );
  AND2_X1 U11253 ( .A1(n13198), .A2(n13278), .ZN(n13207) );
  INV_X1 U11254 ( .A(n19133), .ZN(n19136) );
  INV_X1 U11255 ( .A(n12084), .ZN(n19053) );
  AND2_X1 U11256 ( .A1(n11964), .A2(n11957), .ZN(n19116) );
  AND2_X1 U11257 ( .A1(n16315), .A2(n11152), .ZN(n11151) );
  INV_X1 U11258 ( .A(n12079), .ZN(n10961) );
  NAND2_X1 U11259 ( .A1(n13187), .A2(n13186), .ZN(n13198) );
  OR2_X1 U11260 ( .A1(n15464), .A2(n15457), .ZN(n15459) );
  AND2_X1 U11261 ( .A1(n11962), .A2(n11960), .ZN(n12185) );
  NAND2_X1 U11262 ( .A1(n13768), .A2(n13767), .ZN(n13920) );
  AND2_X1 U11263 ( .A1(n18499), .A2(n13944), .ZN(n11964) );
  AND2_X1 U11264 ( .A1(n13944), .A2(n11138), .ZN(n11961) );
  NAND2_X1 U11265 ( .A1(n13763), .A2(n13762), .ZN(n13768) );
  NOR2_X2 U11266 ( .A1(n21112), .A2(n21126), .ZN(n20949) );
  NOR2_X1 U11267 ( .A1(n18036), .A2(n11945), .ZN(n11963) );
  AND2_X1 U11268 ( .A1(n18427), .A2(n18036), .ZN(n11957) );
  OAI21_X1 U11269 ( .B1(n18036), .B2(n14032), .A(n13727), .ZN(n13846) );
  OR2_X1 U11270 ( .A1(n15484), .A2(n15483), .ZN(n15486) );
  XNOR2_X1 U11271 ( .A(n11934), .B(n11933), .ZN(n13838) );
  NOR2_X1 U11272 ( .A1(n18036), .A2(n11944), .ZN(n11960) );
  OR2_X1 U11273 ( .A1(n21199), .A2(n14261), .ZN(n14709) );
  NAND2_X2 U11274 ( .A1(n19892), .A2(n15511), .ZN(n15509) );
  NAND2_X2 U11275 ( .A1(n11940), .A2(n11938), .ZN(n18036) );
  NAND2_X1 U11276 ( .A1(n11216), .A2(n13124), .ZN(n14070) );
  OR2_X2 U11278 ( .A1(n13557), .A2(n12978), .ZN(n13603) );
  AND2_X1 U11279 ( .A1(n11927), .A2(n11895), .ZN(n11933) );
  OR2_X1 U11280 ( .A1(n11937), .A2(n11936), .ZN(n11938) );
  AOI21_X1 U11281 ( .B1(n11906), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11867), .ZN(n11891) );
  INV_X2 U11282 ( .A(n12703), .ZN(n15223) );
  OR2_X1 U11283 ( .A1(n12460), .A2(n12457), .ZN(n14082) );
  NOR2_X1 U11284 ( .A1(n20078), .A2(n20030), .ZN(n20077) );
  AOI21_X1 U11285 ( .B1(n11930), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11890), .ZN(n11892) );
  NOR2_X1 U11286 ( .A1(n14097), .A2(n11191), .ZN(n14257) );
  XNOR2_X1 U11287 ( .A(n11156), .B(n13033), .ZN(n21749) );
  NAND2_X1 U11288 ( .A1(n13075), .A2(n13074), .ZN(n13076) );
  NAND2_X1 U11289 ( .A1(n12983), .A2(n13035), .ZN(n12994) );
  INV_X2 U11290 ( .A(n15821), .ZN(n19586) );
  AOI22_X1 U11291 ( .A1(n13987), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12407), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11897) );
  INV_X2 U11292 ( .A(n20030), .ZN(n20080) );
  NAND2_X1 U11293 ( .A1(n11397), .A2(n11118), .ZN(n13034) );
  AND2_X1 U11294 ( .A1(n11302), .A2(n13024), .ZN(n11301) );
  CLKBUF_X1 U11295 ( .A(n12376), .Z(n13711) );
  NAND3_X1 U11296 ( .A1(n11877), .A2(n11876), .A3(n11903), .ZN(n11908) );
  OR2_X1 U11297 ( .A1(n12434), .A2(n18021), .ZN(n11914) );
  AND2_X1 U11298 ( .A1(n12993), .A2(n13446), .ZN(n11118) );
  AOI21_X1 U11299 ( .B1(n11248), .B2(n11249), .A(n11500), .ZN(n11502) );
  AOI21_X1 U11300 ( .B1(n13021), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11305), 
        .ZN(n11304) );
  AND2_X1 U11301 ( .A1(n11635), .A2(n11504), .ZN(n11507) );
  NOR2_X1 U11302 ( .A1(n17131), .A2(n11680), .ZN(n11617) );
  CLKBUF_X1 U11303 ( .A(n11854), .Z(n13750) );
  XNOR2_X1 U11304 ( .A(n11499), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11248) );
  AOI21_X1 U11305 ( .B1(n18898), .B2(n18807), .A(n20710), .ZN(n11696) );
  NAND2_X1 U11306 ( .A1(n11115), .A2(n12979), .ZN(n12991) );
  INV_X1 U11307 ( .A(n11880), .ZN(n12438) );
  NOR2_X1 U11308 ( .A1(n11639), .A2(n20570), .ZN(n11504) );
  NAND2_X1 U11309 ( .A1(n11498), .A2(n11639), .ZN(n11499) );
  AND2_X1 U11310 ( .A1(n11859), .A2(n11864), .ZN(n12401) );
  NOR2_X1 U11311 ( .A1(n17910), .A2(n17916), .ZN(n17909) );
  INV_X1 U11312 ( .A(n11682), .ZN(n20586) );
  INV_X1 U11313 ( .A(n12985), .ZN(n15291) );
  CLKBUF_X1 U11314 ( .A(n11862), .Z(n13740) );
  OR2_X1 U11315 ( .A1(n13441), .A2(n21716), .ZN(n13313) );
  MUX2_X1 U11316 ( .A(n12912), .B(n12960), .S(n12965), .Z(n12913) );
  OR2_X1 U11317 ( .A1(n13442), .A2(n13342), .ZN(n13695) );
  NAND2_X1 U11318 ( .A1(n11448), .A2(n20698), .ZN(n11639) );
  NAND2_X1 U11319 ( .A1(n20703), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17916) );
  INV_X1 U11320 ( .A(n12967), .ZN(n13674) );
  AND2_X2 U11321 ( .A1(n12135), .A2(n12134), .ZN(n15212) );
  CLKBUF_X1 U11322 ( .A(n12980), .Z(n13441) );
  NAND3_X1 U11323 ( .A1(n11536), .A2(n11535), .A3(n11534), .ZN(n20520) );
  CLKBUF_X1 U11324 ( .A(n11872), .Z(n11873) );
  CLKBUF_X1 U11325 ( .A(n14524), .Z(n19291) );
  INV_X1 U11326 ( .A(n14272), .ZN(n21716) );
  XNOR2_X1 U11327 ( .A(n20698), .B(n11497), .ZN(n17910) );
  OR3_X2 U11328 ( .A1(n11124), .A2(n11584), .A3(n11585), .ZN(n11609) );
  INV_X2 U11329 ( .A(U212), .ZN(n10962) );
  OR2_X1 U11330 ( .A1(n13017), .A2(n13016), .ZN(n13054) );
  OR2_X1 U11331 ( .A1(n13006), .A2(n13005), .ZN(n13206) );
  NOR2_X1 U11332 ( .A1(n13315), .A2(n21898), .ZN(n14656) );
  NAND2_X2 U11333 ( .A1(U214), .A2(n19972), .ZN(n20013) );
  NAND2_X2 U11334 ( .A1(n11802), .A2(n11801), .ZN(n11858) );
  NAND4_X1 U11335 ( .A1(n12834), .A2(n12833), .A3(n12832), .A4(n12831), .ZN(
        n12855) );
  NAND2_X1 U11336 ( .A1(n11849), .A2(n13958), .ZN(n11850) );
  AND4_X1 U11337 ( .A1(n12847), .A2(n12846), .A3(n12845), .A4(n12844), .ZN(
        n12853) );
  NAND2_X1 U11338 ( .A1(n12911), .A2(n11396), .ZN(n12965) );
  AND4_X1 U11339 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12936) );
  AND4_X1 U11340 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12959) );
  BUF_X2 U11341 ( .A(n12901), .Z(n15144) );
  AND4_X1 U11342 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12873) );
  AND4_X1 U11343 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11770) );
  AND4_X1 U11344 ( .A1(n12863), .A2(n12862), .A3(n12861), .A4(n12860), .ZN(
        n12874) );
  AND4_X1 U11345 ( .A1(n12838), .A2(n12837), .A3(n12836), .A4(n12835), .ZN(
        n12843) );
  AND4_X1 U11346 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12934) );
  AND4_X1 U11347 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n13958), .ZN(
        n11756) );
  AND4_X1 U11348 ( .A1(n12859), .A2(n12858), .A3(n12857), .A4(n12856), .ZN(
        n12875) );
  AND4_X1 U11349 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12935) );
  AND4_X1 U11350 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12933) );
  AND2_X2 U11351 ( .A1(n21872), .A2(n13776), .ZN(n19952) );
  AND4_X1 U11352 ( .A1(n12879), .A2(n12878), .A3(n12877), .A4(n12876), .ZN(
        n12897) );
  AND4_X1 U11353 ( .A1(n12905), .A2(n12904), .A3(n12903), .A4(n12902), .ZN(
        n12911) );
  AND4_X1 U11354 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n12895) );
  AND4_X1 U11355 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12852) );
  AND4_X1 U11356 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  AND4_X1 U11357 ( .A1(n12825), .A2(n12824), .A3(n12823), .A4(n12822), .ZN(
        n12834) );
  AND4_X1 U11358 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12872) );
  AND2_X1 U11359 ( .A1(n12829), .A2(n12828), .ZN(n12832) );
  NAND2_X2 U11360 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17128), .ZN(n17124) );
  NAND2_X2 U11361 ( .A1(n20082), .A2(n17520), .ZN(n21105) );
  NAND2_X2 U11362 ( .A1(n17128), .A2(n21682), .ZN(n17125) );
  CLKBUF_X1 U11363 ( .A(n18386), .Z(n18371) );
  BUF_X4 U11364 ( .A(n11434), .Z(n17491) );
  BUF_X2 U11365 ( .A(n13044), .Z(n12999) );
  INV_X2 U11366 ( .A(n10959), .ZN(n10963) );
  AND2_X2 U11367 ( .A1(n16036), .A2(n13958), .ZN(n15866) );
  AND2_X1 U11368 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  BUF_X2 U11369 ( .A(n14411), .Z(n15100) );
  INV_X2 U11370 ( .A(n18890), .ZN(U215) );
  AND4_X1 U11371 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        n12956) );
  INV_X4 U11372 ( .A(n17354), .ZN(n10965) );
  AND2_X2 U11373 ( .A1(n11213), .A2(n14063), .ZN(n12901) );
  OR2_X1 U11374 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20729), .ZN(
        n20739) );
  AND2_X1 U11375 ( .A1(n12826), .A2(n14055), .ZN(n12906) );
  AOI22_X1 U11376 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12822) );
  INV_X2 U11377 ( .A(n19722), .ZN(n19776) );
  AND2_X1 U11378 ( .A1(n20918), .A2(n20915), .ZN(n10969) );
  AND2_X1 U11379 ( .A1(n11274), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11975) );
  AND2_X2 U11380 ( .A1(n12366), .A2(n12168), .ZN(n11988) );
  NAND2_X1 U11381 ( .A1(n20761), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20740) );
  AND2_X2 U11382 ( .A1(n14063), .A2(n14055), .ZN(n12951) );
  AND2_X2 U11383 ( .A1(n14063), .A2(n12830), .ZN(n13045) );
  NOR2_X2 U11384 ( .A1(n21659), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22319) );
  INV_X1 U11385 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13985) );
  AND2_X1 U11386 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12366) );
  INV_X1 U11387 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12820) );
  AND2_X1 U11388 ( .A1(n12814), .A2(n11227), .ZN(n10967) );
  AND2_X1 U11389 ( .A1(n11226), .A2(n11227), .ZN(n10968) );
  OR2_X1 U11390 ( .A1(n16269), .A2(n15190), .ZN(n16246) );
  NAND3_X1 U11391 ( .A1(n17794), .A2(n10969), .A3(n17554), .ZN(n11245) );
  BUF_X4 U11392 ( .A(n11578), .Z(n17300) );
  BUF_X4 U11393 ( .A(n11578), .Z(n17482) );
  NOR2_X2 U11394 ( .A1(n14252), .A2(n14253), .ZN(n14421) );
  NAND2_X1 U11395 ( .A1(n15327), .A2(n15328), .ZN(n15314) );
  NAND2_X2 U11396 ( .A1(n11765), .A2(n11764), .ZN(n11861) );
  NAND2_X2 U11397 ( .A1(n12309), .A2(n11228), .ZN(n12310) );
  NAND2_X2 U11398 ( .A1(n15199), .A2(n15198), .ZN(n16231) );
  AND2_X2 U11399 ( .A1(n14704), .A2(n14703), .ZN(n10970) );
  AND2_X4 U11400 ( .A1(n17006), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16399) );
  NAND2_X1 U11401 ( .A1(n16339), .A2(n12812), .ZN(n16532) );
  NOR2_X4 U11402 ( .A1(n17007), .A2(n16642), .ZN(n17006) );
  AND2_X1 U11403 ( .A1(n11759), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11763) );
  INV_X2 U11404 ( .A(n11078), .ZN(n12354) );
  NAND2_X2 U11405 ( .A1(n11776), .A2(n11775), .ZN(n11078) );
  NAND4_X2 U11406 ( .A1(n20695), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n20583), .ZN(n20688) );
  XNOR2_X1 U11407 ( .A(n10971), .B(n19959), .ZN(n21380) );
  INV_X1 U11408 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10971) );
  INV_X2 U11409 ( .A(n11758), .ZN(n10972) );
  INV_X2 U11410 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12168) );
  INV_X2 U11411 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11752) );
  AND2_X4 U11412 ( .A1(n11975), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10973) );
  NAND3_X1 U11413 ( .A1(n20752), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n11406), .ZN(n17354) );
  XNOR2_X2 U11414 ( .A(n12799), .B(n12800), .ZN(n12791) );
  BUF_X4 U11415 ( .A(n11592), .Z(n10974) );
  NOR2_X1 U11416 ( .A1(n11404), .A2(n20741), .ZN(n11592) );
  CLKBUF_X2 U11417 ( .A(n11482), .Z(n10975) );
  NOR3_X1 U11418 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11405), .ZN(n11482) );
  AOI21_X2 U11419 ( .B1(n10980), .B2(n13278), .A(n13103), .ZN(n16955) );
  AND2_X2 U11420 ( .A1(n12964), .A2(n12977), .ZN(n13308) );
  AND2_X2 U11421 ( .A1(n12819), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14042) );
  NAND2_X2 U11422 ( .A1(n13038), .A2(n13037), .ZN(n21730) );
  NOR2_X1 U11424 ( .A1(n20089), .A2(n11081), .ZN(n11435) );
  INV_X2 U11425 ( .A(n17261), .ZN(n10976) );
  OR2_X1 U11426 ( .A1(n11405), .A2(n11403), .ZN(n17261) );
  NAND2_X2 U11427 ( .A1(n12963), .A2(n12966), .ZN(n12969) );
  INV_X2 U11428 ( .A(n12855), .ZN(n12963) );
  AND2_X1 U11429 ( .A1(n12826), .A2(n14055), .ZN(n10977) );
  AND2_X1 U11430 ( .A1(n12826), .A2(n14055), .ZN(n10978) );
  NOR2_X4 U11431 ( .A1(n20741), .A2(n20089), .ZN(n11434) );
  NAND2_X1 U11432 ( .A1(n20712), .A2(n11406), .ZN(n20089) );
  AND2_X2 U11433 ( .A1(n12826), .A2(n14042), .ZN(n13080) );
  NAND2_X4 U11434 ( .A1(n13207), .A2(n11162), .ZN(n13221) );
  INV_X1 U11435 ( .A(n13065), .ZN(n13033) );
  NAND2_X2 U11436 ( .A1(n13061), .A2(n13060), .ZN(n13059) );
  NAND2_X2 U11437 ( .A1(n13777), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13778) );
  XNOR2_X2 U11438 ( .A(n13062), .B(n13059), .ZN(n13777) );
  NAND2_X2 U11439 ( .A1(n11310), .A2(n11307), .ZN(n13224) );
  NAND2_X2 U11440 ( .A1(n15692), .A2(n11311), .ZN(n11310) );
  AND2_X2 U11441 ( .A1(n14042), .A2(n13698), .ZN(n13039) );
  OR2_X2 U11442 ( .A1(n12984), .A2(n12961), .ZN(n13323) );
  AND2_X2 U11443 ( .A1(n15454), .A2(n15456), .ZN(n15432) );
  NOR2_X2 U11444 ( .A1(n15365), .A2(n15462), .ZN(n15454) );
  NAND2_X2 U11445 ( .A1(n15173), .A2(n13213), .ZN(n15692) );
  OAI21_X2 U11446 ( .B1(n13671), .B2(n13148), .A(n13027), .ZN(n13791) );
  NAND3_X2 U11447 ( .A1(n12898), .A2(n13435), .A3(n15511), .ZN(n12972) );
  INV_X2 U11448 ( .A(n12969), .ZN(n12898) );
  NOR2_X2 U11449 ( .A1(n15352), .A2(n15353), .ZN(n15341) );
  XNOR2_X2 U11450 ( .A(n12994), .B(n13034), .ZN(n13673) );
  AOI211_X2 U11451 ( .C1(n19946), .C2(n15610), .A(n15609), .B(n15608), .ZN(
        n15611) );
  OAI21_X2 U11453 ( .B1(n15327), .B2(n15328), .A(n15314), .ZN(n15607) );
  AND2_X2 U11454 ( .A1(n15341), .A2(n15340), .ZN(n15327) );
  AND2_X1 U11455 ( .A1(n14055), .A2(n12827), .ZN(n10982) );
  AND2_X4 U11456 ( .A1(n14055), .A2(n12827), .ZN(n10983) );
  AND2_X1 U11457 ( .A1(n12966), .A2(n12978), .ZN(n13278) );
  NAND2_X1 U11458 ( .A1(n12462), .A2(n12461), .ZN(n11330) );
  INV_X1 U11459 ( .A(n14082), .ZN(n12462) );
  INV_X1 U11460 ( .A(n14163), .ZN(n11329) );
  NAND2_X1 U11461 ( .A1(n12970), .A2(n12966), .ZN(n12973) );
  AND2_X1 U11462 ( .A1(n13748), .A2(n13747), .ZN(n12452) );
  NAND2_X1 U11463 ( .A1(n11018), .A2(n12353), .ZN(n11852) );
  NOR2_X1 U11464 ( .A1(n15315), .A2(n11242), .ZN(n11241) );
  INV_X1 U11465 ( .A(n15328), .ZN(n11242) );
  INV_X1 U11466 ( .A(n15494), .ZN(n11187) );
  INV_X1 U11467 ( .A(n11195), .ZN(n11194) );
  OR2_X1 U11468 ( .A1(n14096), .A2(n11196), .ZN(n11195) );
  INV_X1 U11469 ( .A(n14146), .ZN(n11196) );
  NAND2_X1 U11470 ( .A1(n13684), .A2(n13390), .ZN(n13420) );
  AND3_X1 U11471 ( .A1(n12970), .A2(n12963), .A3(n15511), .ZN(n12977) );
  NAND2_X1 U11472 ( .A1(n14272), .A2(n12854), .ZN(n13423) );
  NAND2_X1 U11473 ( .A1(n13325), .A2(n11220), .ZN(n11219) );
  NAND2_X1 U11474 ( .A1(n21915), .A2(n11221), .ZN(n11220) );
  XNOR2_X1 U11475 ( .A(n12665), .B(n12666), .ZN(n12662) );
  AND2_X1 U11476 ( .A1(n13728), .A2(n13740), .ZN(n15990) );
  AND2_X1 U11477 ( .A1(n11291), .A2(n14785), .ZN(n11290) );
  INV_X1 U11478 ( .A(n13833), .ZN(n11332) );
  NAND2_X1 U11479 ( .A1(n11896), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11883) );
  AND2_X1 U11480 ( .A1(n16987), .A2(n11030), .ZN(n11357) );
  INV_X1 U11481 ( .A(n15269), .ZN(n12648) );
  AOI221_X1 U11482 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12332), 
        .C1(n14020), .C2(n12332), .A(n12331), .ZN(n12391) );
  NOR2_X1 U11483 ( .A1(n11404), .A2(n11256), .ZN(n11433) );
  NAND2_X1 U11484 ( .A1(n21143), .A2(n20761), .ZN(n11256) );
  INV_X1 U11485 ( .A(n17665), .ZN(n11524) );
  AND2_X1 U11486 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11513), .ZN(
        n11514) );
  OR2_X1 U11487 ( .A1(n11404), .A2(n11403), .ZN(n11377) );
  NOR2_X1 U11488 ( .A1(n13208), .A2(n21614), .ZN(n11162) );
  AND2_X1 U11489 ( .A1(n16094), .A2(n11046), .ZN(n16055) );
  NOR2_X1 U11490 ( .A1(n11325), .A2(n14206), .ZN(n11324) );
  INV_X1 U11491 ( .A(n14546), .ZN(n11325) );
  INV_X1 U11492 ( .A(n12711), .ZN(n15227) );
  AND2_X1 U11493 ( .A1(n11858), .A2(n19183), .ZN(n12437) );
  NAND2_X1 U11494 ( .A1(n11322), .A2(n14215), .ZN(n11321) );
  INV_X1 U11495 ( .A(n14523), .ZN(n11322) );
  AND2_X1 U11496 ( .A1(n12400), .A2(n18535), .ZN(n12815) );
  AND2_X1 U11497 ( .A1(n14018), .A2(n18535), .ZN(n18538) );
  NAND2_X1 U11498 ( .A1(n18383), .A2(n17021), .ZN(n16226) );
  OR2_X1 U11499 ( .A1(n20935), .A2(n11073), .ZN(n11072) );
  INV_X1 U11500 ( .A(n20936), .ZN(n11075) );
  NAND2_X1 U11501 ( .A1(n21102), .A2(n20937), .ZN(n11074) );
  NAND2_X1 U11502 ( .A1(n11957), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11141) );
  AND2_X2 U11503 ( .A1(n11111), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12826) );
  AOI22_X1 U11504 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15896), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U11505 ( .A1(n12405), .A2(n11349), .ZN(n12382) );
  INV_X1 U11506 ( .A(n11350), .ZN(n11349) );
  OAI21_X1 U11507 ( .B1(n13749), .B2(n12379), .A(n11860), .ZN(n11350) );
  NAND2_X1 U11508 ( .A1(n12147), .A2(n12146), .ZN(n12149) );
  AOI21_X1 U11509 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21153), .A(
        n11662), .ZN(n11663) );
  NOR2_X1 U11510 ( .A1(n11667), .A2(n11666), .ZN(n11662) );
  INV_X1 U11511 ( .A(n13189), .ZN(n13187) );
  NAND2_X1 U11512 ( .A1(n12971), .A2(n11398), .ZN(n11293) );
  AND2_X1 U11513 ( .A1(n12969), .A2(n12970), .ZN(n12971) );
  AOI22_X1 U11514 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12825) );
  AND2_X1 U11515 ( .A1(n14272), .A2(n13435), .ZN(n13078) );
  NAND2_X1 U11516 ( .A1(n11204), .A2(n12343), .ZN(n12386) );
  NAND2_X1 U11517 ( .A1(n12138), .A2(n11146), .ZN(n11204) );
  NAND2_X1 U11518 ( .A1(n11871), .A2(n11870), .ZN(n11880) );
  NAND2_X1 U11519 ( .A1(n11342), .A2(n12660), .ZN(n11341) );
  NOR2_X1 U11520 ( .A1(n16147), .A2(n11343), .ZN(n11342) );
  OR2_X1 U11521 ( .A1(n12799), .A2(n12801), .ZN(n12806) );
  INV_X1 U11522 ( .A(n12800), .ZN(n12801) );
  AND2_X1 U11523 ( .A1(n13728), .A2(n19597), .ZN(n11136) );
  NAND2_X1 U11524 ( .A1(n11078), .A2(n11872), .ZN(n11857) );
  NOR2_X1 U11525 ( .A1(n12009), .A2(n12008), .ZN(n12774) );
  INV_X1 U11526 ( .A(n20566), .ZN(n11635) );
  NOR2_X1 U11527 ( .A1(n20586), .A2(n18725), .ZN(n11625) );
  NOR2_X1 U11528 ( .A1(n11238), .A2(n14459), .ZN(n11237) );
  INV_X1 U11529 ( .A(n14493), .ZN(n11238) );
  NAND2_X1 U11530 ( .A1(n15432), .A2(n15052), .ZN(n15352) );
  AND2_X1 U11531 ( .A1(n15051), .A2(n15433), .ZN(n15052) );
  AND2_X1 U11532 ( .A1(n15442), .A2(n15450), .ZN(n15433) );
  INV_X1 U11533 ( .A(n19940), .ZN(n11309) );
  NAND2_X1 U11534 ( .A1(n11314), .A2(n11382), .ZN(n11308) );
  INV_X1 U11535 ( .A(n11313), .ZN(n11314) );
  INV_X1 U11536 ( .A(n15158), .ZN(n15127) );
  AND2_X1 U11537 ( .A1(n11237), .A2(n11234), .ZN(n11233) );
  INV_X1 U11538 ( .A(n14714), .ZN(n11234) );
  NAND2_X1 U11539 ( .A1(n11236), .A2(n11235), .ZN(n14680) );
  NAND2_X1 U11540 ( .A1(n11165), .A2(n13132), .ZN(n13172) );
  AND2_X1 U11541 ( .A1(n14070), .A2(n13151), .ZN(n11165) );
  INV_X1 U11542 ( .A(n14144), .ZN(n11215) );
  OR2_X1 U11543 ( .A1(n15511), .A2(n21898), .ZN(n15087) );
  NAND2_X1 U11544 ( .A1(n11200), .A2(n13415), .ZN(n11199) );
  INV_X1 U11545 ( .A(n15452), .ZN(n11200) );
  INV_X1 U11546 ( .A(n15443), .ZN(n11201) );
  INV_X1 U11547 ( .A(n14790), .ZN(n11188) );
  AND2_X1 U11548 ( .A1(n13104), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U11549 ( .A1(n13348), .A2(n13684), .ZN(n13429) );
  INV_X1 U11550 ( .A(n11114), .ZN(n11115) );
  OAI21_X1 U11551 ( .B1(n13442), .B2(n22202), .A(n21195), .ZN(n11114) );
  NAND2_X1 U11552 ( .A1(n11304), .A2(n11306), .ZN(n11302) );
  NAND2_X1 U11553 ( .A1(n13092), .A2(n13759), .ZN(n13107) );
  AND2_X1 U11554 ( .A1(n13078), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U11555 ( .A1(n11117), .A2(n13035), .ZN(n13036) );
  OR2_X1 U11556 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21897), .ZN(
        n13255) );
  NOR3_X1 U11557 ( .A1(n12304), .A2(n11002), .A3(n11211), .ZN(n12327) );
  OR2_X1 U11558 ( .A1(n12303), .A2(n12324), .ZN(n11211) );
  AND2_X1 U11559 ( .A1(n12260), .A2(n11035), .ZN(n12256) );
  INV_X1 U11560 ( .A(n12254), .ZN(n11210) );
  NOR2_X1 U11561 ( .A1(n12235), .A2(n12234), .ZN(n12240) );
  NOR2_X1 U11562 ( .A1(n12226), .A2(n11209), .ZN(n11208) );
  INV_X1 U11563 ( .A(n12218), .ZN(n11209) );
  NAND2_X1 U11564 ( .A1(n12219), .A2(n10986), .ZN(n12233) );
  AND2_X1 U11565 ( .A1(n11044), .A2(n11267), .ZN(n11266) );
  INV_X1 U11566 ( .A(n12756), .ZN(n11267) );
  NOR2_X1 U11567 ( .A1(n12402), .A2(n12420), .ZN(n11886) );
  AND2_X2 U11568 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11981) );
  NOR2_X1 U11569 ( .A1(n14766), .A2(n11292), .ZN(n11291) );
  INV_X1 U11570 ( .A(n14522), .ZN(n11292) );
  INV_X1 U11571 ( .A(n15990), .ZN(n15931) );
  NOR2_X1 U11572 ( .A1(n11155), .A2(n16313), .ZN(n11154) );
  INV_X1 U11573 ( .A(n16312), .ZN(n11155) );
  NAND2_X1 U11574 ( .A1(n12219), .A2(n12218), .ZN(n15210) );
  NOR2_X1 U11575 ( .A1(n18342), .A2(n15212), .ZN(n15189) );
  AND2_X1 U11576 ( .A1(n18317), .A2(n11337), .ZN(n12321) );
  NAND2_X1 U11577 ( .A1(n11126), .A2(n11128), .ZN(n12308) );
  INV_X1 U11578 ( .A(n11129), .ZN(n11128) );
  NAND2_X1 U11579 ( .A1(n12297), .A2(n11127), .ZN(n11126) );
  NOR2_X1 U11580 ( .A1(n11056), .A2(n11228), .ZN(n11227) );
  AND2_X1 U11581 ( .A1(n16350), .A2(n12259), .ZN(n16322) );
  AND2_X1 U11582 ( .A1(n14236), .A2(n14198), .ZN(n11273) );
  OR2_X1 U11583 ( .A1(n18106), .A2(n15212), .ZN(n12231) );
  NAND2_X1 U11584 ( .A1(n11367), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11366) );
  INV_X1 U11585 ( .A(n12790), .ZN(n11367) );
  NAND2_X1 U11586 ( .A1(n11360), .A2(n12113), .ZN(n11351) );
  XNOR2_X1 U11587 ( .A(n12447), .B(n12452), .ZN(n13809) );
  OR2_X1 U11588 ( .A1(n12452), .A2(n12451), .ZN(n12456) );
  NAND2_X1 U11589 ( .A1(n13843), .A2(n13842), .ZN(n13867) );
  OAI21_X1 U11590 ( .B1(n13944), .B2(n14032), .A(n13860), .ZN(n13863) );
  NAND2_X1 U11591 ( .A1(n13863), .A2(n13862), .ZN(n13871) );
  NOR2_X1 U11592 ( .A1(n11853), .A2(n11852), .ZN(n11879) );
  NAND2_X1 U11593 ( .A1(n11961), .A2(n11965), .ZN(n12079) );
  NOR2_X1 U11594 ( .A1(n20740), .A2(n20089), .ZN(n11449) );
  NOR2_X1 U11595 ( .A1(n20761), .A2(n20729), .ZN(n11441) );
  NOR2_X1 U11596 ( .A1(n20446), .A2(n11095), .ZN(n11094) );
  NOR2_X1 U11597 ( .A1(n20096), .A2(n11092), .ZN(n11091) );
  INV_X1 U11598 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11092) );
  OAI21_X1 U11599 ( .B1(n11695), .B2(n20586), .A(n11683), .ZN(n11612) );
  NAND2_X1 U11600 ( .A1(n11245), .A2(n17708), .ZN(n11522) );
  NAND2_X1 U11601 ( .A1(n11612), .A2(n11688), .ZN(n11626) );
  NOR2_X1 U11602 ( .A1(n20558), .A2(n11512), .ZN(n11515) );
  NAND2_X1 U11603 ( .A1(n17863), .A2(n11649), .ZN(n11651) );
  NAND2_X1 U11604 ( .A1(n17892), .A2(n11645), .ZN(n11647) );
  NOR2_X1 U11605 ( .A1(n11609), .A2(n11682), .ZN(n11687) );
  AOI22_X1 U11606 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n21147), .B2(n11406), .ZN(
        n11678) );
  NOR2_X1 U11607 ( .A1(n20597), .A2(n18766), .ZN(n11688) );
  NAND2_X1 U11608 ( .A1(n11611), .A2(n11617), .ZN(n20746) );
  AND2_X1 U11609 ( .A1(n14709), .A2(n14273), .ZN(n14282) );
  OR2_X1 U11610 ( .A1(n13682), .A2(n13681), .ZN(n13824) );
  INV_X1 U11611 ( .A(n15087), .ZN(n15165) );
  INV_X1 U11612 ( .A(n15257), .ZN(n11240) );
  OR2_X1 U11613 ( .A1(n15134), .A2(n15133), .ZN(n15160) );
  NAND2_X1 U11614 ( .A1(n15045), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15048) );
  AND2_X1 U11615 ( .A1(n15432), .A2(n15450), .ZN(n15448) );
  NAND2_X1 U11616 ( .A1(n14421), .A2(n14420), .ZN(n14457) );
  INV_X1 U11617 ( .A(n14423), .ZN(n14420) );
  INV_X1 U11618 ( .A(n13203), .ZN(n13204) );
  INV_X1 U11619 ( .A(n15244), .ZN(n15592) );
  NAND2_X1 U11620 ( .A1(n13226), .A2(n13221), .ZN(n15627) );
  NAND2_X1 U11621 ( .A1(n11313), .A2(n11312), .ZN(n11311) );
  NAND2_X1 U11622 ( .A1(n11315), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11312) );
  NAND2_X1 U11623 ( .A1(n13221), .A2(n11157), .ZN(n11159) );
  NAND2_X1 U11624 ( .A1(n11158), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11157) );
  INV_X1 U11625 ( .A(n13215), .ZN(n11158) );
  OR2_X1 U11626 ( .A1(n13193), .A2(n21262), .ZN(n13194) );
  NAND2_X1 U11627 ( .A1(n11194), .A2(n11192), .ZN(n11191) );
  NOR2_X1 U11628 ( .A1(n19880), .A2(n19886), .ZN(n11192) );
  NAND2_X1 U11629 ( .A1(n11105), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13150) );
  AND2_X1 U11630 ( .A1(n13457), .A2(n13451), .ZN(n21206) );
  OR2_X1 U11631 ( .A1(n15203), .A2(n15202), .ZN(n15209) );
  NAND2_X1 U11632 ( .A1(n15201), .A2(n15200), .ZN(n15203) );
  AND2_X1 U11633 ( .A1(n12327), .A2(n12326), .ZN(n15201) );
  NOR2_X1 U11634 ( .A1(n16155), .A2(n16147), .ZN(n16149) );
  OR2_X1 U11635 ( .A1(n12302), .A2(n12301), .ZN(n12304) );
  AND2_X1 U11636 ( .A1(n12499), .A2(n12498), .ZN(n13833) );
  AOI21_X1 U11637 ( .B1(n13799), .B2(n11336), .A(n11335), .ZN(n11334) );
  INV_X1 U11638 ( .A(n13821), .ZN(n11335) );
  AND2_X1 U11639 ( .A1(n12155), .A2(n12154), .ZN(n12219) );
  AND2_X1 U11640 ( .A1(n16094), .A2(n11266), .ZN(n16065) );
  NOR2_X1 U11641 ( .A1(n14535), .A2(n14534), .ZN(n14582) );
  OAI21_X1 U11642 ( .B1(n16010), .B2(n11281), .A(n11277), .ZN(n11287) );
  INV_X1 U11643 ( .A(n11282), .ZN(n11281) );
  INV_X1 U11644 ( .A(n16053), .ZN(n11278) );
  NAND2_X1 U11645 ( .A1(n11275), .A2(n15913), .ZN(n16093) );
  OR2_X1 U11646 ( .A1(n13875), .A2(n13876), .ZN(n13928) );
  NOR2_X1 U11647 ( .A1(n12125), .A2(n12124), .ZN(n12135) );
  AND2_X1 U11648 ( .A1(n18355), .A2(n11337), .ZN(n16243) );
  OAI21_X1 U11649 ( .B1(n16263), .B2(n15197), .A(n15189), .ZN(n16242) );
  NAND2_X1 U11650 ( .A1(n12618), .A2(n16207), .ZN(n11319) );
  OR2_X1 U11651 ( .A1(n14431), .A2(n14430), .ZN(n14496) );
  NAND2_X1 U11652 ( .A1(n14126), .A2(n14153), .ZN(n14184) );
  NAND2_X1 U11653 ( .A1(n12239), .A2(n12238), .ZN(n16311) );
  NAND2_X1 U11654 ( .A1(n12635), .A2(n11337), .ZN(n11336) );
  OR2_X1 U11655 ( .A1(n13875), .A2(n11261), .ZN(n14105) );
  OR2_X1 U11656 ( .A1(n11263), .A2(n11262), .ZN(n11261) );
  INV_X1 U11657 ( .A(n13907), .ZN(n11262) );
  NOR2_X1 U11658 ( .A1(n13875), .A2(n11263), .ZN(n13929) );
  AND2_X1 U11659 ( .A1(n14545), .A2(n12476), .ZN(n13800) );
  OR2_X1 U11660 ( .A1(n12788), .A2(n12787), .ZN(n12789) );
  AND2_X1 U11661 ( .A1(n12471), .A2(n12470), .ZN(n14206) );
  AND2_X1 U11662 ( .A1(n13848), .A2(n13847), .ZN(n13849) );
  XNOR2_X1 U11663 ( .A(n13867), .B(n13865), .ZN(n13850) );
  NAND2_X1 U11664 ( .A1(n13733), .A2(n13732), .ZN(n13848) );
  OR2_X1 U11665 ( .A1(n12355), .A2(n12352), .ZN(n14335) );
  NAND2_X1 U11666 ( .A1(n19198), .A2(n19142), .ZN(n19193) );
  AND2_X1 U11667 ( .A1(n19219), .A2(n19200), .ZN(n19215) );
  AOI21_X1 U11668 ( .B1(n19036), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n13500), 
        .ZN(n19044) );
  INV_X1 U11669 ( .A(n19219), .ZN(n19594) );
  NOR2_X1 U11670 ( .A1(n20411), .A2(n20482), .ZN(n20412) );
  INV_X1 U11671 ( .A(n11547), .ZN(n17492) );
  NAND2_X1 U11672 ( .A1(n21143), .A2(n20761), .ZN(n11081) );
  NOR2_X1 U11673 ( .A1(n17745), .A2(n20481), .ZN(n17744) );
  NAND2_X1 U11674 ( .A1(n17691), .A2(n17692), .ZN(n17690) );
  NOR2_X1 U11675 ( .A1(n17670), .A2(n17655), .ZN(n17713) );
  INV_X1 U11676 ( .A(n17668), .ZN(n11246) );
  NOR2_X1 U11677 ( .A1(n17622), .A2(n17604), .ZN(n17637) );
  NAND2_X1 U11678 ( .A1(n17540), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17622) );
  NOR2_X1 U11679 ( .A1(n17855), .A2(n20159), .ZN(n17830) );
  INV_X1 U11680 ( .A(n17909), .ZN(n11247) );
  AOI211_X1 U11681 ( .C1(n17481), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n11533), .B(n11532), .ZN(n11534) );
  OAI21_X1 U11682 ( .B1(n20879), .B2(n17534), .A(n20945), .ZN(n20770) );
  NAND2_X1 U11683 ( .A1(n11258), .A2(n11257), .ZN(n17852) );
  NAND2_X1 U11684 ( .A1(n11511), .A2(n11259), .ZN(n11257) );
  NAND2_X1 U11685 ( .A1(n17862), .A2(n11015), .ZN(n11258) );
  INV_X2 U11686 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21898) );
  XNOR2_X1 U11687 ( .A(n13433), .B(n13432), .ZN(n15424) );
  NAND2_X1 U11688 ( .A1(n15344), .A2(n11053), .ZN(n11184) );
  NAND2_X1 U11689 ( .A1(n13236), .A2(n11112), .ZN(n15172) );
  INV_X1 U11690 ( .A(n11113), .ZN(n11112) );
  OR2_X1 U11691 ( .A1(n19967), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21373) );
  AND2_X1 U11692 ( .A1(n13457), .A2(n13327), .ZN(n21393) );
  INV_X1 U11693 ( .A(n21393), .ZN(n21353) );
  AND3_X1 U11694 ( .A1(n16714), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18535) );
  OR2_X1 U11695 ( .A1(n18538), .A2(n13525), .ZN(n17018) );
  AND2_X1 U11696 ( .A1(n17018), .A2(n16713), .ZN(n17021) );
  INV_X1 U11697 ( .A(n17024), .ZN(n17035) );
  XNOR2_X1 U11698 ( .A(n15229), .B(n15228), .ZN(n18403) );
  XNOR2_X1 U11699 ( .A(n16119), .B(n15270), .ZN(n18994) );
  INV_X1 U11700 ( .A(n11318), .ZN(n11317) );
  AOI21_X1 U11701 ( .B1(n18382), .B2(n18466), .A(n16448), .ZN(n16449) );
  OR2_X1 U11702 ( .A1(n16447), .A2(n16446), .ZN(n16448) );
  XNOR2_X1 U11703 ( .A(n16048), .B(n16058), .ZN(n18383) );
  INV_X1 U11704 ( .A(n16357), .ZN(n18249) );
  XNOR2_X1 U11705 ( .A(n16353), .B(n11045), .ZN(n16581) );
  INV_X1 U11706 ( .A(n18494), .ZN(n18481) );
  INV_X1 U11707 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19146) );
  INV_X1 U11708 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19183) );
  NAND2_X1 U11709 ( .A1(n14335), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16694) );
  NAND2_X1 U11710 ( .A1(n20016), .A2(n20521), .ZN(n20088) );
  OAI21_X1 U11711 ( .B1(n20362), .B2(n20482), .A(n11097), .ZN(n20386) );
  AOI21_X1 U11712 ( .B1(n20387), .B2(n11099), .A(n11098), .ZN(n11097) );
  INV_X1 U11713 ( .A(n20363), .ZN(n11099) );
  INV_X1 U11714 ( .A(n20382), .ZN(n11098) );
  AND2_X1 U11715 ( .A1(n11714), .A2(n21105), .ZN(n11119) );
  NAND2_X1 U11716 ( .A1(n11121), .A2(n20998), .ZN(n11120) );
  NAND2_X1 U11717 ( .A1(n11251), .A2(n11253), .ZN(n11122) );
  NAND2_X1 U11718 ( .A1(n20770), .A2(n17596), .ZN(n20938) );
  AND2_X1 U11719 ( .A1(n20939), .A2(n21120), .ZN(n11070) );
  NAND2_X1 U11720 ( .A1(n20767), .A2(n11076), .ZN(n20935) );
  AND2_X1 U11721 ( .A1(n21041), .A2(n20768), .ZN(n11076) );
  NAND2_X1 U11722 ( .A1(n11733), .A2(n20847), .ZN(n21110) );
  INV_X1 U11723 ( .A(n16302), .ZN(n11130) );
  AOI22_X1 U11724 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12031), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12033) );
  OAI21_X1 U11725 ( .B1(n11143), .B2(n11142), .A(n11141), .ZN(n11140) );
  NOR2_X1 U11726 ( .A1(n11678), .A2(n11669), .ZN(n11661) );
  NAND2_X1 U11727 ( .A1(n13219), .A2(n13218), .ZN(n13220) );
  NOR2_X1 U11728 ( .A1(n15673), .A2(n19933), .ZN(n13218) );
  INV_X1 U11729 ( .A(n15670), .ZN(n13219) );
  OR2_X1 U11730 ( .A1(n13183), .A2(n13182), .ZN(n13200) );
  OR2_X1 U11731 ( .A1(n13162), .A2(n13161), .ZN(n13190) );
  INV_X1 U11732 ( .A(n13265), .ZN(n11221) );
  INV_X1 U11733 ( .A(n13021), .ZN(n11306) );
  INV_X1 U11734 ( .A(n13026), .ZN(n11305) );
  AND2_X1 U11735 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12900) );
  AND2_X2 U11736 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14055) );
  AND2_X1 U11737 ( .A1(n11752), .A2(n13958), .ZN(n15891) );
  AND2_X1 U11738 ( .A1(n12440), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13728) );
  NOR2_X1 U11739 ( .A1(n12420), .A2(n18022), .ZN(n11903) );
  INV_X1 U11740 ( .A(n16282), .ZN(n12319) );
  INV_X1 U11741 ( .A(n16265), .ZN(n12320) );
  NOR2_X1 U11742 ( .A1(n11130), .A2(n11135), .ZN(n11127) );
  OAI21_X1 U11743 ( .B1(n11009), .B2(n11130), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U11744 ( .A1(n11394), .A2(n11393), .ZN(n12112) );
  INV_X1 U11745 ( .A(n14524), .ZN(n11870) );
  OR2_X1 U11746 ( .A1(n12027), .A2(n12026), .ZN(n12138) );
  NAND2_X1 U11747 ( .A1(n11148), .A2(n11149), .ZN(n11145) );
  NOR2_X1 U11748 ( .A1(n13749), .A2(n11878), .ZN(n11149) );
  NAND2_X1 U11749 ( .A1(n11084), .A2(n11878), .ZN(n11147) );
  OAI21_X1 U11750 ( .B1(n13740), .B2(n11870), .A(n11860), .ZN(n11363) );
  NOR2_X1 U11751 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  INV_X1 U11752 ( .A(n12149), .ZN(n12151) );
  NAND2_X1 U11753 ( .A1(n13737), .A2(n18036), .ZN(n11143) );
  AND3_X1 U11754 ( .A1(n12384), .A2(n12383), .A3(n12410), .ZN(n12404) );
  NAND2_X1 U11755 ( .A1(n12377), .A2(n11860), .ZN(n12378) );
  NAND2_X1 U11756 ( .A1(n11507), .A2(n11632), .ZN(n11512) );
  INV_X1 U11757 ( .A(n20698), .ZN(n11627) );
  NAND2_X1 U11758 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U11759 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11403) );
  AND2_X1 U11760 ( .A1(n13254), .A2(n13239), .ZN(n13249) );
  AND2_X1 U11761 ( .A1(n12974), .A2(n22104), .ZN(n13680) );
  AOI22_X1 U11762 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12842) );
  INV_X1 U11763 ( .A(n15473), .ZN(n11229) );
  AND2_X1 U11764 ( .A1(n15482), .A2(n15378), .ZN(n11230) );
  INV_X1 U11765 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14662) );
  NOR2_X1 U11766 ( .A1(n15319), .A2(n11183), .ZN(n11182) );
  INV_X1 U11767 ( .A(n15331), .ZN(n11183) );
  OAI21_X1 U11768 ( .B1(n11108), .B2(n11110), .A(n11107), .ZN(n13226) );
  INV_X1 U11769 ( .A(n11310), .ZN(n11108) );
  INV_X1 U11770 ( .A(n13220), .ZN(n11315) );
  INV_X1 U11771 ( .A(n19901), .ZN(n11299) );
  NOR2_X1 U11772 ( .A1(n11299), .A2(n11298), .ZN(n11297) );
  INV_X1 U11773 ( .A(n19894), .ZN(n11298) );
  OR2_X1 U11774 ( .A1(n13142), .A2(n13141), .ZN(n13165) );
  OR2_X1 U11775 ( .A1(n13090), .A2(n13089), .ZN(n13125) );
  OR2_X1 U11776 ( .A1(n13429), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13331) );
  AND2_X1 U11777 ( .A1(n13680), .A2(n12985), .ZN(n13692) );
  NAND2_X1 U11778 ( .A1(n12986), .A2(n13056), .ZN(n12980) );
  OR2_X1 U11779 ( .A1(n13123), .A2(n13122), .ZN(n13145) );
  NOR2_X1 U11780 ( .A1(n12986), .A2(n12965), .ZN(n12974) );
  AOI22_X1 U11781 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12923), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U11782 ( .A1(n12941), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12831) );
  INV_X1 U11783 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21853) );
  NAND2_X1 U11784 ( .A1(n13079), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13279) );
  INV_X1 U11785 ( .A(n13078), .ZN(n13079) );
  INV_X1 U11786 ( .A(n13269), .ZN(n13294) );
  AND2_X1 U11787 ( .A1(n11347), .A2(n16173), .ZN(n11346) );
  AND2_X1 U11788 ( .A1(n12256), .A2(n12251), .ZN(n12279) );
  AND2_X1 U11789 ( .A1(n12260), .A2(n12261), .ZN(n12272) );
  NOR2_X1 U11790 ( .A1(n12175), .A2(n12174), .ZN(n12164) );
  OAI21_X1 U11791 ( .B1(n12386), .B2(n15204), .A(n11203), .ZN(n12174) );
  NAND2_X1 U11792 ( .A1(n15204), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11203) );
  INV_X1 U11793 ( .A(n11280), .ZN(n11279) );
  INV_X1 U11794 ( .A(n15895), .ZN(n16033) );
  CLKBUF_X1 U11795 ( .A(n15897), .Z(n16019) );
  INV_X1 U11796 ( .A(n16071), .ZN(n11284) );
  INV_X1 U11797 ( .A(n11858), .ZN(n13749) );
  NOR2_X1 U11798 ( .A1(n18295), .A2(n11169), .ZN(n11168) );
  INV_X1 U11799 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11169) );
  INV_X1 U11800 ( .A(n16391), .ZN(n16383) );
  NAND2_X1 U11801 ( .A1(n11154), .A2(n16422), .ZN(n11152) );
  NAND2_X1 U11802 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16401), .ZN(
        n16391) );
  NOR2_X1 U11803 ( .A1(n17019), .A2(n16403), .ZN(n16401) );
  NOR2_X1 U11804 ( .A1(n18140), .A2(n11172), .ZN(n11171) );
  INV_X1 U11805 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11172) );
  NOR2_X1 U11806 ( .A1(n18083), .A2(n11177), .ZN(n11176) );
  AND2_X1 U11807 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U11808 ( .A1(n14030), .A2(n10989), .ZN(n11915) );
  NAND2_X1 U11809 ( .A1(n11340), .A2(n16126), .ZN(n11339) );
  INV_X1 U11810 ( .A(n11341), .ZN(n11340) );
  NAND2_X1 U11811 ( .A1(n11986), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14571) );
  NAND2_X1 U11812 ( .A1(n15973), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14569) );
  INV_X1 U11813 ( .A(n16076), .ZN(n11268) );
  NAND2_X1 U11814 ( .A1(n16562), .A2(n11345), .ZN(n16167) );
  AND2_X1 U11815 ( .A1(n11346), .A2(n12653), .ZN(n11345) );
  NOR2_X1 U11816 ( .A1(n11354), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11132) );
  INV_X1 U11817 ( .A(n16525), .ZN(n11354) );
  INV_X1 U11818 ( .A(n18296), .ZN(n12307) );
  AND2_X1 U11819 ( .A1(n16376), .A2(n16375), .ZN(n16320) );
  NOR2_X1 U11820 ( .A1(n16995), .A2(n16668), .ZN(n11371) );
  NAND2_X1 U11821 ( .A1(n11265), .A2(n11264), .ZN(n11263) );
  INV_X1 U11822 ( .A(n13927), .ZN(n11264) );
  INV_X1 U11823 ( .A(n13876), .ZN(n11265) );
  OR2_X1 U11824 ( .A1(n12213), .A2(n12212), .ZN(n12475) );
  AND2_X1 U11825 ( .A1(n11366), .A2(n12795), .ZN(n11365) );
  NAND2_X1 U11826 ( .A1(n11929), .A2(n11928), .ZN(n12665) );
  NAND2_X1 U11827 ( .A1(n12164), .A2(n12163), .ZN(n12165) );
  NAND2_X1 U11828 ( .A1(n11926), .A2(n11925), .ZN(n11934) );
  OAI21_X1 U11829 ( .B1(n12401), .B2(n11865), .A(n12374), .ZN(n12434) );
  NAND2_X1 U11830 ( .A1(n11860), .A2(n12440), .ZN(n11865) );
  INV_X1 U11831 ( .A(n11872), .ZN(n11862) );
  AND2_X1 U11832 ( .A1(n12450), .A2(n12449), .ZN(n13808) );
  OR2_X1 U11833 ( .A1(n12056), .A2(n12055), .ZN(n12463) );
  NAND2_X1 U11834 ( .A1(n12376), .A2(n11882), .ZN(n11896) );
  CLKBUF_X1 U11835 ( .A(n12366), .Z(n12367) );
  NAND2_X1 U11836 ( .A1(n11966), .A2(n11965), .ZN(n12086) );
  NAND3_X1 U11837 ( .A1(n11390), .A2(n11774), .A3(n11773), .ZN(n11775) );
  NAND2_X1 U11838 ( .A1(n11770), .A2(n13958), .ZN(n11776) );
  NOR2_X1 U11839 ( .A1(n17535), .A2(n21071), .ZN(n17597) );
  AND2_X1 U11840 ( .A1(n17561), .A2(n17530), .ZN(n17537) );
  OR2_X1 U11841 ( .A1(n17845), .A2(n20850), .ZN(n11656) );
  INV_X1 U11842 ( .A(n11692), .ZN(n11616) );
  OAI21_X1 U11843 ( .B1(n11623), .B2(n21135), .A(n21165), .ZN(n11621) );
  INV_X1 U11844 ( .A(n20752), .ZN(n20109) );
  OAI21_X1 U11845 ( .B1(n11676), .B2(n11674), .A(n11677), .ZN(n21134) );
  AND2_X1 U11846 ( .A1(n14403), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14442) );
  NAND2_X1 U11847 ( .A1(n13918), .A2(n13917), .ZN(n14087) );
  INV_X1 U11848 ( .A(n13921), .ZN(n13918) );
  INV_X1 U11849 ( .A(n13920), .ZN(n13917) );
  NAND2_X1 U11850 ( .A1(n13069), .A2(n13068), .ZN(n13077) );
  NAND2_X1 U11851 ( .A1(n13070), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13075) );
  AND2_X1 U11852 ( .A1(n14118), .A2(n15293), .ZN(n19780) );
  INV_X1 U11853 ( .A(n13670), .ZN(n13624) );
  NAND2_X1 U11854 ( .A1(n15327), .A2(n11241), .ZN(n15317) );
  AND2_X1 U11855 ( .A1(n15610), .A2(n15161), .ZN(n15112) );
  NAND2_X1 U11856 ( .A1(n14264), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15090) );
  INV_X1 U11857 ( .A(n15069), .ZN(n14264) );
  OR2_X1 U11858 ( .A1(n15090), .A2(n15089), .ZN(n15111) );
  NAND2_X1 U11859 ( .A1(n14263), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15027) );
  OR2_X1 U11860 ( .A1(n15027), .A2(n15026), .ZN(n15069) );
  AND2_X1 U11861 ( .A1(n14262), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15045) );
  AND2_X1 U11862 ( .A1(n15050), .A2(n15049), .ZN(n15450) );
  AND2_X1 U11863 ( .A1(n14979), .A2(n14978), .ZN(n15456) );
  NOR2_X1 U11864 ( .A1(n14944), .A2(n15656), .ZN(n14961) );
  NAND2_X1 U11865 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n14961), .ZN(
        n14977) );
  CLKBUF_X1 U11866 ( .A(n15365), .Z(n15461) );
  AND2_X1 U11867 ( .A1(n14897), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14928) );
  NAND2_X1 U11868 ( .A1(n14928), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14944) );
  NOR2_X1 U11869 ( .A1(n14882), .A2(n15383), .ZN(n14897) );
  NOR2_X1 U11870 ( .A1(n14847), .A2(n14848), .ZN(n14866) );
  NAND2_X1 U11871 ( .A1(n14686), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14847) );
  NOR2_X1 U11872 ( .A1(n14661), .A2(n14662), .ZN(n14686) );
  NOR2_X2 U11873 ( .A1(n14457), .A2(n11231), .ZN(n14704) );
  NAND2_X1 U11874 ( .A1(n11232), .A2(n11031), .ZN(n11231) );
  OR2_X1 U11875 ( .A1(n11235), .A2(n11233), .ZN(n11232) );
  NOR2_X1 U11876 ( .A1(n14475), .A2(n14474), .ZN(n14631) );
  NAND2_X1 U11877 ( .A1(n14631), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14630) );
  NAND2_X1 U11878 ( .A1(n14442), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14475) );
  INV_X1 U11879 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14474) );
  AND2_X1 U11880 ( .A1(n14419), .A2(n14418), .ZN(n14423) );
  NOR2_X1 U11881 ( .A1(n14246), .A2(n14245), .ZN(n14403) );
  INV_X1 U11882 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14245) );
  AOI21_X1 U11883 ( .B1(n14251), .B2(n14656), .A(n14250), .ZN(n14253) );
  INV_X1 U11884 ( .A(n14218), .ZN(n14219) );
  NAND2_X1 U11885 ( .A1(n14219), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14246) );
  NAND2_X1 U11886 ( .A1(n14223), .A2(n14222), .ZN(n14225) );
  INV_X1 U11887 ( .A(n14187), .ZN(n14188) );
  NAND2_X1 U11888 ( .A1(n14188), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14218) );
  NOR2_X1 U11889 ( .A1(n14193), .A2(n14143), .ZN(n11214) );
  NAND2_X1 U11890 ( .A1(n14135), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14187) );
  NAND2_X1 U11891 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14089) );
  NOR2_X1 U11892 ( .A1(n14089), .A2(n14088), .ZN(n14135) );
  INV_X1 U11893 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14088) );
  NOR2_X1 U11894 ( .A1(n15354), .A2(n15345), .ZN(n15344) );
  OR3_X1 U11895 ( .A1(n11201), .A2(n15355), .A3(n11199), .ZN(n11198) );
  NOR3_X1 U11896 ( .A1(n15459), .A2(n11201), .A3(n15452), .ZN(n15445) );
  NOR2_X1 U11897 ( .A1(n15459), .A2(n15452), .ZN(n15451) );
  NAND2_X1 U11898 ( .A1(n15463), .A2(n13401), .ZN(n15464) );
  AND2_X1 U11899 ( .A1(n15477), .A2(n15372), .ZN(n15463) );
  NOR2_X1 U11900 ( .A1(n15486), .A2(n15476), .ZN(n15477) );
  NAND2_X1 U11901 ( .A1(n14791), .A2(n10999), .ZN(n15484) );
  INV_X1 U11902 ( .A(n15385), .ZN(n11186) );
  AND2_X1 U11903 ( .A1(n15692), .A2(n11315), .ZN(n19941) );
  AND2_X1 U11904 ( .A1(n13386), .A2(n13385), .ZN(n15494) );
  NAND2_X1 U11905 ( .A1(n14791), .A2(n11024), .ZN(n15506) );
  NAND2_X1 U11906 ( .A1(n14791), .A2(n14790), .ZN(n15504) );
  NAND2_X1 U11907 ( .A1(n13221), .A2(n13215), .ZN(n15695) );
  NAND2_X1 U11908 ( .A1(n13221), .A2(n13214), .ZN(n19925) );
  OR2_X1 U11909 ( .A1(n14798), .A2(n13369), .ZN(n14799) );
  NAND2_X1 U11910 ( .A1(n11294), .A2(n11295), .ZN(n15175) );
  AOI21_X1 U11911 ( .B1(n15182), .B2(n11296), .A(n11013), .ZN(n11295) );
  INV_X1 U11912 ( .A(n13205), .ZN(n11296) );
  XNOR2_X1 U11913 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15174) );
  OR2_X1 U11914 ( .A1(n14462), .A2(n14461), .ZN(n14798) );
  NAND2_X1 U11915 ( .A1(n14425), .A2(n14424), .ZN(n14462) );
  AND2_X1 U11916 ( .A1(n14257), .A2(n14256), .ZN(n14425) );
  NAND2_X1 U11917 ( .A1(n11103), .A2(n11102), .ZN(n19907) );
  INV_X1 U11918 ( .A(n11104), .ZN(n11103) );
  NAND2_X1 U11919 ( .A1(n19895), .A2(n11297), .ZN(n11102) );
  OAI21_X1 U11920 ( .B1(n13150), .B2(n11299), .A(n13171), .ZN(n11104) );
  AND2_X1 U11921 ( .A1(n13354), .A2(n13353), .ZN(n19880) );
  OR2_X1 U11922 ( .A1(n14097), .A2(n11190), .ZN(n19884) );
  NAND2_X1 U11923 ( .A1(n11194), .A2(n11193), .ZN(n11190) );
  OR2_X1 U11924 ( .A1(n14097), .A2(n11195), .ZN(n19887) );
  NOR2_X1 U11925 ( .A1(n14097), .A2(n14096), .ZN(n14147) );
  AND2_X1 U11926 ( .A1(n13453), .A2(n21367), .ZN(n21333) );
  AND2_X1 U11927 ( .A1(n13339), .A2(n13338), .ZN(n13922) );
  NAND2_X1 U11928 ( .A1(n13341), .A2(n13340), .ZN(n14097) );
  INV_X1 U11929 ( .A(n13922), .ZN(n13340) );
  INV_X1 U11930 ( .A(n11180), .ZN(n13341) );
  INV_X1 U11931 ( .A(n13684), .ZN(n13770) );
  CLKBUF_X1 U11932 ( .A(n13062), .Z(n13792) );
  NAND2_X1 U11933 ( .A1(n13692), .A2(n13674), .ZN(n13436) );
  AND2_X1 U11934 ( .A1(n13322), .A2(n19965), .ZN(n13457) );
  NAND2_X1 U11935 ( .A1(n13423), .A2(n13390), .ZN(n13687) );
  NAND2_X1 U11936 ( .A1(n13093), .A2(n13099), .ZN(n13759) );
  NAND2_X1 U11937 ( .A1(n13108), .A2(n11217), .ZN(n13131) );
  INV_X1 U11938 ( .A(n13107), .ZN(n11217) );
  OR2_X1 U11939 ( .A1(n21802), .A2(n10980), .ZN(n21753) );
  AND2_X1 U11940 ( .A1(n10980), .A2(n14071), .ZN(n21792) );
  OR2_X1 U11941 ( .A1(n14068), .A2(n13672), .ZN(n21819) );
  NOR2_X1 U11942 ( .A1(n12885), .A2(n12884), .ZN(n12896) );
  INV_X1 U11943 ( .A(n12966), .ZN(n22104) );
  AND2_X1 U11944 ( .A1(n14068), .A2(n21707), .ZN(n21791) );
  AND2_X1 U11945 ( .A1(n14068), .A2(n13672), .ZN(n21876) );
  NAND2_X1 U11946 ( .A1(n19952), .A2(n21712), .ZN(n22205) );
  INV_X1 U11947 ( .A(n13279), .ZN(n13305) );
  INV_X1 U11948 ( .A(n13297), .ZN(n13301) );
  AOI21_X1 U11949 ( .B1(n13247), .B2(n13246), .A(n13245), .ZN(n13304) );
  INV_X1 U11950 ( .A(n13321), .ZN(n16762) );
  INV_X1 U11951 ( .A(n13715), .ZN(n18021) );
  INV_X2 U11952 ( .A(n19291), .ZN(n15204) );
  OR2_X1 U11953 ( .A1(n15201), .A2(n12328), .ZN(n18342) );
  NOR2_X1 U11954 ( .A1(n11348), .A2(n16180), .ZN(n11347) );
  INV_X1 U11955 ( .A(n16190), .ZN(n11348) );
  OR2_X1 U11956 ( .A1(n12299), .A2(n12298), .ZN(n12302) );
  NAND2_X1 U11957 ( .A1(n12279), .A2(n12278), .ZN(n12299) );
  NAND2_X1 U11958 ( .A1(n16205), .A2(n16583), .ZN(n16585) );
  NAND2_X1 U11959 ( .A1(n12260), .A2(n10997), .ZN(n12255) );
  AND2_X1 U11960 ( .A1(n16383), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16385) );
  NAND2_X1 U11961 ( .A1(n16383), .A2(n10994), .ZN(n16367) );
  NAND2_X1 U11962 ( .A1(n12260), .A2(n10993), .ZN(n12276) );
  OR2_X1 U11963 ( .A1(n12268), .A2(n12266), .ZN(n12264) );
  NOR2_X2 U11964 ( .A1(n12264), .A2(n12263), .ZN(n12260) );
  NAND2_X1 U11965 ( .A1(n11392), .A2(n12241), .ZN(n12268) );
  AND2_X1 U11966 ( .A1(n10986), .A2(n11043), .ZN(n11207) );
  AND2_X1 U11967 ( .A1(n15204), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12234) );
  AND2_X1 U11968 ( .A1(n12539), .A2(n12538), .ZN(n13884) );
  AND2_X1 U11969 ( .A1(n12219), .A2(n11208), .ZN(n12228) );
  NOR2_X1 U11970 ( .A1(n12165), .A2(n12159), .ZN(n12155) );
  CLKBUF_X1 U11971 ( .A(n18257), .Z(n18385) );
  OR2_X1 U11972 ( .A1(n14014), .A2(n18532), .ZN(n13508) );
  INV_X1 U11973 ( .A(n14105), .ZN(n12691) );
  AND2_X1 U11974 ( .A1(n13935), .A2(n11054), .ZN(n11288) );
  INV_X1 U11975 ( .A(n16052), .ZN(n11286) );
  AOI21_X1 U11976 ( .B1(n16009), .B2(n11284), .A(n11283), .ZN(n11282) );
  INV_X1 U11977 ( .A(n16062), .ZN(n11283) );
  AND2_X1 U11978 ( .A1(n11290), .A2(n14828), .ZN(n11289) );
  INV_X1 U11979 ( .A(n14180), .ZN(n14526) );
  OR2_X1 U11980 ( .A1(n14767), .A2(n14764), .ZN(n14602) );
  AND2_X1 U11981 ( .A1(n10992), .A2(n13836), .ZN(n11331) );
  AND2_X1 U11982 ( .A1(n13871), .A2(n13870), .ZN(n13872) );
  AND2_X1 U11983 ( .A1(n19597), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13715) );
  AND2_X1 U11984 ( .A1(n13714), .A2(n21669), .ZN(n17076) );
  INV_X1 U11985 ( .A(n15271), .ZN(n11225) );
  XNOR2_X1 U11986 ( .A(n11179), .B(n11178), .ZN(n15811) );
  INV_X1 U11987 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U11988 ( .A1(n16221), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U11989 ( .A1(n16255), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16247) );
  AND2_X1 U11990 ( .A1(n16273), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16255) );
  NAND2_X1 U11991 ( .A1(n17030), .A2(n11167), .ZN(n16284) );
  AND2_X1 U11992 ( .A1(n10995), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11167) );
  NOR2_X1 U11993 ( .A1(n16284), .A2(n16272), .ZN(n16273) );
  NAND2_X1 U11994 ( .A1(n17030), .A2(n10995), .ZN(n16295) );
  NAND2_X1 U11995 ( .A1(n17030), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17029) );
  NOR2_X1 U11996 ( .A1(n16344), .A2(n16334), .ZN(n17030) );
  INV_X1 U11997 ( .A(n16318), .ZN(n16394) );
  OR2_X1 U11998 ( .A1(n14496), .A2(n14495), .ZN(n14535) );
  NAND2_X1 U11999 ( .A1(n17020), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17019) );
  AND2_X1 U12000 ( .A1(n16985), .A2(n11170), .ZN(n17020) );
  AND2_X1 U12001 ( .A1(n10987), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U12002 ( .A1(n16311), .A2(n11154), .ZN(n16406) );
  NAND2_X1 U12003 ( .A1(n16985), .A2(n10987), .ZN(n17004) );
  INV_X1 U12004 ( .A(n16433), .ZN(n16985) );
  NAND2_X1 U12005 ( .A1(n16985), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16984) );
  NAND2_X1 U12006 ( .A1(n11175), .A2(n11173), .ZN(n16433) );
  NOR2_X1 U12007 ( .A1(n10985), .A2(n11174), .ZN(n11173) );
  NAND2_X1 U12008 ( .A1(n11175), .A2(n11176), .ZN(n16975) );
  NOR2_X1 U12009 ( .A1(n16966), .A2(n10985), .ZN(n16974) );
  INV_X1 U12010 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18083) );
  NOR2_X1 U12011 ( .A1(n16966), .A2(n18083), .ZN(n14729) );
  NAND2_X1 U12012 ( .A1(n14357), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14395) );
  INV_X1 U12013 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14396) );
  NOR2_X1 U12014 ( .A1(n14395), .A2(n14396), .ZN(n16967) );
  NAND2_X1 U12015 ( .A1(n11206), .A2(n11205), .ZN(n18395) );
  NAND2_X1 U12016 ( .A1(n15211), .A2(n19291), .ZN(n11205) );
  OAI21_X1 U12017 ( .B1(n15209), .B2(P2_EBX_REG_30__SCAN_IN), .A(n15204), .ZN(
        n11206) );
  OR2_X1 U12018 ( .A1(n16492), .A2(n12813), .ZN(n16457) );
  NAND2_X1 U12019 ( .A1(n10967), .A2(n11226), .ZN(n16269) );
  NOR2_X1 U12020 ( .A1(n12321), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16282) );
  NOR2_X1 U12021 ( .A1(n16532), .A2(n11056), .ZN(n16306) );
  INV_X1 U12022 ( .A(n11132), .ZN(n11131) );
  NAND2_X1 U12023 ( .A1(n16311), .A2(n12249), .ZN(n12285) );
  OR2_X1 U12024 ( .A1(n18262), .A2(n15212), .ZN(n16324) );
  NOR2_X1 U12025 ( .A1(n14580), .A2(n11269), .ZN(n14742) );
  INV_X1 U12026 ( .A(n14604), .ZN(n11271) );
  INV_X1 U12027 ( .A(n14803), .ZN(n11270) );
  NAND2_X1 U12028 ( .A1(n16351), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16352) );
  AND2_X1 U12029 ( .A1(n12639), .A2(n12638), .ZN(n14523) );
  INV_X1 U12030 ( .A(n14215), .ZN(n11320) );
  AND2_X1 U12031 ( .A1(n11028), .A2(n14328), .ZN(n11272) );
  NAND2_X1 U12032 ( .A1(n13882), .A2(n13948), .ZN(n14127) );
  AND2_X1 U12033 ( .A1(n12577), .A2(n12576), .ZN(n14128) );
  CLKBUF_X1 U12034 ( .A(n16339), .Z(n16432) );
  INV_X1 U12035 ( .A(n16979), .ZN(n11358) );
  XNOR2_X1 U12036 ( .A(n12807), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16976) );
  AND2_X1 U12037 ( .A1(n12231), .A2(n12230), .ZN(n16979) );
  OR2_X1 U12038 ( .A1(n18094), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14724) );
  NAND2_X1 U12039 ( .A1(n12794), .A2(n11366), .ZN(n12796) );
  NOR2_X1 U12040 ( .A1(n11326), .A2(n14206), .ZN(n11323) );
  INV_X1 U12041 ( .A(n13938), .ZN(n12676) );
  OAI21_X1 U12043 ( .B1(n15269), .B2(n11137), .A(n12446), .ZN(n13747) );
  AOI21_X1 U12044 ( .B1(n18427), .B2(n13837), .A(n13731), .ZN(n13732) );
  INV_X1 U12045 ( .A(n18385), .ZN(n18246) );
  NAND2_X1 U12046 ( .A1(n11961), .A2(n11960), .ZN(n19203) );
  NAND2_X1 U12047 ( .A1(n11962), .A2(n11963), .ZN(n19064) );
  INV_X1 U12048 ( .A(n12086), .ZN(n14344) );
  OR2_X1 U12049 ( .A1(n19035), .A2(n18038), .ZN(n19192) );
  OR2_X1 U12050 ( .A1(n19035), .A2(n19034), .ZN(n19182) );
  NAND3_X1 U12051 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14526), .A3(n19215), 
        .ZN(n19602) );
  NAND3_X1 U12052 ( .A1(n16187), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19215), 
        .ZN(n19600) );
  INV_X1 U12053 ( .A(n19602), .ZN(n19593) );
  INV_X1 U12054 ( .A(n19600), .ZN(n19592) );
  INV_X1 U12055 ( .A(n19354), .ZN(n19596) );
  NAND2_X1 U12056 ( .A1(n19170), .A2(n19085), .ZN(n19051) );
  NAND2_X1 U12057 ( .A1(n19035), .A2(n18038), .ZN(n19143) );
  AND2_X1 U12058 ( .A1(n12371), .A2(n17044), .ZN(n18520) );
  NOR3_X2 U12059 ( .A1(n11626), .A2(n11609), .A3(n11619), .ZN(n11610) );
  INV_X1 U12060 ( .A(n21134), .ZN(n21130) );
  AOI21_X1 U12061 ( .B1(n20411), .B2(n11100), .A(n20482), .ZN(n20434) );
  INV_X1 U12062 ( .A(n20413), .ZN(n11100) );
  NOR2_X1 U12063 ( .A1(n20434), .A2(n20435), .ZN(n20441) );
  NAND2_X1 U12064 ( .A1(n20400), .A2(n11388), .ZN(n20401) );
  NAND2_X1 U12065 ( .A1(n20386), .A2(n20387), .ZN(n20400) );
  OAI21_X1 U12066 ( .B1(n20524), .B2(n20523), .A(n21164), .ZN(n20527) );
  INV_X1 U12067 ( .A(n20527), .ZN(n20596) );
  NOR2_X1 U12068 ( .A1(n20027), .A2(n16705), .ZN(n17973) );
  NAND2_X1 U12069 ( .A1(n20520), .A2(n11610), .ZN(n20028) );
  NAND2_X1 U12070 ( .A1(n21130), .A2(n21649), .ZN(n20029) );
  NAND2_X1 U12071 ( .A1(n17744), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17723) );
  NAND2_X1 U12072 ( .A1(n17713), .A2(n11003), .ZN(n17745) );
  NAND2_X1 U12073 ( .A1(n17713), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17712) );
  INV_X1 U12074 ( .A(n17670), .ZN(n17671) );
  NAND2_X1 U12075 ( .A1(n17637), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17670) );
  NAND2_X1 U12076 ( .A1(n17751), .A2(n10998), .ZN(n17541) );
  NAND2_X1 U12077 ( .A1(n17751), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17528) );
  NAND2_X1 U12078 ( .A1(n17776), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21061) );
  NAND2_X1 U12079 ( .A1(n17571), .A2(n11725), .ZN(n17550) );
  INV_X1 U12080 ( .A(n20280), .ZN(n11725) );
  NOR2_X1 U12081 ( .A1(n20213), .A2(n20231), .ZN(n17571) );
  INV_X1 U12082 ( .A(n20250), .ZN(n17771) );
  NOR4_X1 U12083 ( .A1(n20185), .A2(n20174), .A3(n20201), .A4(n20220), .ZN(
        n17770) );
  NOR2_X1 U12084 ( .A1(n17553), .A2(n20858), .ZN(n17786) );
  NAND2_X1 U12085 ( .A1(n11101), .A2(n11017), .ZN(n17855) );
  INV_X1 U12086 ( .A(n17891), .ZN(n11101) );
  INV_X1 U12087 ( .A(n17918), .ZN(n17875) );
  NAND2_X1 U12088 ( .A1(n17690), .A2(n20798), .ZN(n11700) );
  NOR2_X1 U12089 ( .A1(n20981), .A2(n20980), .ZN(n11252) );
  NAND2_X1 U12090 ( .A1(n20798), .A2(n17793), .ZN(n11253) );
  NOR2_X1 U12091 ( .A1(n17618), .A2(n11523), .ZN(n17667) );
  OR2_X1 U12092 ( .A1(n21061), .A2(n17595), .ZN(n20765) );
  NOR2_X1 U12093 ( .A1(n17618), .A2(n17537), .ZN(n17535) );
  NAND2_X1 U12094 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17764), .ZN(
        n20920) );
  INV_X1 U12095 ( .A(n21061), .ZN(n21018) );
  NOR2_X1 U12096 ( .A1(n17777), .A2(n20918), .ZN(n17776) );
  NOR2_X1 U12097 ( .A1(n20918), .A2(n17765), .ZN(n17764) );
  INV_X1 U12098 ( .A(n16707), .ZN(n20021) );
  INV_X1 U12099 ( .A(n20931), .ZN(n21103) );
  NOR2_X1 U12100 ( .A1(n17840), .A2(n11518), .ZN(n17828) );
  NAND2_X1 U12101 ( .A1(n17856), .A2(n11652), .ZN(n17846) );
  NOR2_X1 U12102 ( .A1(n17846), .A2(n17847), .ZN(n17845) );
  NAND2_X1 U12103 ( .A1(n17882), .A2(n11648), .ZN(n17864) );
  NAND2_X1 U12104 ( .A1(n17864), .A2(n17865), .ZN(n17863) );
  INV_X1 U12105 ( .A(n11509), .ZN(n11508) );
  AND2_X1 U12106 ( .A1(n17862), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17868) );
  OR2_X1 U12107 ( .A1(n17877), .A2(n20819), .ZN(n17882) );
  NAND2_X1 U12108 ( .A1(n20792), .A2(n11644), .ZN(n17893) );
  XNOR2_X1 U12109 ( .A(n11637), .B(n11501), .ZN(n17894) );
  NAND2_X1 U12110 ( .A1(n17893), .A2(n17894), .ZN(n17892) );
  NOR2_X1 U12111 ( .A1(n17890), .A2(n17889), .ZN(n17888) );
  INV_X1 U12112 ( .A(n21132), .ZN(n20798) );
  INV_X1 U12113 ( .A(n20995), .ZN(n21125) );
  NOR2_X1 U12114 ( .A1(n11598), .A2(n11597), .ZN(n11682) );
  AND2_X1 U12115 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20742) );
  INV_X1 U12116 ( .A(n20742), .ZN(n20720) );
  INV_X1 U12117 ( .A(n20746), .ZN(n11123) );
  INV_X1 U12118 ( .A(n21094), .ZN(n21126) );
  INV_X1 U12119 ( .A(n20721), .ZN(n20713) );
  NAND3_X1 U12120 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16697) );
  INV_X1 U12121 ( .A(n20520), .ZN(n20084) );
  NOR2_X2 U12122 ( .A1(n11608), .A2(n11607), .ZN(n18807) );
  NOR2_X1 U12123 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18567), .ZN(n18895) );
  NOR2_X1 U12124 ( .A1(n11557), .A2(n11556), .ZN(n18766) );
  NOR2_X1 U12125 ( .A1(n11577), .A2(n11576), .ZN(n18725) );
  INV_X1 U12126 ( .A(n11609), .ZN(n20585) );
  INV_X1 U12127 ( .A(n18895), .ZN(n18765) );
  AND2_X1 U12128 ( .A1(n15291), .A2(n13342), .ZN(n13517) );
  INV_X1 U12129 ( .A(n21507), .ZN(n21596) );
  AND2_X1 U12130 ( .A1(n14709), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21553) );
  INV_X1 U12131 ( .A(n21605), .ZN(n21592) );
  OR2_X1 U12132 ( .A1(n21588), .A2(n14269), .ZN(n21428) );
  AND2_X1 U12133 ( .A1(n14282), .A2(n14281), .ZN(n21597) );
  AND2_X1 U12134 ( .A1(n13686), .A2(n13685), .ZN(n19892) );
  INV_X1 U12135 ( .A(n19888), .ZN(n15497) );
  INV_X1 U12136 ( .A(n15511), .ZN(n22202) );
  INV_X1 U12137 ( .A(n15304), .ZN(n15517) );
  INV_X1 U12138 ( .A(n15597), .ZN(n15522) );
  INV_X1 U12139 ( .A(n15510), .ZN(n15580) );
  AND2_X1 U12140 ( .A1(n15238), .A2(n21712), .ZN(n15581) );
  OR2_X1 U12141 ( .A1(n15239), .A2(n13828), .ZN(n15585) );
  BUF_X1 U12142 ( .A(n19802), .Z(n19813) );
  BUF_X1 U12143 ( .A(n19797), .Z(n21200) );
  NOR2_X1 U12144 ( .A1(n19780), .A2(n21200), .ZN(n19802) );
  XNOR2_X1 U12145 ( .A(n14267), .B(n14266), .ZN(n15169) );
  OR2_X1 U12146 ( .A1(n15160), .A2(n15260), .ZN(n14267) );
  INV_X1 U12147 ( .A(n15166), .ZN(n11243) );
  AND2_X1 U12148 ( .A1(n14718), .A2(n14717), .ZN(n19930) );
  CLKBUF_X1 U12149 ( .A(n14457), .Z(n14458) );
  NAND2_X1 U12150 ( .A1(n19911), .A2(n13205), .ZN(n15183) );
  INV_X1 U12151 ( .A(n21610), .ZN(n19961) );
  OR2_X1 U12152 ( .A1(n16749), .A2(n21631), .ZN(n21610) );
  NOR2_X1 U12153 ( .A1(n15245), .A2(n15592), .ZN(n15246) );
  NAND2_X1 U12154 ( .A1(n13227), .A2(n13228), .ZN(n15619) );
  OAI21_X1 U12155 ( .B1(n11310), .B2(n11055), .A(n11109), .ZN(n15646) );
  AND2_X1 U12156 ( .A1(n15698), .A2(n11159), .ZN(n15682) );
  NAND2_X1 U12157 ( .A1(n19899), .A2(n19901), .ZN(n19900) );
  INV_X1 U12158 ( .A(n11106), .ZN(n14229) );
  INV_X1 U12159 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21864) );
  CLKBUF_X1 U12160 ( .A(n21872), .Z(n21908) );
  INV_X1 U12161 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16765) );
  AND2_X1 U12162 ( .A1(n21623), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15801) );
  NOR2_X1 U12163 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15797) );
  OR2_X1 U12164 ( .A1(n21753), .A2(n21841), .ZN(n22230) );
  INV_X1 U12165 ( .A(n22230), .ZN(n22239) );
  INV_X1 U12166 ( .A(n22178), .ZN(n22275) );
  AND2_X1 U12167 ( .A1(n21877), .A2(n21873), .ZN(n22304) );
  AND2_X1 U12168 ( .A1(n21877), .A2(n21791), .ZN(n22314) );
  NOR2_X1 U12169 ( .A1(n13508), .A2(n13499), .ZN(n15824) );
  NAND2_X1 U12170 ( .A1(n18358), .A2(n18385), .ZN(n18360) );
  NAND2_X1 U12171 ( .A1(n18360), .A2(n18359), .ZN(n18369) );
  OR2_X1 U12172 ( .A1(n15265), .A2(n12661), .ZN(n18353) );
  NAND2_X1 U12173 ( .A1(n18332), .A2(n18385), .ZN(n18334) );
  NAND2_X1 U12174 ( .A1(n18334), .A2(n18333), .ZN(n18348) );
  NAND2_X1 U12175 ( .A1(n12313), .A2(n12312), .ZN(n12318) );
  NAND2_X1 U12176 ( .A1(n11166), .A2(n18303), .ZN(n18310) );
  NAND2_X1 U12177 ( .A1(n11333), .A2(n11334), .ZN(n13832) );
  INV_X1 U12178 ( .A(n18378), .ZN(n18396) );
  OR2_X1 U12179 ( .A1(n19591), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n18283) );
  INV_X1 U12180 ( .A(n18193), .ZN(n18260) );
  INV_X1 U12181 ( .A(n18340), .ZN(n18402) );
  NOR2_X1 U12182 ( .A1(n18516), .A2(n18246), .ZN(n18393) );
  OR2_X1 U12183 ( .A1(n16058), .A2(n16057), .ZN(n16233) );
  OR2_X1 U12184 ( .A1(n16055), .A2(n16066), .ZN(n16248) );
  OR2_X1 U12185 ( .A1(n12555), .A2(n12554), .ZN(n14195) );
  OR2_X1 U12186 ( .A1(n12516), .A2(n12515), .ZN(n14156) );
  NAND2_X1 U12187 ( .A1(n13936), .A2(n13935), .ZN(n13934) );
  AND2_X1 U12188 ( .A1(n13736), .A2(n18535), .ZN(n16112) );
  XNOR2_X1 U12189 ( .A(n11285), .B(n16045), .ZN(n16124) );
  NAND2_X1 U12190 ( .A1(n11287), .A2(n11286), .ZN(n11285) );
  INV_X1 U12191 ( .A(n19474), .ZN(n18995) );
  AND2_X1 U12192 ( .A1(n19468), .A2(n19467), .ZN(n19287) );
  NAND2_X1 U12193 ( .A1(n13746), .A2(n18535), .ZN(n19465) );
  CLKBUF_X1 U12195 ( .A(n17096), .Z(n17108) );
  NOR2_X1 U12196 ( .A1(n17076), .A2(n17108), .ZN(n17095) );
  INV_X1 U12197 ( .A(n18999), .ZN(n19589) );
  NAND2_X1 U12198 ( .A1(n18403), .A2(n17021), .ZN(n15233) );
  NOR2_X1 U12199 ( .A1(n16608), .A2(n11374), .ZN(n11372) );
  AND2_X1 U12200 ( .A1(n16399), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16400) );
  INV_X1 U12201 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15836) );
  INV_X1 U12202 ( .A(n17014), .ZN(n17032) );
  INV_X1 U12203 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13531) );
  INV_X1 U12204 ( .A(n17018), .ZN(n17031) );
  INV_X1 U12205 ( .A(n16233), .ZN(n18368) );
  INV_X1 U12206 ( .A(n16248), .ZN(n18357) );
  NAND2_X1 U12207 ( .A1(n16242), .A2(n15190), .ZN(n11082) );
  NOR3_X1 U12208 ( .A1(n14184), .A2(n11321), .A3(n14183), .ZN(n16208) );
  NAND2_X1 U12209 ( .A1(n16399), .A2(n11373), .ZN(n16598) );
  NAND2_X1 U12210 ( .A1(n16311), .A2(n16312), .ZN(n17001) );
  NAND2_X1 U12211 ( .A1(n16432), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16994) );
  OAI21_X1 U12212 ( .B1(n13800), .B2(n13799), .A(n11336), .ZN(n13822) );
  CLKBUF_X1 U12213 ( .A(n14608), .Z(n14609) );
  NAND2_X1 U12214 ( .A1(n11370), .A2(n11368), .ZN(n14540) );
  NAND2_X1 U12215 ( .A1(n12793), .A2(n12790), .ZN(n11370) );
  OR2_X1 U12216 ( .A1(n12793), .A2(n12790), .ZN(n11368) );
  INV_X1 U12217 ( .A(n18450), .ZN(n18501) );
  INV_X1 U12218 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19164) );
  INV_X1 U12219 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19179) );
  INV_X1 U12220 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19160) );
  OR2_X1 U12221 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  INV_X1 U12222 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19159) );
  NAND2_X1 U12223 ( .A1(n19170), .A2(n19142), .ZN(n19083) );
  AND2_X1 U12224 ( .A1(n11330), .A2(n11327), .ZN(n14164) );
  INV_X1 U12225 ( .A(n12460), .ZN(n11327) );
  INV_X1 U12226 ( .A(n19198), .ZN(n19170) );
  INV_X1 U12227 ( .A(n19034), .ZN(n18038) );
  NAND2_X1 U12228 ( .A1(n13848), .A2(n13734), .ZN(n19035) );
  OR2_X1 U12229 ( .A1(n13733), .A2(n13732), .ZN(n13734) );
  XNOR2_X1 U12230 ( .A(n13943), .B(n13942), .ZN(n19198) );
  OAI21_X1 U12231 ( .B1(n19270), .B2(n19220), .A(n19219), .ZN(n19716) );
  OR2_X1 U12232 ( .A1(n19193), .A2(n19143), .ZN(n19686) );
  OR2_X1 U12233 ( .A1(n19131), .A2(n19182), .ZN(n19670) );
  NOR2_X1 U12234 ( .A1(n19131), .A2(n19167), .ZN(n19657) );
  NAND2_X1 U12235 ( .A1(n19101), .A2(n19100), .ZN(n19651) );
  OAI22_X1 U12236 ( .A1(n19077), .A2(n19074), .B1(n19215), .B2(n19073), .ZN(
        n19636) );
  AOI21_X1 U12237 ( .B1(n19357), .B2(n19219), .A(n19045), .ZN(n19611) );
  INV_X1 U12238 ( .A(n19709), .ZN(n19702) );
  AND2_X1 U12239 ( .A1(n16011), .A2(n19596), .ZN(n19573) );
  INV_X1 U12240 ( .A(n19231), .ZN(n19604) );
  INV_X1 U12241 ( .A(n19211), .ZN(n19197) );
  INV_X1 U12242 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16714) );
  NOR2_X1 U12243 ( .A1(n21129), .A2(n20027), .ZN(n20016) );
  INV_X1 U12244 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20082) );
  INV_X1 U12245 ( .A(n20494), .ZN(n11090) );
  OR2_X1 U12246 ( .A1(n20483), .A2(n20482), .ZN(n20493) );
  INV_X1 U12247 ( .A(n20491), .ZN(n11087) );
  NOR2_X1 U12248 ( .A1(n20459), .A2(n20482), .ZN(n20460) );
  NOR2_X1 U12249 ( .A1(n20412), .A2(n20413), .ZN(n20433) );
  NAND2_X1 U12250 ( .A1(n20380), .A2(n20387), .ZN(n20381) );
  NAND2_X1 U12251 ( .A1(n20362), .A2(n20363), .ZN(n20380) );
  INV_X1 U12252 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20220) );
  INV_X1 U12253 ( .A(n20409), .ZN(n20500) );
  INV_X1 U12254 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21139) );
  INV_X1 U12255 ( .A(n20515), .ZN(n20490) );
  INV_X1 U12256 ( .A(n20514), .ZN(n20431) );
  NOR2_X2 U12257 ( .A1(n21176), .A2(n20431), .ZN(n20409) );
  NAND4_X1 U12258 ( .A1(n21105), .A2(n20090), .A3(n21173), .A4(n21185), .ZN(
        n20514) );
  INV_X1 U12259 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17353) );
  AOI211_X1 U12260 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11564), .B(n11563), .ZN(n11565) );
  NOR2_X1 U12261 ( .A1(n20661), .A2(n20626), .ZN(n20632) );
  NOR2_X1 U12262 ( .A1(n20625), .A2(n20667), .ZN(n20662) );
  NAND2_X1 U12263 ( .A1(n20662), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20661) );
  NOR2_X1 U12264 ( .A1(n20607), .A2(n20612), .ZN(n20606) );
  NOR3_X1 U12265 ( .A1(n20625), .A2(n20675), .A3(n20584), .ZN(n20616) );
  INV_X1 U12266 ( .A(n20631), .ZN(n20674) );
  INV_X1 U12267 ( .A(n20672), .ZN(n20673) );
  NOR2_X1 U12268 ( .A1(n20536), .A2(n20542), .ZN(n20540) );
  NOR2_X1 U12269 ( .A1(n11412), .A2(n11411), .ZN(n20558) );
  NOR2_X1 U12270 ( .A1(n20526), .A2(n20557), .ZN(n20560) );
  NOR2_X1 U12271 ( .A1(n20525), .A2(n20565), .ZN(n20568) );
  NOR2_X1 U12272 ( .A1(n11432), .A2(n11431), .ZN(n20579) );
  NAND2_X1 U12273 ( .A1(n20625), .A2(n20596), .ZN(n20700) );
  INV_X1 U12274 ( .A(n20691), .ZN(n20704) );
  INV_X1 U12275 ( .A(n20573), .ZN(n20705) );
  CLKBUF_X1 U12276 ( .A(n21177), .Z(n17990) );
  NOR3_X1 U12278 ( .A1(n21188), .A2(n20029), .A3(n20028), .ZN(n20071) );
  INV_X1 U12280 ( .A(n20765), .ZN(n17651) );
  INV_X1 U12281 ( .A(n17637), .ZN(n17600) );
  AOI21_X1 U12282 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17636), .A(
        n18894), .ZN(n17680) );
  NOR2_X1 U12283 ( .A1(n17550), .A2(n17564), .ZN(n17751) );
  NAND3_X1 U12284 ( .A1(n21644), .A2(n17918), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17755) );
  INV_X1 U12285 ( .A(n17821), .ZN(n17806) );
  INV_X1 U12286 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20201) );
  INV_X1 U12287 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20159) );
  AND3_X1 U12288 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20128) );
  INV_X1 U12289 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17884) );
  NAND2_X1 U12290 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17891) );
  OR2_X1 U12291 ( .A1(n18765), .A2(n18609), .ZN(n18893) );
  INV_X1 U12292 ( .A(n11249), .ZN(n17902) );
  INV_X1 U12293 ( .A(n11248), .ZN(n17901) );
  AND2_X1 U12294 ( .A1(n11248), .A2(n11249), .ZN(n17900) );
  INV_X1 U12295 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20096) );
  INV_X1 U12296 ( .A(n17922), .ZN(n17912) );
  NAND2_X1 U12297 ( .A1(n17755), .A2(n17754), .ZN(n17911) );
  XNOR2_X1 U12298 ( .A(n11723), .B(n20716), .ZN(n11737) );
  NAND2_X1 U12299 ( .A1(n11722), .A2(n11007), .ZN(n11723) );
  OR3_X2 U12300 ( .A1(n17738), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U12301 ( .A1(n21016), .A2(n20978), .ZN(n20981) );
  NOR2_X1 U12302 ( .A1(n11721), .A2(n11701), .ZN(n17699) );
  NOR2_X1 U12303 ( .A1(n20938), .A2(n20942), .ZN(n21016) );
  INV_X1 U12304 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21153) );
  NAND2_X1 U12305 ( .A1(n20742), .A2(n21143), .ZN(n20729) );
  BUF_X1 U12306 ( .A(n18564), .Z(n18890) );
  OAI21_X1 U12307 ( .B1(n15172), .B2(n21353), .A(n11160), .ZN(P1_U3000) );
  INV_X1 U12308 ( .A(n11161), .ZN(n11160) );
  OAI21_X1 U12309 ( .B1(n15424), .B2(n21399), .A(n13473), .ZN(n11161) );
  NAND2_X1 U12310 ( .A1(n16226), .A2(n16225), .ZN(n16227) );
  OAI21_X1 U12311 ( .B1(n16581), .B2(n17014), .A(n11019), .ZN(P2_U2995) );
  NAND2_X1 U12312 ( .A1(n18994), .A2(n18466), .ZN(n11316) );
  NAND2_X1 U12313 ( .A1(n16450), .A2(n16449), .ZN(n16451) );
  NAND2_X1 U12314 ( .A1(n11088), .A2(n11086), .ZN(P3_U2641) );
  NAND2_X1 U12315 ( .A1(n11089), .A2(n20488), .ZN(n11088) );
  NOR4_X1 U12316 ( .A1(n11008), .A2(n20507), .A3(n20487), .A4(n11087), .ZN(
        n11086) );
  XNOR2_X1 U12317 ( .A(n20493), .B(n11090), .ZN(n11089) );
  NOR2_X1 U12318 ( .A1(n11716), .A2(n11006), .ZN(n11717) );
  NAND2_X1 U12319 ( .A1(n11120), .A2(n11119), .ZN(n11718) );
  AOI21_X1 U12320 ( .B1(n11072), .B2(n11071), .A(n11070), .ZN(n20941) );
  AOI21_X1 U12321 ( .B1(n20938), .B2(n20942), .A(n20997), .ZN(n11071) );
  NOR2_X1 U12322 ( .A1(n20712), .A2(n20755), .ZN(n11461) );
  CLKBUF_X3 U12323 ( .A(n11461), .Z(n17457) );
  INV_X1 U12324 ( .A(n11930), .ZN(n12703) );
  OR3_X1 U12325 ( .A1(n14184), .A2(n14183), .A3(n11320), .ZN(n10984) );
  AND2_X1 U12326 ( .A1(n15492), .A2(n11025), .ZN(n15364) );
  NAND2_X1 U12327 ( .A1(n12914), .A2(n12913), .ZN(n12984) );
  NAND2_X1 U12328 ( .A1(n11236), .A2(n11237), .ZN(n14678) );
  NAND2_X1 U12329 ( .A1(n15492), .A2(n11230), .ZN(n15472) );
  NAND2_X1 U12330 ( .A1(n11176), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10985) );
  AND2_X1 U12331 ( .A1(n11208), .A2(n12227), .ZN(n10986) );
  AND2_X1 U12332 ( .A1(n11171), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10987) );
  NAND2_X1 U12333 ( .A1(n14521), .A2(n14522), .ZN(n14767) );
  AND2_X1 U12334 ( .A1(n11356), .A2(n11030), .ZN(n16988) );
  AND2_X1 U12335 ( .A1(n15182), .A2(n19912), .ZN(n10988) );
  AND2_X1 U12336 ( .A1(n11136), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10989) );
  NOR2_X1 U12337 ( .A1(n15197), .A2(n15189), .ZN(n10990) );
  AND2_X1 U12338 ( .A1(n16562), .A2(n11347), .ZN(n10991) );
  AND2_X1 U12339 ( .A1(n11334), .A2(n11332), .ZN(n10992) );
  OAI21_X1 U12340 ( .B1(n13294), .B2(n13144), .A(n13143), .ZN(n13151) );
  NAND2_X1 U12341 ( .A1(n11330), .A2(n11328), .ZN(n14165) );
  AND2_X1 U12342 ( .A1(n12270), .A2(n12261), .ZN(n10993) );
  AND2_X1 U12343 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U12344 ( .A1(n12691), .A2(n12690), .ZN(n14107) );
  AND2_X1 U12345 ( .A1(n11168), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10995) );
  AND2_X1 U12346 ( .A1(n11024), .A2(n11187), .ZN(n10996) );
  AND2_X1 U12347 ( .A1(n10993), .A2(n11042), .ZN(n10997) );
  AND2_X1 U12348 ( .A1(n11091), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10998) );
  AND2_X1 U12349 ( .A1(n10996), .A2(n11186), .ZN(n10999) );
  AND2_X1 U12350 ( .A1(n14195), .A2(n11389), .ZN(n11000) );
  AND2_X1 U12351 ( .A1(n10994), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11001) );
  OR2_X1 U12352 ( .A1(n12316), .A2(n11212), .ZN(n11002) );
  AND2_X1 U12353 ( .A1(n11094), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11003) );
  AND2_X2 U12354 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U12355 ( .A1(n11351), .A2(n12799), .ZN(n12790) );
  AND2_X2 U12356 ( .A1(n16018), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12003) );
  NAND2_X1 U12357 ( .A1(n11226), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16305) );
  NAND2_X1 U12358 ( .A1(n16562), .A2(n16190), .ZN(n16179) );
  NAND2_X1 U12359 ( .A1(n12311), .A2(n12310), .ZN(n16264) );
  BUF_X1 U12360 ( .A(n12743), .Z(n12752) );
  NAND2_X1 U12361 ( .A1(n16094), .A2(n16088), .ZN(n16075) );
  AOI21_X1 U12362 ( .B1(n13807), .B2(n12456), .A(n12455), .ZN(n12460) );
  OR2_X1 U12363 ( .A1(n16010), .A2(n16009), .ZN(n11004) );
  AND4_X1 U12364 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n11005) );
  INV_X1 U12365 ( .A(n11255), .ZN(n11701) );
  NOR3_X1 U12366 ( .A1(n11715), .A2(n21110), .A3(n17692), .ZN(n11006) );
  OR3_X1 U12367 ( .A1(n17737), .A2(n21007), .A3(n21008), .ZN(n11007) );
  NOR2_X1 U12368 ( .A1(n20492), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11008) );
  AOI21_X1 U12369 ( .B1(n14141), .B2(n14656), .A(n14140), .ZN(n14143) );
  NAND2_X1 U12370 ( .A1(n12297), .A2(n11134), .ZN(n11133) );
  NAND2_X1 U12371 ( .A1(n13226), .A2(n15647), .ZN(n15599) );
  INV_X1 U12372 ( .A(n11360), .ZN(n12115) );
  AND2_X1 U12373 ( .A1(n11356), .A2(n11358), .ZN(n16430) );
  NAND2_X1 U12374 ( .A1(n12297), .A2(n12296), .ZN(n16524) );
  NAND2_X1 U12375 ( .A1(n11133), .A2(n11131), .ZN(n16300) );
  NAND2_X1 U12376 ( .A1(n11300), .A2(n13228), .ZN(n15612) );
  NOR2_X1 U12377 ( .A1(n16301), .A2(n11132), .ZN(n11009) );
  AND2_X1 U12378 ( .A1(n13864), .A2(n13871), .ZN(n13942) );
  AND2_X1 U12379 ( .A1(n16055), .A2(n16056), .ZN(n16058) );
  INV_X1 U12380 ( .A(n11636), .ZN(n20570) );
  NAND2_X1 U12381 ( .A1(n16395), .A2(n16394), .ZN(n16374) );
  OAI22_X1 U12382 ( .A1(n15612), .A2(n13229), .B1(n13212), .B2(n15724), .ZN(
        n15589) );
  INV_X1 U12383 ( .A(n12402), .ZN(n11146) );
  AND2_X1 U12384 ( .A1(n12416), .A2(n11856), .ZN(n11918) );
  AND3_X1 U12385 ( .A1(n11317), .A2(n15278), .A3(n11316), .ZN(n11010) );
  AND2_X1 U12386 ( .A1(n12320), .A2(n12319), .ZN(n11011) );
  INV_X1 U12387 ( .A(n12239), .ZN(n16423) );
  OR2_X1 U12388 ( .A1(n20698), .A2(n11497), .ZN(n11012) );
  AND2_X1 U12389 ( .A1(n13211), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11013) );
  OR2_X1 U12390 ( .A1(n16525), .A2(n11355), .ZN(n11014) );
  AND2_X1 U12391 ( .A1(n11259), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U12392 ( .A1(n13130), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11016) );
  INV_X2 U12393 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13958) );
  AND2_X1 U12394 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11017) );
  AND3_X1 U12395 ( .A1(n14524), .A2(n11858), .A3(n11078), .ZN(n11018) );
  NAND2_X1 U12396 ( .A1(n11085), .A2(n16302), .ZN(n16291) );
  INV_X1 U12397 ( .A(n20387), .ZN(n20482) );
  AND2_X1 U12398 ( .A1(n16362), .A2(n16361), .ZN(n11019) );
  INV_X1 U12399 ( .A(n11110), .ZN(n11109) );
  OAI21_X1 U12400 ( .B1(n11307), .B2(n11055), .A(n13221), .ZN(n11110) );
  NOR2_X1 U12401 ( .A1(n16155), .A2(n11339), .ZN(n11338) );
  NAND3_X1 U12402 ( .A1(n13985), .A2(n11752), .A3(n11352), .ZN(n11783) );
  BUF_X1 U12403 ( .A(n15896), .Z(n16018) );
  AND2_X1 U12404 ( .A1(n11145), .A2(n11147), .ZN(n11020) );
  INV_X1 U12405 ( .A(n11135), .ZN(n11134) );
  NAND2_X1 U12406 ( .A1(n12296), .A2(n11014), .ZN(n11135) );
  INV_X1 U12407 ( .A(n11143), .ZN(n11965) );
  OR3_X1 U12408 ( .A1(n12790), .A2(n12800), .A3(n14548), .ZN(n11021) );
  AND3_X1 U12409 ( .A1(n12311), .A2(n12310), .A3(n11011), .ZN(n16263) );
  INV_X2 U12410 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21143) );
  NAND2_X1 U12411 ( .A1(n11303), .A2(n11301), .ZN(n13093) );
  AND2_X1 U12412 ( .A1(n12223), .A2(n11080), .ZN(n11022) );
  AOI22_X1 U12413 ( .A1(n15811), .A2(n18022), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n15216), .ZN(n18257) );
  INV_X1 U12414 ( .A(n16115), .ZN(n16082) );
  AND2_X1 U12415 ( .A1(n13308), .A2(n14272), .ZN(n13325) );
  INV_X1 U12416 ( .A(n11860), .ZN(n12353) );
  NAND2_X1 U12417 ( .A1(n14239), .A2(n11000), .ZN(n14435) );
  INV_X1 U12418 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U12419 ( .A1(n14239), .A2(n14195), .ZN(n14301) );
  AND2_X1 U12420 ( .A1(n16985), .A2(n11171), .ZN(n11023) );
  NOR2_X1 U12421 ( .A1(n15503), .A2(n11188), .ZN(n11024) );
  NOR3_X1 U12422 ( .A1(n14184), .A2(n11319), .A3(n11321), .ZN(n16205) );
  AND2_X1 U12423 ( .A1(n11214), .A2(n11215), .ZN(n14224) );
  NAND2_X1 U12424 ( .A1(n14224), .A2(n14225), .ZN(n14252) );
  AND2_X1 U12425 ( .A1(n11229), .A2(n11230), .ZN(n11025) );
  INV_X1 U12426 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11111) );
  AND2_X1 U12427 ( .A1(n15864), .A2(n16108), .ZN(n16098) );
  AND2_X1 U12428 ( .A1(n17751), .A2(n11091), .ZN(n11026) );
  AND2_X1 U12429 ( .A1(n17708), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11027) );
  AND2_X1 U12430 ( .A1(n14237), .A2(n11273), .ZN(n14196) );
  AND2_X1 U12431 ( .A1(n14498), .A2(n14500), .ZN(n14521) );
  NOR2_X1 U12432 ( .A1(n14457), .A2(n14459), .ZN(n14492) );
  NAND2_X1 U12433 ( .A1(n16967), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16966) );
  INV_X1 U12434 ( .A(n16966), .ZN(n11175) );
  AND2_X1 U12435 ( .A1(n11273), .A2(n14300), .ZN(n11028) );
  OR2_X1 U12436 ( .A1(n14580), .A2(n14604), .ZN(n11029) );
  NAND2_X1 U12437 ( .A1(n19913), .A2(n19912), .ZN(n19911) );
  AND2_X1 U12438 ( .A1(n11358), .A2(n16429), .ZN(n11030) );
  NAND2_X1 U12439 ( .A1(n15183), .A2(n15182), .ZN(n15181) );
  NAND2_X1 U12440 ( .A1(n19893), .A2(n13150), .ZN(n19899) );
  AND2_X1 U12441 ( .A1(n14679), .A2(n14715), .ZN(n11031) );
  NOR3_X1 U12442 ( .A1(n14580), .A2(n14604), .A3(n14803), .ZN(n14743) );
  NOR2_X1 U12443 ( .A1(n15459), .A2(n11198), .ZN(n11202) );
  INV_X1 U12444 ( .A(n19886), .ZN(n11193) );
  INV_X1 U12445 ( .A(n11197), .ZN(n15437) );
  NOR3_X1 U12446 ( .A1(n15459), .A2(n11199), .A3(n11201), .ZN(n11197) );
  AND2_X1 U12447 ( .A1(n14521), .A2(n11289), .ZN(n15864) );
  NAND2_X1 U12448 ( .A1(n14521), .A2(n11290), .ZN(n14827) );
  INV_X1 U12449 ( .A(n14457), .ZN(n11236) );
  AND2_X1 U12450 ( .A1(n14524), .A2(n12441), .ZN(n12635) );
  AND2_X1 U12451 ( .A1(n14521), .A2(n11291), .ZN(n14786) );
  INV_X1 U12452 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18107) );
  OR2_X1 U12453 ( .A1(n11804), .A2(n13749), .ZN(n11032) );
  OAI21_X1 U12454 ( .B1(n13294), .B2(n13164), .A(n13163), .ZN(n13173) );
  NAND2_X1 U12455 ( .A1(n13232), .A2(n13706), .ZN(n11033) );
  AND2_X1 U12456 ( .A1(n15492), .A2(n15378), .ZN(n15379) );
  NAND2_X1 U12457 ( .A1(n16562), .A2(n11346), .ZN(n16164) );
  AND2_X1 U12458 ( .A1(n11241), .A2(n11240), .ZN(n11034) );
  AND2_X1 U12459 ( .A1(n10997), .A2(n11210), .ZN(n11035) );
  OR2_X1 U12460 ( .A1(n12077), .A2(n12076), .ZN(n12466) );
  AND2_X1 U12461 ( .A1(n11025), .A2(n11385), .ZN(n11036) );
  AND2_X1 U12462 ( .A1(n11288), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11037) );
  AND2_X1 U12463 ( .A1(n13173), .A2(n13151), .ZN(n11038) );
  INV_X1 U12464 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U12465 ( .A1(n13873), .A2(n13872), .ZN(n13936) );
  NAND2_X1 U12466 ( .A1(n13800), .A2(n11336), .ZN(n11333) );
  AND2_X1 U12467 ( .A1(n13936), .A2(n11288), .ZN(n14108) );
  AND2_X1 U12468 ( .A1(n11323), .A2(n11330), .ZN(n14207) );
  AND2_X1 U12469 ( .A1(n11877), .A2(n11876), .ZN(n13967) );
  AND2_X1 U12470 ( .A1(n17030), .A2(n11168), .ZN(n11039) );
  NOR2_X1 U12471 ( .A1(n13883), .A2(n13884), .ZN(n13882) );
  AND2_X1 U12472 ( .A1(n17713), .A2(n11094), .ZN(n11040) );
  AND2_X1 U12473 ( .A1(n11333), .A2(n10992), .ZN(n13831) );
  AND2_X1 U12474 ( .A1(n14237), .A2(n14236), .ZN(n14197) );
  AND2_X1 U12475 ( .A1(n14237), .A2(n11028), .ZN(n14298) );
  NOR2_X1 U12476 ( .A1(n14184), .A2(n14183), .ZN(n14185) );
  AND2_X1 U12477 ( .A1(n16383), .A2(n11001), .ZN(n11041) );
  NAND2_X1 U12478 ( .A1(n15204), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11042) );
  NAND2_X1 U12479 ( .A1(n15204), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11043) );
  NOR2_X1 U12480 ( .A1(n16247), .A2(n16235), .ZN(n16221) );
  AND2_X1 U12481 ( .A1(n16088), .A2(n11268), .ZN(n11044) );
  AND2_X1 U12482 ( .A1(n16350), .A2(n16349), .ZN(n11045) );
  NOR2_X1 U12483 ( .A1(n17541), .A2(n20355), .ZN(n17540) );
  AND2_X1 U12484 ( .A1(n11266), .A2(n16064), .ZN(n11046) );
  NOR2_X1 U12485 ( .A1(n17868), .A2(n11511), .ZN(n11047) );
  AND2_X1 U12486 ( .A1(n14434), .A2(n14437), .ZN(n11048) );
  INV_X1 U12487 ( .A(n11328), .ZN(n11326) );
  NOR2_X1 U12488 ( .A1(n12460), .A2(n11329), .ZN(n11328) );
  NAND2_X1 U12489 ( .A1(n14791), .A2(n10996), .ZN(n11189) );
  AND2_X1 U12490 ( .A1(n13936), .A2(n11037), .ZN(n11049) );
  INV_X1 U12491 ( .A(n20997), .ZN(n21093) );
  NOR2_X1 U12492 ( .A1(n17692), .A2(n17708), .ZN(n11050) );
  AND2_X1 U12493 ( .A1(n11000), .A2(n11048), .ZN(n11051) );
  AND2_X1 U12494 ( .A1(n11001), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11052) );
  INV_X1 U12495 ( .A(n15237), .ZN(n21712) );
  NAND2_X1 U12496 ( .A1(n11247), .A2(n11012), .ZN(n11249) );
  NAND2_X1 U12497 ( .A1(n11515), .A2(n11733), .ZN(n17708) );
  INV_X1 U12498 ( .A(n13838), .ZN(n11138) );
  INV_X1 U12499 ( .A(n12312), .ZN(n11212) );
  INV_X1 U12500 ( .A(n14633), .ZN(n11239) );
  INV_X1 U12501 ( .A(n12660), .ZN(n11344) );
  AND2_X1 U12502 ( .A1(n11182), .A2(n15249), .ZN(n11053) );
  AND2_X1 U12503 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U12504 ( .A1(n15780), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11055) );
  OR2_X1 U12505 ( .A1(n16515), .A2(n11355), .ZN(n11056) );
  INV_X1 U12506 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11228) );
  INV_X1 U12507 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11177) );
  INV_X1 U12508 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11174) );
  INV_X1 U12509 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11095) );
  INV_X1 U12510 ( .A(n11374), .ZN(n11373) );
  NAND2_X1 U12511 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11374) );
  INV_X1 U12512 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11142) );
  INV_X2 U12513 ( .A(n22319), .ZN(n11057) );
  AOI211_X1 U12514 ( .C1(n16211), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        n16123) );
  OAI22_X2 U12515 ( .A1(n21961), .A2(n22207), .B1(n21960), .B2(n22205), .ZN(
        n21997) );
  INV_X1 U12516 ( .A(n22140), .ZN(n11058) );
  INV_X1 U12517 ( .A(n11058), .ZN(n11059) );
  OAI22_X2 U12518 ( .A1(n21914), .A2(n22207), .B1(n21913), .B2(n22205), .ZN(
        n21950) );
  INV_X1 U12519 ( .A(n21955), .ZN(n11060) );
  INV_X1 U12520 ( .A(n11060), .ZN(n11061) );
  INV_X1 U12521 ( .A(n22097), .ZN(n11062) );
  INV_X1 U12522 ( .A(n11062), .ZN(n11063) );
  INV_X1 U12523 ( .A(n22194), .ZN(n11064) );
  INV_X1 U12524 ( .A(n11064), .ZN(n11065) );
  INV_X1 U12525 ( .A(n22303), .ZN(n11066) );
  INV_X1 U12526 ( .A(n11066), .ZN(n11067) );
  INV_X1 U12527 ( .A(n21889), .ZN(n11068) );
  INV_X1 U12528 ( .A(n11068), .ZN(n11069) );
  NOR2_X1 U12529 ( .A1(n21177), .A2(n17973), .ZN(n17982) );
  OAI22_X2 U12530 ( .A1(n22011), .A2(n22207), .B1(n22010), .B2(n22205), .ZN(
        n22050) );
  NOR3_X2 U12531 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21896), .ZN(n22249) );
  INV_X2 U12532 ( .A(n18001), .ZN(n18008) );
  NOR2_X2 U12533 ( .A1(n19354), .A2(n11077), .ZN(n19396) );
  NAND3_X1 U12534 ( .A1(n11075), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11074), .ZN(n11073) );
  CLKBUF_X1 U12535 ( .A(n11078), .Z(n11077) );
  AND3_X1 U12536 ( .A1(n11862), .A2(n11078), .A3(n11861), .ZN(n11863) );
  NAND2_X1 U12537 ( .A1(n12420), .A2(n11077), .ZN(n12412) );
  NAND2_X1 U12538 ( .A1(n12380), .A2(n11077), .ZN(n12381) );
  MUX2_X1 U12539 ( .A(n12380), .B(n11854), .S(n12354), .Z(n11804) );
  NAND2_X1 U12540 ( .A1(n12224), .A2(n12223), .ZN(n14727) );
  NAND2_X1 U12541 ( .A1(n11079), .A2(n14724), .ZN(n16978) );
  NAND2_X1 U12542 ( .A1(n12224), .A2(n11022), .ZN(n11079) );
  INV_X1 U12543 ( .A(n14725), .ZN(n11080) );
  XNOR2_X1 U12544 ( .A(n11638), .B(n20570), .ZN(n11637) );
  NAND2_X1 U12545 ( .A1(n20794), .A2(n20793), .ZN(n20792) );
  INV_X2 U12546 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11406) );
  INV_X4 U12547 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20712) );
  INV_X1 U12548 ( .A(n11656), .ZN(n11653) );
  NAND2_X1 U12549 ( .A1(n11934), .A2(n11933), .ZN(n11083) );
  XNOR2_X2 U12550 ( .A(n12664), .B(n12662), .ZN(n13944) );
  NAND3_X1 U12551 ( .A1(n12414), .A2(n12758), .A3(n11084), .ZN(n13744) );
  INV_X1 U12553 ( .A(n16291), .ZN(n12309) );
  NAND2_X1 U12554 ( .A1(n11133), .A2(n11009), .ZN(n11085) );
  NAND2_X1 U12555 ( .A1(n14353), .A2(n15212), .ZN(n12167) );
  OR2_X2 U12556 ( .A1(n11496), .A2(n11495), .ZN(n20703) );
  INV_X1 U12557 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11093) );
  INV_X1 U12558 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11096) );
  XNOR2_X2 U12559 ( .A(n11105), .B(n21248), .ZN(n19895) );
  NAND2_X2 U12560 ( .A1(n11106), .A2(n11016), .ZN(n11105) );
  OR2_X2 U12561 ( .A1(n14228), .A2(n14230), .ZN(n11106) );
  NOR2_X2 U12562 ( .A1(n16954), .A2(n13105), .ZN(n13129) );
  NOR2_X2 U12563 ( .A1(n16953), .A2(n16955), .ZN(n16954) );
  AND2_X4 U12564 ( .A1(n12830), .A2(n12826), .ZN(n12946) );
  OAI21_X2 U12565 ( .B1(n15588), .B2(n13237), .A(n11033), .ZN(n11113) );
  NOR2_X2 U12566 ( .A1(n15589), .A2(n15590), .ZN(n15588) );
  NAND3_X1 U12567 ( .A1(n12981), .A2(n11381), .A3(n12991), .ZN(n12982) );
  INV_X2 U12568 ( .A(n12978), .ZN(n21915) );
  NAND2_X1 U12569 ( .A1(n11116), .A2(n13053), .ZN(n13092) );
  NAND3_X1 U12570 ( .A1(n21730), .A2(n13069), .A3(n21614), .ZN(n11116) );
  NAND2_X1 U12571 ( .A1(n21730), .A2(n13069), .ZN(n21805) );
  NAND3_X1 U12572 ( .A1(n13070), .A2(n13034), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11117) );
  NAND2_X2 U12573 ( .A1(n13028), .A2(n13065), .ZN(n13070) );
  NAND3_X1 U12574 ( .A1(n11250), .A2(n11122), .A3(n21093), .ZN(n11121) );
  NAND2_X2 U12575 ( .A1(n20747), .A2(n11123), .ZN(n20721) );
  INV_X2 U12576 ( .A(n20748), .ZN(n20747) );
  OR2_X2 U12577 ( .A1(n20738), .A2(n20751), .ZN(n20748) );
  NOR2_X2 U12578 ( .A1(n20586), .A2(n20585), .ZN(n20710) );
  NAND3_X1 U12579 ( .A1(n11586), .A2(n11587), .A3(n11125), .ZN(n11124) );
  NAND2_X1 U12580 ( .A1(n20798), .A2(n20554), .ZN(n20993) );
  AND2_X2 U12581 ( .A1(n21129), .A2(n11622), .ZN(n20931) );
  NOR2_X2 U12582 ( .A1(n14840), .A2(n11621), .ZN(n21129) );
  NAND2_X2 U12583 ( .A1(n14030), .A2(n11136), .ZN(n12707) );
  AND2_X2 U12584 ( .A1(n11359), .A2(n11357), .ZN(n12239) );
  NOR2_X2 U12585 ( .A1(n13944), .A2(n11138), .ZN(n11966) );
  NAND3_X1 U12586 ( .A1(n11139), .A2(n12061), .A3(n12466), .ZN(n11360) );
  INV_X1 U12587 ( .A(n12161), .ZN(n11139) );
  AND2_X1 U12588 ( .A1(n11964), .A2(n11965), .ZN(n19152) );
  AND2_X1 U12589 ( .A1(n11964), .A2(n11140), .ZN(n11958) );
  NAND2_X1 U12590 ( .A1(n11918), .A2(n11144), .ZN(n11150) );
  NAND3_X1 U12591 ( .A1(n11145), .A2(n11146), .A3(n11147), .ZN(n11144) );
  INV_X1 U12592 ( .A(n11804), .ZN(n11148) );
  NAND2_X1 U12593 ( .A1(n11150), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11866) );
  OAI21_X1 U12594 ( .B1(n12239), .B2(n11153), .A(n11151), .ZN(n16317) );
  INV_X1 U12595 ( .A(n11154), .ZN(n11153) );
  NAND2_X1 U12596 ( .A1(n13036), .A2(n21749), .ZN(n13069) );
  NAND2_X1 U12597 ( .A1(n13032), .A2(n13031), .ZN(n11156) );
  NAND3_X1 U12598 ( .A1(n15698), .A2(n13216), .A3(n11159), .ZN(n15670) );
  OAI21_X2 U12599 ( .B1(n15599), .B2(n15601), .A(n13212), .ZN(n13228) );
  INV_X1 U12600 ( .A(n11382), .ZN(n11164) );
  NAND3_X1 U12601 ( .A1(n13132), .A2(n14070), .A3(n11038), .ZN(n13189) );
  NAND2_X1 U12602 ( .A1(n13132), .A2(n14070), .ZN(n13152) );
  OAI211_X1 U12603 ( .C1(n11166), .C2(n18303), .A(n18310), .B(n18386), .ZN(
        n18304) );
  NAND2_X1 U12604 ( .A1(n18301), .A2(n18385), .ZN(n11166) );
  NAND2_X1 U12605 ( .A1(n16383), .A2(n11052), .ZN(n16344) );
  NAND2_X1 U12606 ( .A1(n11180), .A2(n13922), .ZN(n13923) );
  NAND2_X1 U12607 ( .A1(n13771), .A2(n13334), .ZN(n11180) );
  NAND2_X1 U12608 ( .A1(n15344), .A2(n11182), .ZN(n11185) );
  NAND2_X1 U12609 ( .A1(n11185), .A2(n13390), .ZN(n11181) );
  NAND2_X1 U12610 ( .A1(n15344), .A2(n15331), .ZN(n15333) );
  NAND2_X1 U12611 ( .A1(n11184), .A2(n11181), .ZN(n13433) );
  INV_X1 U12612 ( .A(n11185), .ZN(n15318) );
  INV_X1 U12613 ( .A(n11189), .ZN(n15495) );
  INV_X1 U12614 ( .A(n11202), .ZN(n15354) );
  NAND2_X1 U12615 ( .A1(n12219), .A2(n11207), .ZN(n12235) );
  NOR2_X1 U12616 ( .A1(n12304), .A2(n12303), .ZN(n12313) );
  OR3_X1 U12617 ( .A1(n12304), .A2(n11002), .A3(n12303), .ZN(n12325) );
  AND2_X2 U12618 ( .A1(n11213), .A2(n13698), .ZN(n13044) );
  AND2_X2 U12619 ( .A1(n12827), .A2(n11213), .ZN(n14411) );
  AND2_X2 U12620 ( .A1(n12820), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11213) );
  NAND2_X1 U12621 ( .A1(n11215), .A2(n14142), .ZN(n14192) );
  AOI21_X1 U12622 ( .B1(n14191), .B2(n14656), .A(n14190), .ZN(n14193) );
  NAND3_X1 U12623 ( .A1(n12162), .A2(n12785), .A3(n14352), .ZN(n12783) );
  NAND2_X1 U12624 ( .A1(n21802), .A2(n14656), .ZN(n14095) );
  NAND2_X1 U12625 ( .A1(n21804), .A2(n21614), .ZN(n11216) );
  NAND3_X1 U12626 ( .A1(n13323), .A2(n11219), .A3(n13436), .ZN(n11218) );
  OAI21_X1 U12627 ( .B1(n16246), .B2(n11223), .A(n11222), .ZN(n15279) );
  OR2_X1 U12628 ( .A1(n11224), .A2(n15216), .ZN(n11223) );
  NAND2_X1 U12629 ( .A1(n11225), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11224) );
  OAI21_X1 U12630 ( .B1(n15279), .B2(n18494), .A(n11378), .ZN(n11318) );
  INV_X1 U12631 ( .A(n16532), .ZN(n11226) );
  NAND2_X1 U12632 ( .A1(n15492), .A2(n11036), .ZN(n15365) );
  AND2_X1 U12633 ( .A1(n11237), .A2(n14633), .ZN(n11235) );
  NAND2_X1 U12634 ( .A1(n15327), .A2(n11034), .ZN(n11244) );
  INV_X1 U12635 ( .A(n11244), .ZN(n15256) );
  NOR2_X2 U12636 ( .A1(n17826), .A2(n11027), .ZN(n17794) );
  NAND2_X1 U12637 ( .A1(n17691), .A2(n11251), .ZN(n11250) );
  AOI21_X1 U12638 ( .B1(n11050), .B2(n20798), .A(n11252), .ZN(n11251) );
  NAND2_X1 U12639 ( .A1(n11526), .A2(n20980), .ZN(n11715) );
  INV_X1 U12640 ( .A(n11526), .ZN(n11254) );
  INV_X1 U12641 ( .A(n11715), .ZN(n11721) );
  NAND3_X1 U12642 ( .A1(n11255), .A2(n11715), .A3(n17793), .ZN(n17698) );
  XNOR2_X1 U12643 ( .A(n11510), .B(n11508), .ZN(n17862) );
  INV_X1 U12644 ( .A(n17853), .ZN(n11259) );
  AND2_X4 U12645 ( .A1(n11260), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15897) );
  NOR2_X1 U12646 ( .A1(n13970), .A2(n11260), .ZN(n13971) );
  NAND2_X1 U12647 ( .A1(n16094), .A2(n11044), .ZN(n16078) );
  NAND3_X1 U12648 ( .A1(n11271), .A2(n14744), .A3(n11270), .ZN(n11269) );
  NAND2_X1 U12649 ( .A1(n14237), .A2(n11272), .ZN(n14431) );
  INV_X1 U12650 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11274) );
  AND2_X4 U12651 ( .A1(n11975), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11987) );
  NAND2_X1 U12652 ( .A1(n16098), .A2(n16099), .ZN(n11275) );
  NAND2_X1 U12653 ( .A1(n16010), .A2(n16009), .ZN(n16069) );
  NAND2_X1 U12654 ( .A1(n11276), .A2(n11282), .ZN(n16051) );
  NAND2_X1 U12655 ( .A1(n16010), .A2(n11280), .ZN(n11276) );
  AOI21_X1 U12656 ( .B1(n11279), .B2(n11282), .A(n11278), .ZN(n11277) );
  OR2_X1 U12657 ( .A1(n16009), .A2(n11284), .ZN(n11280) );
  NAND2_X1 U12658 ( .A1(n11293), .A2(n12972), .ZN(n12976) );
  NAND3_X1 U12659 ( .A1(n12972), .A2(n11293), .A3(n12978), .ZN(n12992) );
  AND2_X1 U12660 ( .A1(n13318), .A2(n11293), .ZN(n13438) );
  NAND2_X1 U12661 ( .A1(n19913), .A2(n10988), .ZN(n11294) );
  NAND2_X1 U12662 ( .A1(n19895), .A2(n19894), .ZN(n19893) );
  NAND2_X1 U12663 ( .A1(n13227), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11300) );
  NAND2_X1 U12664 ( .A1(n13673), .A2(n11304), .ZN(n11303) );
  INV_X1 U12665 ( .A(n15692), .ZN(n15681) );
  NAND3_X1 U12666 ( .A1(n11328), .A2(n11324), .A3(n11330), .ZN(n14545) );
  NAND2_X1 U12667 ( .A1(n11333), .A2(n11331), .ZN(n13883) );
  NOR2_X1 U12668 ( .A1(n16155), .A2(n11341), .ZN(n16134) );
  INV_X1 U12669 ( .A(n11338), .ZN(n16125) );
  NOR3_X1 U12670 ( .A1(n16155), .A2(n16147), .A3(n11344), .ZN(n15265) );
  INV_X1 U12671 ( .A(n16133), .ZN(n11343) );
  NAND3_X1 U12672 ( .A1(n11351), .A2(n12799), .A3(n15212), .ZN(n12158) );
  NAND4_X1 U12673 ( .A1(n12311), .A2(n11011), .A3(n15192), .A4(n12310), .ZN(
        n11353) );
  NAND2_X1 U12674 ( .A1(n11353), .A2(n15193), .ZN(n15196) );
  INV_X1 U12675 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U12676 ( .A1(n16978), .A2(n12232), .ZN(n11359) );
  CLKBUF_X1 U12677 ( .A(n11359), .Z(n11356) );
  NAND2_X1 U12678 ( .A1(n11361), .A2(n12379), .ZN(n12416) );
  NAND2_X1 U12679 ( .A1(n11364), .A2(n11362), .ZN(n11361) );
  NAND2_X1 U12680 ( .A1(n11363), .A2(n11852), .ZN(n11362) );
  INV_X1 U12681 ( .A(n11853), .ZN(n11364) );
  NAND2_X1 U12682 ( .A1(n12794), .A2(n11365), .ZN(n11369) );
  NAND2_X1 U12683 ( .A1(n14608), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U12684 ( .A1(n16339), .A2(n11371), .ZN(n16416) );
  NAND2_X2 U12685 ( .A1(n16399), .A2(n11372), .ZN(n16380) );
  OAI21_X2 U12686 ( .B1(n13077), .B2(n13076), .A(n13661), .ZN(n21850) );
  AND2_X1 U12687 ( .A1(n11908), .A2(n11907), .ZN(n11909) );
  INV_X1 U12688 ( .A(n11885), .ZN(n14030) );
  NAND2_X1 U12689 ( .A1(n12354), .A2(n11858), .ZN(n11868) );
  OAI211_X1 U12690 ( .C1(n12707), .C2(n14356), .A(n11932), .B(n11931), .ZN(
        n12666) );
  OAI211_X1 U12691 ( .C1(n12707), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        n11890) );
  NAND2_X1 U12692 ( .A1(n11879), .A2(n12379), .ZN(n12376) );
  NAND2_X1 U12693 ( .A1(n12158), .A2(n18069), .ZN(n12182) );
  AOI22_X1 U12694 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U12695 ( .A1(n12783), .A2(n12782), .ZN(n12787) );
  NAND2_X1 U12696 ( .A1(n13838), .A2(n13837), .ZN(n13843) );
  AND2_X1 U12697 ( .A1(n15967), .A2(n15990), .ZN(n11375) );
  OR2_X1 U12698 ( .A1(n16091), .A2(n15952), .ZN(n11376) );
  NOR2_X1 U12699 ( .A1(n13557), .A2(n13556), .ZN(n13669) );
  INV_X1 U12700 ( .A(n11450), .ZN(n11547) );
  NOR2_X1 U12701 ( .A1(n15277), .A2(n15276), .ZN(n11378) );
  INV_X1 U12702 ( .A(n15364), .ZN(n15475) );
  NOR2_X1 U12703 ( .A1(n14196), .A2(n14199), .ZN(n11379) );
  AND3_X1 U12704 ( .A1(n11493), .A2(n11492), .A3(n11491), .ZN(n11380) );
  INV_X1 U12705 ( .A(n17636), .ZN(n17754) );
  NOR2_X1 U12706 ( .A1(n17917), .A2(n17875), .ZN(n17636) );
  INV_X1 U12707 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14020) );
  OR2_X1 U12708 ( .A1(n12495), .A2(n12494), .ZN(n14109) );
  AND3_X1 U12709 ( .A1(n12976), .A2(n13695), .A3(n12975), .ZN(n11381) );
  OR2_X1 U12710 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11382) );
  INV_X1 U12711 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11497) );
  OR2_X1 U12712 ( .A1(n11745), .A2(n17785), .ZN(n11383) );
  INV_X2 U12713 ( .A(n17517), .ZN(n17513) );
  OAI21_X1 U12714 ( .B1(n13210), .B2(n13209), .A(n13221), .ZN(n13211) );
  BUF_X4 U12715 ( .A(n11441), .Z(n17475) );
  OR2_X1 U12716 ( .A1(n15874), .A2(n12018), .ZN(n11384) );
  INV_X1 U12717 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13106) );
  AND2_X1 U12718 ( .A1(n14946), .A2(n14945), .ZN(n11385) );
  NAND2_X1 U12719 ( .A1(n15204), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11386) );
  INV_X1 U12720 ( .A(n15968), .ZN(n16011) );
  INV_X1 U12721 ( .A(n14081), .ZN(n12461) );
  INV_X1 U12722 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11501) );
  AND2_X1 U12723 ( .A1(n13212), .A2(n15723), .ZN(n11387) );
  OR2_X1 U12724 ( .A1(n20482), .A2(n20399), .ZN(n11388) );
  OR2_X1 U12725 ( .A1(n12573), .A2(n12572), .ZN(n11389) );
  AND3_X1 U12726 ( .A1(n11772), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11771), .ZN(n11390) );
  INV_X1 U12727 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21614) );
  AND2_X1 U12728 ( .A1(n16216), .A2(n16230), .ZN(n11391) );
  AND2_X1 U12729 ( .A1(n12240), .A2(n11386), .ZN(n11392) );
  AND4_X1 U12730 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n11393) );
  NAND2_X1 U12731 ( .A1(n11962), .A2(n11957), .ZN(n12085) );
  AND4_X1 U12732 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n11394) );
  AND2_X2 U12733 ( .A1(n14055), .A2(n13698), .ZN(n12928) );
  NAND2_X1 U12734 ( .A1(n13026), .A2(n13025), .ZN(n11395) );
  AND4_X1 U12735 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n11396) );
  AND3_X1 U12736 ( .A1(n13450), .A2(n12992), .A3(n12991), .ZN(n11397) );
  NAND2_X1 U12737 ( .A1(n12986), .A2(n12978), .ZN(n13342) );
  AND2_X1 U12738 ( .A1(n12968), .A2(n15511), .ZN(n11398) );
  OR2_X1 U12739 ( .A1(n12085), .A2(n11941), .ZN(n11942) );
  NAND2_X1 U12740 ( .A1(n13020), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U12741 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11841) );
  OR2_X1 U12742 ( .A1(n13252), .A2(n13268), .ZN(n13254) );
  INV_X1 U12743 ( .A(n15273), .ZN(n15274) );
  INV_X1 U12744 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15190) );
  INV_X1 U12745 ( .A(n11838), .ZN(n11843) );
  XNOR2_X1 U12746 ( .A(n11872), .B(n11861), .ZN(n12380) );
  INV_X1 U12747 ( .A(n13188), .ZN(n13186) );
  AND2_X1 U12748 ( .A1(n13185), .A2(n13184), .ZN(n13188) );
  OR2_X1 U12749 ( .A1(n13052), .A2(n13051), .ZN(n13094) );
  AOI22_X1 U12750 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11759) );
  NOR2_X1 U12751 ( .A1(n11857), .A2(n11858), .ZN(n11803) );
  OR2_X1 U12752 ( .A1(n12015), .A2(n12624), .ZN(n12127) );
  INV_X1 U12753 ( .A(n15048), .ZN(n14263) );
  OR2_X1 U12754 ( .A1(n21623), .A2(n21915), .ZN(n13647) );
  AND2_X1 U12755 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12885) );
  AND2_X1 U12756 ( .A1(n19146), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12337) );
  INV_X1 U12757 ( .A(n16422), .ZN(n12238) );
  XNOR2_X1 U12758 ( .A(n12182), .B(n14548), .ZN(n14541) );
  AND2_X1 U12759 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11505), .ZN(
        n11506) );
  OR2_X1 U12760 ( .A1(n15595), .A2(n14136), .ZN(n15136) );
  INV_X1 U12761 ( .A(n14977), .ZN(n14262) );
  NAND2_X1 U12762 ( .A1(n14646), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14661) );
  NAND2_X1 U12763 ( .A1(n14217), .A2(n14656), .ZN(n14223) );
  NAND2_X1 U12764 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13213) );
  NAND2_X1 U12765 ( .A1(n13070), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13113) );
  AOI21_X1 U12766 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19159), .A(
        n12152), .ZN(n12332) );
  OR2_X1 U12767 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  AND2_X1 U12768 ( .A1(n15969), .A2(n11375), .ZN(n15970) );
  INV_X1 U12769 ( .A(n12806), .ZN(n12808) );
  INV_X1 U12770 ( .A(n19203), .ZN(n12078) );
  NAND2_X1 U12771 ( .A1(n17771), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20280) );
  INV_X1 U12772 ( .A(n11613), .ZN(n11611) );
  AOI21_X1 U12773 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21147), .A(
        n11661), .ZN(n11667) );
  AND2_X1 U12774 ( .A1(n21898), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15164) );
  NAND2_X1 U12775 ( .A1(n15793), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15158) );
  INV_X1 U12776 ( .A(n15502), .ZN(n14865) );
  INV_X1 U12777 ( .A(n14136), .ZN(n15161) );
  NAND2_X1 U12778 ( .A1(n15612), .A2(n15242), .ZN(n15243) );
  AND2_X1 U12779 ( .A1(n15627), .A2(n15600), .ZN(n13227) );
  NAND2_X1 U12780 ( .A1(n15669), .A2(n15671), .ZN(n19940) );
  NAND2_X1 U12781 ( .A1(n13113), .A2(n13112), .ZN(n21764) );
  INV_X1 U12782 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21827) );
  INV_X1 U12783 ( .A(n21863), .ZN(n21895) );
  INV_X1 U12784 ( .A(n16101), .ZN(n12742) );
  INV_X1 U12785 ( .A(n14106), .ZN(n12690) );
  OR2_X1 U12786 ( .A1(n12109), .A2(n12108), .ZN(n12472) );
  AND2_X1 U12787 ( .A1(n16407), .A2(n12291), .ZN(n16316) );
  NOR2_X1 U12788 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  INV_X1 U12789 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15216) );
  AND3_X1 U12790 ( .A1(n11860), .A2(n19410), .A3(n11858), .ZN(n11864) );
  OR2_X1 U12791 ( .A1(n12406), .A2(n12405), .ZN(n13957) );
  OR2_X2 U12792 ( .A1(n11896), .A2(n12433), .ZN(n13987) );
  INV_X1 U12793 ( .A(n19109), .ZN(n19104) );
  INV_X1 U12794 ( .A(n19064), .ZN(n19061) );
  NOR2_X1 U12795 ( .A1(n20712), .A2(n16697), .ZN(n11450) );
  NOR2_X1 U12796 ( .A1(n11624), .A2(n20528), .ZN(n11686) );
  INV_X1 U12797 ( .A(n20558), .ZN(n11630) );
  NOR2_X1 U12798 ( .A1(n21072), .A2(n20784), .ZN(n20810) );
  OR2_X1 U12799 ( .A1(n11668), .A2(n11675), .ZN(n11676) );
  AND2_X1 U12800 ( .A1(n13263), .A2(n13262), .ZN(n15288) );
  INV_X1 U12801 ( .A(n21597), .ZN(n21580) );
  AND2_X1 U12802 ( .A1(n15169), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U12803 ( .A1(n14282), .A2(n14280), .ZN(n21544) );
  OR2_X1 U12804 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  OR2_X1 U12805 ( .A1(n15030), .A2(n15029), .ZN(n15434) );
  NAND2_X1 U12806 ( .A1(n14866), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14882) );
  INV_X1 U12807 ( .A(n14630), .ZN(n14646) );
  XOR2_X1 U12808 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n15673) );
  AND2_X1 U12809 ( .A1(n21333), .A2(n21256), .ZN(n21389) );
  NAND2_X1 U12810 ( .A1(n13457), .A2(n15282), .ZN(n21256) );
  OR2_X1 U12811 ( .A1(n21753), .A2(n21822), .ZN(n22221) );
  OR2_X1 U12812 ( .A1(n21842), .A2(n21819), .ZN(n22178) );
  AOI21_X1 U12813 ( .B1(n21196), .B2(n21615), .A(n15801), .ZN(n21715) );
  INV_X1 U12814 ( .A(n21903), .ZN(n21869) );
  OR3_X1 U12815 ( .A1(n21859), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n21715), 
        .ZN(n22203) );
  INV_X1 U12816 ( .A(n18380), .ZN(n18394) );
  NAND2_X1 U12817 ( .A1(n18396), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18340) );
  NAND2_X1 U12818 ( .A1(n13850), .A2(n13849), .ZN(n13869) );
  INV_X1 U12819 ( .A(n15952), .ZN(n15949) );
  NAND2_X1 U12820 ( .A1(n13495), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n14180)
         );
  NAND2_X1 U12821 ( .A1(n18403), .A2(n18500), .ZN(n15278) );
  OR2_X1 U12822 ( .A1(n12322), .A2(n16497), .ZN(n16280) );
  AND2_X1 U12823 ( .A1(n18270), .A2(n12294), .ZN(n16329) );
  INV_X1 U12824 ( .A(n13957), .ZN(n14005) );
  INV_X1 U12825 ( .A(n19664), .ZN(n19557) );
  NAND2_X1 U12826 ( .A1(n13869), .A2(n13851), .ZN(n19142) );
  OR2_X1 U12827 ( .A1(n19051), .A2(n19167), .ZN(n19608) );
  NOR2_X1 U12828 ( .A1(n20746), .A2(n18807), .ZN(n11689) );
  NOR2_X1 U12829 ( .A1(n11626), .A2(n20724), .ZN(n17133) );
  INV_X1 U12830 ( .A(n20920), .ZN(n21017) );
  INV_X1 U12831 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20231) );
  AND2_X1 U12832 ( .A1(n17708), .A2(n17828), .ZN(n17553) );
  AND2_X1 U12833 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  NAND2_X1 U12834 ( .A1(n20021), .A2(n17133), .ZN(n21094) );
  INV_X1 U12835 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21147) );
  AND2_X1 U12836 ( .A1(n13307), .A2(n13306), .ZN(n21623) );
  INV_X1 U12837 ( .A(n21529), .ZN(n21519) );
  AND2_X1 U12838 ( .A1(n14709), .A2(n14268), .ZN(n21588) );
  INV_X1 U12839 ( .A(n21544), .ZN(n21436) );
  AND2_X1 U12840 ( .A1(n14282), .A2(n14277), .ZN(n21605) );
  AND2_X1 U12841 ( .A1(n19892), .A2(n22202), .ZN(n19888) );
  NAND2_X1 U12842 ( .A1(n13827), .A2(n19965), .ZN(n15239) );
  INV_X1 U12844 ( .A(n19923), .ZN(n19955) );
  AND2_X1 U12845 ( .A1(n19923), .A2(n13783), .ZN(n19946) );
  INV_X1 U12846 ( .A(n21389), .ZN(n21337) );
  NOR2_X1 U12847 ( .A1(n21333), .A2(n21388), .ZN(n21265) );
  INV_X1 U12848 ( .A(n21256), .ZN(n21314) );
  AND2_X1 U12849 ( .A1(n13457), .A2(n13437), .ZN(n21382) );
  INV_X1 U12850 ( .A(n21725), .ZN(n22215) );
  INV_X1 U12851 ( .A(n22221), .ZN(n22232) );
  OAI21_X1 U12852 ( .B1(n22238), .B2(n21770), .A(n21887), .ZN(n22240) );
  AND2_X1 U12853 ( .A1(n21792), .A2(n21873), .ZN(n22250) );
  AND2_X1 U12854 ( .A1(n21792), .A2(n21876), .ZN(n22257) );
  INV_X1 U12855 ( .A(n22261), .ZN(n22264) );
  INV_X1 U12856 ( .A(n22286), .ZN(n22276) );
  INV_X1 U12857 ( .A(n21846), .ZN(n22289) );
  NOR2_X1 U12858 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21715), .ZN(n22199) );
  INV_X1 U12859 ( .A(n21763), .ZN(n21845) );
  AND2_X1 U12860 ( .A1(n16765), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13321) );
  INV_X1 U12861 ( .A(n16072), .ZN(n18347) );
  AND2_X1 U12862 ( .A1(n15824), .A2(n15818), .ZN(n18380) );
  AND2_X1 U12863 ( .A1(n16965), .A2(n15815), .ZN(n18405) );
  INV_X1 U12864 ( .A(n18283), .ZN(n18404) );
  OR2_X1 U12865 ( .A1(n14602), .A2(n14763), .ZN(n14805) );
  AND2_X1 U12866 ( .A1(n14529), .A2(n14527), .ZN(n18996) );
  NOR2_X1 U12867 ( .A1(n13552), .A2(n19586), .ZN(n19587) );
  AND2_X1 U12868 ( .A1(n17018), .A2(n13537), .ZN(n17005) );
  INV_X1 U12869 ( .A(n18422), .ZN(n18460) );
  INV_X1 U12870 ( .A(n13500), .ZN(n19200) );
  OAI21_X2 U12871 ( .B1(n16694), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14337), 
        .ZN(n19219) );
  INV_X1 U12872 ( .A(n19142), .ZN(n19085) );
  NAND2_X1 U12873 ( .A1(n19223), .A2(n19222), .ZN(n19715) );
  INV_X1 U12874 ( .A(n19686), .ZN(n19679) );
  OAI21_X1 U12875 ( .B1(n19155), .B2(n19154), .A(n19153), .ZN(n19680) );
  NAND2_X1 U12876 ( .A1(n19198), .A2(n19085), .ZN(n19131) );
  INV_X1 U12877 ( .A(n19641), .ZN(n19634) );
  OAI21_X1 U12878 ( .B1(n19077), .B2(n19076), .A(n19075), .ZN(n19635) );
  NAND2_X1 U12879 ( .A1(n19035), .A2(n19034), .ZN(n19167) );
  INV_X1 U12880 ( .A(n19620), .ZN(n19610) );
  INV_X1 U12881 ( .A(n19523), .ZN(n19519) );
  INV_X1 U12882 ( .A(n19336), .ZN(n19332) );
  INV_X1 U12883 ( .A(n19608), .ZN(n19603) );
  INV_X1 U12884 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18022) );
  INV_X1 U12885 ( .A(n20445), .ZN(n20468) );
  NOR2_X2 U12886 ( .A1(n21166), .A2(n20088), .ZN(n20445) );
  NOR2_X1 U12887 ( .A1(n20387), .A2(n21173), .ZN(n20281) );
  INV_X1 U12888 ( .A(n17519), .ZN(n17506) );
  NOR2_X1 U12889 ( .A1(n11546), .A2(n11545), .ZN(n18898) );
  NAND2_X1 U12890 ( .A1(n20685), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20675) );
  NOR3_X1 U12891 ( .A1(n20625), .A2(n20699), .A3(n20576), .ZN(n20575) );
  NAND2_X1 U12892 ( .A1(n20709), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n20699) );
  INV_X1 U12893 ( .A(n18898), .ZN(n20521) );
  INV_X1 U12894 ( .A(n17755), .ZN(n17747) );
  NAND2_X1 U12895 ( .A1(n11658), .A2(n17822), .ZN(n20869) );
  OAI21_X1 U12896 ( .B1(n20738), .B2(n20723), .A(n11620), .ZN(n20946) );
  INV_X1 U12897 ( .A(n21110), .ZN(n21120) );
  NOR2_X1 U12898 ( .A1(n20849), .A2(n20848), .ZN(n20877) );
  INV_X1 U12899 ( .A(n21022), .ZN(n21006) );
  NOR2_X1 U12900 ( .A1(n20997), .A2(n21132), .ZN(n20847) );
  INV_X1 U12901 ( .A(n20736), .ZN(n21178) );
  INV_X1 U12902 ( .A(n14526), .ZN(n16187) );
  NAND2_X1 U12903 ( .A1(n21623), .A2(n13504), .ZN(n13557) );
  INV_X1 U12904 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21881) );
  AND2_X1 U12905 ( .A1(n15358), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15351) );
  INV_X1 U12906 ( .A(n21588), .ZN(n21602) );
  INV_X1 U12907 ( .A(n19930), .ZN(n21493) );
  INV_X1 U12908 ( .A(n19780), .ZN(n19815) );
  OR2_X1 U12909 ( .A1(n13640), .A2(n21915), .ZN(n13670) );
  OAI21_X1 U12910 ( .B1(n15448), .B2(n15442), .A(n15441), .ZN(n21585) );
  NAND2_X1 U12911 ( .A1(n21610), .A2(n13781), .ZN(n19923) );
  INV_X1 U12912 ( .A(n19946), .ZN(n19964) );
  INV_X1 U12913 ( .A(n21382), .ZN(n21399) );
  INV_X1 U12914 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21897) );
  OR2_X1 U12915 ( .A1(n21753), .A2(n21819), .ZN(n22219) );
  INV_X1 U12916 ( .A(n21752), .ZN(n22236) );
  NAND2_X1 U12917 ( .A1(n21792), .A2(n21845), .ZN(n22248) );
  NAND2_X1 U12918 ( .A1(n21803), .A2(n21845), .ZN(n22273) );
  OR2_X1 U12919 ( .A1(n21842), .A2(n21822), .ZN(n22286) );
  NAND2_X1 U12920 ( .A1(n21877), .A2(n21845), .ZN(n22300) );
  NAND2_X1 U12921 ( .A1(n21877), .A2(n21876), .ZN(n22318) );
  INV_X1 U12922 ( .A(n21634), .ZN(n21636) );
  NOR2_X1 U12923 ( .A1(n13508), .A2(n13507), .ZN(n16965) );
  INV_X1 U12924 ( .A(n18405), .ZN(n18354) );
  OR2_X1 U12925 ( .A1(n13846), .A2(n13741), .ZN(n19034) );
  INV_X1 U12926 ( .A(n19465), .ZN(n19278) );
  OR2_X1 U12927 ( .A1(n19465), .A2(n13750), .ZN(n19468) );
  INV_X1 U12928 ( .A(n17076), .ZN(n17110) );
  INV_X1 U12929 ( .A(n17005), .ZN(n17042) );
  INV_X1 U12930 ( .A(n17021), .ZN(n17038) );
  NAND2_X1 U12931 ( .A1(n12815), .A2(n13998), .ZN(n18450) );
  INV_X1 U12932 ( .A(n16695), .ZN(n16690) );
  OR2_X1 U12933 ( .A1(n19193), .A2(n19192), .ZN(n19711) );
  OR2_X1 U12934 ( .A1(n19193), .A2(n19167), .ZN(n19700) );
  NOR2_X1 U12935 ( .A1(n19166), .A2(n19165), .ZN(n19693) );
  AOI21_X1 U12936 ( .B1(n19151), .B2(n19154), .A(n19149), .ZN(n19684) );
  OR2_X1 U12937 ( .A1(n19131), .A2(n19192), .ZN(n19677) );
  INV_X1 U12938 ( .A(n19657), .ZN(n19668) );
  OR2_X1 U12939 ( .A1(n19131), .A2(n19143), .ZN(n19661) );
  OR2_X1 U12940 ( .A1(n19083), .A2(n19192), .ZN(n19649) );
  OR2_X1 U12941 ( .A1(n19083), .A2(n19182), .ZN(n19641) );
  OR2_X1 U12942 ( .A1(n19083), .A2(n19167), .ZN(n19639) );
  AOI22_X1 U12943 ( .A1(n14342), .A2(n14341), .B1(n14340), .B2(n14339), .ZN(
        n19626) );
  OR2_X1 U12944 ( .A1(n19051), .A2(n19182), .ZN(n19620) );
  OAI21_X1 U12945 ( .B1(n19044), .B2(n19040), .A(n19039), .ZN(n19614) );
  OR2_X1 U12946 ( .A1(n19051), .A2(n19143), .ZN(n19719) );
  INV_X1 U12947 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21685) );
  INV_X1 U12948 ( .A(n20516), .ZN(n20498) );
  INV_X1 U12949 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20174) );
  NAND3_X1 U12950 ( .A1(n11567), .A2(n11566), .A3(n11565), .ZN(n20625) );
  INV_X1 U12951 ( .A(n17429), .ZN(n17443) );
  NOR2_X1 U12952 ( .A1(n20346), .A2(n17472), .ZN(n17490) );
  INV_X1 U12953 ( .A(n20700), .ZN(n20686) );
  NOR2_X1 U12954 ( .A1(n20581), .A2(n20553), .ZN(n20552) );
  NOR2_X1 U12955 ( .A1(n11422), .A2(n11421), .ZN(n20566) );
  NAND2_X1 U12956 ( .A1(n20710), .A2(n20596), .ZN(n20691) );
  INV_X1 U12957 ( .A(n17973), .ZN(n17972) );
  NAND2_X1 U12958 ( .A1(n17806), .A2(n21058), .ZN(n17753) );
  NAND2_X1 U12959 ( .A1(n11733), .A2(n17912), .ZN(n17810) );
  INV_X1 U12960 ( .A(n17911), .ZN(n17895) );
  INV_X1 U12961 ( .A(n11705), .ZN(n20997) );
  INV_X1 U12962 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21144) );
  INV_X1 U12963 ( .A(n21647), .ZN(n16702) );
  NAND2_X1 U12964 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20769) );
  INV_X1 U12965 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20937) );
  NOR2_X1 U12966 ( .A1(n20769), .A2(n20937), .ZN(n17596) );
  NAND2_X1 U12967 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17596), .ZN(
        n11707) );
  INV_X1 U12968 ( .A(n11707), .ZN(n20932) );
  NAND2_X1 U12969 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n20932), .ZN(
        n17668) );
  AOI22_X1 U12970 ( .A1(n17435), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11402) );
  AND2_X2 U12971 ( .A1(n20712), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n20752) );
  NAND2_X2 U12972 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21143), .ZN(
        n20741) );
  AOI22_X1 U12973 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U12974 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11400) );
  NAND3_X1 U12975 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n20761), .ZN(n20755) );
  INV_X2 U12976 ( .A(n20739), .ZN(n17474) );
  AOI22_X1 U12977 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U12978 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11412) );
  AOI22_X1 U12979 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11410) );
  INV_X2 U12980 ( .A(n11377), .ZN(n17498) );
  INV_X1 U12981 ( .A(n11435), .ZN(n11484) );
  AOI22_X1 U12982 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U12983 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11408) );
  NOR3_X4 U12984 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11406), .A3(
        n20109), .ZN(n11578) );
  AOI22_X1 U12985 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U12986 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11411) );
  AOI22_X1 U12987 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U12988 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U12989 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U12990 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U12991 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11422) );
  INV_X2 U12992 ( .A(n11377), .ZN(n17481) );
  AOI22_X1 U12993 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U12994 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U12995 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U12996 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11417) );
  NAND4_X1 U12997 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(
        n11421) );
  AOI22_X1 U12998 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U12999 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U13000 ( .A1(n11441), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U13001 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11423) );
  NAND4_X1 U13002 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11432) );
  AOI22_X1 U13003 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11449), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U13004 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U13005 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U13006 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11427) );
  NAND4_X1 U13007 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11431) );
  INV_X1 U13008 ( .A(n20579), .ZN(n11448) );
  AOI22_X1 U13009 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17462), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U13010 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n10974), .ZN(n11438) );
  AOI22_X1 U13011 ( .A1(n11483), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17498), .ZN(n11437) );
  AOI22_X1 U13012 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10960), .B1(
        n11578), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11436) );
  NAND4_X1 U13013 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11447) );
  AOI22_X1 U13014 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17499), .B1(
        n10952), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U13015 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U13016 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17220), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10948), .ZN(n11443) );
  AOI22_X1 U13017 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11441), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n11450), .ZN(n11442) );
  NAND4_X1 U13018 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  OR2_X2 U13019 ( .A1(n11447), .A2(n11446), .ZN(n20698) );
  AOI22_X1 U13020 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U13021 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11459) );
  INV_X1 U13022 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U13023 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11451) );
  OAI21_X1 U13024 ( .B1(n11547), .B2(n17342), .A(n11451), .ZN(n11457) );
  AOI22_X1 U13025 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U13026 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U13027 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U13028 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U13029 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11456) );
  AOI211_X1 U13030 ( .C1(n17475), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n11457), .B(n11456), .ZN(n11458) );
  NAND3_X1 U13031 ( .A1(n11460), .A2(n11459), .A3(n11458), .ZN(n11636) );
  AOI22_X1 U13032 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U13033 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U13034 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11462) );
  OAI21_X1 U13035 ( .B1(n11547), .B2(n17353), .A(n11462), .ZN(n11468) );
  AOI22_X1 U13036 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U13037 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U13038 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U13039 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U13040 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11467) );
  AOI211_X1 U13041 ( .C1(n11441), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11468), .B(n11467), .ZN(n11469) );
  NAND3_X1 U13042 ( .A1(n11471), .A2(n11470), .A3(n11469), .ZN(n11632) );
  AOI22_X1 U13043 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U13044 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11480) );
  INV_X1 U13045 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17157) );
  AOI22_X1 U13046 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11472) );
  OAI21_X1 U13047 ( .B1(n11547), .B2(n17157), .A(n11472), .ZN(n11478) );
  AOI22_X1 U13048 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U13049 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11578), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U13050 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U13051 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11473) );
  NAND4_X1 U13052 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11477) );
  AOI211_X1 U13053 ( .C1(n17475), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n11478), .B(n11477), .ZN(n11479) );
  NAND3_X1 U13054 ( .A1(n11481), .A2(n11480), .A3(n11479), .ZN(n11733) );
  INV_X1 U13055 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21090) );
  INV_X1 U13056 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U13057 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U13058 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U13059 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U13060 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11485) );
  NAND4_X1 U13061 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11496) );
  INV_X1 U13062 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U13063 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11489) );
  OAI21_X1 U13064 ( .B1(n11547), .B2(n17143), .A(n11489), .ZN(n11490) );
  INV_X1 U13065 ( .A(n11490), .ZN(n11494) );
  AOI22_X1 U13066 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U13067 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U13068 ( .A1(n11441), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U13069 ( .A1(n11494), .A2(n11380), .ZN(n11495) );
  INV_X1 U13070 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20801) );
  NAND2_X1 U13071 ( .A1(n20579), .A2(n11627), .ZN(n11498) );
  NOR2_X1 U13072 ( .A1(n20801), .A2(n11499), .ZN(n11500) );
  XNOR2_X1 U13073 ( .A(n11502), .B(n11501), .ZN(n17890) );
  XNOR2_X1 U13074 ( .A(n20570), .B(n11639), .ZN(n17889) );
  NOR2_X1 U13075 ( .A1(n11502), .A2(n11501), .ZN(n11503) );
  NOR2_X1 U13076 ( .A1(n17888), .A2(n11503), .ZN(n17880) );
  INV_X1 U13077 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20819) );
  XOR2_X1 U13078 ( .A(n11635), .B(n11504), .Z(n11505) );
  XOR2_X1 U13079 ( .A(n20819), .B(n11505), .Z(n17879) );
  NOR2_X1 U13080 ( .A1(n17880), .A2(n17879), .ZN(n17878) );
  NOR2_X1 U13081 ( .A1(n17878), .A2(n11506), .ZN(n11510) );
  INV_X1 U13082 ( .A(n11632), .ZN(n20561) );
  XOR2_X1 U13083 ( .A(n20561), .B(n11507), .Z(n11509) );
  NOR2_X1 U13084 ( .A1(n11510), .A2(n11509), .ZN(n11511) );
  INV_X1 U13085 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20849) );
  XNOR2_X1 U13086 ( .A(n11630), .B(n11512), .ZN(n11513) );
  XOR2_X1 U13087 ( .A(n20849), .B(n11513), .Z(n17853) );
  NOR2_X2 U13088 ( .A1(n17852), .A2(n11514), .ZN(n11516) );
  OAI21_X1 U13089 ( .B1(n11515), .B2(n11733), .A(n17708), .ZN(n11517) );
  XNOR2_X1 U13090 ( .A(n11516), .B(n11517), .ZN(n17841) );
  NOR2_X1 U13091 ( .A1(n20850), .A2(n17841), .ZN(n17840) );
  NOR2_X1 U13092 ( .A1(n11516), .A2(n11517), .ZN(n11518) );
  NAND2_X1 U13093 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17708), .ZN(
        n11519) );
  OAI21_X1 U13094 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17708), .A(
        n11519), .ZN(n17827) );
  INV_X1 U13095 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20918) );
  NAND2_X1 U13096 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20880) );
  INV_X1 U13097 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20899) );
  INV_X1 U13098 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20875) );
  NOR3_X1 U13099 ( .A1(n20880), .A2(n20899), .A3(n20875), .ZN(n20900) );
  NAND2_X1 U13100 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20900), .ZN(
        n20919) );
  INV_X1 U13101 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20915) );
  NOR3_X1 U13102 ( .A1(n20918), .A2(n20919), .A3(n20915), .ZN(n21058) );
  INV_X1 U13103 ( .A(n21058), .ZN(n11704) );
  NOR2_X1 U13104 ( .A1(n17794), .A2(n11704), .ZN(n11520) );
  INV_X1 U13105 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21115) );
  INV_X1 U13106 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20874) );
  NAND2_X1 U13107 ( .A1(n21115), .A2(n20874), .ZN(n17807) );
  NOR2_X1 U13108 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17807), .ZN(
        n17578) );
  NAND2_X1 U13109 ( .A1(n17578), .A2(n20899), .ZN(n17585) );
  NOR2_X1 U13110 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17585), .ZN(
        n17554) );
  OAI221_X1 U13111 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17708), 
        .C1(n21090), .C2(n11520), .A(n11522), .ZN(n17757) );
  NOR2_X1 U13112 ( .A1(n17757), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17756) );
  INV_X1 U13113 ( .A(n17708), .ZN(n17793) );
  NOR2_X2 U13114 ( .A1(n17756), .A2(n17793), .ZN(n17618) );
  INV_X1 U13115 ( .A(n11520), .ZN(n11521) );
  NAND2_X1 U13116 ( .A1(n11522), .A2(n11521), .ZN(n17561) );
  NAND2_X1 U13117 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21065) );
  INV_X1 U13118 ( .A(n21065), .ZN(n17530) );
  INV_X1 U13119 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21071) );
  NOR2_X1 U13120 ( .A1(n21065), .A2(n21071), .ZN(n17626) );
  INV_X1 U13121 ( .A(n17626), .ZN(n11660) );
  NOR2_X1 U13122 ( .A1(n11660), .A2(n17668), .ZN(n21019) );
  NAND2_X1 U13123 ( .A1(n17708), .A2(n21071), .ZN(n17619) );
  INV_X1 U13124 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21048) );
  INV_X1 U13125 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21053) );
  NAND2_X1 U13126 ( .A1(n21048), .A2(n21053), .ZN(n21051) );
  OR3_X1 U13127 ( .A1(n17619), .A2(n21051), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17598) );
  NOR2_X1 U13128 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17598), .ZN(
        n17645) );
  INV_X1 U13129 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U13130 ( .A1(n21019), .A2(n17561), .B1(n17645), .B2(n17650), .ZN(
        n11523) );
  INV_X1 U13131 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17666) );
  AND2_X2 U13132 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17660), .ZN(
        n17709) );
  INV_X1 U13133 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20962) );
  INV_X1 U13134 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20963) );
  NAND3_X1 U13135 ( .A1(n11524), .A2(n20962), .A3(n20963), .ZN(n11525) );
  AOI22_X2 U13136 ( .A1(n17709), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n17708), .B2(n11525), .ZN(n11526) );
  INV_X1 U13137 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20980) );
  NAND2_X1 U13138 ( .A1(n11715), .A2(n17698), .ZN(n17691) );
  NOR2_X1 U13139 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17793), .ZN(
        n11720) );
  AOI21_X1 U13140 ( .B1(n17793), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11720), .ZN(n17692) );
  AOI22_X1 U13141 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U13142 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11535) );
  INV_X1 U13143 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U13144 ( .A1(n17300), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11527) );
  OAI21_X1 U13145 ( .B1(n11484), .B2(n17514), .A(n11527), .ZN(n11533) );
  AOI22_X1 U13146 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U13147 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10952), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U13148 ( .A1(n10948), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U13149 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11528) );
  NAND4_X1 U13150 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11532) );
  AOI22_X1 U13151 ( .A1(n17435), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U13152 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U13153 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11538) );
  INV_X2 U13154 ( .A(n11547), .ZN(n17378) );
  AOI22_X1 U13155 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11537) );
  NAND4_X1 U13156 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11546) );
  AOI22_X1 U13157 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U13158 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U13159 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U13160 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11541) );
  NAND4_X1 U13161 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11545) );
  NAND2_X1 U13162 ( .A1(n18898), .A2(n20520), .ZN(n11623) );
  AOI22_X1 U13163 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13164 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U13165 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U13166 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U13167 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11557) );
  AOI22_X1 U13168 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U13169 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11554) );
  INV_X2 U13170 ( .A(n11484), .ZN(n17444) );
  AOI22_X1 U13171 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U13172 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U13173 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11556) );
  AOI22_X1 U13174 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U13175 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U13176 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11558) );
  OAI21_X1 U13177 ( .B1(n11484), .B2(n17157), .A(n11558), .ZN(n11564) );
  AOI22_X1 U13178 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U13179 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U13180 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U13181 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U13182 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11563) );
  NAND3_X1 U13183 ( .A1(n18898), .A2(n18766), .A3(n20625), .ZN(n11613) );
  AOI22_X1 U13184 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U13185 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13186 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13187 ( .A1(n10948), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U13188 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11577) );
  AOI22_X1 U13189 ( .A1(n10974), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13190 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U13191 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U13192 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U13193 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  INV_X1 U13194 ( .A(n18725), .ZN(n17131) );
  AOI22_X1 U13195 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U13196 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13197 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11579) );
  OAI21_X1 U13198 ( .B1(n11484), .B2(n17353), .A(n11579), .ZN(n11585) );
  AOI22_X1 U13199 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U13200 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U13201 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U13202 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U13203 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  AOI22_X1 U13204 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U13205 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U13206 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U13207 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U13208 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11598) );
  AOI22_X1 U13209 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U13210 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13211 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U13212 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11593) );
  NAND4_X1 U13213 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11597) );
  NAND2_X1 U13214 ( .A1(n11609), .A2(n20586), .ZN(n11680) );
  AOI22_X1 U13215 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U13216 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U13217 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13218 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U13219 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11608) );
  AOI22_X1 U13220 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13221 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U13222 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13223 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U13224 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  NAND2_X1 U13225 ( .A1(n18807), .A2(n18725), .ZN(n11695) );
  NAND2_X1 U13226 ( .A1(n11609), .A2(n18807), .ZN(n11683) );
  NOR3_X4 U13227 ( .A1(n11687), .A2(n11696), .A3(n11625), .ZN(n11619) );
  NOR2_X2 U13228 ( .A1(n11689), .A2(n11610), .ZN(n21135) );
  NAND2_X1 U13229 ( .A1(n20084), .A2(n11610), .ZN(n21165) );
  INV_X1 U13230 ( .A(n11621), .ZN(n14838) );
  NAND2_X1 U13231 ( .A1(n18807), .A2(n11623), .ZN(n11692) );
  NAND3_X1 U13232 ( .A1(n11611), .A2(n11687), .A3(n11616), .ZN(n11622) );
  NAND2_X1 U13233 ( .A1(n18807), .A2(n18766), .ZN(n20723) );
  NAND2_X1 U13234 ( .A1(n20521), .A2(n20084), .ZN(n11624) );
  NOR2_X1 U13235 ( .A1(n20597), .A2(n20710), .ZN(n20528) );
  INV_X1 U13236 ( .A(n11612), .ZN(n11614) );
  OAI21_X1 U13237 ( .B1(n18766), .B2(n11614), .A(n11613), .ZN(n11615) );
  OAI221_X1 U13238 ( .B1(n11617), .B2(n11616), .C1(n11617), .C2(n11680), .A(
        n11615), .ZN(n11618) );
  INV_X1 U13239 ( .A(n11620), .ZN(n20751) );
  NAND2_X1 U13240 ( .A1(n11624), .A2(n11623), .ZN(n16707) );
  INV_X1 U13241 ( .A(n11625), .ZN(n20724) );
  INV_X1 U13242 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20942) );
  INV_X1 U13243 ( .A(n11733), .ZN(n20554) );
  INV_X1 U13244 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20858) );
  INV_X1 U13245 ( .A(n20703), .ZN(n11640) );
  OAI21_X1 U13246 ( .B1(n11627), .B2(n11640), .A(n20579), .ZN(n11638) );
  AND2_X1 U13247 ( .A1(n11636), .A2(n11638), .ZN(n11634) );
  NAND2_X1 U13248 ( .A1(n11634), .A2(n11635), .ZN(n11631) );
  NOR2_X1 U13249 ( .A1(n20561), .A2(n11631), .ZN(n11629) );
  NAND2_X1 U13250 ( .A1(n11629), .A2(n11630), .ZN(n11628) );
  NOR2_X1 U13251 ( .A1(n20554), .A2(n11628), .ZN(n11657) );
  XOR2_X1 U13252 ( .A(n20554), .B(n11628), .Z(n17847) );
  XOR2_X1 U13253 ( .A(n11630), .B(n11629), .Z(n11650) );
  XNOR2_X1 U13254 ( .A(n11632), .B(n11631), .ZN(n11633) );
  NAND2_X1 U13255 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11633), .ZN(
        n11649) );
  XOR2_X1 U13256 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11633), .Z(
        n17865) );
  XOR2_X1 U13257 ( .A(n11635), .B(n11634), .Z(n11646) );
  NAND2_X1 U13258 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11637), .ZN(
        n11645) );
  OAI21_X1 U13259 ( .B1(n11640), .B2(n11639), .A(n11638), .ZN(n11641) );
  NAND2_X1 U13260 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11641), .ZN(
        n11644) );
  XNOR2_X1 U13261 ( .A(n20801), .B(n11641), .ZN(n20794) );
  AOI21_X1 U13262 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20698), .A(
        n20703), .ZN(n11643) );
  INV_X1 U13263 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20886) );
  NOR2_X1 U13264 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20698), .ZN(
        n11642) );
  AOI221_X1 U13265 ( .B1(n20703), .B2(n20698), .C1(n11643), .C2(n20886), .A(
        n11642), .ZN(n20793) );
  NAND2_X1 U13266 ( .A1(n11646), .A2(n11647), .ZN(n11648) );
  XNOR2_X1 U13267 ( .A(n11647), .B(n11646), .ZN(n17877) );
  NAND2_X1 U13268 ( .A1(n11650), .A2(n11651), .ZN(n11652) );
  XOR2_X1 U13269 ( .A(n11651), .B(n11650), .Z(n17857) );
  NAND2_X1 U13270 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17857), .ZN(
        n17856) );
  NAND2_X1 U13271 ( .A1(n11657), .A2(n11653), .ZN(n11658) );
  NAND2_X1 U13272 ( .A1(n17847), .A2(n17846), .ZN(n11655) );
  NAND2_X1 U13273 ( .A1(n11657), .A2(n11656), .ZN(n11654) );
  OAI211_X1 U13274 ( .C1(n11657), .C2(n11656), .A(n11655), .B(n11654), .ZN(
        n17823) );
  NAND2_X1 U13275 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17823), .ZN(
        n17822) );
  AOI22_X1 U13276 ( .A1(n21063), .A2(n17786), .B1(n21125), .B2(n20869), .ZN(
        n20879) );
  NAND2_X1 U13277 ( .A1(n21058), .A2(n17626), .ZN(n17534) );
  NOR2_X1 U13278 ( .A1(n20858), .A2(n20850), .ZN(n20878) );
  INV_X1 U13279 ( .A(n20878), .ZN(n17552) );
  AOI21_X1 U13280 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20813) );
  INV_X1 U13281 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20833) );
  NOR3_X1 U13282 ( .A1(n20819), .A2(n11501), .A3(n20833), .ZN(n20836) );
  INV_X1 U13283 ( .A(n20836), .ZN(n11659) );
  NOR2_X1 U13284 ( .A1(n20813), .A2(n11659), .ZN(n20826) );
  NAND2_X1 U13285 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20826), .ZN(
        n20851) );
  NOR2_X1 U13286 ( .A1(n17552), .A2(n20851), .ZN(n20887) );
  NAND2_X1 U13287 ( .A1(n21058), .A2(n20887), .ZN(n21064) );
  NOR2_X1 U13288 ( .A1(n11660), .A2(n21064), .ZN(n11706) );
  INV_X1 U13289 ( .A(n21112), .ZN(n21072) );
  NOR2_X1 U13290 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21103), .ZN(
        n20784) );
  NAND3_X1 U13291 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20836), .ZN(n20827) );
  NOR2_X1 U13292 ( .A1(n20849), .A2(n20827), .ZN(n20853) );
  NAND2_X1 U13293 ( .A1(n20878), .A2(n20853), .ZN(n21113) );
  NOR2_X1 U13294 ( .A1(n17534), .A2(n21113), .ZN(n20933) );
  AOI22_X1 U13295 ( .A1(n21126), .A2(n11706), .B1(n20810), .B2(n20933), .ZN(
        n20945) );
  NAND3_X1 U13296 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20968) );
  NOR2_X1 U13297 ( .A1(n20962), .A2(n20968), .ZN(n20978) );
  NAND2_X1 U13298 ( .A1(n21144), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11669) );
  AOI22_X1 U13299 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n21153), .B2(n21143), .ZN(
        n11666) );
  AOI22_X1 U13300 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21139), .B1(
        n11663), .B2(n20761), .ZN(n11670) );
  INV_X1 U13301 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21156) );
  NOR2_X1 U13302 ( .A1(n11663), .A2(n20761), .ZN(n11671) );
  NAND2_X1 U13303 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21139), .ZN(
        n11664) );
  OAI22_X1 U13304 ( .A1(n11670), .A2(n21156), .B1(n11671), .B2(n11664), .ZN(
        n11668) );
  INV_X1 U13305 ( .A(n11668), .ZN(n11665) );
  OAI211_X1 U13306 ( .C1(n21144), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11669), .B(n11665), .ZN(n11679) );
  XNOR2_X1 U13307 ( .A(n11667), .B(n11666), .ZN(n11675) );
  XNOR2_X1 U13308 ( .A(n11669), .B(n11678), .ZN(n11674) );
  OAI21_X1 U13309 ( .B1(n21156), .B2(n11671), .A(n11670), .ZN(n11672) );
  OAI21_X1 U13310 ( .B1(n21139), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n11672), .ZN(n11673) );
  INV_X1 U13311 ( .A(n11673), .ZN(n11677) );
  OAI21_X1 U13312 ( .B1(n11679), .B2(n11675), .A(n21130), .ZN(n11719) );
  INV_X1 U13313 ( .A(n11719), .ZN(n21131) );
  NAND2_X1 U13314 ( .A1(n21131), .A2(n20520), .ZN(n11681) );
  OAI211_X1 U13315 ( .C1(n11679), .C2(n11678), .A(n11677), .B(n11676), .ZN(
        n14839) );
  OAI22_X1 U13316 ( .A1(n11682), .A2(n11681), .B1(n14839), .B2(n11680), .ZN(
        n11698) );
  INV_X1 U13317 ( .A(n11683), .ZN(n11685) );
  INV_X1 U13318 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21689) );
  NAND2_X1 U13319 ( .A1(n21689), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18012) );
  INV_X2 U13320 ( .A(n18012), .ZN(n18006) );
  INV_X1 U13321 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21698) );
  NOR2_X1 U13322 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n21698), .ZN(n21695) );
  NOR2_X1 U13323 ( .A1(n21698), .A2(n18012), .ZN(n18003) );
  INV_X2 U13324 ( .A(n18003), .ZN(n18005) );
  OAI21_X1 U13325 ( .B1(n18006), .B2(n21695), .A(n18005), .ZN(n20085) );
  OAI21_X1 U13326 ( .B1(n18807), .B2(n20520), .A(n20085), .ZN(n11684) );
  AOI21_X1 U13327 ( .B1(n18807), .B2(n20520), .A(n11684), .ZN(n21133) );
  NAND2_X1 U13328 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21649) );
  NOR3_X1 U13329 ( .A1(n11685), .A2(n21133), .A3(n20029), .ZN(n11697) );
  INV_X1 U13330 ( .A(n11686), .ZN(n11694) );
  INV_X1 U13331 ( .A(n11687), .ZN(n17130) );
  OAI211_X1 U13332 ( .C1(n20710), .C2(n18725), .A(n11688), .B(n17130), .ZN(
        n11691) );
  INV_X1 U13333 ( .A(n11689), .ZN(n11690) );
  OAI21_X1 U13334 ( .B1(n11692), .B2(n11691), .A(n11690), .ZN(n11693) );
  OAI211_X1 U13335 ( .C1(n11696), .C2(n11695), .A(n11694), .B(n11693), .ZN(
        n14842) );
  AOI211_X1 U13336 ( .C1(n18807), .C2(n11698), .A(n11697), .B(n14842), .ZN(
        n11699) );
  NOR2_X1 U13337 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20082), .ZN(n21169) );
  NAND2_X1 U13338 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21169), .ZN(n21188) );
  AOI221_X1 U13339 ( .B1(n18725), .B2(n11699), .C1(n14839), .C2(n11699), .A(
        n21188), .ZN(n11705) );
  OAI21_X1 U13340 ( .B1(n11700), .B2(n20554), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11702) );
  NAND3_X1 U13341 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17793), .A3(
        n11701), .ZN(n17737) );
  NAND2_X1 U13342 ( .A1(n11702), .A2(n17737), .ZN(n11713) );
  NAND2_X1 U13343 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17728) );
  INV_X1 U13344 ( .A(n20919), .ZN(n11703) );
  NAND2_X1 U13345 ( .A1(n17786), .A2(n11703), .ZN(n17765) );
  NAND2_X1 U13346 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n20978), .ZN(
        n17688) );
  NAND2_X1 U13347 ( .A1(n17626), .A2(n17596), .ZN(n17595) );
  NOR2_X1 U13348 ( .A1(n17688), .A2(n17595), .ZN(n17731) );
  NAND2_X1 U13349 ( .A1(n21017), .A2(n17731), .ZN(n20976) );
  NOR2_X1 U13350 ( .A1(n17728), .A2(n20976), .ZN(n20991) );
  OR2_X1 U13351 ( .A1(n20991), .A2(n20993), .ZN(n11711) );
  NAND2_X1 U13352 ( .A1(n11703), .A2(n20869), .ZN(n17777) );
  NOR2_X1 U13353 ( .A1(n17728), .A2(n17688), .ZN(n11740) );
  NAND2_X1 U13354 ( .A1(n17651), .A2(n11740), .ZN(n20988) );
  NOR2_X1 U13355 ( .A1(n11704), .A2(n21113), .ZN(n21060) );
  INV_X1 U13356 ( .A(n17731), .ZN(n17701) );
  NOR2_X1 U13357 ( .A1(n20980), .A2(n17701), .ZN(n17689) );
  NAND2_X1 U13358 ( .A1(n21060), .A2(n17689), .ZN(n11741) );
  INV_X1 U13359 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n17919) );
  INV_X1 U13360 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20081) );
  NAND2_X1 U13361 ( .A1(n17919), .A2(n20081), .ZN(n20022) );
  NOR2_X1 U13362 ( .A1(n20022), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17520) );
  NAND2_X1 U13363 ( .A1(n21105), .A2(n20997), .ZN(n21022) );
  INV_X1 U13364 ( .A(n11706), .ZN(n20764) );
  OAI21_X1 U13365 ( .B1(n20764), .B2(n11707), .A(n21126), .ZN(n21025) );
  OAI21_X1 U13366 ( .B1(n20978), .B2(n21094), .A(n21025), .ZN(n20975) );
  AOI221_X1 U13367 ( .B1(n20886), .B2(n20946), .C1(n11741), .C2(n20946), .A(
        n20975), .ZN(n11743) );
  OAI21_X1 U13368 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21094), .A(
        n11743), .ZN(n21002) );
  AOI211_X1 U13369 ( .C1(n21103), .C2(n11741), .A(n21006), .B(n21002), .ZN(
        n11708) );
  INV_X1 U13370 ( .A(n11708), .ZN(n11709) );
  AOI21_X1 U13371 ( .B1(n20988), .B2(n21125), .A(n11709), .ZN(n11710) );
  NAND2_X1 U13372 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  INV_X1 U13373 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20466) );
  NOR2_X1 U13374 ( .A1(n21105), .A2(n20466), .ZN(n11716) );
  NAND2_X1 U13375 ( .A1(n11718), .A2(n11717), .ZN(P3_U2834) );
  INV_X1 U13376 ( .A(n21188), .ZN(n21164) );
  NAND2_X1 U13378 ( .A1(n11721), .A2(n11720), .ZN(n17738) );
  INV_X1 U13379 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21007) );
  INV_X1 U13380 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21008) );
  INV_X1 U13381 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20716) );
  NAND2_X1 U13382 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11739) );
  NOR2_X1 U13383 ( .A1(n11739), .A2(n20988), .ZN(n11724) );
  XNOR2_X1 U13384 ( .A(n20716), .B(n11724), .ZN(n11736) );
  AOI22_X1 U13385 ( .A1(n17837), .A2(n11737), .B1(n17908), .B2(n11736), .ZN(
        n11735) );
  INV_X1 U13386 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20501) );
  INV_X1 U13387 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20185) );
  NAND2_X1 U13388 ( .A1(n17770), .A2(n17830), .ZN(n20213) );
  NAND2_X1 U13389 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20250) );
  NAND2_X1 U13390 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17564) );
  INV_X1 U13391 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20355) );
  NAND2_X1 U13392 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17604) );
  INV_X1 U13393 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n20398) );
  NAND2_X1 U13394 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17655) );
  INV_X1 U13395 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20446) );
  INV_X1 U13396 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20481) );
  XOR2_X2 U13397 ( .A(n20501), .B(n17723), .Z(n20387) );
  INV_X1 U13398 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21644) );
  INV_X1 U13399 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21176) );
  NAND2_X1 U13400 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17523) );
  NAND2_X1 U13401 ( .A1(n21176), .A2(n17523), .ZN(n20018) );
  INV_X1 U13402 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18007) );
  NOR2_X1 U13403 ( .A1(n21105), .A2(n18007), .ZN(n11738) );
  OR2_X1 U13404 ( .A1(n17528), .A2(n11093), .ZN(n17539) );
  NOR2_X1 U13405 ( .A1(n20355), .A2(n17539), .ZN(n17623) );
  NAND2_X1 U13406 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17623), .ZN(
        n17603) );
  NOR2_X1 U13407 ( .A1(n17604), .A2(n17603), .ZN(n17641) );
  NAND2_X1 U13408 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17641), .ZN(
        n17654) );
  NOR2_X1 U13409 ( .A1(n17655), .A2(n17654), .ZN(n17711) );
  NAND2_X1 U13410 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17711), .ZN(
        n17682) );
  NOR2_X1 U13411 ( .A1(n20446), .A2(n17682), .ZN(n17684) );
  NAND2_X1 U13412 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17684), .ZN(
        n17734) );
  NOR2_X1 U13413 ( .A1(n20481), .A2(n17734), .ZN(n11726) );
  NAND2_X1 U13414 ( .A1(n20082), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17917) );
  NAND2_X1 U13415 ( .A1(n21139), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20736) );
  AOI21_X1 U13416 ( .B1(n20022), .B2(n17523), .A(n21178), .ZN(n18567) );
  NAND3_X1 U13417 ( .A1(n20081), .A2(n21176), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18609) );
  INV_X2 U13418 ( .A(n18893), .ZN(n18894) );
  INV_X1 U13419 ( .A(n17680), .ZN(n17683) );
  NAND2_X1 U13420 ( .A1(n11726), .A2(n17683), .ZN(n17725) );
  XNOR2_X1 U13421 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11729) );
  NOR2_X1 U13422 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17754), .ZN(
        n17746) );
  INV_X1 U13423 ( .A(n11726), .ZN(n11727) );
  INV_X1 U13424 ( .A(n17917), .ZN(n17635) );
  AOI22_X1 U13425 ( .A1(n18894), .A2(n11727), .B1(n17635), .B2(n17745), .ZN(
        n11728) );
  NAND2_X1 U13426 ( .A1(n11728), .A2(n17918), .ZN(n17736) );
  NOR2_X1 U13427 ( .A1(n17746), .A2(n17736), .ZN(n17724) );
  OAI22_X1 U13428 ( .A1(n17725), .A2(n11729), .B1(n17724), .B2(n20501), .ZN(
        n11730) );
  AOI211_X1 U13429 ( .C1(n20387), .C2(n17747), .A(n11738), .B(n11730), .ZN(
        n11734) );
  INV_X1 U13430 ( .A(n11739), .ZN(n11731) );
  NAND2_X1 U13431 ( .A1(n20991), .A2(n11731), .ZN(n11732) );
  XNOR2_X1 U13432 ( .A(n20716), .B(n11732), .ZN(n11745) );
  INV_X1 U13433 ( .A(n17836), .ZN(n17785) );
  NAND3_X1 U13434 ( .A1(n11735), .A2(n11734), .A3(n11383), .ZN(P3_U2799) );
  NAND2_X1 U13435 ( .A1(n21093), .A2(n21125), .ZN(n20953) );
  INV_X1 U13436 ( .A(n20953), .ZN(n20965) );
  AOI22_X1 U13437 ( .A1(n21120), .A2(n11737), .B1(n20965), .B2(n11736), .ZN(
        n11751) );
  AOI21_X1 U13438 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21006), .A(
        n11738), .ZN(n11750) );
  NOR2_X1 U13439 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n11739), .ZN(
        n11747) );
  INV_X1 U13440 ( .A(n17596), .ZN(n20944) );
  INV_X1 U13441 ( .A(n11740), .ZN(n17741) );
  NOR3_X1 U13442 ( .A1(n20945), .A2(n20944), .A3(n17741), .ZN(n20990) );
  INV_X1 U13443 ( .A(n20949), .ZN(n21085) );
  INV_X1 U13444 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20998) );
  OAI21_X1 U13445 ( .B1(n20998), .B2(n11741), .A(n21103), .ZN(n20999) );
  OAI21_X1 U13446 ( .B1(n17728), .B2(n21008), .A(n21085), .ZN(n11742) );
  NAND4_X1 U13447 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n11743), .A3(
        n20999), .A4(n11742), .ZN(n21011) );
  NAND3_X1 U13448 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21085), .A3(
        n21011), .ZN(n11744) );
  OAI21_X1 U13449 ( .B1(n11745), .B2(n20993), .A(n11744), .ZN(n11746) );
  AOI21_X1 U13450 ( .B1(n11747), .B2(n20990), .A(n11746), .ZN(n11748) );
  OR2_X1 U13451 ( .A1(n11748), .A2(n20997), .ZN(n11749) );
  NAND3_X1 U13452 ( .A1(n11751), .A2(n11750), .A3(n11749), .ZN(P3_U2831) );
  AOI22_X1 U13453 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U13454 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11755) );
  AND2_X4 U13455 ( .A1(n13975), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11974) );
  AOI22_X1 U13456 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11754) );
  NAND2_X2 U13457 ( .A1(n11981), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11758) );
  INV_X2 U13458 ( .A(n11758), .ZN(n11825) );
  AOI22_X1 U13459 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U13460 ( .A1(n11757), .A2(n11756), .ZN(n11765) );
  AOI22_X1 U13461 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U13462 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U13463 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11760) );
  NAND4_X1 U13464 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11764) );
  INV_X2 U13465 ( .A(n11861), .ZN(n14524) );
  AOI22_X1 U13466 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U13467 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11768) );
  AND2_X4 U13468 ( .A1(n11981), .A2(n13952), .ZN(n15973) );
  AOI22_X1 U13469 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U13470 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U13471 ( .A1(n15897), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13472 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15896), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U13473 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U13474 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11777) );
  AND2_X1 U13475 ( .A1(n11778), .A2(n11777), .ZN(n11781) );
  AOI22_X1 U13476 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U13477 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11779) );
  NAND3_X1 U13478 ( .A1(n11781), .A2(n11780), .A3(n11779), .ZN(n11782) );
  NAND2_X1 U13479 ( .A1(n11782), .A2(n13958), .ZN(n11790) );
  INV_X2 U13480 ( .A(n11783), .ZN(n15896) );
  AOI22_X1 U13481 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U13482 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U13483 ( .A1(n15897), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U13484 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U13485 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11788) );
  NAND2_X1 U13486 ( .A1(n11788), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11789) );
  NAND2_X2 U13487 ( .A1(n11790), .A2(n11789), .ZN(n11872) );
  AOI22_X1 U13488 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10973), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U13489 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U13490 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U13491 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U13492 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11795) );
  NAND2_X1 U13493 ( .A1(n11795), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11802) );
  AOI22_X1 U13494 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U13495 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U13496 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U13497 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U13498 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  NAND2_X1 U13499 ( .A1(n11800), .A2(n13958), .ZN(n11801) );
  NAND2_X1 U13500 ( .A1(n11870), .A2(n11803), .ZN(n11855) );
  AOI22_X1 U13501 ( .A1(n15897), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U13502 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13503 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U13504 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11805) );
  NAND4_X1 U13505 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11814) );
  AOI22_X1 U13506 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U13507 ( .A1(n15897), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U13508 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U13509 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11809) );
  NAND4_X1 U13510 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n11813) );
  MUX2_X2 U13511 ( .A(n11814), .B(n11813), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19410) );
  AOI22_X1 U13512 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U13513 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U13514 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U13515 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11815) );
  NAND4_X1 U13516 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11824) );
  AOI22_X1 U13517 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U13518 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U13519 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U13520 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11819) );
  NAND4_X1 U13521 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11823) );
  MUX2_X2 U13522 ( .A(n11824), .B(n11823), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19597) );
  AOI22_X1 U13523 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U13524 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U13525 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U13526 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U13527 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11835) );
  AOI22_X1 U13528 ( .A1(n15897), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11974), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U13529 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U13530 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U13531 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U13532 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11834) );
  MUX2_X2 U13533 ( .A(n11835), .B(n11834), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12440) );
  NAND2_X2 U13534 ( .A1(n19597), .A2(n12440), .ZN(n12402) );
  NAND2_X1 U13535 ( .A1(n11868), .A2(n11857), .ZN(n11837) );
  NAND2_X1 U13536 ( .A1(n11854), .A2(n19410), .ZN(n11836) );
  NAND2_X1 U13537 ( .A1(n11837), .A2(n11836), .ZN(n11853) );
  AOI22_X1 U13538 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13539 ( .A1(n10972), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U13540 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11839) );
  NAND3_X1 U13541 ( .A1(n11841), .A2(n11840), .A3(n11839), .ZN(n11842) );
  NOR2_X1 U13542 ( .A1(n11843), .A2(n11842), .ZN(n11844) );
  NAND2_X1 U13543 ( .A1(n11844), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11851) );
  AOI22_X1 U13544 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15897), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U13545 ( .A1(n11974), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U13546 ( .A1(n15896), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U13547 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11845) );
  NAND2_X2 U13548 ( .A1(n11851), .A2(n11850), .ZN(n11860) );
  NAND3_X1 U13549 ( .A1(n11855), .A2(n11871), .A3(n11854), .ZN(n11917) );
  NAND2_X1 U13550 ( .A1(n11917), .A2(n12379), .ZN(n11856) );
  NOR2_X1 U13551 ( .A1(n11857), .A2(n11870), .ZN(n11859) );
  NAND2_X1 U13552 ( .A1(n11864), .A2(n11863), .ZN(n11885) );
  NAND2_X2 U13553 ( .A1(n11866), .A2(n11914), .ZN(n11906) );
  OAI21_X1 U13554 ( .B1(n19160), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16714), 
        .ZN(n11867) );
  NAND2_X1 U13555 ( .A1(n13715), .A2(n11871), .ZN(n11884) );
  NAND2_X1 U13556 ( .A1(n11871), .A2(n12379), .ZN(n12413) );
  NAND2_X1 U13557 ( .A1(n12402), .A2(n12413), .ZN(n12411) );
  INV_X1 U13558 ( .A(n11868), .ZN(n11869) );
  NOR2_X1 U13559 ( .A1(n11880), .A2(n11873), .ZN(n11875) );
  INV_X1 U13560 ( .A(n11854), .ZN(n11874) );
  AND2_X1 U13561 ( .A1(n12379), .A2(n11858), .ZN(n11881) );
  NAND4_X1 U13562 ( .A1(n12758), .A2(n12438), .A3(n11881), .A4(n11873), .ZN(
        n11882) );
  OAI211_X2 U13563 ( .C1(n12374), .C2(n11884), .A(n11908), .B(n11883), .ZN(
        n11930) );
  INV_X1 U13564 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n11889) );
  AND2_X4 U13565 ( .A1(n12422), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U13566 ( .A1(n12743), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U13567 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U13568 ( .A1(n11891), .A2(n11892), .ZN(n11927) );
  INV_X1 U13569 ( .A(n11891), .ZN(n11894) );
  INV_X1 U13570 ( .A(n11892), .ZN(n11893) );
  NAND2_X1 U13571 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  NAND2_X1 U13572 ( .A1(n11906), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11898) );
  NOR2_X1 U13573 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U13574 ( .A1(n11898), .A2(n11897), .ZN(n11922) );
  INV_X1 U13575 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U13576 ( .A1(n12743), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11900) );
  NAND2_X1 U13577 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11899) );
  OAI211_X1 U13578 ( .C1(n12707), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11902) );
  AOI21_X2 U13579 ( .B1(n11930), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11902), .ZN(n11923) );
  XNOR2_X1 U13580 ( .A(n11922), .B(n11923), .ZN(n11939) );
  INV_X1 U13581 ( .A(n11903), .ZN(n11904) );
  NOR2_X1 U13582 ( .A1(n11904), .A2(n12402), .ZN(n11905) );
  OAI22_X1 U13583 ( .A1(n11906), .A2(n11905), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12752), .ZN(n11910) );
  NAND2_X1 U13584 ( .A1(n12407), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U13585 ( .A1(n11910), .A2(n11909), .ZN(n11937) );
  NAND2_X1 U13586 ( .A1(n12743), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11913) );
  INV_X1 U13587 ( .A(n12407), .ZN(n18510) );
  NAND2_X1 U13588 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11911) );
  AND2_X1 U13589 ( .A1(n18510), .A2(n11911), .ZN(n11912) );
  NAND4_X1 U13590 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  AOI21_X1 U13591 ( .B1(n11930), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11916), .ZN(n11921) );
  NAND2_X1 U13592 ( .A1(n11020), .A2(n11917), .ZN(n12421) );
  AOI21_X1 U13593 ( .B1(n12421), .B2(n11918), .A(n18022), .ZN(n11919) );
  INV_X1 U13594 ( .A(n11919), .ZN(n11920) );
  NAND2_X1 U13595 ( .A1(n11921), .A2(n11920), .ZN(n11936) );
  NAND2_X1 U13596 ( .A1(n11937), .A2(n11936), .ZN(n11935) );
  NAND2_X1 U13597 ( .A1(n11939), .A2(n11935), .ZN(n11926) );
  INV_X1 U13598 ( .A(n11922), .ZN(n11924) );
  NAND2_X1 U13599 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  NAND2_X1 U13600 ( .A1(n11906), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U13601 ( .A1(n12407), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11928) );
  INV_X1 U13602 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U13603 ( .A1(n11930), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11932) );
  AOI22_X1 U13604 ( .A1(n12752), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U13605 ( .A1(n11964), .A2(n11960), .ZN(n19133) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11943) );
  NOR2_X2 U13607 ( .A1(n13944), .A2(n18499), .ZN(n11962) );
  XNOR2_X2 U13608 ( .A(n11940), .B(n11944), .ZN(n18427) );
  INV_X1 U13609 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11941) );
  OAI211_X1 U13610 ( .C1(n19133), .C2(n11943), .A(n11942), .B(n16011), .ZN(
        n11948) );
  INV_X1 U13611 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14568) );
  INV_X1 U13612 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11946) );
  INV_X1 U13613 ( .A(n11944), .ZN(n11945) );
  NAND2_X2 U13614 ( .A1(n11961), .A2(n11963), .ZN(n19161) );
  NOR2_X1 U13615 ( .A1(n11948), .A2(n11947), .ZN(n11973) );
  INV_X1 U13616 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14565) );
  INV_X1 U13617 ( .A(n19027), .ZN(n11950) );
  INV_X1 U13618 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11949) );
  INV_X1 U13619 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11952) );
  INV_X1 U13620 ( .A(n18427), .ZN(n13737) );
  INV_X1 U13621 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11951) );
  OAI22_X1 U13622 ( .A1(n11952), .A2(n12079), .B1(n19080), .B2(n11951), .ZN(
        n11953) );
  INV_X1 U13623 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U13624 ( .A1(n11961), .A2(n11957), .ZN(n12036) );
  INV_X1 U13625 ( .A(n12087), .ZN(n11956) );
  INV_X1 U13626 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11955) );
  OAI22_X1 U13627 ( .A1(n14570), .A2(n12036), .B1(n11956), .B2(n11955), .ZN(
        n11959) );
  NOR2_X1 U13628 ( .A1(n11959), .A2(n11958), .ZN(n11971) );
  INV_X1 U13629 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12510) );
  INV_X1 U13630 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12505) );
  OAI22_X1 U13631 ( .A1(n12510), .A2(n19203), .B1(n19064), .B2(n12505), .ZN(
        n11969) );
  INV_X1 U13632 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U13633 ( .A1(n11964), .A2(n11963), .ZN(n19109) );
  INV_X1 U13634 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14562) );
  OAI22_X1 U13635 ( .A1(n11967), .A2(n19109), .B1(n12086), .B2(n14562), .ZN(
        n11968) );
  NOR2_X1 U13636 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND4_X1 U13637 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n12029) );
  INV_X1 U13638 ( .A(n11974), .ZN(n15895) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U13640 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11977) );
  NAND2_X1 U13641 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11976) );
  OAI211_X1 U13642 ( .C1(n15874), .C2(n11978), .A(n11977), .B(n11976), .ZN(
        n11985) );
  NAND2_X1 U13643 ( .A1(n11979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12015) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12485) );
  AND2_X1 U13645 ( .A1(n13985), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11980) );
  NAND2_X1 U13646 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11983) );
  INV_X1 U13647 ( .A(n11981), .ZN(n13953) );
  INV_X1 U13648 ( .A(n13953), .ZN(n13970) );
  NAND2_X1 U13649 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11982) );
  OAI211_X1 U13650 ( .C1(n12015), .C2(n12485), .A(n11983), .B(n11982), .ZN(
        n11984) );
  NOR2_X1 U13651 ( .A1(n11985), .A2(n11984), .ZN(n11997) );
  AOI22_X1 U13652 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11996) );
  AND2_X2 U13653 ( .A1(n10973), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12126) );
  AOI22_X1 U13654 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11991) );
  AND2_X2 U13655 ( .A1(n11987), .A2(n13958), .ZN(n11998) );
  AOI22_X1 U13656 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11990) );
  AND2_X2 U13657 ( .A1(n16036), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12092) );
  AOI22_X1 U13658 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11989) );
  NAND3_X1 U13659 ( .A1(n11991), .A2(n11990), .A3(n11989), .ZN(n11994) );
  INV_X1 U13660 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11992) );
  INV_X1 U13661 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14509) );
  OAI22_X1 U13662 ( .A1(n11992), .A2(n14571), .B1(n14569), .B2(n14509), .ZN(
        n11993) );
  NAND3_X1 U13663 ( .A1(n11997), .A2(n11996), .A3(n11995), .ZN(n13535) );
  INV_X1 U13664 ( .A(n13535), .ZN(n12010) );
  AOI22_X1 U13665 ( .A1(n15865), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15884), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U13666 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15883), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12001) );
  INV_X1 U13667 ( .A(n12015), .ZN(n12609) );
  AOI22_X1 U13668 ( .A1(n12609), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12000) );
  INV_X1 U13669 ( .A(n15874), .ZN(n12602) );
  AOI22_X1 U13670 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12602), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U13671 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12009) );
  AOI22_X1 U13672 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15875), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U13673 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15876), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U13674 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U13675 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12092), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12004) );
  NAND4_X1 U13676 ( .A1(n12007), .A2(n12006), .A3(n12005), .A4(n12004), .ZN(
        n12008) );
  NOR2_X1 U13677 ( .A1(n12010), .A2(n12774), .ZN(n12011) );
  NAND2_X1 U13678 ( .A1(n15968), .A2(n12011), .ZN(n12777) );
  AOI22_X1 U13679 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U13680 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U13681 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12012) );
  NAND3_X1 U13682 ( .A1(n12014), .A2(n12013), .A3(n12012), .ZN(n12027) );
  INV_X1 U13683 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U13684 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12017) );
  NAND2_X1 U13685 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12016) );
  OAI211_X1 U13686 ( .C1(n12015), .C2(n12523), .A(n12017), .B(n12016), .ZN(
        n12022) );
  NAND2_X1 U13687 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12020) );
  NAND2_X1 U13688 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12019) );
  INV_X1 U13689 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12018) );
  NAND3_X1 U13690 ( .A1(n12020), .A2(n12019), .A3(n11384), .ZN(n12021) );
  NOR2_X1 U13691 ( .A1(n12022), .A2(n12021), .ZN(n12025) );
  AOI22_X1 U13692 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U13693 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15883), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12023) );
  NAND3_X1 U13694 ( .A1(n12025), .A2(n12024), .A3(n12023), .ZN(n12026) );
  INV_X1 U13695 ( .A(n12138), .ZN(n12776) );
  NAND2_X1 U13696 ( .A1(n12777), .A2(n12776), .ZN(n12028) );
  NAND2_X1 U13697 ( .A1(n12029), .A2(n12028), .ZN(n12161) );
  INV_X1 U13698 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12545) );
  INV_X1 U13699 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14751) );
  OAI22_X1 U13700 ( .A1(n12545), .A2(n19064), .B1(n12086), .B2(n14751), .ZN(
        n12030) );
  INV_X1 U13701 ( .A(n12030), .ZN(n12035) );
  AOI22_X1 U13702 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12084), .B1(
        n12185), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12034) );
  INV_X1 U13703 ( .A(n12085), .ZN(n12031) );
  AOI22_X1 U13704 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19027), .B1(
        n12078), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U13705 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12060) );
  AOI22_X1 U13706 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19152), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U13707 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19104), .B1(
        n19184), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U13708 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12059) );
  AOI22_X1 U13709 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U13710 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U13711 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12041) );
  NAND3_X1 U13712 ( .A1(n12043), .A2(n12042), .A3(n12041), .ZN(n12056) );
  INV_X1 U13713 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12046) );
  NAND2_X1 U13714 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12045) );
  NAND2_X1 U13715 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12044) );
  OAI211_X1 U13716 ( .C1(n15874), .C2(n12046), .A(n12045), .B(n12044), .ZN(
        n12050) );
  NAND2_X1 U13717 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U13718 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12047) );
  OAI211_X1 U13719 ( .C1(n12015), .C2(n12545), .A(n12048), .B(n12047), .ZN(
        n12049) );
  NOR2_X1 U13720 ( .A1(n12050), .A2(n12049), .ZN(n12054) );
  AOI22_X1 U13721 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12053) );
  INV_X1 U13722 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13861) );
  OAI22_X1 U13723 ( .A1(n14571), .A2(n13861), .B1(n14569), .B2(n14751), .ZN(
        n12051) );
  INV_X1 U13724 ( .A(n12051), .ZN(n12052) );
  NAND3_X1 U13725 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12055) );
  INV_X1 U13726 ( .A(n12463), .ZN(n12057) );
  NAND2_X1 U13727 ( .A1(n12057), .A2(n15968), .ZN(n12058) );
  INV_X1 U13728 ( .A(n12160), .ZN(n12061) );
  AOI22_X1 U13729 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13730 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U13731 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12062) );
  NAND3_X1 U13732 ( .A1(n12064), .A2(n12063), .A3(n12062), .ZN(n12077) );
  INV_X1 U13733 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U13734 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12066) );
  NAND2_X1 U13735 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12065) );
  OAI211_X1 U13736 ( .C1(n15874), .C2(n12067), .A(n12066), .B(n12065), .ZN(
        n12071) );
  INV_X1 U13737 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U13738 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12069) );
  NAND2_X1 U13739 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12068) );
  OAI211_X1 U13740 ( .C1(n12015), .C2(n12562), .A(n12069), .B(n12068), .ZN(
        n12070) );
  NOR2_X1 U13741 ( .A1(n12071), .A2(n12070), .ZN(n12075) );
  AOI22_X1 U13742 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U13743 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12073) );
  NAND2_X1 U13744 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12072) );
  NAND4_X1 U13745 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12076) );
  INV_X1 U13746 ( .A(n12466), .ZN(n12784) );
  AOI22_X1 U13747 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12078), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19061), .B1(
        n19027), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13749 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19152), .B1(
        n19116), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U13750 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19136), .B1(
        n12191), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13751 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n12084), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U13752 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14344), .B1(
        n12185), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19184), .B1(
        n19104), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U13754 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n12087), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U13755 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U13756 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U13757 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12093) );
  NAND3_X1 U13758 ( .A1(n12095), .A2(n12094), .A3(n12093), .ZN(n12109) );
  INV_X1 U13759 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U13760 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12097) );
  NAND2_X1 U13761 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12096) );
  OAI211_X1 U13762 ( .C1(n15874), .C2(n12098), .A(n12097), .B(n12096), .ZN(
        n12102) );
  INV_X1 U13763 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12583) );
  NAND2_X1 U13764 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U13765 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12099) );
  OAI211_X1 U13766 ( .C1(n12015), .C2(n12583), .A(n12100), .B(n12099), .ZN(
        n12101) );
  NOR2_X1 U13767 ( .A1(n12102), .A2(n12101), .ZN(n12107) );
  AOI22_X1 U13768 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12106) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12103) );
  INV_X1 U13770 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14815) );
  OAI22_X1 U13771 ( .A1(n12103), .A2(n14571), .B1(n14569), .B2(n14815), .ZN(
        n12104) );
  INV_X1 U13772 ( .A(n12104), .ZN(n12105) );
  NAND3_X1 U13773 ( .A1(n12107), .A2(n12106), .A3(n12105), .ZN(n12108) );
  INV_X1 U13774 ( .A(n12472), .ZN(n12110) );
  NAND2_X1 U13775 ( .A1(n12110), .A2(n15968), .ZN(n12111) );
  INV_X1 U13776 ( .A(n12114), .ZN(n12113) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n15870), .B1(
        n15875), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n15871), .B1(
        n15876), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U13779 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12117) );
  NAND2_X1 U13780 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12116) );
  NAND4_X1 U13781 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  NAND2_X1 U13782 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U13783 ( .A1(n15882), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U13784 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U13785 ( .A1(n15866), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12120) );
  NAND4_X1 U13786 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  NAND2_X1 U13787 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U13788 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U13789 ( .A1(n15865), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12128) );
  INV_X1 U13790 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12624) );
  NAND4_X1 U13791 ( .A1(n12130), .A2(n12129), .A3(n12128), .A4(n12127), .ZN(
        n12133) );
  INV_X1 U13792 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12131) );
  INV_X1 U13793 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19060) );
  OAI22_X1 U13794 ( .A1(n12131), .A2(n14571), .B1(n14569), .B2(n19060), .ZN(
        n12132) );
  NOR2_X1 U13795 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  INV_X1 U13796 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12136) );
  INV_X1 U13797 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13742) );
  NAND2_X1 U13798 ( .A1(n12136), .A2(n13742), .ZN(n12137) );
  MUX2_X1 U13799 ( .A(n12774), .B(n12137), .S(n15204), .Z(n12175) );
  XNOR2_X1 U13800 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U13801 ( .A1(n12387), .A2(n12337), .ZN(n12140) );
  NAND2_X1 U13802 ( .A1(n19179), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U13803 ( .A1(n12140), .A2(n12139), .ZN(n12144) );
  INV_X1 U13804 ( .A(n12144), .ZN(n12142) );
  XNOR2_X1 U13805 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12143) );
  INV_X1 U13806 ( .A(n12143), .ZN(n12141) );
  NAND2_X1 U13807 ( .A1(n12142), .A2(n12141), .ZN(n12145) );
  NAND2_X1 U13808 ( .A1(n12144), .A2(n12143), .ZN(n12147) );
  AND2_X1 U13809 ( .A1(n12145), .A2(n12147), .ZN(n12358) );
  NAND2_X1 U13810 ( .A1(n12402), .A2(n12358), .ZN(n12343) );
  NAND2_X1 U13811 ( .A1(n19160), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12146) );
  XNOR2_X1 U13812 ( .A(n13958), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12150) );
  XNOR2_X1 U13813 ( .A(n12149), .B(n12150), .ZN(n12359) );
  MUX2_X1 U13814 ( .A(n12463), .B(n12359), .S(n12402), .Z(n12334) );
  INV_X1 U13815 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12148) );
  MUX2_X1 U13816 ( .A(n12334), .B(n12148), .S(n15204), .Z(n12163) );
  NAND3_X1 U13817 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12332), .A3(
        n14020), .ZN(n12360) );
  MUX2_X1 U13818 ( .A(n12360), .B(n12466), .S(n11146), .Z(n12335) );
  INV_X1 U13819 ( .A(n12335), .ZN(n12153) );
  MUX2_X1 U13820 ( .A(n12153), .B(P2_EBX_REG_4__SCAN_IN), .S(n15204), .Z(
        n12159) );
  INV_X1 U13821 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18081) );
  MUX2_X1 U13822 ( .A(n12472), .B(n18081), .S(n15204), .Z(n12154) );
  INV_X1 U13823 ( .A(n12219), .ZN(n12157) );
  OR2_X1 U13824 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  NAND2_X1 U13825 ( .A1(n12157), .A2(n12156), .ZN(n18069) );
  INV_X1 U13826 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14548) );
  XNOR2_X1 U13827 ( .A(n12165), .B(n12159), .ZN(n18056) );
  INV_X1 U13828 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14544) );
  OR2_X1 U13829 ( .A1(n12164), .A2(n12163), .ZN(n12166) );
  NAND2_X1 U13830 ( .A1(n12166), .A2(n12165), .ZN(n15819) );
  NAND2_X1 U13831 ( .A1(n12167), .A2(n15819), .ZN(n14382) );
  INV_X1 U13832 ( .A(n12337), .ZN(n12170) );
  NAND2_X1 U13833 ( .A1(n12168), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12169) );
  NAND2_X1 U13834 ( .A1(n12170), .A2(n12169), .ZN(n12363) );
  INV_X1 U13835 ( .A(n12363), .ZN(n12339) );
  MUX2_X1 U13836 ( .A(n13535), .B(n12339), .S(n12402), .Z(n12388) );
  MUX2_X1 U13837 ( .A(n12388), .B(P2_EBX_REG_0__SCAN_IN), .S(n15204), .Z(
        n18030) );
  AND2_X1 U13838 ( .A1(n18030), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12173) );
  NAND3_X1 U13839 ( .A1(n15204), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U13840 ( .A1(n12175), .A2(n12171), .ZN(n18043) );
  INV_X1 U13841 ( .A(n18043), .ZN(n12172) );
  NOR2_X1 U13842 ( .A1(n12173), .A2(n12172), .ZN(n13521) );
  AND2_X1 U13843 ( .A1(n12173), .A2(n12172), .ZN(n13520) );
  NOR2_X1 U13844 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13520), .ZN(
        n13519) );
  NOR2_X1 U13845 ( .A1(n13521), .A2(n13519), .ZN(n13596) );
  XNOR2_X1 U13846 ( .A(n12175), .B(n12174), .ZN(n15838) );
  XNOR2_X1 U13847 ( .A(n15838), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13594) );
  INV_X1 U13848 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18508) );
  NOR2_X1 U13849 ( .A1(n15838), .A2(n18508), .ZN(n12176) );
  AOI21_X1 U13850 ( .B1(n13596), .B2(n13594), .A(n12176), .ZN(n14354) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14365) );
  AND2_X1 U13852 ( .A1(n18056), .A2(n14544), .ZN(n12178) );
  AOI21_X1 U13853 ( .B1(n14354), .B2(n14365), .A(n12178), .ZN(n12177) );
  NAND2_X1 U13854 ( .A1(n14382), .A2(n12177), .ZN(n12181) );
  INV_X1 U13855 ( .A(n14354), .ZN(n14383) );
  INV_X1 U13856 ( .A(n12178), .ZN(n12179) );
  NAND3_X1 U13857 ( .A1(n14383), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12179), .ZN(n12180) );
  OAI211_X1 U13858 ( .C1(n18056), .C2(n14544), .A(n12181), .B(n12180), .ZN(
        n14542) );
  NAND2_X1 U13859 ( .A1(n14541), .A2(n14542), .ZN(n12184) );
  NAND2_X1 U13860 ( .A1(n12182), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12183) );
  NAND2_X1 U13861 ( .A1(n12184), .A2(n12183), .ZN(n14611) );
  AOI22_X1 U13862 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12031), .B1(
        n10961), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U13863 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12084), .B1(
        n12185), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19027), .B1(
        n12078), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13865 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19061), .B1(
        n14344), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U13866 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12197) );
  AOI22_X1 U13867 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19104), .B1(
        n19184), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U13868 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19152), .B1(
        n12087), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19116), .B1(
        n12190), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U13870 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19136), .B1(
        n12191), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U13871 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12196) );
  AOI22_X1 U13872 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13873 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12200) );
  NAND2_X1 U13874 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U13875 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12198) );
  NAND4_X1 U13876 ( .A1(n12201), .A2(n12200), .A3(n12199), .A4(n12198), .ZN(
        n12213) );
  INV_X1 U13877 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12204) );
  NAND2_X1 U13878 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12203) );
  NAND2_X1 U13879 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12202) );
  OAI211_X1 U13880 ( .C1(n15874), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        n12208) );
  INV_X1 U13881 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U13882 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12206) );
  NAND2_X1 U13883 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12205) );
  OAI211_X1 U13884 ( .C1(n12015), .C2(n16017), .A(n12206), .B(n12205), .ZN(
        n12207) );
  NOR2_X1 U13885 ( .A1(n12208), .A2(n12207), .ZN(n12211) );
  AOI22_X1 U13886 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15883), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U13887 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12209) );
  NAND3_X1 U13888 ( .A1(n12211), .A2(n12210), .A3(n12209), .ZN(n12212) );
  INV_X1 U13889 ( .A(n12475), .ZN(n12214) );
  NAND2_X1 U13890 ( .A1(n12214), .A2(n15968), .ZN(n12215) );
  NAND2_X1 U13891 ( .A1(n12791), .A2(n15212), .ZN(n12220) );
  INV_X1 U13892 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12217) );
  MUX2_X1 U13893 ( .A(n12475), .B(n12217), .S(n15204), .Z(n12218) );
  OAI21_X1 U13894 ( .B1(n12219), .B2(n12218), .A(n15210), .ZN(n18082) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U13896 ( .A1(n14611), .A2(n14610), .ZN(n12224) );
  NAND2_X1 U13897 ( .A1(n12222), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12223) );
  MUX2_X1 U13898 ( .A(n15212), .B(P2_EBX_REG_7__SCAN_IN), .S(n15204), .Z(
        n12226) );
  INV_X1 U13899 ( .A(n12226), .ZN(n12225) );
  XNOR2_X1 U13900 ( .A(n15210), .B(n12225), .ZN(n18094) );
  AND2_X1 U13901 ( .A1(n18094), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14725) );
  NAND2_X1 U13902 ( .A1(n15204), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12227) );
  OR2_X1 U13903 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  NAND2_X1 U13904 ( .A1(n12233), .A2(n12229), .ZN(n18106) );
  INV_X1 U13905 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12230) );
  NOR2_X1 U13906 ( .A1(n12231), .A2(n12230), .ZN(n16980) );
  NAND2_X1 U13907 ( .A1(n16980), .A2(n14724), .ZN(n12232) );
  XNOR2_X1 U13908 ( .A(n12233), .B(n11043), .ZN(n18121) );
  NAND2_X1 U13909 ( .A1(n18121), .A2(n11337), .ZN(n12246) );
  INV_X1 U13910 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16668) );
  NAND2_X1 U13911 ( .A1(n12246), .A2(n16668), .ZN(n16429) );
  INV_X1 U13912 ( .A(n12240), .ZN(n12237) );
  NAND2_X1 U13913 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  NAND2_X1 U13914 ( .A1(n12237), .A2(n12236), .ZN(n18130) );
  INV_X1 U13915 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16995) );
  OAI21_X1 U13916 ( .B1(n18130), .B2(n15212), .A(n16995), .ZN(n16987) );
  XNOR2_X1 U13917 ( .A(n12237), .B(n11386), .ZN(n18143) );
  AOI21_X1 U13918 ( .B1(n18143), .B2(n11337), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16422) );
  NAND2_X1 U13919 ( .A1(n15204), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12241) );
  OR2_X1 U13920 ( .A1(n11392), .A2(n12241), .ZN(n12242) );
  NAND2_X1 U13921 ( .A1(n12268), .A2(n12242), .ZN(n18156) );
  INV_X1 U13922 ( .A(n18156), .ZN(n12244) );
  INV_X1 U13923 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12702) );
  NOR2_X1 U13924 ( .A1(n15212), .A2(n12702), .ZN(n12243) );
  NAND2_X1 U13925 ( .A1(n12244), .A2(n12243), .ZN(n16998) );
  INV_X1 U13926 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16659) );
  NOR2_X1 U13927 ( .A1(n15212), .A2(n16659), .ZN(n12245) );
  NAND2_X1 U13928 ( .A1(n18143), .A2(n12245), .ZN(n16420) );
  OR2_X1 U13929 ( .A1(n12246), .A2(n16668), .ZN(n16989) );
  INV_X1 U13930 ( .A(n18130), .ZN(n12248) );
  NOR2_X1 U13931 ( .A1(n15212), .A2(n16995), .ZN(n12247) );
  NAND2_X1 U13932 ( .A1(n12248), .A2(n12247), .ZN(n16986) );
  AND4_X1 U13933 ( .A1(n16998), .A2(n16420), .A3(n16989), .A4(n16986), .ZN(
        n12249) );
  AND2_X1 U13934 ( .A1(n15204), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12266) );
  AND2_X1 U13935 ( .A1(n15204), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12263) );
  NAND2_X1 U13936 ( .A1(n15204), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U13937 ( .A1(n15204), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12270) );
  AND2_X1 U13938 ( .A1(n15204), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12254) );
  NAND2_X1 U13939 ( .A1(n15204), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U13940 ( .A1(n15204), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12278) );
  AND2_X1 U13941 ( .A1(n15204), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12298) );
  INV_X1 U13942 ( .A(n12298), .ZN(n12250) );
  XNOR2_X1 U13943 ( .A(n12299), .B(n12250), .ZN(n18270) );
  AOI21_X1 U13944 ( .B1(n18270), .B2(n11337), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16328) );
  INV_X1 U13945 ( .A(n12251), .ZN(n12252) );
  XNOR2_X1 U13946 ( .A(n12256), .B(n12252), .ZN(n18239) );
  NAND2_X1 U13947 ( .A1(n18239), .A2(n11337), .ZN(n12253) );
  INV_X1 U13948 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16576) );
  NAND2_X1 U13949 ( .A1(n12253), .A2(n16576), .ZN(n16350) );
  AND2_X1 U13950 ( .A1(n12255), .A2(n12254), .ZN(n12257) );
  OR2_X1 U13951 ( .A1(n12257), .A2(n12256), .ZN(n18232) );
  INV_X1 U13952 ( .A(n18232), .ZN(n12258) );
  NAND2_X1 U13953 ( .A1(n12258), .A2(n11337), .ZN(n16363) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16588) );
  NAND2_X1 U13955 ( .A1(n16363), .A2(n16588), .ZN(n12259) );
  NOR2_X1 U13956 ( .A1(n12260), .A2(n12261), .ZN(n12262) );
  OR2_X1 U13957 ( .A1(n12272), .A2(n12262), .ZN(n18194) );
  NOR2_X1 U13958 ( .A1(n18194), .A2(n15212), .ZN(n12289) );
  OR2_X1 U13959 ( .A1(n12289), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16405) );
  AND2_X1 U13960 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  OR2_X1 U13961 ( .A1(n12265), .A2(n12260), .ZN(n18182) );
  NOR2_X1 U13962 ( .A1(n18182), .A2(n15212), .ZN(n12290) );
  OR2_X1 U13963 ( .A1(n12290), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16409) );
  INV_X1 U13964 ( .A(n12266), .ZN(n12267) );
  XNOR2_X1 U13965 ( .A(n12268), .B(n12267), .ZN(n18165) );
  NAND2_X1 U13966 ( .A1(n18165), .A2(n11337), .ZN(n12269) );
  INV_X1 U13967 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18457) );
  NAND2_X1 U13968 ( .A1(n12269), .A2(n18457), .ZN(n16638) );
  OAI21_X1 U13969 ( .B1(n18156), .B2(n15212), .A(n12702), .ZN(n16999) );
  NAND4_X1 U13970 ( .A1(n16405), .A2(n16409), .A3(n16638), .A4(n16999), .ZN(
        n16314) );
  INV_X1 U13971 ( .A(n12270), .ZN(n12271) );
  XNOR2_X1 U13972 ( .A(n12272), .B(n12271), .ZN(n18207) );
  NAND2_X1 U13973 ( .A1(n18207), .A2(n11337), .ZN(n12273) );
  INV_X1 U13974 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16622) );
  NAND2_X1 U13975 ( .A1(n12273), .A2(n16622), .ZN(n12275) );
  NOR2_X1 U13976 ( .A1(n15212), .A2(n16622), .ZN(n12274) );
  NAND2_X1 U13977 ( .A1(n18207), .A2(n12274), .ZN(n16375) );
  NAND2_X1 U13978 ( .A1(n12275), .A2(n16375), .ZN(n16318) );
  NOR2_X1 U13979 ( .A1(n16314), .A2(n16318), .ZN(n12282) );
  XNOR2_X1 U13980 ( .A(n12276), .B(n11042), .ZN(n18217) );
  NAND2_X1 U13981 ( .A1(n18217), .A2(n11337), .ZN(n12277) );
  INV_X1 U13982 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16608) );
  NAND2_X1 U13983 ( .A1(n12277), .A2(n16608), .ZN(n16377) );
  OR2_X1 U13984 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  NAND2_X1 U13985 ( .A1(n12299), .A2(n12280), .ZN(n18262) );
  INV_X1 U13986 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16558) );
  NAND2_X1 U13987 ( .A1(n16324), .A2(n16558), .ZN(n12281) );
  NAND4_X1 U13988 ( .A1(n16322), .A2(n12282), .A3(n16377), .A4(n12281), .ZN(
        n12283) );
  NOR2_X1 U13989 ( .A1(n16328), .A2(n12283), .ZN(n12284) );
  NAND2_X1 U13990 ( .A1(n12285), .A2(n12284), .ZN(n12297) );
  INV_X1 U13991 ( .A(n16363), .ZN(n12286) );
  NAND2_X1 U13992 ( .A1(n12286), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16321) );
  NOR2_X1 U13993 ( .A1(n15212), .A2(n16608), .ZN(n12287) );
  NAND2_X1 U13994 ( .A1(n18217), .A2(n12287), .ZN(n16376) );
  NOR2_X1 U13995 ( .A1(n15212), .A2(n18457), .ZN(n12288) );
  NAND2_X1 U13996 ( .A1(n18165), .A2(n12288), .ZN(n16407) );
  NAND2_X1 U13997 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12289), .ZN(
        n16404) );
  NAND2_X1 U13998 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n12290), .ZN(
        n16408) );
  AND2_X1 U13999 ( .A1(n16404), .A2(n16408), .ZN(n12291) );
  AND3_X1 U14000 ( .A1(n16321), .A2(n16320), .A3(n16316), .ZN(n12293) );
  NOR2_X1 U14001 ( .A1(n15212), .A2(n16576), .ZN(n12292) );
  NAND2_X1 U14002 ( .A1(n18239), .A2(n12292), .ZN(n16349) );
  OAI211_X1 U14003 ( .C1(n16324), .C2(n16558), .A(n12293), .B(n16349), .ZN(
        n12295) );
  INV_X1 U14004 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16537) );
  NOR2_X1 U14005 ( .A1(n15212), .A2(n16537), .ZN(n12294) );
  NOR2_X1 U14006 ( .A1(n12295), .A2(n16329), .ZN(n12296) );
  AND2_X1 U14007 ( .A1(n15204), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12301) );
  INV_X1 U14008 ( .A(n12301), .ZN(n12300) );
  XNOR2_X1 U14009 ( .A(n12302), .B(n12300), .ZN(n18281) );
  NAND2_X1 U14010 ( .A1(n18281), .A2(n11337), .ZN(n16525) );
  AND2_X1 U14011 ( .A1(n15204), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12303) );
  AND2_X1 U14012 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  OR2_X1 U14013 ( .A1(n12305), .A2(n12313), .ZN(n18296) );
  AOI21_X1 U14014 ( .B1(n12307), .B2(n11337), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16301) );
  INV_X1 U14015 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16515) );
  NOR2_X1 U14016 ( .A1(n15212), .A2(n16515), .ZN(n12306) );
  NAND2_X1 U14017 ( .A1(n12307), .A2(n12306), .ZN(n16302) );
  NAND2_X1 U14018 ( .A1(n15204), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12312) );
  XNOR2_X1 U14019 ( .A(n12313), .B(n11212), .ZN(n18307) );
  NAND2_X1 U14020 ( .A1(n18307), .A2(n11337), .ZN(n16292) );
  NAND2_X1 U14021 ( .A1(n12308), .A2(n16292), .ZN(n12311) );
  AND2_X1 U14022 ( .A1(n15204), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12324) );
  AND2_X1 U14023 ( .A1(n15204), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12316) );
  XOR2_X1 U14024 ( .A(n12324), .B(n12325), .Z(n18328) );
  INV_X1 U14025 ( .A(n18328), .ZN(n12314) );
  NOR2_X1 U14026 ( .A1(n12314), .A2(n15212), .ZN(n12315) );
  NAND3_X1 U14027 ( .A1(n18328), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11337), .ZN(n12323) );
  OAI21_X1 U14028 ( .B1(n12315), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12323), .ZN(n16265) );
  INV_X1 U14029 ( .A(n12316), .ZN(n12317) );
  XNOR2_X1 U14030 ( .A(n12318), .B(n12317), .ZN(n18317) );
  INV_X1 U14031 ( .A(n12321), .ZN(n12322) );
  INV_X1 U14032 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16497) );
  NAND2_X1 U14033 ( .A1(n12323), .A2(n16280), .ZN(n15197) );
  NAND2_X1 U14034 ( .A1(n15204), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12326) );
  NOR2_X1 U14035 ( .A1(n12327), .A2(n12326), .ZN(n12328) );
  NAND2_X1 U14036 ( .A1(n12329), .A2(n16242), .ZN(n12330) );
  XNOR2_X1 U14037 ( .A(n12330), .B(n15190), .ZN(n16262) );
  INV_X1 U14038 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16717) );
  NOR2_X1 U14039 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16717), .ZN(
        n12331) );
  NOR2_X1 U14040 ( .A1(n12360), .A2(n12402), .ZN(n12333) );
  OR2_X1 U14041 ( .A1(n12391), .A2(n12333), .ZN(n12350) );
  NAND2_X1 U14042 ( .A1(n12335), .A2(n12334), .ZN(n12390) );
  INV_X1 U14043 ( .A(n12358), .ZN(n12342) );
  NAND2_X1 U14044 ( .A1(n12339), .A2(n12387), .ZN(n12336) );
  NAND2_X1 U14045 ( .A1(n11146), .A2(n12336), .ZN(n12341) );
  XNOR2_X1 U14046 ( .A(n12387), .B(n12337), .ZN(n12361) );
  INV_X1 U14047 ( .A(n12361), .ZN(n12338) );
  OAI211_X1 U14048 ( .C1(n16011), .C2(n12339), .A(n12379), .B(n12338), .ZN(
        n12340) );
  OAI211_X1 U14049 ( .C1(n12413), .C2(n12342), .A(n12341), .B(n12340), .ZN(
        n12347) );
  OAI21_X1 U14050 ( .B1(n13715), .B2(n15968), .A(n12342), .ZN(n12344) );
  NAND2_X1 U14051 ( .A1(n12344), .A2(n12343), .ZN(n12346) );
  INV_X1 U14052 ( .A(n12359), .ZN(n12345) );
  AOI21_X1 U14053 ( .B1(n12347), .B2(n12346), .A(n12345), .ZN(n12348) );
  AOI21_X1 U14054 ( .B1(n12390), .B2(n12402), .A(n12348), .ZN(n12349) );
  NOR2_X1 U14055 ( .A1(n12350), .A2(n12349), .ZN(n12351) );
  MUX2_X1 U14056 ( .A(n14020), .B(n12351), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12355) );
  AND2_X1 U14057 ( .A1(n12391), .A2(n13715), .ZN(n12352) );
  NAND2_X1 U14058 ( .A1(n14335), .A2(n16011), .ZN(n13713) );
  NAND2_X1 U14059 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18527) );
  INV_X1 U14060 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21682) );
  NOR2_X1 U14061 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n16709) );
  INV_X1 U14062 ( .A(n16709), .ZN(n21679) );
  NAND2_X1 U14063 ( .A1(n21685), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21666) );
  INV_X2 U14064 ( .A(n21666), .ZN(n17128) );
  OAI21_X1 U14065 ( .B1(n21682), .B2(n21679), .A(n17125), .ZN(n21669) );
  NAND2_X1 U14066 ( .A1(n18527), .A2(n21669), .ZN(n14028) );
  INV_X1 U14067 ( .A(n14028), .ZN(n14009) );
  NAND2_X1 U14068 ( .A1(n12353), .A2(n14009), .ZN(n12399) );
  OAI21_X1 U14069 ( .B1(n12355), .B2(n19597), .A(n12354), .ZN(n12356) );
  INV_X1 U14070 ( .A(n12356), .ZN(n12357) );
  NAND2_X1 U14071 ( .A1(n12357), .A2(n13713), .ZN(n12398) );
  NAND3_X1 U14072 ( .A1(n12360), .A2(n12359), .A3(n12358), .ZN(n12364) );
  NOR2_X1 U14073 ( .A1(n12364), .A2(n12361), .ZN(n12362) );
  OR2_X1 U14074 ( .A1(n12391), .A2(n12362), .ZN(n14014) );
  OAI21_X1 U14075 ( .B1(n12364), .B2(n12363), .A(n16714), .ZN(n12365) );
  OR2_X1 U14076 ( .A1(n14014), .A2(n12365), .ZN(n12371) );
  NAND2_X1 U14077 ( .A1(n12367), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U14078 ( .A1(n12368), .A2(n14020), .ZN(n13548) );
  INV_X1 U14079 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12369) );
  OAI21_X1 U14080 ( .B1(n12126), .B2(n13548), .A(n12369), .ZN(n12370) );
  NAND2_X1 U14081 ( .A1(n12370), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17044) );
  NAND2_X1 U14082 ( .A1(n12401), .A2(n16011), .ZN(n12372) );
  NOR2_X1 U14083 ( .A1(n18520), .A2(n12372), .ZN(n12396) );
  MUX2_X1 U14084 ( .A(n14030), .B(n12353), .S(n15968), .Z(n12373) );
  NAND2_X1 U14085 ( .A1(n12373), .A2(n18527), .ZN(n12394) );
  OR2_X1 U14086 ( .A1(n12374), .A2(n14028), .ZN(n12375) );
  OR2_X1 U14087 ( .A1(n14014), .A2(n12375), .ZN(n12385) );
  NAND2_X1 U14088 ( .A1(n13750), .A2(n12354), .ZN(n12377) );
  NAND2_X1 U14089 ( .A1(n13711), .A2(n12378), .ZN(n12384) );
  OR2_X1 U14090 ( .A1(n11868), .A2(n16011), .ZN(n12405) );
  AND3_X1 U14091 ( .A1(n12382), .A2(n12420), .A3(n12381), .ZN(n12383) );
  AND2_X1 U14092 ( .A1(n15968), .A2(n19597), .ZN(n14029) );
  OAI21_X1 U14093 ( .B1(n12380), .B2(n13749), .A(n14029), .ZN(n12410) );
  AND2_X1 U14094 ( .A1(n12385), .A2(n12404), .ZN(n13544) );
  AOI21_X1 U14095 ( .B1(n12388), .B2(n12387), .A(n12386), .ZN(n12389) );
  NOR2_X1 U14096 ( .A1(n12390), .A2(n12389), .ZN(n12392) );
  OR2_X1 U14097 ( .A1(n12392), .A2(n12391), .ZN(n13999) );
  INV_X1 U14098 ( .A(n13999), .ZN(n12393) );
  AND2_X1 U14099 ( .A1(n12401), .A2(n14029), .ZN(n14000) );
  NAND2_X1 U14100 ( .A1(n12393), .A2(n14000), .ZN(n13522) );
  OAI211_X1 U14101 ( .C1(n14014), .C2(n12394), .A(n13544), .B(n13522), .ZN(
        n12395) );
  NOR2_X1 U14102 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  OAI211_X1 U14103 ( .C1(n13713), .C2(n12399), .A(n12398), .B(n12397), .ZN(
        n12400) );
  INV_X1 U14104 ( .A(n12401), .ZN(n12403) );
  OR2_X1 U14105 ( .A1(n12403), .A2(n12402), .ZN(n13523) );
  INV_X1 U14106 ( .A(n13523), .ZN(n13998) );
  INV_X1 U14107 ( .A(n12404), .ZN(n12406) );
  NAND2_X1 U14108 ( .A1(n12815), .A2(n14005), .ZN(n18495) );
  INV_X1 U14109 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18435) );
  INV_X1 U14110 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18418) );
  OAI21_X1 U14111 ( .B1(n18435), .B2(n18418), .A(n18508), .ZN(n18488) );
  INV_X1 U14112 ( .A(n12815), .ZN(n12408) );
  NAND2_X1 U14113 ( .A1(n19164), .A2(n19183), .ZN(n13500) );
  NAND2_X1 U14114 ( .A1(n19200), .A2(n12407), .ZN(n18240) );
  INV_X1 U14115 ( .A(n18240), .ZN(n18072) );
  INV_X1 U14116 ( .A(n18072), .ZN(n18475) );
  NAND2_X1 U14117 ( .A1(n12408), .A2(n18475), .ZN(n18509) );
  OAI21_X1 U14118 ( .B1(n18495), .B2(n18488), .A(n18509), .ZN(n14364) );
  INV_X1 U14119 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18474) );
  NAND4_X1 U14120 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14616) );
  NOR3_X1 U14121 ( .A1(n12230), .A2(n18474), .A3(n14616), .ZN(n12765) );
  NOR2_X1 U14122 ( .A1(n18495), .A2(n12765), .ZN(n12409) );
  NOR2_X1 U14123 ( .A1(n14364), .A2(n12409), .ZN(n16555) );
  NAND2_X1 U14124 ( .A1(n11032), .A2(n16011), .ZN(n13969) );
  NAND2_X1 U14125 ( .A1(n13969), .A2(n12410), .ZN(n12418) );
  INV_X1 U14126 ( .A(n12411), .ZN(n13512) );
  AOI22_X1 U14127 ( .A1(n13512), .A2(n12412), .B1(n19597), .B2(n12353), .ZN(
        n12415) );
  INV_X1 U14128 ( .A(n12413), .ZN(n12414) );
  NAND3_X1 U14129 ( .A1(n12416), .A2(n12415), .A3(n13744), .ZN(n12417) );
  AOI21_X1 U14130 ( .B1(n12418), .B2(n19410), .A(n12417), .ZN(n12419) );
  OAI21_X1 U14131 ( .B1(n12421), .B2(n12420), .A(n12419), .ZN(n13989) );
  INV_X1 U14132 ( .A(n13989), .ZN(n13949) );
  INV_X1 U14133 ( .A(n12422), .ZN(n13950) );
  NAND2_X1 U14134 ( .A1(n13949), .A2(n13950), .ZN(n12423) );
  NAND2_X1 U14135 ( .A1(n12815), .A2(n12423), .ZN(n18489) );
  INV_X1 U14136 ( .A(n18489), .ZN(n12762) );
  NAND2_X1 U14137 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18428) );
  NOR2_X1 U14138 ( .A1(n18508), .A2(n18428), .ZN(n18486) );
  NAND2_X1 U14139 ( .A1(n12765), .A2(n18486), .ZN(n16549) );
  NAND2_X1 U14140 ( .A1(n12762), .A2(n16549), .ZN(n12424) );
  NAND2_X1 U14141 ( .A1(n16555), .A2(n12424), .ZN(n18459) );
  AND2_X1 U14142 ( .A1(n18495), .A2(n18489), .ZN(n18422) );
  OR2_X1 U14143 ( .A1(n18459), .A2(n18460), .ZN(n16653) );
  NAND2_X1 U14144 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16563) );
  NOR2_X1 U14145 ( .A1(n16563), .A2(n16558), .ZN(n12428) );
  INV_X1 U14146 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16629) );
  NAND2_X1 U14147 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16642) );
  INV_X1 U14148 ( .A(n16642), .ZN(n12427) );
  NAND3_X1 U14149 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18461) );
  INV_X1 U14150 ( .A(n18461), .ZN(n12425) );
  AND2_X1 U14151 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n12425), .ZN(
        n12426) );
  NAND2_X1 U14152 ( .A1(n12427), .A2(n12426), .ZN(n16626) );
  NOR2_X1 U14153 ( .A1(n16629), .A2(n16626), .ZN(n16602) );
  AND3_X1 U14154 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16602), .ZN(n16556) );
  AND2_X1 U14155 ( .A1(n12428), .A2(n16556), .ZN(n16536) );
  NAND2_X1 U14156 ( .A1(n16536), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12811) );
  OR2_X1 U14157 ( .A1(n18459), .A2(n12811), .ZN(n12429) );
  NAND2_X1 U14158 ( .A1(n16653), .A2(n12429), .ZN(n16514) );
  AND2_X1 U14159 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12761) );
  OAI21_X1 U14160 ( .B1(n18422), .B2(n12761), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12430) );
  INV_X1 U14161 ( .A(n12430), .ZN(n12431) );
  NAND2_X1 U14162 ( .A1(n16514), .A2(n12431), .ZN(n16504) );
  NAND2_X1 U14163 ( .A1(n16504), .A2(n16653), .ZN(n16498) );
  NAND2_X1 U14164 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U14165 ( .A1(n16653), .A2(n12813), .ZN(n12432) );
  NAND2_X1 U14166 ( .A1(n16498), .A2(n12432), .ZN(n16455) );
  INV_X1 U14167 ( .A(n12433), .ZN(n13499) );
  NAND2_X1 U14168 ( .A1(n13711), .A2(n13499), .ZN(n14012) );
  NAND2_X1 U14169 ( .A1(n14012), .A2(n16011), .ZN(n12435) );
  NAND2_X1 U14170 ( .A1(n12434), .A2(n13967), .ZN(n13956) );
  NAND2_X1 U14171 ( .A1(n12435), .A2(n13956), .ZN(n12436) );
  NAND2_X1 U14172 ( .A1(n12815), .A2(n12436), .ZN(n18490) );
  NOR2_X1 U14173 ( .A1(n11858), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U14174 ( .A1(n12458), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12439) );
  OAI21_X1 U14175 ( .B1(n15269), .B2(n11901), .A(n12439), .ZN(n12451) );
  INV_X1 U14176 ( .A(n12451), .ZN(n12447) );
  INV_X1 U14177 ( .A(n12467), .ZN(n12647) );
  OR2_X1 U14178 ( .A1(n12647), .A2(n13750), .ZN(n12454) );
  MUX2_X1 U14179 ( .A(n11858), .B(n19146), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12443) );
  NOR2_X1 U14180 ( .A1(n12440), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U14181 ( .A1(n12635), .A2(n13535), .ZN(n12442) );
  NAND3_X1 U14182 ( .A1(n12454), .A2(n12443), .A3(n12442), .ZN(n13748) );
  INV_X1 U14183 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U14184 ( .A1(n12440), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12444) );
  OAI211_X1 U14185 ( .C1(n11858), .C2(n13754), .A(n12444), .B(n19183), .ZN(
        n12445) );
  INV_X1 U14186 ( .A(n12445), .ZN(n12446) );
  INV_X1 U14187 ( .A(n12635), .ZN(n12478) );
  OR2_X1 U14188 ( .A1(n12774), .A2(n12478), .ZN(n12450) );
  NAND2_X1 U14189 ( .A1(n13750), .A2(n11858), .ZN(n12448) );
  MUX2_X1 U14190 ( .A(n12448), .B(n19179), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12449) );
  NAND2_X1 U14191 ( .A1(n13809), .A2(n13808), .ZN(n13807) );
  NAND2_X1 U14192 ( .A1(n12635), .A2(n12138), .ZN(n12453) );
  OAI211_X1 U14193 ( .C1(n19183), .C2(n19160), .A(n12454), .B(n12453), .ZN(
        n12455) );
  AND3_X1 U14194 ( .A1(n13807), .A2(n12456), .A3(n12455), .ZN(n12457) );
  INV_X1 U14195 ( .A(n12458), .ZN(n12646) );
  INV_X2 U14196 ( .A(n12646), .ZN(n12595) );
  AOI22_X1 U14197 ( .A1(n12595), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12459) );
  OAI21_X1 U14198 ( .B1(n15269), .B2(n11889), .A(n12459), .ZN(n14081) );
  AOI22_X1 U14199 ( .A1(n12635), .A2(n12463), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U14200 ( .A1(n12595), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12464) );
  OAI211_X1 U14201 ( .C1(n14356), .C2(n15269), .A(n12465), .B(n12464), .ZN(
        n14163) );
  NAND2_X1 U14202 ( .A1(n12635), .A2(n12466), .ZN(n12469) );
  AOI22_X1 U14203 ( .A1(n12595), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12468) );
  AND2_X1 U14204 ( .A1(n12469), .A2(n12468), .ZN(n12471) );
  NAND2_X1 U14205 ( .A1(n12648), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U14206 ( .A1(n12648), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12635), 
        .B2(n12472), .ZN(n12474) );
  AOI22_X1 U14207 ( .A1(n12595), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12473) );
  NAND2_X1 U14208 ( .A1(n12474), .A2(n12473), .ZN(n14546) );
  NAND2_X1 U14209 ( .A1(n12475), .A2(n12635), .ZN(n12476) );
  INV_X1 U14210 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17088) );
  OAI22_X1 U14211 ( .A1(n12646), .A2(n17088), .B1(n12647), .B2(n12221), .ZN(
        n12477) );
  AOI21_X1 U14212 ( .B1(n12648), .B2(P2_REIP_REG_6__SCAN_IN), .A(n12477), .ZN(
        n13799) );
  INV_X1 U14213 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U14214 ( .A1(n12595), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12479) );
  OAI21_X1 U14215 ( .B1(n15269), .B2(n18096), .A(n12479), .ZN(n13821) );
  AOI22_X1 U14216 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U14217 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U14218 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12480) );
  NAND3_X1 U14219 ( .A1(n12482), .A2(n12481), .A3(n12480), .ZN(n12495) );
  NAND2_X1 U14220 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12484) );
  NAND2_X1 U14221 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12483) );
  OAI211_X1 U14222 ( .C1(n15874), .C2(n12485), .A(n12484), .B(n12483), .ZN(
        n12489) );
  NAND2_X1 U14223 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12487) );
  NAND2_X1 U14224 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12486) );
  OAI211_X1 U14225 ( .C1(n12015), .C2(n14509), .A(n12487), .B(n12486), .ZN(
        n12488) );
  NOR2_X1 U14226 ( .A1(n12489), .A2(n12488), .ZN(n12493) );
  AOI22_X1 U14227 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U14228 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12491) );
  NAND2_X1 U14229 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12490) );
  NAND4_X1 U14230 ( .A1(n12493), .A2(n12492), .A3(n12491), .A4(n12490), .ZN(
        n12494) );
  NAND2_X1 U14231 ( .A1(n12635), .A2(n14109), .ZN(n12497) );
  AOI22_X1 U14232 ( .A1(n12595), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12496) );
  AND2_X1 U14233 ( .A1(n12497), .A2(n12496), .ZN(n12499) );
  NAND2_X1 U14234 ( .A1(n12648), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12498) );
  INV_X1 U14235 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U14236 ( .A1(n12595), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12467), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U14237 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U14238 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U14239 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12500) );
  NAND3_X1 U14240 ( .A1(n12502), .A2(n12501), .A3(n12500), .ZN(n12516) );
  NAND2_X1 U14241 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12504) );
  NAND2_X1 U14242 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12503) );
  OAI211_X1 U14243 ( .C1(n15874), .C2(n12505), .A(n12504), .B(n12503), .ZN(
        n12509) );
  NAND2_X1 U14244 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12507) );
  NAND2_X1 U14245 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12506) );
  OAI211_X1 U14246 ( .C1(n12015), .C2(n14562), .A(n12507), .B(n12506), .ZN(
        n12508) );
  NOR2_X1 U14247 ( .A1(n12509), .A2(n12508), .ZN(n12514) );
  AOI22_X1 U14248 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12513) );
  OAI22_X1 U14249 ( .A1(n14571), .A2(n12510), .B1(n14569), .B2(n14565), .ZN(
        n12511) );
  INV_X1 U14250 ( .A(n12511), .ZN(n12512) );
  NAND3_X1 U14251 ( .A1(n12514), .A2(n12513), .A3(n12512), .ZN(n12515) );
  NAND2_X1 U14252 ( .A1(n12635), .A2(n14156), .ZN(n12517) );
  OAI211_X1 U14253 ( .C1(n15269), .C2(n12694), .A(n12518), .B(n12517), .ZN(
        n13836) );
  AOI22_X1 U14254 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15884), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U14255 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12520) );
  AOI22_X1 U14256 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15876), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12519) );
  AND2_X1 U14257 ( .A1(n12520), .A2(n12519), .ZN(n12527) );
  NAND2_X1 U14258 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12522) );
  NAND2_X1 U14259 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12521) );
  OAI211_X1 U14260 ( .C1(n15874), .C2(n12523), .A(n12522), .B(n12521), .ZN(
        n12524) );
  INV_X1 U14261 ( .A(n12524), .ZN(n12526) );
  AOI22_X1 U14262 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12525) );
  NAND4_X1 U14263 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n12534) );
  AOI22_X1 U14264 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12609), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U14265 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U14266 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12530) );
  NAND2_X1 U14267 ( .A1(n15865), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12529) );
  NAND4_X1 U14268 ( .A1(n12532), .A2(n12531), .A3(n12530), .A4(n12529), .ZN(
        n12533) );
  NOR2_X1 U14269 ( .A1(n12534), .A2(n12533), .ZN(n14241) );
  INV_X1 U14270 ( .A(n14241), .ZN(n12535) );
  NAND2_X1 U14271 ( .A1(n12635), .A2(n12535), .ZN(n12537) );
  AOI22_X1 U14272 ( .A1(n12595), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12536) );
  AND2_X1 U14273 ( .A1(n12537), .A2(n12536), .ZN(n12539) );
  NAND2_X1 U14274 ( .A1(n12648), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12538) );
  INV_X1 U14275 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U14276 ( .A1(n12595), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U14277 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U14278 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U14279 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12540) );
  NAND3_X1 U14280 ( .A1(n12542), .A2(n12541), .A3(n12540), .ZN(n12555) );
  NAND2_X1 U14281 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12544) );
  NAND2_X1 U14282 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12543) );
  OAI211_X1 U14283 ( .C1(n15874), .C2(n12545), .A(n12544), .B(n12543), .ZN(
        n12549) );
  NAND2_X1 U14284 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U14285 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12546) );
  OAI211_X1 U14286 ( .C1(n12015), .C2(n14751), .A(n12547), .B(n12546), .ZN(
        n12548) );
  NOR2_X1 U14287 ( .A1(n12549), .A2(n12548), .ZN(n12553) );
  AOI22_X1 U14288 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U14289 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12551) );
  NAND2_X1 U14290 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12550) );
  NAND4_X1 U14291 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  NAND2_X1 U14292 ( .A1(n12635), .A2(n14195), .ZN(n12556) );
  OAI211_X1 U14293 ( .C1(n15269), .C2(n16417), .A(n12557), .B(n12556), .ZN(
        n13948) );
  AOI22_X1 U14294 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15883), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U14295 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12559) );
  AOI22_X1 U14296 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15875), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12558) );
  AND2_X1 U14297 ( .A1(n12559), .A2(n12558), .ZN(n12566) );
  NAND2_X1 U14298 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U14299 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12560) );
  OAI211_X1 U14300 ( .C1(n15874), .C2(n12562), .A(n12561), .B(n12560), .ZN(
        n12563) );
  INV_X1 U14301 ( .A(n12563), .ZN(n12565) );
  AOI22_X1 U14302 ( .A1(n15882), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12092), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12564) );
  NAND4_X1 U14303 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n12573) );
  AOI22_X1 U14304 ( .A1(n15865), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12609), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U14305 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U14306 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12569) );
  NAND2_X1 U14307 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12568) );
  NAND4_X1 U14308 ( .A1(n12571), .A2(n12570), .A3(n12569), .A4(n12568), .ZN(
        n12572) );
  NAND2_X1 U14309 ( .A1(n12635), .A2(n11389), .ZN(n12575) );
  AOI22_X1 U14310 ( .A1(n12595), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12574) );
  AND2_X1 U14311 ( .A1(n12575), .A2(n12574), .ZN(n12577) );
  NAND2_X1 U14312 ( .A1(n12648), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U14313 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U14314 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U14315 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12578) );
  NAND3_X1 U14316 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(n12594) );
  NAND2_X1 U14317 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U14318 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12581) );
  OAI211_X1 U14319 ( .C1(n15874), .C2(n12583), .A(n12582), .B(n12581), .ZN(
        n12587) );
  NAND2_X1 U14320 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12585) );
  NAND2_X1 U14321 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12584) );
  OAI211_X1 U14322 ( .C1(n12015), .C2(n14815), .A(n12585), .B(n12584), .ZN(
        n12586) );
  NOR2_X1 U14323 ( .A1(n12587), .A2(n12586), .ZN(n12592) );
  AOI22_X1 U14324 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12591) );
  INV_X1 U14325 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12588) );
  INV_X1 U14326 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14818) );
  OAI22_X1 U14327 ( .A1(n12588), .A2(n14571), .B1(n14569), .B2(n14818), .ZN(
        n12589) );
  INV_X1 U14328 ( .A(n12589), .ZN(n12590) );
  NAND3_X1 U14329 ( .A1(n12592), .A2(n12591), .A3(n12590), .ZN(n12593) );
  OR2_X1 U14330 ( .A1(n12594), .A2(n12593), .ZN(n14434) );
  AOI22_X1 U14331 ( .A1(n12648), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n12635), 
        .B2(n14434), .ZN(n12597) );
  AOI22_X1 U14332 ( .A1(n12595), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U14333 ( .A1(n12597), .A2(n12596), .ZN(n14153) );
  INV_X1 U14334 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U14335 ( .A1(n12595), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U14336 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15875), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U14337 ( .A1(n14809), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12598) );
  AND2_X1 U14338 ( .A1(n12599), .A2(n12598), .ZN(n12608) );
  AOI22_X1 U14339 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15876), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U14340 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12600) );
  AND2_X1 U14341 ( .A1(n12601), .A2(n12600), .ZN(n12607) );
  AOI22_X1 U14342 ( .A1(n12602), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12606) );
  INV_X1 U14343 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12603) );
  INV_X1 U14344 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15855) );
  OAI22_X1 U14345 ( .A1(n14571), .A2(n12603), .B1(n14569), .B2(n15855), .ZN(
        n12604) );
  INV_X1 U14346 ( .A(n12604), .ZN(n12605) );
  NAND4_X1 U14347 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        n12615) );
  AOI22_X1 U14348 ( .A1(n15865), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12609), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U14349 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U14350 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U14351 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12610) );
  NAND4_X1 U14352 ( .A1(n12613), .A2(n12612), .A3(n12611), .A4(n12610), .ZN(
        n12614) );
  OR2_X1 U14353 ( .A1(n12615), .A2(n12614), .ZN(n14437) );
  NAND2_X1 U14354 ( .A1(n12635), .A2(n14437), .ZN(n12616) );
  OAI211_X1 U14355 ( .C1(n15269), .C2(n12714), .A(n12617), .B(n12616), .ZN(
        n12618) );
  INV_X1 U14356 ( .A(n12618), .ZN(n14183) );
  INV_X1 U14357 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U14358 ( .A1(n12595), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U14359 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U14360 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U14361 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12092), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12619) );
  NAND3_X1 U14362 ( .A1(n12621), .A2(n12620), .A3(n12619), .ZN(n12634) );
  NAND2_X1 U14363 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12623) );
  NAND2_X1 U14364 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12622) );
  OAI211_X1 U14365 ( .C1(n15874), .C2(n12624), .A(n12623), .B(n12622), .ZN(
        n12628) );
  NAND2_X1 U14366 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12626) );
  NAND2_X1 U14367 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12625) );
  OAI211_X1 U14368 ( .C1(n12015), .C2(n19060), .A(n12626), .B(n12625), .ZN(
        n12627) );
  NOR2_X1 U14369 ( .A1(n12628), .A2(n12627), .ZN(n12632) );
  AOI22_X1 U14370 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12631) );
  NAND2_X1 U14371 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12630) );
  NAND2_X1 U14372 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12629) );
  NAND4_X1 U14373 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12633) );
  OR2_X1 U14374 ( .A1(n12634), .A2(n12633), .ZN(n14500) );
  NAND2_X1 U14375 ( .A1(n12635), .A2(n14500), .ZN(n12636) );
  OAI211_X1 U14376 ( .C1(n15269), .C2(n18191), .A(n12637), .B(n12636), .ZN(
        n14215) );
  NAND2_X1 U14377 ( .A1(n12648), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U14378 ( .A1(n12595), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12638) );
  INV_X1 U14379 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18219) );
  AOI22_X1 U14380 ( .A1(n12595), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12640) );
  OAI21_X1 U14381 ( .B1(n15269), .B2(n18219), .A(n12640), .ZN(n16207) );
  INV_X1 U14382 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U14383 ( .A1(n12595), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12641) );
  OAI21_X1 U14384 ( .B1(n15269), .B2(n17117), .A(n12641), .ZN(n16583) );
  NAND2_X1 U14385 ( .A1(n12648), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U14386 ( .A1(n12595), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12642) );
  AND2_X1 U14387 ( .A1(n12643), .A2(n12642), .ZN(n16197) );
  NAND2_X1 U14388 ( .A1(n12648), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U14389 ( .A1(n12595), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12644) );
  AND2_X1 U14390 ( .A1(n12645), .A2(n12644), .ZN(n16559) );
  NOR2_X4 U14391 ( .A1(n16560), .A2(n16559), .ZN(n16562) );
  INV_X1 U14392 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13891) );
  INV_X1 U14393 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17118) );
  OAI222_X1 U14394 ( .A1(n12647), .A2(n16537), .B1(n12646), .B2(n13891), .C1(
        n15269), .C2(n17118), .ZN(n16190) );
  NAND2_X1 U14395 ( .A1(n12648), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U14396 ( .A1(n12595), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12649) );
  AND2_X1 U14397 ( .A1(n12650), .A2(n12649), .ZN(n16180) );
  INV_X1 U14398 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18294) );
  AOI22_X1 U14399 ( .A1(n12595), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12651) );
  OAI21_X1 U14400 ( .B1(n15269), .B2(n18294), .A(n12651), .ZN(n16173) );
  INV_X1 U14401 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U14402 ( .A1(n12595), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12652) );
  OAI21_X1 U14403 ( .B1(n15269), .B2(n17119), .A(n12652), .ZN(n12653) );
  INV_X1 U14404 ( .A(n12653), .ZN(n16165) );
  INV_X1 U14405 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U14406 ( .A1(n12595), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12654) );
  OAI21_X1 U14407 ( .B1(n15269), .B2(n17120), .A(n12654), .ZN(n16156) );
  INV_X1 U14408 ( .A(n16156), .ZN(n12655) );
  INV_X1 U14409 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16275) );
  AOI22_X1 U14410 ( .A1(n12595), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12656) );
  OAI21_X1 U14411 ( .B1(n15269), .B2(n16275), .A(n12656), .ZN(n12657) );
  INV_X1 U14412 ( .A(n12657), .ZN(n16147) );
  INV_X1 U14413 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U14414 ( .A1(n12595), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12659) );
  OAI21_X1 U14415 ( .B1(n15269), .B2(n18339), .A(n12659), .ZN(n12660) );
  NOR2_X1 U14416 ( .A1(n16149), .A2(n12660), .ZN(n12661) );
  INV_X1 U14417 ( .A(n12662), .ZN(n12663) );
  NAND2_X1 U14418 ( .A1(n12664), .A2(n12663), .ZN(n12670) );
  INV_X1 U14419 ( .A(n12665), .ZN(n12668) );
  INV_X1 U14420 ( .A(n12666), .ZN(n12667) );
  NAND2_X1 U14421 ( .A1(n12668), .A2(n12667), .ZN(n12669) );
  NAND2_X1 U14422 ( .A1(n12670), .A2(n12669), .ZN(n13938) );
  INV_X1 U14423 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U14424 ( .A1(n15224), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U14425 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12671) );
  OAI211_X1 U14426 ( .C1(n12707), .C2(n12673), .A(n12672), .B(n12671), .ZN(
        n12674) );
  AOI21_X1 U14427 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12674), .ZN(n13937) );
  INV_X1 U14428 ( .A(n13937), .ZN(n12675) );
  NAND2_X1 U14429 ( .A1(n12676), .A2(n12675), .ZN(n13875) );
  INV_X1 U14430 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U14431 ( .A1(n15224), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U14432 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12677) );
  OAI211_X1 U14433 ( .C1(n12707), .C2(n14547), .A(n12678), .B(n12677), .ZN(
        n12679) );
  AOI21_X1 U14434 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12679), .ZN(n13876) );
  INV_X1 U14435 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U14436 ( .A1(n12743), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U14437 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12680) );
  OAI211_X1 U14438 ( .C1(n12707), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        n12683) );
  AOI21_X1 U14439 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12683), .ZN(n13927) );
  NAND2_X1 U14440 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12685) );
  AOI22_X1 U14441 ( .A1(n15224), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12684) );
  OAI211_X1 U14442 ( .C1(n12707), .C2(n18096), .A(n12685), .B(n12684), .ZN(
        n13907) );
  INV_X1 U14443 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U14444 ( .A1(n15224), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U14445 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12686) );
  OAI211_X1 U14446 ( .C1(n12707), .C2(n12688), .A(n12687), .B(n12686), .ZN(
        n12689) );
  AOI21_X1 U14447 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12689), .ZN(n14106) );
  NAND2_X1 U14448 ( .A1(n12752), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U14449 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12692) );
  OAI211_X1 U14450 ( .C1(n12707), .C2(n12694), .A(n12693), .B(n12692), .ZN(
        n12695) );
  AOI21_X1 U14451 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12695), .ZN(n14158) );
  INV_X1 U14452 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n18437) );
  NAND2_X1 U14453 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12697) );
  AOI22_X1 U14454 ( .A1(n15224), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12696) );
  OAI211_X1 U14455 ( .C1(n12707), .C2(n18437), .A(n12697), .B(n12696), .ZN(
        n14236) );
  NAND2_X1 U14456 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12699) );
  AOI22_X1 U14457 ( .A1(n15224), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12698) );
  OAI211_X1 U14458 ( .C1(n12707), .C2(n16417), .A(n12699), .B(n12698), .ZN(
        n14198) );
  AOI22_X1 U14459 ( .A1(n12743), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12701) );
  INV_X1 U14460 ( .A(n12707), .ZN(n12711) );
  NAND2_X1 U14461 ( .A1(n12711), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12700) );
  OAI211_X1 U14462 ( .C1(n12703), .C2(n12702), .A(n12701), .B(n12700), .ZN(
        n14300) );
  NAND2_X1 U14463 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12710) );
  INV_X1 U14464 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12706) );
  NAND2_X1 U14465 ( .A1(n15224), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U14466 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12704) );
  OAI211_X1 U14467 ( .C1(n12707), .C2(n12706), .A(n12705), .B(n12704), .ZN(
        n12708) );
  INV_X1 U14468 ( .A(n12708), .ZN(n12709) );
  NAND2_X1 U14469 ( .A1(n12710), .A2(n12709), .ZN(n14328) );
  NAND2_X1 U14470 ( .A1(n15224), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U14471 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12712) );
  OAI211_X1 U14472 ( .C1(n15227), .C2(n12714), .A(n12713), .B(n12712), .ZN(
        n12715) );
  AOI21_X1 U14473 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12715), .ZN(n14430) );
  NAND2_X1 U14474 ( .A1(n12752), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U14475 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12716) );
  OAI211_X1 U14476 ( .C1(n15227), .C2(n18191), .A(n12717), .B(n12716), .ZN(
        n12718) );
  AOI21_X1 U14477 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12718), .ZN(n14495) );
  INV_X1 U14478 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U14479 ( .A1(n15224), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U14480 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12719) );
  OAI211_X1 U14481 ( .C1(n15227), .C2(n12721), .A(n12720), .B(n12719), .ZN(
        n12722) );
  AOI21_X1 U14482 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12722), .ZN(n14534) );
  NAND2_X1 U14483 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12724) );
  AOI22_X1 U14484 ( .A1(n15224), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12723) );
  OAI211_X1 U14485 ( .C1(n15227), .C2(n18219), .A(n12724), .B(n12723), .ZN(
        n14581) );
  NAND2_X1 U14486 ( .A1(n14582), .A2(n14581), .ZN(n14580) );
  NAND2_X1 U14487 ( .A1(n12743), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U14488 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12725) );
  OAI211_X1 U14489 ( .C1(n15227), .C2(n17117), .A(n12726), .B(n12725), .ZN(
        n12727) );
  AOI21_X1 U14490 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12727), .ZN(n14604) );
  INV_X1 U14491 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18242) );
  NAND2_X1 U14492 ( .A1(n15224), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U14493 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12728) );
  OAI211_X1 U14494 ( .C1(n15227), .C2(n18242), .A(n12729), .B(n12728), .ZN(
        n12730) );
  AOI21_X1 U14495 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12730), .ZN(n14803) );
  INV_X1 U14496 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16342) );
  NAND2_X1 U14497 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12732) );
  AOI22_X1 U14498 ( .A1(n15224), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12731) );
  OAI211_X1 U14499 ( .C1(n15227), .C2(n16342), .A(n12732), .B(n12731), .ZN(
        n14744) );
  NAND2_X1 U14500 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12734) );
  AOI22_X1 U14501 ( .A1(n12752), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12733) );
  OAI211_X1 U14502 ( .C1(n15227), .C2(n17118), .A(n12734), .B(n12733), .ZN(
        n14831) );
  NAND2_X1 U14503 ( .A1(n14742), .A2(n14831), .ZN(n14830) );
  INV_X1 U14504 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U14505 ( .A1(n15224), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U14506 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12735) );
  OAI211_X1 U14507 ( .C1(n15227), .C2(n12737), .A(n12736), .B(n12735), .ZN(
        n12738) );
  AOI21_X1 U14508 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12738), .ZN(n16109) );
  NAND2_X1 U14509 ( .A1(n15224), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U14510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12739) );
  OAI211_X1 U14511 ( .C1(n15227), .C2(n18294), .A(n12740), .B(n12739), .ZN(
        n12741) );
  AOI21_X1 U14512 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12741), .ZN(n16101) );
  NAND2_X1 U14513 ( .A1(n12743), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U14514 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12744) );
  OAI211_X1 U14515 ( .C1(n15227), .C2(n17119), .A(n12745), .B(n12744), .ZN(
        n12746) );
  AOI21_X1 U14516 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12746), .ZN(n16095) );
  NAND2_X1 U14517 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12748) );
  AOI22_X1 U14518 ( .A1(n15224), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12747) );
  OAI211_X1 U14519 ( .C1(n15227), .C2(n17120), .A(n12748), .B(n12747), .ZN(
        n16088) );
  NAND2_X1 U14520 ( .A1(n15224), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U14521 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12749) );
  OAI211_X1 U14522 ( .C1(n15227), .C2(n16275), .A(n12750), .B(n12749), .ZN(
        n12751) );
  AOI21_X1 U14523 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12751), .ZN(n16076) );
  NAND2_X1 U14524 ( .A1(n12752), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U14525 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12753) );
  OAI211_X1 U14526 ( .C1(n15227), .C2(n18339), .A(n12754), .B(n12753), .ZN(
        n12755) );
  AOI21_X1 U14527 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12755), .ZN(n12756) );
  AND2_X1 U14528 ( .A1(n16078), .A2(n12756), .ZN(n12757) );
  OR2_X1 U14529 ( .A1(n12757), .A2(n16065), .ZN(n16072) );
  NAND2_X1 U14530 ( .A1(n13987), .A2(n15968), .ZN(n12759) );
  NAND2_X1 U14531 ( .A1(n13967), .A2(n12758), .ZN(n13951) );
  NAND2_X1 U14532 ( .A1(n12759), .A2(n13951), .ZN(n12760) );
  AND2_X2 U14533 ( .A1(n12815), .A2(n12760), .ZN(n18500) );
  NAND2_X1 U14534 ( .A1(n18347), .A2(n18500), .ZN(n12770) );
  INV_X1 U14535 ( .A(n12761), .ZN(n12767) );
  INV_X1 U14536 ( .A(n18495), .ZN(n16548) );
  NAND2_X1 U14537 ( .A1(n16548), .A2(n18488), .ZN(n12764) );
  NAND2_X1 U14538 ( .A1(n12762), .A2(n18486), .ZN(n12763) );
  NAND2_X1 U14539 ( .A1(n12764), .A2(n12763), .ZN(n14612) );
  NAND2_X1 U14540 ( .A1(n14612), .A2(n12765), .ZN(n16651) );
  NOR2_X1 U14541 ( .A1(n12811), .A2(n16651), .ZN(n16529) );
  INV_X1 U14542 ( .A(n16529), .ZN(n12766) );
  NOR2_X1 U14543 ( .A1(n12767), .A2(n12766), .ZN(n16505) );
  NAND2_X1 U14544 ( .A1(n16505), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16492) );
  NOR2_X1 U14545 ( .A1(n16457), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12768) );
  NOR2_X1 U14546 ( .A1(n18240), .A2(n18339), .ZN(n16257) );
  NOR2_X1 U14547 ( .A1(n12768), .A2(n16257), .ZN(n12769) );
  OAI211_X1 U14548 ( .C1(n18490), .C2(n18353), .A(n12770), .B(n12769), .ZN(
        n12771) );
  AOI21_X1 U14549 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16455), .A(
        n12771), .ZN(n12817) );
  NOR2_X1 U14550 ( .A1(n18418), .A2(n13535), .ZN(n13534) );
  INV_X1 U14551 ( .A(n12774), .ZN(n12772) );
  NAND2_X1 U14552 ( .A1(n13534), .A2(n12772), .ZN(n12775) );
  NOR2_X1 U14553 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13535), .ZN(
        n12773) );
  XOR2_X1 U14554 ( .A(n12774), .B(n12773), .Z(n13528) );
  NAND2_X1 U14555 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13528), .ZN(
        n13527) );
  NAND2_X1 U14556 ( .A1(n12775), .A2(n13527), .ZN(n12778) );
  XNOR2_X1 U14557 ( .A(n18508), .B(n12778), .ZN(n13598) );
  XNOR2_X1 U14558 ( .A(n12777), .B(n12776), .ZN(n13597) );
  NAND2_X1 U14559 ( .A1(n13598), .A2(n13597), .ZN(n12780) );
  NAND2_X1 U14560 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12778), .ZN(
        n12779) );
  NAND2_X1 U14561 ( .A1(n12780), .A2(n12779), .ZN(n12781) );
  XNOR2_X1 U14562 ( .A(n12781), .B(n14365), .ZN(n14352) );
  NAND2_X1 U14563 ( .A1(n12781), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12782) );
  XNOR2_X1 U14564 ( .A(n12787), .B(n12786), .ZN(n14388) );
  NAND2_X1 U14565 ( .A1(n14388), .A2(n14544), .ZN(n14387) );
  INV_X1 U14566 ( .A(n12786), .ZN(n12788) );
  AND2_X1 U14567 ( .A1(n12790), .A2(n14548), .ZN(n12792) );
  NAND2_X1 U14568 ( .A1(n12796), .A2(n12791), .ZN(n12797) );
  XNOR2_X1 U14569 ( .A(n12806), .B(n15212), .ZN(n12802) );
  XNOR2_X1 U14570 ( .A(n12802), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14722) );
  NAND2_X1 U14571 ( .A1(n14723), .A2(n14722), .ZN(n12805) );
  INV_X1 U14572 ( .A(n12802), .ZN(n12803) );
  NAND2_X1 U14573 ( .A1(n12803), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12804) );
  NAND2_X1 U14574 ( .A1(n12808), .A2(n11337), .ZN(n12807) );
  NAND2_X1 U14575 ( .A1(n16977), .A2(n16976), .ZN(n12810) );
  NAND3_X1 U14576 ( .A1(n12808), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11337), .ZN(n12809) );
  INV_X1 U14577 ( .A(n12811), .ZN(n12812) );
  INV_X1 U14578 ( .A(n12813), .ZN(n12814) );
  INV_X1 U14579 ( .A(n16246), .ZN(n16237) );
  AOI21_X1 U14580 ( .B1(n15190), .B2(n16269), .A(n16237), .ZN(n16260) );
  NAND2_X1 U14581 ( .A1(n12815), .A2(n14000), .ZN(n18494) );
  NAND2_X1 U14582 ( .A1(n16260), .A2(n18481), .ZN(n12816) );
  OAI21_X1 U14583 ( .B1(n16262), .B2(n18450), .A(n12818), .ZN(P2_U3019) );
  INV_X1 U14584 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12821) );
  AND2_X2 U14585 ( .A1(n12821), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12827) );
  AOI22_X1 U14586 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12824) );
  AND2_X4 U14587 ( .A1(n14055), .A2(n12827), .ZN(n13007) );
  AOI22_X1 U14588 ( .A1(n10982), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12823) );
  AND2_X2 U14589 ( .A1(n12827), .A2(n14042), .ZN(n14651) );
  AOI22_X1 U14590 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12829) );
  AND2_X2 U14591 ( .A1(n12827), .A2(n12830), .ZN(n14406) );
  AOI22_X1 U14592 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U14593 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12923), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U14594 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U14595 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U14596 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U14597 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13080), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U14598 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U14599 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12839) );
  NAND2_X2 U14600 ( .A1(n12843), .A2(n11005), .ZN(n15511) );
  AOI22_X1 U14601 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U14602 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U14603 ( .A1(n12923), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U14604 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12906), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U14605 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U14606 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13039), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U14607 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U14608 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12848) );
  INV_X1 U14609 ( .A(n12986), .ZN(n12854) );
  NAND2_X1 U14610 ( .A1(n13674), .A2(n12854), .ZN(n12899) );
  NAND2_X1 U14611 ( .A1(n12923), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12859) );
  NAND2_X1 U14612 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12858) );
  NAND2_X1 U14613 ( .A1(n12941), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12857) );
  NAND2_X1 U14614 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12856) );
  NAND2_X1 U14615 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12863) );
  NAND2_X1 U14616 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12862) );
  NAND2_X1 U14617 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12861) );
  NAND2_X1 U14618 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U14619 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12867) );
  NAND2_X1 U14620 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12866) );
  NAND2_X1 U14621 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12865) );
  NAND2_X1 U14622 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U14623 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U14624 ( .A1(n12946), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U14625 ( .A1(n12906), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12869) );
  NAND2_X1 U14626 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12868) );
  NAND4_X4 U14627 ( .A1(n12875), .A2(n12874), .A3(n12873), .A4(n12872), .ZN(
        n12966) );
  NAND2_X1 U14628 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U14629 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12878) );
  NAND2_X1 U14630 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U14631 ( .A1(n12923), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12876) );
  NAND2_X1 U14632 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12883) );
  NAND2_X1 U14633 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12881) );
  NAND2_X1 U14634 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12880) );
  NAND2_X1 U14635 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  NAND2_X1 U14636 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12889) );
  NAND2_X1 U14637 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12888) );
  NAND2_X1 U14638 ( .A1(n12906), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U14639 ( .A1(n12946), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12886) );
  NAND2_X1 U14640 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12893) );
  NAND2_X1 U14641 ( .A1(n12941), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12892) );
  NAND2_X1 U14642 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12891) );
  NAND2_X1 U14643 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12890) );
  NAND2_X1 U14644 ( .A1(n12899), .A2(n12972), .ZN(n12914) );
  NAND2_X1 U14645 ( .A1(n12966), .A2(n13315), .ZN(n12912) );
  INV_X1 U14646 ( .A(n12973), .ZN(n12960) );
  AOI22_X1 U14647 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12923), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12905) );
  AOI21_X1 U14648 ( .B1(n12951), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n12900), .ZN(n12904) );
  AOI22_X1 U14649 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12928), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U14650 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U14651 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U14652 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13080), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U14653 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10978), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U14654 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U14655 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12918) );
  NAND2_X1 U14656 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12917) );
  NAND2_X1 U14657 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12916) );
  NAND2_X1 U14658 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12915) );
  NAND2_X1 U14659 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12922) );
  NAND2_X1 U14660 ( .A1(n12941), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U14661 ( .A1(n12946), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12920) );
  NAND2_X1 U14662 ( .A1(n12906), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12919) );
  NAND2_X1 U14663 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12927) );
  NAND2_X1 U14664 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12926) );
  NAND2_X1 U14665 ( .A1(n12923), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12925) );
  NAND2_X1 U14666 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12924) );
  NAND2_X1 U14667 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12932) );
  NAND2_X1 U14668 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12931) );
  NAND2_X1 U14669 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12930) );
  NAND2_X1 U14670 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12929) );
  NAND4_X2 U14671 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12978) );
  NAND2_X1 U14672 ( .A1(n12901), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12940) );
  NAND2_X1 U14673 ( .A1(n14411), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12939) );
  NAND2_X1 U14674 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12938) );
  NAND2_X1 U14675 ( .A1(n12923), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12937) );
  NAND2_X1 U14676 ( .A1(n14406), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12945) );
  NAND2_X1 U14677 ( .A1(n12941), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12944) );
  NAND2_X1 U14678 ( .A1(n13080), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12943) );
  NAND2_X1 U14679 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12942) );
  NAND2_X1 U14680 ( .A1(n13039), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12950) );
  NAND2_X1 U14681 ( .A1(n13044), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12949) );
  NAND2_X1 U14682 ( .A1(n10978), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12948) );
  NAND2_X1 U14683 ( .A1(n12946), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12947) );
  NAND2_X1 U14684 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12955) );
  NAND2_X1 U14685 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12954) );
  NAND2_X1 U14686 ( .A1(n12951), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U14687 ( .A1(n12928), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12952) );
  NAND2_X1 U14688 ( .A1(n12985), .A2(n12960), .ZN(n12961) );
  INV_X1 U14689 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n12962) );
  XNOR2_X1 U14690 ( .A(n12962), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13265) );
  NOR2_X1 U14691 ( .A1(n12980), .A2(n12966), .ZN(n12964) );
  NAND2_X1 U14692 ( .A1(n22104), .A2(n13315), .ZN(n12968) );
  INV_X1 U14693 ( .A(n12974), .ZN(n12975) );
  INV_X1 U14694 ( .A(n12977), .ZN(n12979) );
  OAI21_X1 U14695 ( .B1(n12984), .B2(n15291), .A(n13313), .ZN(n12981) );
  NAND2_X1 U14696 ( .A1(n12982), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U14697 ( .A1(n13070), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12983) );
  NAND2_X1 U14698 ( .A1(n15797), .A2(n21614), .ZN(n13780) );
  MUX2_X1 U14699 ( .A(n13780), .B(n13321), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n13035) );
  NAND2_X1 U14700 ( .A1(n12984), .A2(n12985), .ZN(n13446) );
  NAND2_X1 U14701 ( .A1(n12969), .A2(n12986), .ZN(n12989) );
  NAND2_X1 U14702 ( .A1(n21716), .A2(n12978), .ZN(n14275) );
  NAND2_X1 U14703 ( .A1(n12965), .A2(n14272), .ZN(n12987) );
  NAND4_X1 U14704 ( .A1(n14275), .A2(n15797), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n12987), .ZN(n12988) );
  AOI21_X1 U14705 ( .B1(n13517), .B2(n12989), .A(n12988), .ZN(n12993) );
  NAND2_X1 U14706 ( .A1(n12974), .A2(n12963), .ZN(n12990) );
  AND2_X1 U14707 ( .A1(n13695), .A2(n12990), .ZN(n13450) );
  AOI22_X1 U14708 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14709 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15000), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U14710 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14711 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13045), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U14712 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n13006) );
  AOI22_X1 U14713 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U14714 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14716 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14717 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U14718 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13005) );
  NAND2_X1 U14719 ( .A1(n12970), .A2(n13206), .ZN(n13208) );
  INV_X1 U14720 ( .A(n13208), .ZN(n13019) );
  AOI22_X1 U14721 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U14722 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U14723 ( .A1(n15145), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13009) );
  AOI22_X1 U14724 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13008) );
  NAND4_X1 U14725 ( .A1(n13011), .A2(n13010), .A3(n13009), .A4(n13008), .ZN(
        n13017) );
  AOI22_X1 U14726 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U14727 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U14728 ( .A1(n14651), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U14729 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13012) );
  NAND4_X1 U14730 ( .A1(n13015), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13016) );
  INV_X1 U14731 ( .A(n13054), .ZN(n13018) );
  NAND2_X1 U14732 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NOR2_X1 U14733 ( .A1(n13435), .A2(n21614), .ZN(n13095) );
  INV_X1 U14734 ( .A(n13206), .ZN(n13195) );
  NAND3_X1 U14735 ( .A1(n13095), .A2(n13195), .A3(n13054), .ZN(n13026) );
  INV_X1 U14736 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13023) );
  AOI21_X1 U14737 ( .B1(n21716), .B2(n13054), .A(n21614), .ZN(n13022) );
  OAI211_X1 U14738 ( .C1(n13294), .C2(n13023), .A(n13022), .B(n13208), .ZN(
        n13024) );
  INV_X1 U14739 ( .A(n13024), .ZN(n13025) );
  NAND2_X1 U14740 ( .A1(n13093), .A2(n11395), .ZN(n13671) );
  INV_X1 U14741 ( .A(n13278), .ZN(n13148) );
  AND2_X1 U14742 ( .A1(n21716), .A2(n12986), .ZN(n13100) );
  AOI21_X1 U14743 ( .B1(n13018), .B2(n21195), .A(n13100), .ZN(n13027) );
  NAND2_X1 U14744 ( .A1(n13791), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13062) );
  XNOR2_X1 U14745 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21739) );
  NAND2_X1 U14746 ( .A1(n16762), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13066) );
  OAI21_X1 U14747 ( .B1(n13780), .B2(n21739), .A(n13066), .ZN(n13030) );
  INV_X1 U14748 ( .A(n13030), .ZN(n13029) );
  NAND3_X1 U14749 ( .A1(n13065), .A2(n13029), .A3(n13028), .ZN(n13032) );
  OR2_X1 U14750 ( .A1(n13030), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13031) );
  INV_X1 U14751 ( .A(n21749), .ZN(n13038) );
  INV_X1 U14752 ( .A(n13036), .ZN(n13037) );
  AOI22_X1 U14753 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U14754 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U14755 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10963), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U14756 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13040) );
  NAND4_X1 U14757 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13052) );
  AOI22_X1 U14758 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U14759 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U14760 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U14761 ( .A1(n13045), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13047) );
  NAND4_X1 U14762 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13051) );
  NAND2_X1 U14763 ( .A1(n13095), .A2(n13094), .ZN(n13053) );
  OR2_X2 U14764 ( .A1(n13092), .A2(n13148), .ZN(n13061) );
  NAND2_X1 U14765 ( .A1(n13094), .A2(n13054), .ZN(n13127) );
  OAI21_X1 U14766 ( .B1(n13054), .B2(n13094), .A(n13127), .ZN(n13055) );
  INV_X1 U14767 ( .A(n13055), .ZN(n13058) );
  NAND2_X1 U14768 ( .A1(n13056), .A2(n12966), .ZN(n13057) );
  AOI21_X1 U14769 ( .B1(n13058), .B2(n21195), .A(n13057), .ZN(n13060) );
  INV_X1 U14770 ( .A(n13792), .ZN(n13063) );
  NAND2_X1 U14771 ( .A1(n13059), .A2(n13063), .ZN(n13064) );
  NAND2_X1 U14772 ( .A1(n13066), .A2(n12821), .ZN(n13067) );
  NAND2_X1 U14773 ( .A1(n13033), .A2(n13067), .ZN(n13068) );
  INV_X1 U14774 ( .A(n13780), .ZN(n13111) );
  NAND2_X1 U14775 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U14776 ( .A1(n21853), .A2(n13071), .ZN(n13073) );
  NAND2_X1 U14777 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21896) );
  INV_X1 U14778 ( .A(n21896), .ZN(n13072) );
  NAND2_X1 U14779 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13072), .ZN(
        n21893) );
  AND2_X1 U14780 ( .A1(n13073), .A2(n21893), .ZN(n21717) );
  AOI22_X1 U14781 ( .A1(n13111), .A2(n21717), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16762), .ZN(n13074) );
  NAND2_X2 U14782 ( .A1(n13077), .A2(n13076), .ZN(n13661) );
  AOI22_X1 U14783 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14784 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U14785 ( .A1(n15139), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U14786 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13081) );
  NAND4_X1 U14787 ( .A1(n13084), .A2(n13083), .A3(n13082), .A4(n13081), .ZN(
        n13090) );
  AOI22_X1 U14788 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U14789 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U14790 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U14791 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13085) );
  NAND4_X1 U14792 ( .A1(n13088), .A2(n13087), .A3(n13086), .A4(n13085), .ZN(
        n13089) );
  AOI22_X1 U14793 ( .A1(n13269), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13305), .B2(n13125), .ZN(n13091) );
  NAND3_X1 U14794 ( .A1(n21716), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13094), 
        .ZN(n13097) );
  INV_X1 U14795 ( .A(n13095), .ZN(n13096) );
  NAND2_X1 U14796 ( .A1(n13097), .A2(n13096), .ZN(n13098) );
  AOI21_X1 U14797 ( .B1(n13269), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n13098), .ZN(n13099) );
  INV_X1 U14798 ( .A(n21195), .ZN(n16759) );
  XNOR2_X1 U14799 ( .A(n13127), .B(n13125), .ZN(n13102) );
  INV_X1 U14800 ( .A(n13100), .ZN(n13101) );
  OAI21_X1 U14801 ( .B1(n16759), .B2(n13102), .A(n13101), .ZN(n13103) );
  XNOR2_X1 U14802 ( .A(n13129), .B(n13106), .ZN(n14228) );
  INV_X1 U14803 ( .A(n21893), .ZN(n13109) );
  NAND2_X1 U14804 ( .A1(n13109), .A2(n21897), .ZN(n21793) );
  NAND2_X1 U14805 ( .A1(n21893), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13110) );
  NAND2_X1 U14806 ( .A1(n21793), .A2(n13110), .ZN(n21806) );
  AOI22_X1 U14807 ( .A1(n13111), .A2(n21806), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16762), .ZN(n13112) );
  XNOR2_X2 U14808 ( .A(n13661), .B(n21764), .ZN(n21804) );
  AOI22_X1 U14809 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U14810 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U14811 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U14812 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13114) );
  NAND4_X1 U14813 ( .A1(n13117), .A2(n13116), .A3(n13115), .A4(n13114), .ZN(
        n13123) );
  AOI22_X1 U14814 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U14815 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U14816 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U14817 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13118) );
  NAND4_X1 U14818 ( .A1(n13121), .A2(n13120), .A3(n13119), .A4(n13118), .ZN(
        n13122) );
  AOI22_X1 U14819 ( .A1(n13269), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13305), .B2(n13145), .ZN(n13124) );
  INV_X1 U14820 ( .A(n13125), .ZN(n13126) );
  NAND2_X1 U14821 ( .A1(n13127), .A2(n13126), .ZN(n13146) );
  XOR2_X1 U14822 ( .A(n13146), .B(n13145), .Z(n13128) );
  AOI22_X1 U14823 ( .A1(n21802), .A2(n13278), .B1(n21195), .B2(n13128), .ZN(
        n14230) );
  INV_X1 U14824 ( .A(n13129), .ZN(n13130) );
  INV_X1 U14825 ( .A(n13131), .ZN(n13132) );
  INV_X1 U14826 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U14827 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U14828 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U14829 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U14830 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13133) );
  NAND4_X1 U14831 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        n13142) );
  AOI22_X1 U14832 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U14833 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U14834 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U14835 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13137) );
  NAND4_X1 U14836 ( .A1(n13140), .A2(n13139), .A3(n13138), .A4(n13137), .ZN(
        n13141) );
  NAND2_X1 U14837 ( .A1(n13305), .A2(n13165), .ZN(n13143) );
  XNOR2_X1 U14838 ( .A(n13152), .B(n13151), .ZN(n14141) );
  INV_X1 U14839 ( .A(n14141), .ZN(n13149) );
  NAND2_X1 U14840 ( .A1(n13146), .A2(n13145), .ZN(n13167) );
  XOR2_X1 U14841 ( .A(n13167), .B(n13165), .Z(n13147) );
  OAI22_X1 U14842 ( .A1(n13149), .A2(n13148), .B1(n13147), .B2(n16759), .ZN(
        n19894) );
  INV_X1 U14843 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21248) );
  INV_X1 U14844 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U14845 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U14846 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13155) );
  AOI22_X1 U14847 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U14848 ( .A1(n15138), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13153) );
  NAND4_X1 U14849 ( .A1(n13156), .A2(n13155), .A3(n13154), .A4(n13153), .ZN(
        n13162) );
  AOI22_X1 U14850 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U14851 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U14852 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U14853 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13157) );
  NAND4_X1 U14854 ( .A1(n13160), .A2(n13159), .A3(n13158), .A4(n13157), .ZN(
        n13161) );
  NAND2_X1 U14855 ( .A1(n13305), .A2(n13190), .ZN(n13163) );
  INV_X1 U14856 ( .A(n13165), .ZN(n13166) );
  NOR2_X1 U14857 ( .A1(n13167), .A2(n13166), .ZN(n13191) );
  XOR2_X1 U14858 ( .A(n13190), .B(n13191), .Z(n13168) );
  AOI22_X1 U14859 ( .A1(n14191), .A2(n13278), .B1(n21195), .B2(n13168), .ZN(
        n13169) );
  XNOR2_X1 U14860 ( .A(n13169), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19901) );
  INV_X1 U14861 ( .A(n13169), .ZN(n13170) );
  INV_X1 U14862 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21264) );
  NAND2_X1 U14863 ( .A1(n13170), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13171) );
  NAND2_X1 U14864 ( .A1(n13269), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13185) );
  AOI22_X1 U14865 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U14866 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U14867 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U14868 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13174) );
  NAND4_X1 U14869 ( .A1(n13177), .A2(n13176), .A3(n13175), .A4(n13174), .ZN(
        n13183) );
  AOI22_X1 U14870 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U14871 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U14872 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U14873 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13178) );
  NAND4_X1 U14874 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n13182) );
  NAND2_X1 U14875 ( .A1(n13305), .A2(n13200), .ZN(n13184) );
  NAND2_X1 U14876 ( .A1(n13189), .A2(n13188), .ZN(n14217) );
  NAND2_X1 U14877 ( .A1(n13191), .A2(n13190), .ZN(n13199) );
  XNOR2_X1 U14878 ( .A(n13199), .B(n13200), .ZN(n13192) );
  AOI22_X1 U14879 ( .A1(n13207), .A2(n14217), .B1(n21195), .B2(n13192), .ZN(
        n13193) );
  XNOR2_X1 U14880 ( .A(n13193), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19906) );
  NAND2_X1 U14881 ( .A1(n19907), .A2(n19906), .ZN(n19905) );
  INV_X1 U14882 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21262) );
  NAND2_X1 U14883 ( .A1(n19905), .A2(n13194), .ZN(n19913) );
  INV_X1 U14884 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13196) );
  OAI22_X1 U14885 ( .A1(n13294), .A2(n13196), .B1(n13279), .B2(n13195), .ZN(
        n13197) );
  INV_X1 U14886 ( .A(n13199), .ZN(n13201) );
  NAND2_X1 U14887 ( .A1(n13201), .A2(n13200), .ZN(n13210) );
  XNOR2_X1 U14888 ( .A(n13210), .B(n13206), .ZN(n13202) );
  AOI22_X1 U14889 ( .A1(n14251), .A2(n13278), .B1(n21195), .B2(n13202), .ZN(
        n13203) );
  XNOR2_X1 U14890 ( .A(n13203), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19912) );
  INV_X1 U14891 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21284) );
  NAND2_X1 U14892 ( .A1(n21195), .A2(n13206), .ZN(n13209) );
  XOR2_X1 U14893 ( .A(n13211), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(
        n15182) );
  INV_X1 U14894 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21292) );
  INV_X1 U14895 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U14896 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13215) );
  XNOR2_X1 U14897 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15698) );
  INV_X1 U14898 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U14899 ( .A1(n13221), .A2(n13377), .ZN(n13216) );
  INV_X1 U14900 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13217) );
  INV_X1 U14901 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15705) );
  INV_X1 U14902 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21326) );
  NAND2_X1 U14903 ( .A1(n15705), .A2(n21326), .ZN(n13222) );
  NAND2_X1 U14904 ( .A1(n13212), .A2(n13222), .ZN(n15693) );
  NAND2_X1 U14905 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15696) );
  OAI21_X1 U14906 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n13212), .ZN(n13223) );
  NAND2_X1 U14907 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15671) );
  AND3_X1 U14908 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15780) );
  NAND2_X1 U14909 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15626) );
  INV_X1 U14910 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15756) );
  OAI21_X1 U14911 ( .B1(n15626), .B2(n15756), .A(n13221), .ZN(n15600) );
  INV_X1 U14912 ( .A(n13224), .ZN(n15653) );
  OR4_X1 U14913 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U14914 ( .B1(n13224), .B2(n13225), .A(n13212), .ZN(n15647) );
  INV_X1 U14915 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15763) );
  INV_X1 U14916 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13409) );
  NAND3_X1 U14917 ( .A1(n15763), .A2(n15756), .A3(n13409), .ZN(n15601) );
  INV_X1 U14918 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15747) );
  NOR2_X1 U14919 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15723) );
  NOR2_X1 U14920 ( .A1(n13221), .A2(n15723), .ZN(n13229) );
  AND2_X1 U14921 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15724) );
  NOR2_X1 U14922 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15590) );
  NOR2_X1 U14923 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13231) );
  XNOR2_X1 U14924 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13234) );
  INV_X1 U14925 ( .A(n13234), .ZN(n13230) );
  OAI21_X1 U14926 ( .B1(n13231), .B2(n13221), .A(n13230), .ZN(n13237) );
  INV_X1 U14927 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U14928 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15244) );
  NAND2_X1 U14929 ( .A1(n13221), .A2(n15252), .ZN(n13233) );
  OAI211_X1 U14930 ( .C1(n13221), .C2(n15252), .A(n15244), .B(n13233), .ZN(
        n13232) );
  INV_X1 U14931 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13706) );
  AND2_X1 U14932 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  NAND2_X1 U14933 ( .A1(n15588), .A2(n13235), .ZN(n13236) );
  NAND2_X1 U14934 ( .A1(n21827), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13239) );
  NAND2_X1 U14935 ( .A1(n12821), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13238) );
  NAND2_X1 U14936 ( .A1(n13239), .A2(n13238), .ZN(n13252) );
  NAND2_X1 U14937 ( .A1(n21864), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13268) );
  INV_X1 U14938 ( .A(n13249), .ZN(n13242) );
  NAND2_X1 U14939 ( .A1(n21853), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13243) );
  NAND2_X1 U14940 ( .A1(n12819), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13240) );
  NAND2_X1 U14941 ( .A1(n13243), .A2(n13240), .ZN(n13248) );
  INV_X1 U14942 ( .A(n13248), .ZN(n13241) );
  NAND2_X1 U14943 ( .A1(n13242), .A2(n13241), .ZN(n13250) );
  NAND2_X1 U14944 ( .A1(n13250), .A2(n13243), .ZN(n13260) );
  NAND2_X1 U14945 ( .A1(n13260), .A2(n13255), .ZN(n13247) );
  NAND2_X1 U14946 ( .A1(n21897), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13256) );
  INV_X1 U14947 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16769) );
  NAND2_X1 U14948 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16769), .ZN(
        n13244) );
  AND2_X1 U14949 ( .A1(n13256), .A2(n13244), .ZN(n13246) );
  INV_X1 U14950 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U14951 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14054), .ZN(
        n13257) );
  INV_X1 U14952 ( .A(n13257), .ZN(n13245) );
  INV_X1 U14953 ( .A(n13304), .ZN(n13263) );
  NAND2_X1 U14954 ( .A1(n13249), .A2(n13248), .ZN(n13251) );
  AND2_X1 U14955 ( .A1(n13251), .A2(n13250), .ZN(n13290) );
  NAND2_X1 U14956 ( .A1(n13252), .A2(n13268), .ZN(n13253) );
  NAND2_X1 U14957 ( .A1(n13254), .A2(n13253), .ZN(n13280) );
  INV_X1 U14958 ( .A(n13280), .ZN(n13277) );
  NAND2_X1 U14959 ( .A1(n13290), .A2(n13277), .ZN(n13261) );
  AND2_X1 U14960 ( .A1(n13256), .A2(n13255), .ZN(n13259) );
  INV_X1 U14961 ( .A(n13256), .ZN(n13258) );
  OAI22_X1 U14962 ( .A1(n13260), .A2(n13259), .B1(n13258), .B2(n13257), .ZN(
        n13298) );
  OR2_X1 U14963 ( .A1(n13261), .A2(n13298), .ZN(n13262) );
  INV_X1 U14964 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U14965 ( .A1(n13265), .A2(n13264), .ZN(n21657) );
  NAND2_X1 U14966 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21660) );
  INV_X1 U14967 ( .A(n21660), .ZN(n13643) );
  AOI21_X1 U14968 ( .B1(n12978), .B2(n21657), .A(n13643), .ZN(n13266) );
  NAND2_X1 U14969 ( .A1(n15288), .A2(n13266), .ZN(n13312) );
  NAND2_X1 U14970 ( .A1(n11111), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13267) );
  NAND2_X1 U14971 ( .A1(n13268), .A2(n13267), .ZN(n13271) );
  NAND2_X1 U14972 ( .A1(n13269), .A2(n13278), .ZN(n13297) );
  OAI21_X1 U14973 ( .B1(n13279), .B2(n13271), .A(n13297), .ZN(n13275) );
  NAND2_X1 U14974 ( .A1(n22104), .A2(n14272), .ZN(n13270) );
  NAND2_X1 U14975 ( .A1(n13270), .A2(n21915), .ZN(n13289) );
  INV_X1 U14976 ( .A(n13271), .ZN(n13272) );
  OAI211_X1 U14977 ( .C1(n13442), .C2(n21716), .A(n13289), .B(n13272), .ZN(
        n13274) );
  OR2_X1 U14978 ( .A1(n12966), .A2(n21614), .ZN(n13276) );
  NAND3_X1 U14979 ( .A1(n13276), .A2(n21915), .A3(n13280), .ZN(n13273) );
  NAND3_X1 U14980 ( .A1(n13275), .A2(n13274), .A3(n13273), .ZN(n13285) );
  OAI211_X1 U14981 ( .C1(n13279), .C2(n21915), .A(n13277), .B(n13276), .ZN(
        n13283) );
  NAND2_X1 U14982 ( .A1(n13279), .A2(n13278), .ZN(n13281) );
  NAND2_X1 U14983 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  NAND2_X1 U14984 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  NAND2_X1 U14985 ( .A1(n13285), .A2(n13284), .ZN(n13288) );
  NAND2_X1 U14986 ( .A1(n13305), .A2(n13290), .ZN(n13286) );
  OAI211_X1 U14987 ( .C1(n13294), .C2(n13290), .A(n13286), .B(n13289), .ZN(
        n13287) );
  NAND2_X1 U14988 ( .A1(n13288), .A2(n13287), .ZN(n13293) );
  INV_X1 U14989 ( .A(n13289), .ZN(n13291) );
  NAND3_X1 U14990 ( .A1(n13291), .A2(n13305), .A3(n13290), .ZN(n13292) );
  NAND2_X1 U14991 ( .A1(n13293), .A2(n13292), .ZN(n13296) );
  NAND2_X1 U14992 ( .A1(n13294), .A2(n13298), .ZN(n13295) );
  NAND2_X1 U14993 ( .A1(n13296), .A2(n13295), .ZN(n13300) );
  AOI22_X1 U14994 ( .A1(n13301), .A2(n13298), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21614), .ZN(n13299) );
  NAND2_X1 U14995 ( .A1(n13300), .A2(n13299), .ZN(n13303) );
  NAND2_X1 U14996 ( .A1(n13301), .A2(n13304), .ZN(n13302) );
  NAND2_X1 U14997 ( .A1(n13303), .A2(n13302), .ZN(n13307) );
  NAND2_X1 U14998 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  NAND2_X1 U14999 ( .A1(n21915), .A2(n21657), .ZN(n14274) );
  NAND3_X1 U15000 ( .A1(n13308), .A2(n21660), .A3(n14274), .ZN(n13309) );
  NAND3_X1 U15001 ( .A1(n13309), .A2(n14272), .A3(n12967), .ZN(n13310) );
  NAND2_X1 U15002 ( .A1(n21623), .A2(n13310), .ZN(n13311) );
  MUX2_X1 U15003 ( .A(n13312), .B(n13311), .S(n13056), .Z(n13320) );
  OR2_X1 U15004 ( .A1(n13647), .A2(n12972), .ZN(n13319) );
  NOR2_X1 U15005 ( .A1(n12984), .A2(n13442), .ZN(n13452) );
  NAND2_X1 U15006 ( .A1(n13452), .A2(n21716), .ZN(n15287) );
  NOR2_X1 U15007 ( .A1(n12972), .A2(n13441), .ZN(n13700) );
  INV_X1 U15008 ( .A(n13313), .ZN(n13314) );
  OR2_X1 U15009 ( .A1(n13700), .A2(n13314), .ZN(n13317) );
  OR2_X1 U15010 ( .A1(n13442), .A2(n13315), .ZN(n13316) );
  AND2_X1 U15011 ( .A1(n11398), .A2(n13316), .ZN(n13439) );
  NAND2_X1 U15012 ( .A1(n13317), .A2(n13439), .ZN(n13324) );
  AOI21_X1 U15013 ( .B1(n12898), .B2(n12978), .A(n21716), .ZN(n13318) );
  AOI21_X1 U15014 ( .B1(n15287), .B2(n13324), .A(n13438), .ZN(n13654) );
  NAND3_X1 U15015 ( .A1(n13320), .A2(n13319), .A3(n13654), .ZN(n13322) );
  NAND2_X1 U15016 ( .A1(n13321), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21631) );
  INV_X1 U15017 ( .A(n21631), .ZN(n19965) );
  NOR2_X1 U15018 ( .A1(n13324), .A2(n13442), .ZN(n13779) );
  AND2_X1 U15019 ( .A1(n13700), .A2(n12985), .ZN(n13648) );
  NOR2_X1 U15020 ( .A1(n13779), .A2(n13648), .ZN(n15284) );
  NAND2_X1 U15021 ( .A1(n13325), .A2(n12978), .ZN(n13644) );
  OR2_X1 U15022 ( .A1(n13436), .A2(n12970), .ZN(n13326) );
  NAND4_X1 U15023 ( .A1(n13323), .A2(n15284), .A3(n13644), .A4(n13326), .ZN(
        n13327) );
  INV_X1 U15024 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21230) );
  NAND2_X1 U15025 ( .A1(n13423), .A2(n21230), .ZN(n13329) );
  INV_X1 U15026 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U15027 ( .A1(n13684), .A2(n13773), .ZN(n13328) );
  NAND3_X1 U15028 ( .A1(n13329), .A2(n13390), .A3(n13328), .ZN(n13330) );
  NAND2_X1 U15029 ( .A1(n13331), .A2(n13330), .ZN(n13334) );
  NAND2_X1 U15030 ( .A1(n13423), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13333) );
  INV_X1 U15031 ( .A(n13342), .ZN(n13348) );
  INV_X1 U15032 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13691) );
  NAND2_X1 U15033 ( .A1(n13342), .A2(n13691), .ZN(n13332) );
  NAND2_X1 U15034 ( .A1(n13333), .A2(n13332), .ZN(n13688) );
  XNOR2_X1 U15035 ( .A(n13334), .B(n13688), .ZN(n13769) );
  NAND2_X1 U15036 ( .A1(n13769), .A2(n13684), .ZN(n13771) );
  OR2_X1 U15037 ( .A1(n13429), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13339) );
  INV_X1 U15038 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21237) );
  NAND2_X1 U15039 ( .A1(n13423), .A2(n21237), .ZN(n13337) );
  INV_X1 U15040 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U15041 ( .A1(n13684), .A2(n13335), .ZN(n13336) );
  NAND3_X1 U15042 ( .A1(n13337), .A2(n13390), .A3(n13336), .ZN(n13338) );
  MUX2_X1 U15043 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13343) );
  OAI21_X1 U15044 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13687), .A(
        n13343), .ZN(n14096) );
  OR2_X1 U15045 ( .A1(n13429), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U15046 ( .A1(n13342), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13344) );
  NAND2_X1 U15047 ( .A1(n13423), .A2(n13344), .ZN(n13345) );
  OAI21_X1 U15048 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n13770), .A(n13345), .ZN(
        n13346) );
  NAND2_X1 U15049 ( .A1(n13347), .A2(n13346), .ZN(n14146) );
  NAND2_X1 U15050 ( .A1(n13390), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13349) );
  OAI211_X1 U15051 ( .C1(n13770), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13423), .B(
        n13349), .ZN(n13350) );
  OAI21_X1 U15052 ( .B1(n13420), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13350), .ZN(
        n19886) );
  OR2_X1 U15053 ( .A1(n13429), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U15054 ( .A1(n13423), .A2(n21262), .ZN(n13352) );
  INV_X1 U15055 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19883) );
  NAND2_X1 U15056 ( .A1(n13684), .A2(n19883), .ZN(n13351) );
  NAND3_X1 U15057 ( .A1(n13352), .A2(n13390), .A3(n13351), .ZN(n13353) );
  MUX2_X1 U15058 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13355) );
  OAI21_X1 U15059 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13687), .A(
        n13355), .ZN(n13356) );
  INV_X1 U15060 ( .A(n13356), .ZN(n14256) );
  OR2_X1 U15061 ( .A1(n13429), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U15062 ( .A1(n13423), .A2(n21292), .ZN(n13358) );
  INV_X1 U15063 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U15064 ( .A1(n13684), .A2(n14427), .ZN(n13357) );
  NAND3_X1 U15065 ( .A1(n13358), .A2(n13390), .A3(n13357), .ZN(n13359) );
  NAND2_X1 U15066 ( .A1(n13360), .A2(n13359), .ZN(n14424) );
  MUX2_X1 U15067 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13361) );
  OAI21_X1 U15068 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13687), .A(
        n13361), .ZN(n14461) );
  MUX2_X1 U15069 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13362) );
  OAI21_X1 U15070 ( .B1(n13687), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n13362), .ZN(n14796) );
  INV_X1 U15071 ( .A(n14796), .ZN(n13368) );
  OR2_X1 U15072 ( .A1(n13429), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U15073 ( .A1(n13423), .A2(n15705), .ZN(n13365) );
  INV_X1 U15074 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13363) );
  NAND2_X1 U15075 ( .A1(n13684), .A2(n13363), .ZN(n13364) );
  NAND3_X1 U15076 ( .A1(n13365), .A2(n13390), .A3(n13364), .ZN(n13366) );
  NAND2_X1 U15077 ( .A1(n13367), .A2(n13366), .ZN(n14795) );
  NAND2_X1 U15078 ( .A1(n13368), .A2(n14795), .ZN(n13369) );
  MUX2_X1 U15079 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13371) );
  OR2_X1 U15080 ( .A1(n13687), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13370) );
  AND2_X1 U15081 ( .A1(n13371), .A2(n13370), .ZN(n14682) );
  OR2_X1 U15082 ( .A1(n13429), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U15083 ( .A1(n13390), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13372) );
  NAND2_X1 U15084 ( .A1(n13423), .A2(n13372), .ZN(n13373) );
  OAI21_X1 U15085 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n13770), .A(n13373), .ZN(
        n13374) );
  NAND2_X1 U15086 ( .A1(n13375), .A2(n13374), .ZN(n14719) );
  NAND2_X1 U15087 ( .A1(n14682), .A2(n14719), .ZN(n13376) );
  OR2_X1 U15088 ( .A1(n13429), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U15089 ( .A1(n13423), .A2(n13377), .ZN(n13379) );
  INV_X1 U15090 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15392) );
  NAND2_X1 U15091 ( .A1(n13684), .A2(n15392), .ZN(n13378) );
  NAND3_X1 U15092 ( .A1(n13379), .A2(n13390), .A3(n13378), .ZN(n13380) );
  NAND2_X1 U15093 ( .A1(n13381), .A2(n13380), .ZN(n14790) );
  MUX2_X1 U15094 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13382) );
  OAI21_X1 U15095 ( .B1(n13687), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n13382), .ZN(n15503) );
  OR2_X1 U15096 ( .A1(n13429), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n13386) );
  INV_X1 U15097 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21362) );
  NAND2_X1 U15098 ( .A1(n13423), .A2(n21362), .ZN(n13384) );
  INV_X1 U15099 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21508) );
  NAND2_X1 U15100 ( .A1(n13684), .A2(n21508), .ZN(n13383) );
  NAND3_X1 U15101 ( .A1(n13384), .A2(n13390), .A3(n13383), .ZN(n13385) );
  MUX2_X1 U15102 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13387) );
  OAI21_X1 U15103 ( .B1(n13687), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13387), .ZN(n15385) );
  OR2_X1 U15104 ( .A1(n13429), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n13393) );
  INV_X1 U15105 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U15106 ( .A1(n13423), .A2(n13388), .ZN(n13391) );
  INV_X1 U15107 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21521) );
  NAND2_X1 U15108 ( .A1(n13684), .A2(n21521), .ZN(n13389) );
  NAND3_X1 U15109 ( .A1(n13391), .A2(n13390), .A3(n13389), .ZN(n13392) );
  AND2_X1 U15110 ( .A1(n13393), .A2(n13392), .ZN(n15483) );
  NAND2_X1 U15111 ( .A1(n13390), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13394) );
  OAI211_X1 U15112 ( .C1(n13770), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13423), .B(
        n13394), .ZN(n13395) );
  OAI21_X1 U15113 ( .B1(n13420), .B2(P1_EBX_REG_19__SCAN_IN), .A(n13395), .ZN(
        n15476) );
  OR2_X1 U15114 ( .A1(n13429), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n13399) );
  INV_X1 U15115 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19958) );
  NAND2_X1 U15116 ( .A1(n13423), .A2(n19958), .ZN(n13397) );
  INV_X1 U15117 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U15118 ( .A1(n13684), .A2(n15469), .ZN(n13396) );
  NAND3_X1 U15119 ( .A1(n13397), .A2(n13390), .A3(n13396), .ZN(n13398) );
  NAND2_X1 U15120 ( .A1(n13399), .A2(n13398), .ZN(n15372) );
  MUX2_X1 U15121 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13400) );
  OAI21_X1 U15122 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13687), .A(
        n13400), .ZN(n15467) );
  INV_X1 U15123 ( .A(n15467), .ZN(n13401) );
  OR2_X1 U15124 ( .A1(n13429), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13407) );
  INV_X1 U15125 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13402) );
  NAND2_X1 U15126 ( .A1(n13423), .A2(n13402), .ZN(n13405) );
  INV_X1 U15127 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U15128 ( .A1(n13684), .A2(n13403), .ZN(n13404) );
  NAND3_X1 U15129 ( .A1(n13405), .A2(n13390), .A3(n13404), .ZN(n13406) );
  AND2_X1 U15130 ( .A1(n13407), .A2(n13406), .ZN(n15457) );
  MUX2_X1 U15131 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13408) );
  OAI21_X1 U15132 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13687), .A(
        n13408), .ZN(n15452) );
  OR2_X1 U15133 ( .A1(n13429), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U15134 ( .A1(n13423), .A2(n13409), .ZN(n13411) );
  INV_X1 U15135 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21579) );
  NAND2_X1 U15136 ( .A1(n13684), .A2(n21579), .ZN(n13410) );
  NAND3_X1 U15137 ( .A1(n13411), .A2(n13342), .A3(n13410), .ZN(n13412) );
  NAND2_X1 U15138 ( .A1(n13413), .A2(n13412), .ZN(n15443) );
  MUX2_X1 U15139 ( .A(n13420), .B(n13390), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13414) );
  OAI21_X1 U15140 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13687), .A(
        n13414), .ZN(n15439) );
  INV_X1 U15141 ( .A(n15439), .ZN(n13415) );
  OR2_X1 U15142 ( .A1(n13429), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n13419) );
  NAND2_X1 U15143 ( .A1(n13423), .A2(n15747), .ZN(n13417) );
  INV_X1 U15144 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15360) );
  NAND2_X1 U15145 ( .A1(n13684), .A2(n15360), .ZN(n13416) );
  NAND3_X1 U15146 ( .A1(n13417), .A2(n13342), .A3(n13416), .ZN(n13418) );
  AND2_X1 U15147 ( .A1(n13419), .A2(n13418), .ZN(n15355) );
  MUX2_X1 U15148 ( .A(n13420), .B(n13342), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13421) );
  OAI21_X1 U15149 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13687), .A(
        n13421), .ZN(n15345) );
  OR2_X1 U15150 ( .A1(n13429), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13426) );
  INV_X1 U15151 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U15152 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  OAI211_X1 U15153 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13770), .A(n13424), .B(
        n13342), .ZN(n13425) );
  NAND2_X1 U15154 ( .A1(n13426), .A2(n13425), .ZN(n15331) );
  INV_X1 U15155 ( .A(n13687), .ZN(n13428) );
  INV_X1 U15156 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13461) );
  NOR2_X1 U15157 ( .A1(n13770), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13427) );
  AOI21_X1 U15158 ( .B1(n13428), .B2(n13461), .A(n13427), .ZN(n15247) );
  INV_X1 U15159 ( .A(n13429), .ZN(n13430) );
  INV_X1 U15160 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U15161 ( .A1(n15247), .A2(n13342), .B1(n13430), .B2(n15322), .ZN(
        n15319) );
  AND2_X1 U15162 ( .A1(n13770), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13431) );
  AOI21_X1 U15163 ( .B1(n13687), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13431), .ZN(
        n15249) );
  OAI22_X1 U15164 ( .A1(n13687), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n13770), .ZN(n13432) );
  NAND2_X1 U15165 ( .A1(n13308), .A2(n21195), .ZN(n13434) );
  OAI21_X1 U15166 ( .B1(n13436), .B2(n13435), .A(n13434), .ZN(n13437) );
  INV_X1 U15167 ( .A(n13438), .ZN(n13449) );
  INV_X1 U15168 ( .A(n13439), .ZN(n13440) );
  NAND2_X1 U15169 ( .A1(n13440), .A2(n13348), .ZN(n13448) );
  INV_X1 U15170 ( .A(n14275), .ZN(n13699) );
  AOI22_X1 U15171 ( .A1(n13699), .A2(n13442), .B1(n13441), .B2(n14272), .ZN(
        n13445) );
  AND2_X1 U15172 ( .A1(n12967), .A2(n12965), .ZN(n13443) );
  OAI21_X1 U15173 ( .B1(n12974), .B2(n13443), .A(n12978), .ZN(n13444) );
  AND2_X1 U15174 ( .A1(n13445), .A2(n13444), .ZN(n13447) );
  AND4_X1 U15175 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        n13694) );
  OAI21_X1 U15176 ( .B1(n13450), .B2(n14272), .A(n13694), .ZN(n13451) );
  INV_X1 U15177 ( .A(n21206), .ZN(n13453) );
  NAND2_X1 U15178 ( .A1(n13452), .A2(n13699), .ZN(n14039) );
  INV_X1 U15179 ( .A(n14039), .ZN(n15794) );
  NAND2_X1 U15180 ( .A1(n13457), .A2(n15794), .ZN(n21367) );
  NOR2_X1 U15181 ( .A1(n21248), .A2(n13106), .ZN(n21243) );
  NAND3_X1 U15182 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21243), .ZN(n21275) );
  NOR2_X1 U15183 ( .A1(n21264), .A2(n21275), .ZN(n21277) );
  NOR3_X1 U15184 ( .A1(n21292), .A2(n21284), .A3(n21262), .ZN(n21294) );
  NAND2_X1 U15185 ( .A1(n21277), .A2(n21294), .ZN(n21296) );
  NAND2_X1 U15186 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21304) );
  NOR2_X1 U15187 ( .A1(n21296), .A2(n21304), .ZN(n21316) );
  NAND3_X1 U15188 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n21316), .ZN(n21205) );
  INV_X1 U15189 ( .A(n21205), .ZN(n21332) );
  INV_X1 U15190 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13454) );
  NOR3_X1 U15191 ( .A1(n13217), .A2(n21362), .A3(n13454), .ZN(n21342) );
  INV_X1 U15192 ( .A(n21342), .ZN(n13455) );
  NAND2_X1 U15193 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21336) );
  NOR3_X1 U15194 ( .A1(n13388), .A2(n13455), .A3(n21336), .ZN(n15778) );
  AND2_X1 U15195 ( .A1(n21332), .A2(n15778), .ZN(n13463) );
  INV_X1 U15196 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21228) );
  INV_X1 U15197 ( .A(n13457), .ZN(n13456) );
  NOR2_X1 U15198 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21872) );
  NAND2_X1 U15199 ( .A1(n21908), .A2(n16765), .ZN(n19967) );
  AOI22_X1 U15200 ( .A1(n21206), .A2(n21228), .B1(n13456), .B2(n21373), .ZN(
        n21300) );
  OAI21_X1 U15201 ( .B1(n21333), .B2(n13463), .A(n21300), .ZN(n15784) );
  AND2_X1 U15202 ( .A1(n15780), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13464) );
  OAI21_X1 U15203 ( .B1(n21228), .B2(n21230), .A(n21237), .ZN(n21241) );
  NAND2_X1 U15204 ( .A1(n21243), .A2(n21241), .ZN(n21268) );
  NOR2_X1 U15205 ( .A1(n21264), .A2(n21268), .ZN(n21254) );
  NAND2_X1 U15206 ( .A1(n21294), .A2(n21254), .ZN(n21298) );
  NOR2_X1 U15207 ( .A1(n21304), .A2(n21298), .ZN(n15776) );
  NAND2_X1 U15208 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15776), .ZN(
        n21313) );
  NOR2_X1 U15209 ( .A1(n13214), .A2(n21313), .ZN(n21204) );
  NAND2_X1 U15210 ( .A1(n15778), .A2(n21204), .ZN(n15785) );
  NOR2_X1 U15211 ( .A1(n15785), .A2(n15763), .ZN(n13458) );
  AND2_X1 U15212 ( .A1(n13700), .A2(n13684), .ZN(n15282) );
  AOI21_X1 U15213 ( .B1(n13464), .B2(n13458), .A(n21389), .ZN(n13459) );
  NOR2_X1 U15214 ( .A1(n15784), .A2(n13459), .ZN(n15762) );
  INV_X1 U15215 ( .A(n15762), .ZN(n15768) );
  NOR2_X1 U15216 ( .A1(n15768), .A2(n21337), .ZN(n15726) );
  INV_X1 U15217 ( .A(n21333), .ZN(n21297) );
  NAND2_X1 U15218 ( .A1(n21297), .A2(n15626), .ZN(n13460) );
  OAI211_X1 U15219 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n21256), .A(
        n15762), .B(n13460), .ZN(n15743) );
  NAND2_X1 U15220 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13468) );
  NOR2_X1 U15221 ( .A1(n15743), .A2(n13468), .ZN(n15725) );
  AOI21_X1 U15222 ( .B1(n15725), .B2(n15724), .A(n15726), .ZN(n15715) );
  AOI21_X1 U15223 ( .B1(n13461), .B2(n21337), .A(n15715), .ZN(n15253) );
  OAI21_X1 U15224 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15726), .A(
        n15253), .ZN(n13472) );
  INV_X1 U15225 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n16841) );
  NOR2_X1 U15226 ( .A1(n21373), .A2(n16841), .ZN(n15167) );
  INV_X1 U15227 ( .A(n21367), .ZN(n13462) );
  NOR2_X1 U15228 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13462), .ZN(
        n21388) );
  NAND2_X1 U15229 ( .A1(n13463), .A2(n21265), .ZN(n15779) );
  INV_X1 U15230 ( .A(n13464), .ZN(n13465) );
  NOR2_X1 U15231 ( .A1(n15779), .A2(n13465), .ZN(n13467) );
  NOR3_X1 U15232 ( .A1(n21256), .A2(n15785), .A3(n13465), .ZN(n13466) );
  NOR2_X1 U15233 ( .A1(n13467), .A2(n13466), .ZN(n15771) );
  NOR2_X1 U15234 ( .A1(n15771), .A2(n15626), .ZN(n15757) );
  INV_X1 U15235 ( .A(n13468), .ZN(n13469) );
  NAND2_X1 U15236 ( .A1(n15757), .A2(n13469), .ZN(n15738) );
  INV_X1 U15237 ( .A(n15724), .ZN(n13470) );
  NOR2_X1 U15238 ( .A1(n15738), .A2(n13470), .ZN(n15713) );
  AND4_X1 U15239 ( .A1(n15713), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n13706), .ZN(n13471) );
  AOI211_X1 U15240 ( .C1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13472), .A(
        n15167), .B(n13471), .ZN(n13473) );
  NOR4_X1 U15241 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13477) );
  NOR4_X1 U15242 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13476) );
  NOR4_X1 U15243 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13475) );
  NOR4_X1 U15244 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13474) );
  AND4_X1 U15245 ( .A1(n13477), .A2(n13476), .A3(n13475), .A4(n13474), .ZN(
        n13482) );
  NOR4_X1 U15246 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13480) );
  NOR4_X1 U15247 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13479) );
  NOR4_X1 U15248 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13478) );
  INV_X1 U15249 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19817) );
  AND4_X1 U15250 ( .A1(n13480), .A2(n13479), .A3(n13478), .A4(n19817), .ZN(
        n13481) );
  NAND2_X1 U15251 ( .A1(n13482), .A2(n13481), .ZN(n13483) );
  AND2_X2 U15252 ( .A1(n13483), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15237)
         );
  INV_X1 U15253 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20015) );
  INV_X1 U15254 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n16917) );
  NOR4_X1 U15255 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20015), .A4(n16917), .ZN(n13485) );
  NOR4_X1 U15256 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13484) );
  NAND3_X1 U15257 ( .A1(n15237), .A2(n13485), .A3(n13484), .ZN(U214) );
  NOR4_X1 U15258 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13489) );
  NOR4_X1 U15259 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13488) );
  NOR4_X1 U15260 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13487) );
  NOR4_X1 U15261 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13486) );
  AND4_X1 U15262 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        n13494) );
  NOR4_X1 U15263 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13492) );
  NOR4_X1 U15264 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13491) );
  NOR4_X1 U15265 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13490) );
  INV_X1 U15266 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17113) );
  AND4_X1 U15267 ( .A1(n13492), .A2(n13491), .A3(n13490), .A4(n17113), .ZN(
        n13493) );
  NAND2_X1 U15268 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  NOR2_X1 U15269 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13497) );
  NOR4_X1 U15270 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13496) );
  NAND4_X1 U15271 ( .A1(n13497), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13496), .ZN(n13498) );
  OR2_X1 U15272 ( .A1(n16187), .A2(n13498), .ZN(n19972) );
  INV_X2 U15273 ( .A(U214), .ZN(n20006) );
  OR2_X1 U15274 ( .A1(n19972), .A2(n20006), .ZN(U212) );
  NOR2_X1 U15275 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13498), .ZN(n18564)
         );
  INV_X1 U15276 ( .A(n18535), .ZN(n18532) );
  NOR2_X1 U15277 ( .A1(n13508), .A2(n13711), .ZN(n18049) );
  INV_X1 U15278 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13502) );
  INV_X1 U15279 ( .A(n15824), .ZN(n13501) );
  OR2_X1 U15280 ( .A1(n13500), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U15281 ( .C1(n18049), .C2(n13502), .A(n13501), .B(n13509), .ZN(
        P2_U2814) );
  INV_X1 U15282 ( .A(n15288), .ZN(n13503) );
  NOR3_X1 U15283 ( .A1(n15287), .A2(n21631), .A3(n13503), .ZN(n13506) );
  INV_X1 U15284 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13505) );
  AND2_X1 U15285 ( .A1(n13325), .A2(n19965), .ZN(n13504) );
  OAI211_X1 U15286 ( .C1(n13506), .C2(n13505), .A(n13557), .B(n19967), .ZN(
        P1_U2801) );
  INV_X1 U15287 ( .A(n14012), .ZN(n13507) );
  INV_X1 U15288 ( .A(n16965), .ZN(n18018) );
  INV_X1 U15289 ( .A(n13509), .ZN(n13510) );
  OAI21_X1 U15290 ( .B1(n13510), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18018), 
        .ZN(n13511) );
  OAI21_X1 U15291 ( .B1(n13512), .B2(n18018), .A(n13511), .ZN(P2_U3612) );
  NAND2_X1 U15292 ( .A1(n15288), .A2(n21915), .ZN(n13513) );
  OR2_X1 U15293 ( .A1(n15287), .A2(n13513), .ZN(n13645) );
  NOR2_X1 U15294 ( .A1(n14039), .A2(n21631), .ZN(n13514) );
  NAND2_X1 U15295 ( .A1(n21623), .A2(n13514), .ZN(n14117) );
  OAI211_X1 U15296 ( .C1(n13645), .C2(n21631), .A(n13557), .B(n14117), .ZN(
        n21199) );
  INV_X1 U15297 ( .A(n21199), .ZN(n13516) );
  INV_X1 U15298 ( .A(n19967), .ZN(n14464) );
  OAI21_X1 U15299 ( .B1(n14464), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13516), 
        .ZN(n13515) );
  OAI21_X1 U15300 ( .B1(n13517), .B2(n13516), .A(n13515), .ZN(P1_U3487) );
  INV_X1 U15301 ( .A(n13521), .ZN(n13518) );
  AOI222_X1 U15302 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13521), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13520), .C1(n13519), .C2(
        n13518), .ZN(n18423) );
  OAI21_X1 U15303 ( .B1(n18520), .B2(n13523), .A(n13522), .ZN(n14018) );
  NAND2_X1 U15304 ( .A1(n18538), .A2(n16011), .ZN(n17014) );
  NAND2_X1 U15305 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14336) );
  INV_X1 U15306 ( .A(n14336), .ZN(n13524) );
  NOR2_X1 U15307 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13524), .ZN(n17043) );
  AND2_X1 U15308 ( .A1(n17043), .A2(n18022), .ZN(n13525) );
  NAND2_X1 U15309 ( .A1(n18022), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14032) );
  INV_X1 U15310 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21639) );
  NAND2_X1 U15311 ( .A1(n21639), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13526) );
  NAND2_X1 U15312 ( .A1(n14032), .A2(n13526), .ZN(n13537) );
  NAND2_X1 U15313 ( .A1(n18538), .A2(n15968), .ZN(n17024) );
  OAI21_X1 U15314 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13528), .A(
        n13527), .ZN(n18424) );
  INV_X1 U15315 ( .A(n18240), .ZN(n16539) );
  NAND2_X1 U15316 ( .A1(n16539), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n18433) );
  OAI21_X1 U15317 ( .B1(n17024), .B2(n18424), .A(n18433), .ZN(n13530) );
  NOR2_X1 U15318 ( .A1(n17018), .A2(n13531), .ZN(n13529) );
  AOI211_X1 U15319 ( .C1(n17005), .C2(n13531), .A(n13530), .B(n13529), .ZN(
        n13533) );
  AND2_X1 U15320 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16713) );
  NAND2_X1 U15321 ( .A1(n17021), .A2(n18427), .ZN(n13532) );
  OAI211_X1 U15322 ( .C1(n18423), .C2(n17014), .A(n13533), .B(n13532), .ZN(
        P2_U3013) );
  AOI21_X1 U15323 ( .B1(n18418), .B2(n13535), .A(n13534), .ZN(n18414) );
  NOR2_X1 U15324 ( .A1(n18475), .A2(n11137), .ZN(n18413) );
  XNOR2_X1 U15325 ( .A(n18030), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18411) );
  NOR2_X1 U15326 ( .A1(n17014), .A2(n18411), .ZN(n13536) );
  AOI211_X1 U15327 ( .C1(n18414), .C2(n17035), .A(n18413), .B(n13536), .ZN(
        n13539) );
  OAI21_X1 U15328 ( .B1(n17031), .B2(n13537), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13538) );
  OAI211_X1 U15329 ( .C1(n17038), .C2(n18036), .A(n13539), .B(n13538), .ZN(
        P2_U3014) );
  INV_X1 U15330 ( .A(n13713), .ZN(n13541) );
  NOR2_X1 U15331 ( .A1(n13711), .A2(n14028), .ZN(n13540) );
  NAND2_X1 U15332 ( .A1(n13541), .A2(n13540), .ZN(n13545) );
  AND2_X1 U15333 ( .A1(n12411), .A2(n18527), .ZN(n14010) );
  NAND2_X1 U15334 ( .A1(n14012), .A2(n14010), .ZN(n13542) );
  NOR2_X1 U15335 ( .A1(n14014), .A2(n13542), .ZN(n13543) );
  AOI21_X1 U15336 ( .B1(n14335), .B2(n14005), .A(n13543), .ZN(n13745) );
  INV_X1 U15337 ( .A(n14335), .ZN(n14006) );
  INV_X1 U15338 ( .A(n13956), .ZN(n14004) );
  NAND2_X1 U15339 ( .A1(n14006), .A2(n14004), .ZN(n13735) );
  NAND4_X1 U15340 ( .A1(n13545), .A2(n13544), .A3(n13745), .A4(n13735), .ZN(
        n14021) );
  NAND2_X1 U15341 ( .A1(n14021), .A2(n18535), .ZN(n13547) );
  NOR2_X1 U15342 ( .A1(n18022), .A2(n14336), .ZN(n16716) );
  AOI22_X1 U15343 ( .A1(n18022), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(
        P2_FLUSH_REG_SCAN_IN), .B2(n16716), .ZN(n13546) );
  NAND2_X1 U15344 ( .A1(n13547), .A2(n13546), .ZN(n16695) );
  NOR2_X1 U15345 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16687) );
  INV_X1 U15346 ( .A(n16687), .ZN(n18511) );
  INV_X1 U15347 ( .A(n13548), .ZN(n13549) );
  OR3_X1 U15348 ( .A1(n13711), .A2(n13549), .A3(n16011), .ZN(n14015) );
  OR3_X1 U15349 ( .A1(n16690), .A2(n18511), .A3(n14015), .ZN(n13550) );
  OAI21_X1 U15350 ( .B1(n14020), .B2(n16695), .A(n13550), .ZN(P2_U3595) );
  NAND2_X1 U15351 ( .A1(n15824), .A2(n15968), .ZN(n15821) );
  INV_X1 U15352 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17111) );
  AND2_X1 U15353 ( .A1(n16011), .A2(n18527), .ZN(n13551) );
  NAND2_X2 U15354 ( .A1(n15824), .A2(n13551), .ZN(n19591) );
  INV_X1 U15355 ( .A(n19591), .ZN(n13552) );
  INV_X1 U15356 ( .A(n19587), .ZN(n18999) );
  INV_X1 U15357 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13555) );
  INV_X1 U15358 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13666) );
  OR2_X1 U15359 ( .A1(n16187), .A2(n13666), .ZN(n13554) );
  NAND2_X1 U15360 ( .A1(n14180), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13553) );
  AND2_X1 U15361 ( .A1(n13554), .A2(n13553), .ZN(n14216) );
  OAI222_X1 U15362 ( .A1(n15821), .A2(n17111), .B1(n18999), .B2(n13555), .C1(
        n19591), .C2(n14216), .ZN(P2_U2982) );
  INV_X1 U15363 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19801) );
  NOR2_X1 U15364 ( .A1(n21195), .A2(n21660), .ZN(n13556) );
  INV_X2 U15365 ( .A(n13669), .ZN(n13640) );
  INV_X1 U15366 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n19985) );
  NAND2_X1 U15367 ( .A1(n15237), .A2(n19985), .ZN(n13558) );
  OAI21_X1 U15368 ( .B1(n15237), .B2(DATAI_9_), .A(n13558), .ZN(n15537) );
  INV_X1 U15369 ( .A(n15537), .ZN(n13559) );
  NAND2_X1 U15370 ( .A1(n13624), .A2(n13559), .ZN(n13575) );
  NAND2_X1 U15371 ( .A1(n13640), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13560) );
  OAI211_X1 U15372 ( .C1(n19801), .C2(n13603), .A(n13575), .B(n13560), .ZN(
        P1_U2961) );
  INV_X1 U15373 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19808) );
  INV_X1 U15374 ( .A(DATAI_12_), .ZN(n13561) );
  INV_X1 U15375 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14123) );
  MUX2_X1 U15376 ( .A(n13561), .B(n14123), .S(n15237), .Z(n15523) );
  INV_X1 U15377 ( .A(n15523), .ZN(n13562) );
  NAND2_X1 U15378 ( .A1(n13624), .A2(n13562), .ZN(n13631) );
  NAND2_X1 U15379 ( .A1(n13640), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13563) );
  OAI211_X1 U15380 ( .C1(n19808), .C2(n13603), .A(n13631), .B(n13563), .ZN(
        P1_U2964) );
  INV_X1 U15381 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19804) );
  INV_X1 U15382 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n19987) );
  NAND2_X1 U15383 ( .A1(n15237), .A2(n19987), .ZN(n13564) );
  OAI21_X1 U15384 ( .B1(n15237), .B2(DATAI_10_), .A(n13564), .ZN(n15532) );
  INV_X1 U15385 ( .A(n15532), .ZN(n13565) );
  NAND2_X1 U15386 ( .A1(n13624), .A2(n13565), .ZN(n13573) );
  NAND2_X1 U15387 ( .A1(n13640), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13566) );
  OAI211_X1 U15388 ( .C1(n19804), .C2(n13603), .A(n13573), .B(n13566), .ZN(
        P1_U2962) );
  INV_X1 U15389 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14308) );
  INV_X1 U15390 ( .A(DATAI_6_), .ZN(n13568) );
  NAND2_X1 U15391 ( .A1(n15237), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13567) );
  OAI21_X1 U15392 ( .B1(n15237), .B2(n13568), .A(n13567), .ZN(n22149) );
  NAND2_X1 U15393 ( .A1(n13624), .A2(n22149), .ZN(n13593) );
  NAND2_X1 U15394 ( .A1(n13640), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13569) );
  OAI211_X1 U15395 ( .C1(n14308), .C2(n13603), .A(n13593), .B(n13569), .ZN(
        P1_U2943) );
  INV_X1 U15396 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19810) );
  INV_X1 U15397 ( .A(DATAI_13_), .ZN(n16797) );
  INV_X1 U15398 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n19992) );
  MUX2_X1 U15399 ( .A(n16797), .B(n19992), .S(n15237), .Z(n15518) );
  INV_X1 U15400 ( .A(n15518), .ZN(n13570) );
  NAND2_X1 U15401 ( .A1(n13624), .A2(n13570), .ZN(n13621) );
  NAND2_X1 U15402 ( .A1(n13640), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13571) );
  OAI211_X1 U15403 ( .C1(n19810), .C2(n13603), .A(n13621), .B(n13571), .ZN(
        P1_U2965) );
  INV_X1 U15404 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U15405 ( .A1(n13640), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13572) );
  OAI211_X1 U15406 ( .C1(n14318), .C2(n13603), .A(n13573), .B(n13572), .ZN(
        P1_U2947) );
  INV_X1 U15407 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U15408 ( .A1(n13640), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13574) );
  OAI211_X1 U15409 ( .C1(n14314), .C2(n13603), .A(n13575), .B(n13574), .ZN(
        P1_U2946) );
  INV_X1 U15410 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19799) );
  INV_X1 U15411 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n19983) );
  NAND2_X1 U15412 ( .A1(n15237), .A2(n19983), .ZN(n13576) );
  OAI21_X1 U15413 ( .B1(n15237), .B2(DATAI_8_), .A(n13576), .ZN(n15541) );
  INV_X1 U15414 ( .A(n15541), .ZN(n13577) );
  NAND2_X1 U15415 ( .A1(n13624), .A2(n13577), .ZN(n13583) );
  NAND2_X1 U15416 ( .A1(n13640), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13578) );
  OAI211_X1 U15417 ( .C1(n19799), .C2(n13603), .A(n13583), .B(n13578), .ZN(
        P1_U2960) );
  INV_X1 U15418 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14297) );
  INV_X1 U15419 ( .A(DATAI_7_), .ZN(n13580) );
  NAND2_X1 U15420 ( .A1(n15237), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13579) );
  OAI21_X1 U15421 ( .B1(n15237), .B2(n13580), .A(n13579), .ZN(n22198) );
  NAND2_X1 U15422 ( .A1(n13624), .A2(n22198), .ZN(n13605) );
  NAND2_X1 U15423 ( .A1(n13640), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13581) );
  OAI211_X1 U15424 ( .C1(n14297), .C2(n13603), .A(n13605), .B(n13581), .ZN(
        P1_U2944) );
  INV_X1 U15425 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14306) );
  NAND2_X1 U15426 ( .A1(n13640), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13582) );
  OAI211_X1 U15427 ( .C1(n14306), .C2(n13603), .A(n13583), .B(n13582), .ZN(
        P1_U2945) );
  INV_X1 U15428 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19806) );
  INV_X1 U15429 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n19989) );
  NAND2_X1 U15430 ( .A1(n15237), .A2(n19989), .ZN(n13584) );
  OAI21_X1 U15431 ( .B1(n15237), .B2(DATAI_11_), .A(n13584), .ZN(n15527) );
  INV_X1 U15432 ( .A(n15527), .ZN(n13585) );
  NAND2_X1 U15433 ( .A1(n13624), .A2(n13585), .ZN(n13633) );
  NAND2_X1 U15434 ( .A1(n13640), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13586) );
  OAI211_X1 U15435 ( .C1(n19806), .C2(n13603), .A(n13633), .B(n13586), .ZN(
        P1_U2963) );
  INV_X1 U15436 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19812) );
  INV_X1 U15437 ( .A(DATAI_14_), .ZN(n16796) );
  INV_X1 U15438 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n19994) );
  MUX2_X1 U15439 ( .A(n16796), .B(n19994), .S(n15237), .Z(n15513) );
  INV_X1 U15440 ( .A(n15513), .ZN(n13587) );
  NAND2_X1 U15441 ( .A1(n13624), .A2(n13587), .ZN(n13627) );
  NAND2_X1 U15442 ( .A1(n13640), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13588) );
  OAI211_X1 U15443 ( .C1(n19812), .C2(n13603), .A(n13627), .B(n13588), .ZN(
        P1_U2966) );
  INV_X1 U15444 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19792) );
  INV_X1 U15445 ( .A(DATAI_5_), .ZN(n13590) );
  NAND2_X1 U15446 ( .A1(n15237), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13589) );
  OAI21_X1 U15447 ( .B1(n15237), .B2(n13590), .A(n13589), .ZN(n22101) );
  NAND2_X1 U15448 ( .A1(n13624), .A2(n22101), .ZN(n13629) );
  NAND2_X1 U15449 ( .A1(n13640), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n13591) );
  OAI211_X1 U15450 ( .C1(n19792), .C2(n13603), .A(n13629), .B(n13591), .ZN(
        P1_U2957) );
  INV_X1 U15451 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19794) );
  NAND2_X1 U15452 ( .A1(n13640), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n13592) );
  OAI211_X1 U15453 ( .C1(n19794), .C2(n13603), .A(n13593), .B(n13592), .ZN(
        P1_U2958) );
  INV_X1 U15454 ( .A(n13594), .ZN(n13595) );
  XNOR2_X1 U15455 ( .A(n13596), .B(n13595), .ZN(n18502) );
  NAND2_X1 U15456 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n16539), .ZN(n18506) );
  OAI21_X1 U15457 ( .B1(n17018), .B2(n15836), .A(n18506), .ZN(n13601) );
  AOI21_X1 U15458 ( .B1(n13531), .B2(n15836), .A(n14357), .ZN(n15835) );
  INV_X1 U15459 ( .A(n15835), .ZN(n13599) );
  XNOR2_X1 U15460 ( .A(n13598), .B(n13597), .ZN(n18493) );
  OAI22_X1 U15461 ( .A1(n17042), .A2(n13599), .B1(n17024), .B2(n18493), .ZN(
        n13600) );
  AOI211_X1 U15462 ( .C1(n18502), .C2(n17032), .A(n13601), .B(n13600), .ZN(
        n13602) );
  OAI21_X1 U15463 ( .B1(n11138), .B2(n17038), .A(n13602), .ZN(P2_U3012) );
  INV_X1 U15464 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19796) );
  NAND2_X1 U15465 ( .A1(n13640), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n13604) );
  OAI211_X1 U15466 ( .C1(n19796), .C2(n13603), .A(n13605), .B(n13604), .ZN(
        P1_U2959) );
  INV_X1 U15467 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14122) );
  INV_X1 U15468 ( .A(DATAI_2_), .ZN(n13607) );
  NAND2_X1 U15469 ( .A1(n15237), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13606) );
  OAI21_X1 U15470 ( .B1(n15237), .B2(n13607), .A(n13606), .ZN(n21959) );
  NAND2_X1 U15471 ( .A1(n13624), .A2(n21959), .ZN(n13616) );
  NAND2_X1 U15472 ( .A1(n13640), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13608) );
  OAI211_X1 U15473 ( .C1(n14122), .C2(n13603), .A(n13616), .B(n13608), .ZN(
        P1_U2939) );
  INV_X1 U15474 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19790) );
  INV_X1 U15475 ( .A(DATAI_4_), .ZN(n13610) );
  NAND2_X1 U15476 ( .A1(n15237), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13609) );
  OAI21_X1 U15477 ( .B1(n15237), .B2(n13610), .A(n13609), .ZN(n22054) );
  NAND2_X1 U15478 ( .A1(n13624), .A2(n22054), .ZN(n13635) );
  NAND2_X1 U15479 ( .A1(n13640), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n13611) );
  OAI211_X1 U15480 ( .C1(n19790), .C2(n13603), .A(n13635), .B(n13611), .ZN(
        P1_U2956) );
  INV_X1 U15481 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19788) );
  INV_X1 U15482 ( .A(DATAI_3_), .ZN(n13613) );
  NAND2_X1 U15483 ( .A1(n15237), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13612) );
  OAI21_X1 U15484 ( .B1(n15237), .B2(n13613), .A(n13612), .ZN(n22007) );
  NAND2_X1 U15485 ( .A1(n13624), .A2(n22007), .ZN(n13637) );
  NAND2_X1 U15486 ( .A1(n13640), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n13614) );
  OAI211_X1 U15487 ( .C1(n19788), .C2(n13603), .A(n13637), .B(n13614), .ZN(
        P1_U2955) );
  INV_X1 U15488 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19786) );
  NAND2_X1 U15489 ( .A1(n13640), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n13615) );
  OAI211_X1 U15490 ( .C1(n19786), .C2(n13603), .A(n13616), .B(n13615), .ZN(
        P1_U2954) );
  INV_X1 U15491 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19784) );
  INV_X1 U15492 ( .A(DATAI_1_), .ZN(n13618) );
  NAND2_X1 U15493 ( .A1(n15237), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13617) );
  OAI21_X1 U15494 ( .B1(n15237), .B2(n13618), .A(n13617), .ZN(n21912) );
  NAND2_X1 U15495 ( .A1(n13624), .A2(n21912), .ZN(n13639) );
  NAND2_X1 U15496 ( .A1(n13640), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n13619) );
  OAI211_X1 U15497 ( .C1(n19784), .C2(n13603), .A(n13639), .B(n13619), .ZN(
        P1_U2953) );
  INV_X1 U15498 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14324) );
  NAND2_X1 U15499 ( .A1(n13640), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13620) );
  OAI211_X1 U15500 ( .C1(n14324), .C2(n13603), .A(n13621), .B(n13620), .ZN(
        P1_U2950) );
  INV_X1 U15501 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19782) );
  INV_X1 U15502 ( .A(DATAI_0_), .ZN(n13623) );
  NAND2_X1 U15503 ( .A1(n15237), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13622) );
  OAI21_X1 U15504 ( .B1(n15237), .B2(n13623), .A(n13622), .ZN(n21711) );
  NAND2_X1 U15505 ( .A1(n13624), .A2(n21711), .ZN(n13642) );
  NAND2_X1 U15506 ( .A1(n13640), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n13625) );
  OAI211_X1 U15507 ( .C1(n19782), .C2(n13603), .A(n13642), .B(n13625), .ZN(
        P1_U2952) );
  INV_X1 U15508 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U15509 ( .A1(n13640), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13626) );
  OAI211_X1 U15510 ( .C1(n14316), .C2(n13603), .A(n13627), .B(n13626), .ZN(
        P1_U2951) );
  INV_X1 U15511 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U15512 ( .A1(n13640), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13628) );
  OAI211_X1 U15513 ( .C1(n14320), .C2(n13603), .A(n13629), .B(n13628), .ZN(
        P1_U2942) );
  INV_X1 U15514 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U15515 ( .A1(n13640), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13630) );
  OAI211_X1 U15516 ( .C1(n14312), .C2(n13603), .A(n13631), .B(n13630), .ZN(
        P1_U2949) );
  INV_X1 U15517 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U15518 ( .A1(n13640), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13632) );
  OAI211_X1 U15519 ( .C1(n14310), .C2(n13603), .A(n13633), .B(n13632), .ZN(
        P1_U2948) );
  INV_X1 U15520 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14327) );
  NAND2_X1 U15521 ( .A1(n13640), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13634) );
  OAI211_X1 U15522 ( .C1(n14327), .C2(n13603), .A(n13635), .B(n13634), .ZN(
        P1_U2941) );
  INV_X1 U15523 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U15524 ( .A1(n13640), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13636) );
  OAI211_X1 U15525 ( .C1(n14322), .C2(n13603), .A(n13637), .B(n13636), .ZN(
        P1_U2940) );
  INV_X1 U15526 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U15527 ( .A1(n13640), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13638) );
  OAI211_X1 U15528 ( .C1(n14120), .C2(n13603), .A(n13639), .B(n13638), .ZN(
        P1_U2938) );
  INV_X1 U15529 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U15530 ( .A1(n13640), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13641) );
  OAI211_X1 U15531 ( .C1(n14295), .C2(n13603), .A(n13642), .B(n13641), .ZN(
        P1_U2937) );
  AOI21_X1 U15532 ( .B1(n13645), .B2(n13644), .A(n13643), .ZN(n13646) );
  NAND2_X1 U15533 ( .A1(n13647), .A2(n13646), .ZN(n13650) );
  NAND2_X1 U15534 ( .A1(n21623), .A2(n13648), .ZN(n13649) );
  NAND2_X1 U15535 ( .A1(n13650), .A2(n13649), .ZN(n13826) );
  INV_X1 U15536 ( .A(n15282), .ZN(n13651) );
  OR2_X1 U15537 ( .A1(n21623), .A2(n13651), .ZN(n13656) );
  INV_X1 U15538 ( .A(n21657), .ZN(n15293) );
  INV_X1 U15539 ( .A(n13308), .ZN(n16760) );
  NAND2_X1 U15540 ( .A1(n14039), .A2(n16760), .ZN(n13652) );
  NAND4_X1 U15541 ( .A1(n21623), .A2(n15293), .A3(n21660), .A4(n13652), .ZN(
        n13655) );
  OR2_X1 U15542 ( .A1(n14275), .A2(n12965), .ZN(n13653) );
  NAND4_X1 U15543 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13657) );
  NOR2_X1 U15544 ( .A1(n13826), .A2(n13657), .ZN(n16736) );
  OR2_X1 U15545 ( .A1(n16736), .A2(n21631), .ZN(n13660) );
  NOR2_X1 U15546 ( .A1(n16765), .A2(n21898), .ZN(n14100) );
  NAND2_X1 U15547 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14100), .ZN(n21620) );
  INV_X1 U15548 ( .A(n21620), .ZN(n13658) );
  NAND2_X1 U15549 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13658), .ZN(n13659) );
  NAND2_X1 U15550 ( .A1(n13660), .A2(n13659), .ZN(n13663) );
  AOI21_X1 U15551 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21614), .A(n13663), 
        .ZN(n15809) );
  INV_X1 U15552 ( .A(n15809), .ZN(n13665) );
  INV_X1 U15553 ( .A(n21764), .ZN(n21849) );
  OR2_X1 U15554 ( .A1(n13661), .A2(n21849), .ZN(n13662) );
  XNOR2_X1 U15555 ( .A(n13662), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21412) );
  INV_X1 U15556 ( .A(n13323), .ZN(n14052) );
  NAND4_X1 U15557 ( .A1(n21412), .A2(n15797), .A3(n14052), .A4(n13663), .ZN(
        n13664) );
  OAI21_X1 U15558 ( .B1(n13665), .B2(n14054), .A(n13664), .ZN(P1_U3468) );
  INV_X1 U15559 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19816) );
  INV_X1 U15560 ( .A(DATAI_15_), .ZN(n13667) );
  MUX2_X1 U15561 ( .A(n13667), .B(n13666), .S(n15237), .Z(n15584) );
  INV_X1 U15562 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13668) );
  OAI222_X1 U15563 ( .A1(n13603), .A2(n19816), .B1(n13670), .B2(n15584), .C1(
        n13669), .C2(n13668), .ZN(P1_U2967) );
  BUF_X1 U15564 ( .A(n13671), .Z(n13672) );
  AOI21_X1 U15565 ( .B1(n13672), .B2(n12963), .A(n21898), .ZN(n13679) );
  INV_X1 U15566 ( .A(n13673), .ZN(n21748) );
  NAND2_X1 U15567 ( .A1(n21748), .A2(n14656), .ZN(n13678) );
  AND2_X1 U15568 ( .A1(n13674), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14132) );
  INV_X1 U15569 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13675) );
  OAI22_X1 U15570 ( .A1(n15087), .A2(n19782), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13675), .ZN(n13676) );
  AOI21_X1 U15571 ( .B1(n14132), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13676), .ZN(n13677) );
  NAND2_X1 U15572 ( .A1(n13678), .A2(n13677), .ZN(n13764) );
  NAND2_X1 U15573 ( .A1(n13679), .A2(n13764), .ZN(n13766) );
  OAI21_X1 U15574 ( .B1(n13679), .B2(n13764), .A(n13766), .ZN(n15415) );
  INV_X1 U15575 ( .A(n13700), .ZN(n13683) );
  INV_X1 U15576 ( .A(n13680), .ZN(n13682) );
  NAND3_X1 U15577 ( .A1(n12970), .A2(n22202), .A3(n13315), .ZN(n13681) );
  OAI21_X1 U15578 ( .B1(n21623), .B2(n13683), .A(n13824), .ZN(n13686) );
  AND2_X1 U15579 ( .A1(n13684), .A2(n19965), .ZN(n13685) );
  OR2_X1 U15580 ( .A1(n13687), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13689) );
  AND2_X1 U15581 ( .A1(n13689), .A2(n13688), .ZN(n15418) );
  INV_X1 U15582 ( .A(n15418), .ZN(n13690) );
  OAI222_X1 U15583 ( .A1(n15415), .A2(n15509), .B1(n13691), .B2(n19892), .C1(
        n13690), .C2(n15497), .ZN(P1_U2872) );
  NOR2_X1 U15584 ( .A1(n13692), .A2(n13308), .ZN(n13693) );
  AND2_X1 U15585 ( .A1(n13694), .A2(n13693), .ZN(n13697) );
  AND2_X1 U15586 ( .A1(n13323), .A2(n13695), .ZN(n13696) );
  NAND2_X1 U15587 ( .A1(n13697), .A2(n13696), .ZN(n14050) );
  INV_X1 U15588 ( .A(n14050), .ZN(n15796) );
  OR2_X1 U15589 ( .A1(n21850), .A2(n15796), .ZN(n13705) );
  NAND2_X1 U15590 ( .A1(n13697), .A2(n12974), .ZN(n14047) );
  INV_X1 U15591 ( .A(n14047), .ZN(n13703) );
  XNOR2_X1 U15592 ( .A(n13698), .B(n12819), .ZN(n13707) );
  XNOR2_X1 U15593 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13701) );
  NOR2_X1 U15594 ( .A1(n13699), .A2(n21195), .ZN(n15294) );
  NAND2_X1 U15595 ( .A1(n13700), .A2(n15294), .ZN(n14036) );
  OAI22_X1 U15596 ( .A1(n14039), .A2(n13701), .B1(n13707), .B2(n14036), .ZN(
        n13702) );
  AOI21_X1 U15597 ( .B1(n13703), .B2(n13707), .A(n13702), .ZN(n13704) );
  NAND2_X1 U15598 ( .A1(n13705), .A2(n13704), .ZN(n14051) );
  NOR2_X1 U15599 ( .A1(n16765), .A2(n21228), .ZN(n15799) );
  OAI22_X1 U15600 ( .A1(n21230), .A2(n13706), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15798) );
  INV_X1 U15601 ( .A(n15798), .ZN(n13708) );
  AOI222_X1 U15602 ( .A1(n14051), .A2(n15797), .B1(n15799), .B2(n13708), .C1(
        n13707), .C2(n15801), .ZN(n13710) );
  NAND2_X1 U15603 ( .A1(n15809), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13709) );
  OAI21_X1 U15604 ( .B1(n13710), .B2(n15809), .A(n13709), .ZN(P1_U3472) );
  INV_X1 U15605 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13717) );
  OR2_X1 U15606 ( .A1(n13711), .A2(n18532), .ZN(n13712) );
  OAI21_X1 U15607 ( .B1(n13713), .B2(n13712), .A(n15821), .ZN(n13714) );
  NAND2_X1 U15608 ( .A1(n17076), .A2(n13715), .ZN(n13905) );
  NOR2_X1 U15609 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14336), .ZN(n17096) );
  AOI22_X1 U15610 ( .A1(n17096), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U15611 ( .B1(n13717), .B2(n13905), .A(n13716), .ZN(P2_U2933) );
  INV_X1 U15612 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U15613 ( .A1(n17096), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13718) );
  OAI21_X1 U15614 ( .B1(n13719), .B2(n13905), .A(n13718), .ZN(P2_U2934) );
  OR2_X1 U15615 ( .A1(n13673), .A2(n15796), .ZN(n13721) );
  INV_X1 U15616 ( .A(n12972), .ZN(n15793) );
  NAND2_X1 U15617 ( .A1(n15793), .A2(n11111), .ZN(n13720) );
  NAND2_X1 U15618 ( .A1(n13721), .A2(n13720), .ZN(n16735) );
  INV_X1 U15619 ( .A(n15801), .ZN(n15805) );
  OAI22_X1 U15620 ( .A1(n15805), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16765), .ZN(n13722) );
  AOI21_X1 U15621 ( .B1(n16735), .B2(n15797), .A(n13722), .ZN(n13725) );
  OR2_X1 U15622 ( .A1(n14039), .A2(n11111), .ZN(n16733) );
  INV_X1 U15623 ( .A(n16733), .ZN(n13723) );
  AOI22_X1 U15624 ( .A1(n15809), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n15797), .B2(n13723), .ZN(n13724) );
  OAI21_X1 U15625 ( .B1(n15809), .B2(n13725), .A(n13724), .ZN(P1_U3474) );
  NAND2_X1 U15626 ( .A1(n11873), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U15627 ( .A1(n13726), .A2(n19183), .ZN(n13859) );
  AOI22_X1 U15628 ( .A1(n13859), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19200), .B2(n19146), .ZN(n13727) );
  NAND2_X1 U15629 ( .A1(n15990), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13844) );
  XNOR2_X1 U15630 ( .A(n13846), .B(n13844), .ZN(n13733) );
  INV_X1 U15631 ( .A(n14032), .ZN(n13837) );
  NAND2_X1 U15632 ( .A1(n13859), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13730) );
  NAND2_X1 U15633 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19179), .ZN(
        n19195) );
  INV_X1 U15634 ( .A(n19195), .ZN(n13729) );
  AOI21_X1 U15635 ( .B1(n19146), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13729), .ZN(n19114) );
  OR2_X1 U15636 ( .A1(n19114), .A2(n13500), .ZN(n19180) );
  NAND2_X1 U15637 ( .A1(n13730), .A2(n19180), .ZN(n13731) );
  INV_X1 U15638 ( .A(n19035), .ZN(n19049) );
  NAND2_X1 U15639 ( .A1(n13735), .A2(n13950), .ZN(n13736) );
  NAND2_X1 U15640 ( .A1(n16112), .A2(n11858), .ZN(n16115) );
  MUX2_X1 U15641 ( .A(n12136), .B(n13737), .S(n16112), .Z(n13738) );
  OAI21_X1 U15642 ( .B1(n19049), .B2(n16115), .A(n13738), .ZN(P2_U2886) );
  NAND2_X1 U15643 ( .A1(n16011), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13739) );
  AND4_X1 U15644 ( .A1(n13740), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13739), 
        .A4(n19183), .ZN(n13741) );
  MUX2_X1 U15645 ( .A(n13742), .B(n18036), .S(n16112), .Z(n13743) );
  OAI21_X1 U15646 ( .B1(n19034), .B2(n16115), .A(n13743), .ZN(P2_U2887) );
  NAND2_X1 U15647 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  XNOR2_X1 U15648 ( .A(n13748), .B(n13747), .ZN(n18410) );
  XNOR2_X1 U15649 ( .A(n19034), .B(n18410), .ZN(n13758) );
  NOR2_X1 U15650 ( .A1(n19465), .A2(n13749), .ZN(n14529) );
  NAND2_X1 U15651 ( .A1(n14529), .A2(n13750), .ZN(n19279) );
  INV_X1 U15652 ( .A(n19279), .ZN(n14176) );
  INV_X1 U15653 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13751) );
  OR2_X1 U15654 ( .A1(n16187), .A2(n13751), .ZN(n13753) );
  NAND2_X1 U15655 ( .A1(n16187), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13752) );
  AND2_X1 U15656 ( .A1(n13753), .A2(n13752), .ZN(n19595) );
  INV_X1 U15657 ( .A(n19595), .ZN(n13756) );
  OR2_X1 U15658 ( .A1(n19465), .A2(n11858), .ZN(n19467) );
  OAI22_X1 U15659 ( .A1(n18410), .A2(n19467), .B1(n19278), .B2(n13754), .ZN(
        n13755) );
  AOI21_X1 U15660 ( .B1(n14176), .B2(n13756), .A(n13755), .ZN(n13757) );
  OAI21_X1 U15661 ( .B1(n19468), .B2(n13758), .A(n13757), .ZN(P2_U2919) );
  INV_X1 U15662 ( .A(n13092), .ZN(n13760) );
  XNOR2_X1 U15663 ( .A(n13760), .B(n13759), .ZN(n14068) );
  NAND2_X1 U15664 ( .A1(n14068), .A2(n14656), .ZN(n13763) );
  INV_X1 U15665 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13786) );
  OAI22_X1 U15666 ( .A1(n15087), .A2(n19784), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13786), .ZN(n13761) );
  AOI21_X1 U15667 ( .B1(n14132), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13761), .ZN(n13762) );
  NAND2_X1 U15668 ( .A1(n21898), .A2(n21881), .ZN(n14136) );
  OR2_X1 U15669 ( .A1(n13764), .A2(n14136), .ZN(n13765) );
  NAND2_X1 U15670 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  OAI21_X1 U15671 ( .B1(n13768), .B2(n13767), .A(n13920), .ZN(n15414) );
  INV_X1 U15672 ( .A(n13769), .ZN(n15410) );
  NAND2_X1 U15673 ( .A1(n15410), .A2(n13770), .ZN(n13772) );
  AND2_X1 U15674 ( .A1(n13772), .A2(n13771), .ZN(n21400) );
  OAI22_X1 U15675 ( .A1(n15497), .A2(n21400), .B1(n13773), .B2(n19892), .ZN(
        n13774) );
  INV_X1 U15676 ( .A(n13774), .ZN(n13775) );
  OAI21_X1 U15677 ( .B1(n15414), .B2(n15509), .A(n13775), .ZN(P1_U2871) );
  NOR2_X1 U15678 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16765), .ZN(n21627) );
  NAND2_X1 U15679 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21627), .ZN(n21619) );
  INV_X1 U15680 ( .A(n21619), .ZN(n13776) );
  INV_X1 U15681 ( .A(n19952), .ZN(n15679) );
  OR2_X1 U15682 ( .A1(n13777), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21394) );
  NAND2_X1 U15683 ( .A1(n21623), .A2(n13779), .ZN(n16749) );
  NAND3_X1 U15684 ( .A1(n21394), .A2(n13778), .A3(n19961), .ZN(n13788) );
  INV_X1 U15685 ( .A(n21872), .ZN(n21900) );
  NAND2_X1 U15686 ( .A1(n21900), .A2(n13780), .ZN(n21198) );
  NAND2_X1 U15687 ( .A1(n21198), .A2(n21614), .ZN(n13781) );
  NAND2_X1 U15688 ( .A1(n21614), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16756) );
  NAND2_X1 U15689 ( .A1(n21881), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13782) );
  AND2_X1 U15690 ( .A1(n16756), .A2(n13782), .ZN(n13789) );
  INV_X1 U15691 ( .A(n13789), .ZN(n13783) );
  INV_X1 U15692 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13784) );
  OAI22_X1 U15693 ( .A1(n19923), .A2(n13786), .B1(n21373), .B2(n13784), .ZN(
        n13785) );
  AOI21_X1 U15694 ( .B1(n19946), .B2(n13786), .A(n13785), .ZN(n13787) );
  OAI211_X1 U15695 ( .C1(n15414), .C2(n15679), .A(n13788), .B(n13787), .ZN(
        P1_U2998) );
  NAND2_X1 U15696 ( .A1(n13789), .A2(n19923), .ZN(n13794) );
  AND2_X1 U15697 ( .A1(n13790), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13803) );
  OAI21_X1 U15698 ( .B1(n13791), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13792), .ZN(n13806) );
  NOR2_X1 U15699 ( .A1(n13806), .A2(n21610), .ZN(n13793) );
  AOI211_X1 U15700 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13794), .A(
        n13803), .B(n13793), .ZN(n13795) );
  OAI21_X1 U15701 ( .B1(n15679), .B2(n15415), .A(n13795), .ZN(P1_U2999) );
  INV_X1 U15702 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13796) );
  OR2_X1 U15703 ( .A1(n16187), .A2(n13796), .ZN(n13798) );
  NAND2_X1 U15704 ( .A1(n16187), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13797) );
  AND2_X1 U15705 ( .A1(n13798), .A2(n13797), .ZN(n19230) );
  XNOR2_X1 U15706 ( .A(n13800), .B(n13799), .ZN(n18093) );
  OAI222_X1 U15707 ( .A1(n19279), .A2(n19230), .B1(n18093), .B2(n19287), .C1(
        n17088), .C2(n19278), .ZN(P2_U2913) );
  INV_X1 U15708 ( .A(n21300), .ZN(n21312) );
  AOI21_X1 U15709 ( .B1(n21314), .B2(n21228), .A(n21312), .ZN(n21390) );
  NOR3_X1 U15710 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21314), .A3(
        n21206), .ZN(n13801) );
  AOI21_X1 U15711 ( .B1(n21390), .B2(n21367), .A(n13801), .ZN(n13802) );
  INV_X1 U15712 ( .A(n13802), .ZN(n13805) );
  AOI21_X1 U15713 ( .B1(n21382), .B2(n15418), .A(n13803), .ZN(n13804) );
  OAI211_X1 U15714 ( .C1(n21353), .C2(n13806), .A(n13805), .B(n13804), .ZN(
        P1_U3031) );
  NOR2_X1 U15715 ( .A1(n19034), .A2(n18410), .ZN(n13811) );
  OAI21_X1 U15716 ( .B1(n13809), .B2(n13808), .A(n13807), .ZN(n18046) );
  XNOR2_X1 U15717 ( .A(n19035), .B(n18046), .ZN(n13810) );
  NOR2_X1 U15718 ( .A1(n13810), .A2(n13811), .ZN(n14080) );
  AOI21_X1 U15719 ( .B1(n13811), .B2(n13810), .A(n14080), .ZN(n13817) );
  INV_X1 U15720 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13812) );
  OR2_X1 U15721 ( .A1(n16187), .A2(n13812), .ZN(n13814) );
  NAND2_X1 U15722 ( .A1(n16187), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13813) );
  AND2_X1 U15723 ( .A1(n13814), .A2(n13813), .ZN(n19532) );
  INV_X1 U15724 ( .A(n19532), .ZN(n16210) );
  INV_X1 U15725 ( .A(n18046), .ZN(n18425) );
  INV_X1 U15726 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17079) );
  OAI22_X1 U15727 ( .A1(n18425), .A2(n19467), .B1(n19278), .B2(n17079), .ZN(
        n13815) );
  AOI21_X1 U15728 ( .B1(n14176), .B2(n16210), .A(n13815), .ZN(n13816) );
  OAI21_X1 U15729 ( .B1(n13817), .B2(n19468), .A(n13816), .ZN(P2_U2918) );
  INV_X1 U15730 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13818) );
  OR2_X1 U15731 ( .A1(n16187), .A2(n13818), .ZN(n13820) );
  NAND2_X1 U15732 ( .A1(n16187), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13819) );
  AND2_X1 U15733 ( .A1(n13820), .A2(n13819), .ZN(n19029) );
  XOR2_X1 U15734 ( .A(n13822), .B(n13821), .Z(n18101) );
  INV_X1 U15735 ( .A(n18101), .ZN(n13823) );
  INV_X1 U15736 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17090) );
  OAI222_X1 U15737 ( .A1(n19279), .A2(n19029), .B1(n13823), .B2(n19287), .C1(
        n17090), .C2(n19278), .ZN(P2_U2912) );
  NOR2_X1 U15738 ( .A1(n13824), .A2(n15291), .ZN(n13825) );
  NAND2_X1 U15739 ( .A1(n12969), .A2(n15511), .ZN(n13828) );
  NAND2_X2 U15740 ( .A1(n15553), .A2(n13828), .ZN(n15587) );
  INV_X2 U15741 ( .A(n15239), .ZN(n15553) );
  INV_X1 U15742 ( .A(n21711), .ZN(n15577) );
  OAI222_X1 U15743 ( .A1(n15587), .A2(n15415), .B1(n15553), .B2(n19782), .C1(
        n15585), .C2(n15577), .ZN(P1_U2904) );
  INV_X1 U15744 ( .A(n21912), .ZN(n15572) );
  OAI222_X1 U15745 ( .A1(n15587), .A2(n15414), .B1(n15553), .B2(n19784), .C1(
        n15585), .C2(n15572), .ZN(P1_U2903) );
  OR2_X1 U15746 ( .A1(n14180), .A2(n19983), .ZN(n13830) );
  NAND2_X1 U15747 ( .A1(n14180), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13829) );
  AND2_X1 U15748 ( .A1(n13830), .A2(n13829), .ZN(n19020) );
  AOI21_X1 U15749 ( .B1(n13833), .B2(n13832), .A(n13831), .ZN(n18113) );
  INV_X1 U15750 ( .A(n18113), .ZN(n18476) );
  INV_X1 U15751 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17092) );
  OAI222_X1 U15752 ( .A1(n19279), .A2(n19020), .B1(n18476), .B2(n19287), .C1(
        n17092), .C2(n19278), .ZN(P2_U2911) );
  OR2_X1 U15753 ( .A1(n14180), .A2(n19985), .ZN(n13835) );
  NAND2_X1 U15754 ( .A1(n14180), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13834) );
  AND2_X1 U15755 ( .A1(n13835), .A2(n13834), .ZN(n19017) );
  OAI21_X1 U15756 ( .B1(n13836), .B2(n13831), .A(n13883), .ZN(n18123) );
  INV_X1 U15757 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17094) );
  OAI222_X1 U15758 ( .A1(n19279), .A2(n19017), .B1(n18123), .B2(n19287), .C1(
        n17094), .C2(n19278), .ZN(P2_U2910) );
  AND2_X1 U15759 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19163) );
  NAND2_X1 U15760 ( .A1(n19163), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13856) );
  INV_X1 U15761 ( .A(n19163), .ZN(n13839) );
  NAND2_X1 U15762 ( .A1(n13839), .A2(n19160), .ZN(n13840) );
  NAND2_X1 U15763 ( .A1(n13856), .A2(n13840), .ZN(n14333) );
  NOR2_X1 U15764 ( .A1(n14333), .A2(n13500), .ZN(n13841) );
  AOI21_X1 U15765 ( .B1(n13859), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13841), .ZN(n13842) );
  NAND2_X1 U15766 ( .A1(n15990), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13865) );
  INV_X1 U15767 ( .A(n13844), .ZN(n13845) );
  OR2_X1 U15768 ( .A1(n13846), .A2(n13845), .ZN(n13847) );
  MUX2_X1 U15769 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n18499), .S(n16112), .Z(
        n13852) );
  AOI21_X1 U15770 ( .B1(n19085), .B2(n16082), .A(n13852), .ZN(n13853) );
  INV_X1 U15771 ( .A(n13853), .ZN(P2_U2885) );
  INV_X1 U15772 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U15773 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17107), .B1(n17108), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13854) );
  OAI21_X1 U15774 ( .B1(n13855), .B2(n13905), .A(n13854), .ZN(P2_U2935) );
  AOI21_X1 U15775 ( .B1(n19159), .B2(n13856), .A(n13500), .ZN(n13858) );
  INV_X1 U15776 ( .A(n13856), .ZN(n13857) );
  NAND2_X1 U15777 ( .A1(n13857), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19218) );
  AND2_X1 U15778 ( .A1(n13858), .A2(n19218), .ZN(n14343) );
  AOI21_X1 U15779 ( .B1(n13859), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14343), .ZN(n13860) );
  NOR2_X1 U15780 ( .A1(n15931), .A2(n13861), .ZN(n13862) );
  INV_X1 U15781 ( .A(n13865), .ZN(n13866) );
  NAND2_X1 U15782 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  NAND2_X1 U15783 ( .A1(n13942), .A2(n13943), .ZN(n13873) );
  NAND2_X1 U15784 ( .A1(n11873), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13870) );
  INV_X1 U15785 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13874) );
  NOR2_X1 U15786 ( .A1(n15931), .A2(n13874), .ZN(n13935) );
  XOR2_X1 U15787 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13934), .Z(n13879)
         );
  NAND2_X1 U15788 ( .A1(n13875), .A2(n13876), .ZN(n13877) );
  AND2_X1 U15789 ( .A1(n13928), .A2(n13877), .ZN(n16971) );
  INV_X1 U15790 ( .A(n16971), .ZN(n18076) );
  MUX2_X1 U15791 ( .A(n18076), .B(n18081), .S(n16046), .Z(n13878) );
  OAI21_X1 U15792 ( .B1(n13879), .B2(n16115), .A(n13878), .ZN(P2_U2882) );
  OR2_X1 U15793 ( .A1(n16187), .A2(n19987), .ZN(n13881) );
  NAND2_X1 U15794 ( .A1(n14180), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13880) );
  AND2_X1 U15795 ( .A1(n13881), .A2(n13880), .ZN(n19014) );
  AOI21_X1 U15796 ( .B1(n13884), .B2(n13883), .A(n13882), .ZN(n18136) );
  INV_X1 U15797 ( .A(n18136), .ZN(n18438) );
  INV_X1 U15798 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17098) );
  OAI222_X1 U15799 ( .A1(n19279), .A2(n19014), .B1(n18438), .B2(n19287), .C1(
        n17098), .C2(n19278), .ZN(P2_U2909) );
  INV_X1 U15800 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U15801 ( .A1(n17108), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U15802 ( .B1(n13886), .B2(n13905), .A(n13885), .ZN(P2_U2923) );
  INV_X1 U15803 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U15804 ( .A1(n17108), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13887) );
  OAI21_X1 U15805 ( .B1(n13888), .B2(n13905), .A(n13887), .ZN(P2_U2929) );
  INV_X1 U15806 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U15807 ( .A1(n17108), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13889) );
  OAI21_X1 U15808 ( .B1(n16127), .B2(n13905), .A(n13889), .ZN(P2_U2922) );
  AOI22_X1 U15809 ( .A1(n17108), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13890) );
  OAI21_X1 U15810 ( .B1(n13891), .B2(n13905), .A(n13890), .ZN(P2_U2930) );
  INV_X1 U15811 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U15812 ( .A1(n17108), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13892) );
  OAI21_X1 U15813 ( .B1(n13893), .B2(n13905), .A(n13892), .ZN(P2_U2931) );
  INV_X1 U15814 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16141) );
  AOI22_X1 U15815 ( .A1(n17108), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13894) );
  OAI21_X1 U15816 ( .B1(n16141), .B2(n13905), .A(n13894), .ZN(P2_U2924) );
  INV_X1 U15817 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U15818 ( .A1(n17108), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13895) );
  OAI21_X1 U15819 ( .B1(n16158), .B2(n13905), .A(n13895), .ZN(P2_U2926) );
  INV_X1 U15820 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U15821 ( .A1(n17108), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13896) );
  OAI21_X1 U15822 ( .B1(n13897), .B2(n13905), .A(n13896), .ZN(P2_U2927) );
  INV_X1 U15823 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U15824 ( .A1(n17108), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13898) );
  OAI21_X1 U15825 ( .B1(n13899), .B2(n13905), .A(n13898), .ZN(P2_U2928) );
  INV_X1 U15826 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15827 ( .A1(n17108), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13900) );
  OAI21_X1 U15828 ( .B1(n13901), .B2(n13905), .A(n13900), .ZN(P2_U2925) );
  INV_X1 U15829 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U15830 ( .A1(n17096), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13902) );
  OAI21_X1 U15831 ( .B1(n13903), .B2(n13905), .A(n13902), .ZN(P2_U2932) );
  INV_X1 U15832 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U15833 ( .A1(n17096), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U15834 ( .B1(n13906), .B2(n13905), .A(n13904), .ZN(P2_U2921) );
  XNOR2_X1 U15835 ( .A(n14108), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13911) );
  OR2_X1 U15836 ( .A1(n13929), .A2(n13907), .ZN(n13908) );
  NAND2_X1 U15837 ( .A1(n14105), .A2(n13908), .ZN(n18105) );
  INV_X1 U15838 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13909) );
  MUX2_X1 U15839 ( .A(n18105), .B(n13909), .S(n16046), .Z(n13910) );
  OAI21_X1 U15840 ( .B1(n13911), .B2(n16115), .A(n13910), .ZN(P2_U2880) );
  NAND2_X1 U15841 ( .A1(n10979), .A2(n14656), .ZN(n13915) );
  XNOR2_X1 U15842 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16957) );
  AOI21_X1 U15843 ( .B1(n15161), .B2(n16957), .A(n15164), .ZN(n13912) );
  OAI21_X1 U15844 ( .B1(n15087), .B2(n19786), .A(n13912), .ZN(n13913) );
  AOI21_X1 U15845 ( .B1(n14132), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13913), .ZN(n13914) );
  NAND2_X1 U15846 ( .A1(n13915), .A2(n13914), .ZN(n13916) );
  NAND2_X1 U15847 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14086) );
  NAND2_X1 U15848 ( .A1(n13916), .A2(n14086), .ZN(n13921) );
  INV_X1 U15849 ( .A(n14087), .ZN(n13919) );
  AOI21_X1 U15850 ( .B1(n13921), .B2(n13920), .A(n13919), .ZN(n16959) );
  INV_X1 U15851 ( .A(n16959), .ZN(n13933) );
  AND2_X1 U15852 ( .A1(n14097), .A2(n13923), .ZN(n21233) );
  INV_X1 U15853 ( .A(n19892), .ZN(n15507) );
  AOI22_X1 U15854 ( .A1(n19888), .A2(n21233), .B1(n15507), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U15855 ( .B1(n13933), .B2(n15509), .A(n13924), .ZN(P1_U2870) );
  NOR2_X1 U15856 ( .A1(n13934), .A2(n12103), .ZN(n13926) );
  INV_X1 U15857 ( .A(n14108), .ZN(n13925) );
  OAI211_X1 U15858 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13926), .A(
        n13925), .B(n16082), .ZN(n13932) );
  AND2_X1 U15859 ( .A1(n13928), .A2(n13927), .ZN(n13930) );
  OR2_X1 U15860 ( .A1(n13930), .A2(n13929), .ZN(n14625) );
  INV_X1 U15861 ( .A(n14625), .ZN(n18089) );
  NAND2_X1 U15862 ( .A1(n18089), .A2(n16112), .ZN(n13931) );
  OAI211_X1 U15863 ( .C1(n16112), .C2(n12217), .A(n13932), .B(n13931), .ZN(
        P2_U2881) );
  INV_X1 U15864 ( .A(n21959), .ZN(n15567) );
  OAI222_X1 U15865 ( .A1(n15587), .A2(n13933), .B1(n15553), .B2(n19786), .C1(
        n15585), .C2(n15567), .ZN(P1_U2902) );
  OAI21_X1 U15866 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n19281) );
  NAND2_X1 U15867 ( .A1(n13938), .A2(n13937), .ZN(n13939) );
  NAND2_X1 U15868 ( .A1(n13875), .A2(n13939), .ZN(n18068) );
  NOR2_X1 U15869 ( .A1(n18068), .A2(n16046), .ZN(n13940) );
  AOI21_X1 U15870 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16046), .A(n13940), .ZN(
        n13941) );
  OAI21_X1 U15871 ( .B1(n19281), .B2(n16115), .A(n13941), .ZN(P2_U2883) );
  CLKBUF_X1 U15872 ( .A(n13944), .Z(n15814) );
  MUX2_X1 U15873 ( .A(n12148), .B(n15814), .S(n16112), .Z(n13945) );
  OAI21_X1 U15874 ( .B1(n19198), .B2(n16115), .A(n13945), .ZN(P2_U2884) );
  OR2_X1 U15875 ( .A1(n14180), .A2(n19989), .ZN(n13947) );
  NAND2_X1 U15876 ( .A1(n14180), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13946) );
  AND2_X1 U15877 ( .A1(n13947), .A2(n13946), .ZN(n19011) );
  OAI21_X1 U15878 ( .B1(n13948), .B2(n13882), .A(n14127), .ZN(n16654) );
  INV_X1 U15879 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17100) );
  OAI222_X1 U15880 ( .A1(n19279), .A2(n19011), .B1(n16654), .B2(n19287), .C1(
        n17100), .C2(n19278), .ZN(P2_U2908) );
  OR2_X1 U15881 ( .A1(n15814), .A2(n13949), .ZN(n13964) );
  AND2_X1 U15882 ( .A1(n13951), .A2(n13950), .ZN(n13979) );
  INV_X1 U15883 ( .A(n12367), .ZN(n13976) );
  NAND2_X1 U15884 ( .A1(n13987), .A2(n13976), .ZN(n13954) );
  NAND2_X1 U15885 ( .A1(n13953), .A2(n13952), .ZN(n13974) );
  OAI211_X1 U15886 ( .C1(n11986), .C2(n13979), .A(n13954), .B(n13974), .ZN(
        n13955) );
  INV_X1 U15887 ( .A(n13955), .ZN(n13960) );
  NAND2_X1 U15888 ( .A1(n13957), .A2(n13956), .ZN(n13982) );
  AOI22_X1 U15889 ( .A1(n13982), .A2(n13974), .B1(n12367), .B2(n13987), .ZN(
        n13959) );
  MUX2_X1 U15890 ( .A(n13960), .B(n13959), .S(n13958), .Z(n13962) );
  INV_X1 U15891 ( .A(n15882), .ZN(n13961) );
  AND2_X1 U15892 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  NAND2_X1 U15893 ( .A1(n13964), .A2(n13963), .ZN(n16692) );
  INV_X1 U15894 ( .A(n14021), .ZN(n13965) );
  MUX2_X1 U15895 ( .A(n16692), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13965), .Z(n14024) );
  INV_X1 U15896 ( .A(n14024), .ZN(n13966) );
  OR2_X1 U15897 ( .A1(n13966), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13996) );
  NAND2_X1 U15898 ( .A1(n18427), .A2(n13989), .ZN(n13973) );
  INV_X1 U15899 ( .A(n13967), .ZN(n13968) );
  NAND2_X1 U15900 ( .A1(n13969), .A2(n13968), .ZN(n13986) );
  AOI22_X1 U15901 ( .A1(n11352), .A2(n13987), .B1(n13986), .B2(n13971), .ZN(
        n13972) );
  NAND2_X1 U15902 ( .A1(n13973), .A2(n13972), .ZN(n16681) );
  INV_X1 U15903 ( .A(n16681), .ZN(n13993) );
  NAND2_X1 U15904 ( .A1(n18499), .A2(n13989), .ZN(n13984) );
  NAND2_X1 U15905 ( .A1(n11758), .A2(n13974), .ZN(n13981) );
  INV_X1 U15906 ( .A(n13975), .ZN(n13977) );
  NAND3_X1 U15907 ( .A1(n13987), .A2(n13977), .A3(n13976), .ZN(n13978) );
  OAI21_X1 U15908 ( .B1(n13979), .B2(n13981), .A(n13978), .ZN(n13980) );
  AOI21_X1 U15909 ( .B1(n13982), .B2(n13981), .A(n13980), .ZN(n13983) );
  NAND2_X1 U15910 ( .A1(n13984), .A2(n13983), .ZN(n16688) );
  NOR2_X1 U15911 ( .A1(n19160), .A2(n16688), .ZN(n13992) );
  INV_X1 U15912 ( .A(n18036), .ZN(n18415) );
  MUX2_X1 U15913 ( .A(n13987), .B(n13986), .S(n13985), .Z(n13988) );
  AOI21_X1 U15914 ( .B1(n18415), .B2(n13989), .A(n13988), .ZN(n13990) );
  INV_X1 U15915 ( .A(n13990), .ZN(n16675) );
  AOI211_X1 U15916 ( .C1(n16681), .C2(n19179), .A(n19146), .B(n16675), .ZN(
        n13991) );
  AOI211_X1 U15917 ( .C1(n13993), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13992), .B(n13991), .ZN(n13994) );
  MUX2_X1 U15918 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16688), .S(
        n14021), .Z(n14023) );
  AOI22_X1 U15919 ( .A1(n13994), .A2(n14021), .B1(n19160), .B2(n14023), .ZN(
        n13995) );
  NAND2_X1 U15920 ( .A1(n13996), .A2(n13995), .ZN(n13997) );
  OAI211_X1 U15921 ( .C1(n14024), .C2(n19159), .A(n16717), .B(n13997), .ZN(
        n14026) );
  NAND2_X1 U15922 ( .A1(n18520), .A2(n13998), .ZN(n14002) );
  AOI22_X1 U15923 ( .A1(n14000), .A2(n13999), .B1(n14014), .B2(n14012), .ZN(
        n14001) );
  NAND2_X1 U15924 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  AOI21_X1 U15925 ( .B1(n14004), .B2(n14335), .A(n14003), .ZN(n14008) );
  NAND2_X1 U15926 ( .A1(n14006), .A2(n14005), .ZN(n14007) );
  AND2_X1 U15927 ( .A1(n14008), .A2(n14007), .ZN(n18537) );
  NOR2_X1 U15928 ( .A1(n14010), .A2(n14009), .ZN(n14011) );
  NAND2_X1 U15929 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  OR2_X1 U15930 ( .A1(n14014), .A2(n14013), .ZN(n18534) );
  NOR2_X1 U15931 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14016) );
  OAI21_X1 U15932 ( .B1(n18534), .B2(n14016), .A(n14015), .ZN(n14017) );
  NOR2_X1 U15933 ( .A1(n14018), .A2(n14017), .ZN(n14019) );
  OAI211_X1 U15934 ( .C1(n14021), .C2(n14020), .A(n18537), .B(n14019), .ZN(
        n14022) );
  AOI21_X1 U15935 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14025) );
  AND2_X1 U15936 ( .A1(n14026), .A2(n14025), .ZN(n18533) );
  AND2_X1 U15937 ( .A1(n16714), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14027) );
  NAND2_X1 U15938 ( .A1(n18533), .A2(n14027), .ZN(n14033) );
  NOR2_X1 U15939 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14028), .ZN(n15820) );
  AND2_X1 U15940 ( .A1(n14029), .A2(n15820), .ZN(n15815) );
  AND2_X1 U15941 ( .A1(n14030), .A2(n15815), .ZN(n14031) );
  AOI21_X1 U15942 ( .B1(n14033), .B2(n14032), .A(n14031), .ZN(n18524) );
  OAI21_X1 U15943 ( .B1(n18524), .B2(n18022), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14034) );
  INV_X1 U15944 ( .A(n16716), .ZN(n18519) );
  NAND2_X1 U15945 ( .A1(n14034), .A2(n18519), .ZN(P2_U3593) );
  AND2_X1 U15946 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14035) );
  NOR2_X1 U15947 ( .A1(n14039), .A2(n14035), .ZN(n14041) );
  INV_X1 U15948 ( .A(n14035), .ZN(n14038) );
  NOR2_X1 U15949 ( .A1(n13698), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14037) );
  OAI22_X1 U15950 ( .A1(n14039), .A2(n14038), .B1(n14037), .B2(n14036), .ZN(
        n14040) );
  MUX2_X1 U15951 ( .A(n14041), .B(n14040), .S(n12820), .Z(n14049) );
  INV_X1 U15952 ( .A(n14042), .ZN(n14043) );
  OAI21_X1 U15953 ( .B1(n13698), .B2(n12820), .A(n14043), .ZN(n14044) );
  NOR2_X1 U15954 ( .A1(n14044), .A2(n12999), .ZN(n15806) );
  INV_X1 U15955 ( .A(n13698), .ZN(n14045) );
  NAND2_X1 U15956 ( .A1(n14045), .A2(n14042), .ZN(n14046) );
  OAI21_X1 U15957 ( .B1(n14047), .B2(n15806), .A(n14046), .ZN(n14048) );
  AOI211_X1 U15958 ( .C1(n21804), .C2(n14050), .A(n14049), .B(n14048), .ZN(
        n15808) );
  MUX2_X1 U15959 ( .A(n15808), .B(n12820), .S(n16736), .Z(n16747) );
  MUX2_X1 U15960 ( .A(n14051), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16736), .Z(n16745) );
  NAND2_X1 U15961 ( .A1(n16745), .A2(n16765), .ZN(n14062) );
  AOI21_X1 U15962 ( .B1(n21412), .B2(n14052), .A(n16736), .ZN(n14053) );
  AOI211_X1 U15963 ( .C1(n14054), .C2(n16736), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n14053), .ZN(n14060) );
  NOR2_X1 U15964 ( .A1(n16765), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14056) );
  INV_X1 U15965 ( .A(n14056), .ZN(n14058) );
  INV_X1 U15966 ( .A(n14055), .ZN(n14057) );
  NAND2_X1 U15967 ( .A1(n14056), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14064) );
  OAI21_X1 U15968 ( .B1(n14058), .B2(n14057), .A(n14064), .ZN(n14059) );
  NOR2_X1 U15969 ( .A1(n14060), .A2(n14059), .ZN(n14061) );
  OAI21_X1 U15970 ( .B1(n16747), .B2(n14062), .A(n14061), .ZN(n16753) );
  NAND2_X1 U15971 ( .A1(n14064), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U15972 ( .A1(n16753), .A2(n14065), .ZN(n14101) );
  INV_X1 U15973 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21611) );
  AOI21_X1 U15974 ( .B1(n14101), .B2(n21611), .A(n21620), .ZN(n14066) );
  NAND2_X1 U15975 ( .A1(n16765), .A2(n21898), .ZN(n21196) );
  INV_X1 U15976 ( .A(n14100), .ZN(n21615) );
  OR2_X1 U15977 ( .A1(n14066), .A2(n22199), .ZN(n16768) );
  AND2_X1 U15978 ( .A1(n10980), .A2(n14070), .ZN(n21877) );
  NAND2_X1 U15979 ( .A1(n14068), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21838) );
  INV_X1 U15980 ( .A(n21838), .ZN(n14069) );
  AOI21_X1 U15981 ( .B1(n21877), .B2(n14069), .A(n21900), .ZN(n21905) );
  INV_X1 U15982 ( .A(n21905), .ZN(n14075) );
  INV_X1 U15983 ( .A(n21802), .ZN(n14074) );
  INV_X1 U15984 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21859) );
  NAND2_X1 U15985 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21859), .ZN(n14112) );
  INV_X1 U15986 ( .A(n14070), .ZN(n14071) );
  NOR2_X1 U15987 ( .A1(n21838), .A2(n21900), .ZN(n14072) );
  AND2_X1 U15988 ( .A1(n21792), .A2(n14072), .ZN(n21797) );
  AOI21_X1 U15989 ( .B1(n14112), .B2(n21804), .A(n21797), .ZN(n14073) );
  OAI21_X1 U15990 ( .B1(n14075), .B2(n14074), .A(n14073), .ZN(n14076) );
  NAND2_X1 U15991 ( .A1(n16768), .A2(n14076), .ZN(n14077) );
  OAI21_X1 U15992 ( .B1(n16768), .B2(n21897), .A(n14077), .ZN(P1_U3475) );
  OR2_X1 U15993 ( .A1(n16187), .A2(n19976), .ZN(n14079) );
  NAND2_X1 U15994 ( .A1(n16187), .A2(BUF2_REG_2__SCAN_IN), .ZN(n14078) );
  AND2_X1 U15995 ( .A1(n14079), .A2(n14078), .ZN(n19477) );
  AOI21_X1 U15996 ( .B1(n18425), .B2(n19049), .A(n14080), .ZN(n14168) );
  XNOR2_X1 U15997 ( .A(n14082), .B(n12461), .ZN(n18491) );
  INV_X1 U15998 ( .A(n18491), .ZN(n14167) );
  XNOR2_X1 U15999 ( .A(n14168), .B(n14167), .ZN(n14170) );
  XNOR2_X1 U16000 ( .A(n14170), .B(n19085), .ZN(n14083) );
  INV_X1 U16001 ( .A(n19468), .ZN(n19346) );
  NAND2_X1 U16002 ( .A1(n14083), .A2(n19346), .ZN(n14085) );
  INV_X1 U16003 ( .A(n19467), .ZN(n19345) );
  AOI22_X1 U16004 ( .A1(n19345), .A2(n14167), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19465), .ZN(n14084) );
  OAI211_X1 U16005 ( .C1(n19477), .C2(n19279), .A(n14085), .B(n14084), .ZN(
        P2_U2917) );
  INV_X1 U16006 ( .A(n14089), .ZN(n14091) );
  INV_X1 U16007 ( .A(n14135), .ZN(n14090) );
  OAI21_X1 U16008 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14091), .A(
        n14090), .ZN(n14271) );
  AOI22_X1 U16009 ( .A1(n15161), .A2(n14271), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14092) );
  OAI21_X1 U16010 ( .B1(n15087), .B2(n19788), .A(n14092), .ZN(n14093) );
  AOI21_X1 U16011 ( .B1(n14132), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14093), .ZN(n14094) );
  NAND2_X1 U16012 ( .A1(n14095), .A2(n14094), .ZN(n14130) );
  XOR2_X1 U16013 ( .A(n14131), .B(n14130), .Z(n14233) );
  INV_X1 U16014 ( .A(n14233), .ZN(n14293) );
  INV_X1 U16015 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14099) );
  AND2_X1 U16016 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  NOR2_X1 U16017 ( .A1(n14147), .A2(n14098), .ZN(n21250) );
  INV_X1 U16018 ( .A(n21250), .ZN(n14284) );
  OAI222_X1 U16019 ( .A1(n14293), .A2(n15509), .B1(n19892), .B2(n14099), .C1(
        n14284), .C2(n15497), .ZN(P1_U2869) );
  NAND2_X1 U16020 ( .A1(n14101), .A2(n14100), .ZN(n21624) );
  INV_X1 U16021 ( .A(n21624), .ZN(n14103) );
  INV_X1 U16022 ( .A(n14112), .ZN(n15791) );
  OAI22_X1 U16023 ( .A1(n13672), .A2(n21900), .B1(n13673), .B2(n15791), .ZN(
        n14102) );
  OAI21_X1 U16024 ( .B1(n14103), .B2(n14102), .A(n16768), .ZN(n14104) );
  OAI21_X1 U16025 ( .B1(n16768), .B2(n21864), .A(n14104), .ZN(P1_U3478) );
  OAI21_X1 U16026 ( .B1(n12691), .B2(n12690), .A(n14107), .ZN(n18117) );
  NAND2_X1 U16027 ( .A1(n11049), .A2(n14109), .ZN(n14155) );
  OAI211_X1 U16028 ( .C1(n11049), .C2(n14109), .A(n16082), .B(n14155), .ZN(
        n14111) );
  NAND2_X1 U16029 ( .A1(n16046), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14110) );
  OAI211_X1 U16030 ( .C1(n18117), .C2(n16046), .A(n14111), .B(n14110), .ZN(
        P2_U2879) );
  INV_X1 U16031 ( .A(n22007), .ZN(n15562) );
  OAI222_X1 U16032 ( .A1(n15587), .A2(n14293), .B1(n15553), .B2(n19788), .C1(
        n15585), .C2(n15562), .ZN(P1_U2901) );
  INV_X1 U16033 ( .A(n16768), .ZN(n14116) );
  XNOR2_X1 U16034 ( .A(n10980), .B(n21838), .ZN(n14113) );
  INV_X1 U16035 ( .A(n21850), .ZN(n21710) );
  AOI22_X1 U16036 ( .A1(n14113), .A2(n21908), .B1(n21710), .B2(n14112), .ZN(
        n14115) );
  NAND2_X1 U16037 ( .A1(n14116), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14114) );
  OAI21_X1 U16038 ( .B1(n14116), .B2(n14115), .A(n14114), .ZN(P1_U3476) );
  NAND2_X1 U16039 ( .A1(n13603), .A2(n14117), .ZN(n14118) );
  NAND2_X1 U16040 ( .A1(n19780), .A2(n14272), .ZN(n14326) );
  NOR2_X1 U16041 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21615), .ZN(n19797) );
  AOI22_X1 U16042 ( .A1(n19797), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14119) );
  OAI21_X1 U16043 ( .B1(n14120), .B2(n14326), .A(n14119), .ZN(P1_U2919) );
  AOI22_X1 U16044 ( .A1(n21200), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14121) );
  OAI21_X1 U16045 ( .B1(n14122), .B2(n14326), .A(n14121), .ZN(P1_U2918) );
  OR2_X1 U16046 ( .A1(n14180), .A2(n14123), .ZN(n14125) );
  NAND2_X1 U16047 ( .A1(n14180), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14124) );
  AND2_X1 U16048 ( .A1(n14125), .A2(n14124), .ZN(n19008) );
  AOI21_X1 U16049 ( .B1(n14128), .B2(n14127), .A(n14126), .ZN(n18465) );
  INV_X1 U16050 ( .A(n18465), .ZN(n14129) );
  INV_X1 U16051 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17102) );
  OAI222_X1 U16052 ( .A1(n19279), .A2(n19008), .B1(n14129), .B2(n19287), .C1(
        n17102), .C2(n19278), .ZN(P2_U2907) );
  NAND2_X1 U16053 ( .A1(n14131), .A2(n14130), .ZN(n14144) );
  NAND2_X1 U16054 ( .A1(n14132), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14139) );
  INV_X1 U16055 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14133) );
  AOI21_X1 U16056 ( .B1(n14133), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14134) );
  AOI21_X1 U16057 ( .B1(n15165), .B2(P1_EAX_REG_4__SCAN_IN), .A(n14134), .ZN(
        n14138) );
  OAI21_X1 U16058 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14135), .A(
        n14187), .ZN(n21418) );
  NOR2_X1 U16059 ( .A1(n21418), .A2(n14136), .ZN(n14137) );
  AOI21_X1 U16060 ( .B1(n14139), .B2(n14138), .A(n14137), .ZN(n14140) );
  INV_X1 U16061 ( .A(n14143), .ZN(n14142) );
  NAND2_X1 U16062 ( .A1(n14144), .A2(n14143), .ZN(n14145) );
  AND2_X1 U16063 ( .A1(n14192), .A2(n14145), .ZN(n21404) );
  INV_X1 U16064 ( .A(n21404), .ZN(n14149) );
  INV_X1 U16065 ( .A(n22054), .ZN(n15558) );
  OAI222_X1 U16066 ( .A1(n15587), .A2(n14149), .B1(n15553), .B2(n19790), .C1(
        n15585), .C2(n15558), .ZN(P1_U2900) );
  OR2_X1 U16067 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  NAND2_X1 U16068 ( .A1(n19887), .A2(n14148), .ZN(n21405) );
  INV_X1 U16069 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14150) );
  OAI222_X1 U16070 ( .A1(n21405), .A2(n15497), .B1(n14150), .B2(n19892), .C1(
        n14149), .C2(n15509), .ZN(P1_U2868) );
  OR2_X1 U16071 ( .A1(n16187), .A2(n19992), .ZN(n14152) );
  NAND2_X1 U16072 ( .A1(n14180), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14151) );
  AND2_X1 U16073 ( .A1(n14152), .A2(n14151), .ZN(n19005) );
  INV_X1 U16074 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17104) );
  OAI21_X1 U16075 ( .B1(n14126), .B2(n14153), .A(n14184), .ZN(n18448) );
  OAI222_X1 U16076 ( .A1(n19279), .A2(n19005), .B1(n19278), .B2(n17104), .C1(
        n18448), .C2(n19287), .ZN(P2_U2906) );
  INV_X1 U16077 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14162) );
  INV_X1 U16078 ( .A(n14155), .ZN(n14157) );
  INV_X1 U16079 ( .A(n14156), .ZN(n14154) );
  OAI211_X1 U16080 ( .C1(n14157), .C2(n14156), .A(n16082), .B(n14240), .ZN(
        n14161) );
  AND2_X1 U16081 ( .A1(n14107), .A2(n14158), .ZN(n14159) );
  OR2_X1 U16082 ( .A1(n14159), .A2(n14237), .ZN(n18124) );
  INV_X1 U16083 ( .A(n18124), .ZN(n16671) );
  NAND2_X1 U16084 ( .A1(n16671), .A2(n16112), .ZN(n14160) );
  OAI211_X1 U16085 ( .C1(n16112), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        P2_U2878) );
  OR2_X1 U16086 ( .A1(n14164), .A2(n14163), .ZN(n14166) );
  NAND2_X1 U16087 ( .A1(n14166), .A2(n14165), .ZN(n17056) );
  XNOR2_X1 U16088 ( .A(n19198), .B(n17056), .ZN(n14172) );
  NAND2_X1 U16089 ( .A1(n14168), .A2(n14167), .ZN(n14169) );
  OAI21_X1 U16090 ( .B1(n14170), .B2(n19142), .A(n14169), .ZN(n14171) );
  NOR2_X1 U16091 ( .A1(n14171), .A2(n14172), .ZN(n14211) );
  AOI21_X1 U16092 ( .B1(n14172), .B2(n14171), .A(n14211), .ZN(n14179) );
  INV_X1 U16093 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n14173) );
  OR2_X1 U16094 ( .A1(n16187), .A2(n14173), .ZN(n14175) );
  NAND2_X1 U16095 ( .A1(n14180), .A2(BUF2_REG_3__SCAN_IN), .ZN(n14174) );
  AND2_X1 U16096 ( .A1(n14175), .A2(n14174), .ZN(n19409) );
  INV_X1 U16097 ( .A(n19409), .ZN(n16201) );
  AOI22_X1 U16098 ( .A1(n14176), .A2(n16201), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19465), .ZN(n14178) );
  INV_X1 U16099 ( .A(n17056), .ZN(n14205) );
  NAND2_X1 U16100 ( .A1(n14205), .A2(n19345), .ZN(n14177) );
  OAI211_X1 U16101 ( .C1(n14179), .C2(n19468), .A(n14178), .B(n14177), .ZN(
        P2_U2916) );
  OR2_X1 U16102 ( .A1(n16187), .A2(n19994), .ZN(n14182) );
  NAND2_X1 U16103 ( .A1(n14180), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14181) );
  AND2_X1 U16104 ( .A1(n14182), .A2(n14181), .ZN(n19002) );
  AND2_X1 U16105 ( .A1(n14184), .A2(n14183), .ZN(n14186) );
  OR2_X1 U16106 ( .A1(n14186), .A2(n14185), .ZN(n18184) );
  INV_X1 U16107 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17106) );
  OAI222_X1 U16108 ( .A1(n19279), .A2(n19002), .B1(n18184), .B2(n19287), .C1(
        n17106), .C2(n19278), .ZN(P2_U2905) );
  OAI21_X1 U16109 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14188), .A(
        n14218), .ZN(n21422) );
  AOI22_X1 U16110 ( .A1(n15161), .A2(n21422), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14189) );
  OAI21_X1 U16111 ( .B1(n15087), .B2(n19792), .A(n14189), .ZN(n14190) );
  AOI21_X1 U16112 ( .B1(n14193), .B2(n14192), .A(n14224), .ZN(n21429) );
  INV_X1 U16113 ( .A(n21429), .ZN(n14194) );
  INV_X1 U16114 ( .A(n22101), .ZN(n15554) );
  OAI222_X1 U16115 ( .A1(n15587), .A2(n14194), .B1(n15553), .B2(n19792), .C1(
        n15585), .C2(n15554), .ZN(P1_U2899) );
  INV_X1 U16116 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18141) );
  OAI211_X1 U16117 ( .C1(n14239), .C2(n14195), .A(n14301), .B(n16082), .ZN(
        n14201) );
  NOR2_X1 U16118 ( .A1(n14197), .A2(n14198), .ZN(n14199) );
  NAND2_X1 U16119 ( .A1(n11379), .A2(n16112), .ZN(n14200) );
  OAI211_X1 U16120 ( .C1(n16112), .C2(n18141), .A(n14201), .B(n14200), .ZN(
        P2_U2876) );
  INV_X1 U16121 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n14202) );
  OR2_X1 U16122 ( .A1(n16187), .A2(n14202), .ZN(n14204) );
  NAND2_X1 U16123 ( .A1(n16187), .A2(BUF2_REG_4__SCAN_IN), .ZN(n14203) );
  AND2_X1 U16124 ( .A1(n14204), .A2(n14203), .ZN(n19353) );
  NOR2_X1 U16125 ( .A1(n19170), .A2(n14205), .ZN(n14210) );
  NAND2_X1 U16126 ( .A1(n14206), .A2(n14165), .ZN(n14209) );
  INV_X1 U16127 ( .A(n14207), .ZN(n14208) );
  NAND2_X1 U16128 ( .A1(n14209), .A2(n14208), .ZN(n14391) );
  OAI21_X1 U16129 ( .B1(n14211), .B2(n14210), .A(n14391), .ZN(n19283) );
  XNOR2_X1 U16130 ( .A(n19283), .B(n19281), .ZN(n14212) );
  NAND2_X1 U16131 ( .A1(n14212), .A2(n19346), .ZN(n14214) );
  INV_X1 U16132 ( .A(n14391), .ZN(n18055) );
  AOI22_X1 U16133 ( .A1(n19345), .A2(n18055), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19465), .ZN(n14213) );
  OAI211_X1 U16134 ( .C1(n19353), .C2(n19279), .A(n14214), .B(n14213), .ZN(
        P2_U2915) );
  OAI21_X1 U16135 ( .B1(n14185), .B2(n14215), .A(n10984), .ZN(n18204) );
  OAI222_X1 U16136 ( .A1(n19279), .A2(n14216), .B1(n18204), .B2(n19287), .C1(
        n17111), .C2(n19278), .ZN(P2_U2904) );
  OAI21_X1 U16137 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n14219), .A(
        n14246), .ZN(n21444) );
  AOI22_X1 U16138 ( .A1(n15161), .A2(n21444), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14220) );
  OAI21_X1 U16139 ( .B1(n15087), .B2(n19794), .A(n14220), .ZN(n14221) );
  INV_X1 U16140 ( .A(n14221), .ZN(n14222) );
  OR2_X1 U16141 ( .A1(n14224), .A2(n14225), .ZN(n14226) );
  AND2_X1 U16142 ( .A1(n14252), .A2(n14226), .ZN(n21441) );
  INV_X1 U16143 ( .A(n21441), .ZN(n14227) );
  INV_X1 U16144 ( .A(n22149), .ZN(n15549) );
  OAI222_X1 U16145 ( .A1(n15587), .A2(n14227), .B1(n15553), .B2(n19794), .C1(
        n15585), .C2(n15549), .ZN(P1_U2898) );
  AOI21_X1 U16146 ( .B1(n14228), .B2(n14230), .A(n14229), .ZN(n21249) );
  INV_X1 U16147 ( .A(n21249), .ZN(n14235) );
  AOI22_X1 U16148 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14231) );
  OAI21_X1 U16149 ( .B1(n19964), .B2(n14271), .A(n14231), .ZN(n14232) );
  AOI21_X1 U16150 ( .B1(n14233), .B2(n19952), .A(n14232), .ZN(n14234) );
  OAI21_X1 U16151 ( .B1(n14235), .B2(n21610), .A(n14234), .ZN(P1_U2996) );
  NOR2_X1 U16152 ( .A1(n14237), .A2(n14236), .ZN(n14238) );
  OR2_X1 U16153 ( .A1(n14197), .A2(n14238), .ZN(n18139) );
  NOR2_X1 U16154 ( .A1(n18139), .A2(n16046), .ZN(n14243) );
  AOI211_X1 U16155 ( .C1(n14241), .C2(n14240), .A(n16115), .B(n14239), .ZN(
        n14242) );
  AOI211_X1 U16156 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n16046), .A(n14243), .B(
        n14242), .ZN(n14244) );
  INV_X1 U16157 ( .A(n14244), .ZN(P2_U2877) );
  INV_X1 U16158 ( .A(n14246), .ZN(n14248) );
  INV_X1 U16159 ( .A(n14403), .ZN(n14247) );
  OAI21_X1 U16160 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14248), .A(
        n14247), .ZN(n21449) );
  AOI22_X1 U16161 ( .A1(n15161), .A2(n21449), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14249) );
  OAI21_X1 U16162 ( .B1(n15087), .B2(n19796), .A(n14249), .ZN(n14250) );
  INV_X1 U16163 ( .A(n14421), .ZN(n14422) );
  NAND2_X1 U16164 ( .A1(n14252), .A2(n14253), .ZN(n14254) );
  AND2_X1 U16165 ( .A1(n14422), .A2(n14254), .ZN(n21455) );
  INV_X1 U16166 ( .A(n21455), .ZN(n14259) );
  INV_X1 U16167 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14258) );
  INV_X1 U16168 ( .A(n14425), .ZN(n14255) );
  OAI21_X1 U16169 ( .B1(n14257), .B2(n14256), .A(n14255), .ZN(n21458) );
  OAI222_X1 U16170 ( .A1(n14259), .A2(n15509), .B1(n14258), .B2(n19892), .C1(
        n21458), .C2(n15497), .ZN(P1_U2865) );
  INV_X1 U16171 ( .A(n22198), .ZN(n15545) );
  OAI222_X1 U16172 ( .A1(n15587), .A2(n14259), .B1(n15553), .B2(n19796), .C1(
        n15585), .C2(n15545), .ZN(P1_U2897) );
  MUX2_X1 U16173 ( .A(n15161), .B(n21908), .S(n16765), .Z(n14260) );
  NOR2_X1 U16174 ( .A1(n21859), .A2(n21196), .ZN(n21622) );
  MUX2_X1 U16175 ( .A(n14260), .B(n21622), .S(P1_STATE2_REG_0__SCAN_IN), .Z(
        n14261) );
  INV_X1 U16176 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14848) );
  INV_X1 U16177 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15383) );
  INV_X1 U16178 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15656) );
  INV_X1 U16179 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15026) );
  INV_X1 U16180 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15089) );
  INV_X1 U16181 ( .A(n15111), .ZN(n14265) );
  NAND2_X1 U16182 ( .A1(n14265), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15134) );
  INV_X1 U16183 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15133) );
  INV_X1 U16184 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15260) );
  INV_X1 U16185 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14266) );
  NOR2_X1 U16186 ( .A1(n15169), .A2(n16765), .ZN(n14268) );
  AND3_X1 U16187 ( .A1(n12985), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n14709), 
        .ZN(n14269) );
  INV_X1 U16188 ( .A(n21428), .ZN(n15413) );
  INV_X1 U16189 ( .A(n14271), .ZN(n14291) );
  INV_X1 U16190 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14289) );
  AND2_X1 U16191 ( .A1(n14272), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14273) );
  AND2_X1 U16192 ( .A1(n21660), .A2(n21881), .ZN(n16757) );
  AND2_X1 U16193 ( .A1(n14274), .A2(n16757), .ZN(n14280) );
  INV_X1 U16194 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21231) );
  OAI21_X1 U16195 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21544), .A(n14709), .ZN(
        n15407) );
  AOI21_X1 U16196 ( .B1(n21436), .B2(n21231), .A(n15407), .ZN(n14288) );
  NAND2_X1 U16197 ( .A1(n14289), .A2(n14288), .ZN(n14287) );
  NOR2_X1 U16198 ( .A1(n14275), .A2(n21898), .ZN(n14276) );
  AND2_X1 U16199 ( .A1(n14709), .A2(n14276), .ZN(n21411) );
  NAND2_X1 U16200 ( .A1(n12978), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14278) );
  NOR2_X1 U16201 ( .A1(n14278), .A2(n16757), .ZN(n14277) );
  INV_X1 U16202 ( .A(n14278), .ZN(n14279) );
  NOR2_X1 U16203 ( .A1(n14280), .A2(n14279), .ZN(n14281) );
  AOI22_X1 U16204 ( .A1(n21597), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n21553), .ZN(n14283) );
  OAI21_X1 U16205 ( .B1(n21592), .B2(n14284), .A(n14283), .ZN(n14285) );
  AOI21_X1 U16206 ( .B1(n21411), .B2(n21804), .A(n14285), .ZN(n14286) );
  OAI221_X1 U16207 ( .B1(n14289), .B2(n14288), .C1(n14287), .C2(n21544), .A(
        n14286), .ZN(n14290) );
  AOI21_X1 U16208 ( .B1(n21586), .B2(n14291), .A(n14290), .ZN(n14292) );
  OAI21_X1 U16209 ( .B1(n15413), .B2(n14293), .A(n14292), .ZN(P1_U2837) );
  AOI22_X1 U16210 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19797), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n19813), .ZN(n14294) );
  OAI21_X1 U16211 ( .B1(n14295), .B2(n14326), .A(n14294), .ZN(P1_U2920) );
  AOI22_X1 U16212 ( .A1(n19797), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14296) );
  OAI21_X1 U16213 ( .B1(n14297), .B2(n14326), .A(n14296), .ZN(P1_U2913) );
  INV_X1 U16214 ( .A(n14298), .ZN(n14299) );
  OAI21_X1 U16215 ( .B1(n14196), .B2(n14300), .A(n14299), .ZN(n18162) );
  INV_X1 U16216 ( .A(n14301), .ZN(n14302) );
  OAI211_X1 U16217 ( .C1(n14302), .C2(n11389), .A(n16082), .B(n14435), .ZN(
        n14304) );
  NAND2_X1 U16218 ( .A1(n16046), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14303) );
  OAI211_X1 U16219 ( .C1(n18162), .C2(n16046), .A(n14304), .B(n14303), .ZN(
        P2_U2875) );
  AOI22_X1 U16220 ( .A1(n21200), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14305) );
  OAI21_X1 U16221 ( .B1(n14306), .B2(n14326), .A(n14305), .ZN(P1_U2912) );
  AOI22_X1 U16222 ( .A1(n21200), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14307) );
  OAI21_X1 U16223 ( .B1(n14308), .B2(n14326), .A(n14307), .ZN(P1_U2914) );
  AOI22_X1 U16224 ( .A1(n21200), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14309) );
  OAI21_X1 U16225 ( .B1(n14310), .B2(n14326), .A(n14309), .ZN(P1_U2909) );
  AOI22_X1 U16226 ( .A1(n21200), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14311) );
  OAI21_X1 U16227 ( .B1(n14312), .B2(n14326), .A(n14311), .ZN(P1_U2908) );
  AOI22_X1 U16228 ( .A1(n21200), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14313) );
  OAI21_X1 U16229 ( .B1(n14314), .B2(n14326), .A(n14313), .ZN(P1_U2911) );
  AOI22_X1 U16230 ( .A1(n21200), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U16231 ( .B1(n14316), .B2(n14326), .A(n14315), .ZN(P1_U2906) );
  AOI22_X1 U16232 ( .A1(n21200), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14317) );
  OAI21_X1 U16233 ( .B1(n14318), .B2(n14326), .A(n14317), .ZN(P1_U2910) );
  AOI22_X1 U16234 ( .A1(n21200), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14319) );
  OAI21_X1 U16235 ( .B1(n14320), .B2(n14326), .A(n14319), .ZN(P1_U2915) );
  AOI22_X1 U16236 ( .A1(n21200), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14321) );
  OAI21_X1 U16237 ( .B1(n14322), .B2(n14326), .A(n14321), .ZN(P1_U2917) );
  AOI22_X1 U16238 ( .A1(n21200), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U16239 ( .B1(n14324), .B2(n14326), .A(n14323), .ZN(P1_U2907) );
  AOI22_X1 U16240 ( .A1(n21200), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14325) );
  OAI21_X1 U16241 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(P1_U2916) );
  INV_X1 U16242 ( .A(n14434), .ZN(n14433) );
  XNOR2_X1 U16243 ( .A(n14435), .B(n14433), .ZN(n14332) );
  OR2_X1 U16244 ( .A1(n14328), .A2(n14298), .ZN(n14329) );
  AND2_X1 U16245 ( .A1(n14431), .A2(n14329), .ZN(n18454) );
  INV_X1 U16246 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18164) );
  NOR2_X1 U16247 ( .A1(n16112), .A2(n18164), .ZN(n14330) );
  AOI21_X1 U16248 ( .B1(n16112), .B2(n18454), .A(n14330), .ZN(n14331) );
  OAI21_X1 U16249 ( .B1(n14332), .B2(n16115), .A(n14331), .ZN(P2_U2874) );
  NOR2_X2 U16250 ( .A1(n19083), .A2(n19143), .ZN(n19630) );
  NOR2_X2 U16251 ( .A1(n19192), .A2(n19051), .ZN(n19623) );
  OAI21_X1 U16252 ( .B1(n19630), .B2(n19623), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14342) );
  INV_X1 U16253 ( .A(n19114), .ZN(n14334) );
  NOR2_X1 U16254 ( .A1(n14334), .A2(n14333), .ZN(n19145) );
  NAND2_X1 U16255 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19145), .ZN(
        n14341) );
  NAND3_X1 U16256 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19179), .ZN(n19050) );
  NOR2_X1 U16257 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19050), .ZN(
        n19621) );
  AOI21_X1 U16258 ( .B1(n16714), .B2(n19164), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18528) );
  AND2_X1 U16259 ( .A1(n14336), .A2(n18528), .ZN(n14338) );
  INV_X1 U16260 ( .A(n14338), .ZN(n14337) );
  AOI21_X1 U16261 ( .B1(n19621), .B2(n19219), .A(n19215), .ZN(n14340) );
  NAND2_X1 U16262 ( .A1(n19183), .A2(n14338), .ZN(n19202) );
  INV_X1 U16263 ( .A(n19202), .ZN(n19216) );
  NAND2_X1 U16264 ( .A1(n14344), .A2(n19216), .ZN(n14339) );
  AOI22_X1 U16265 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19592), .ZN(n19585) );
  INV_X1 U16266 ( .A(n19585), .ZN(n19574) );
  AOI22_X2 U16267 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19592), .ZN(n19580) );
  INV_X1 U16268 ( .A(n19580), .ZN(n19552) );
  AOI22_X1 U16269 ( .A1(n19630), .A2(n19574), .B1(n19623), .B2(n19552), .ZN(
        n14349) );
  INV_X1 U16270 ( .A(n14343), .ZN(n14347) );
  INV_X1 U16271 ( .A(n19145), .ZN(n14346) );
  OAI21_X1 U16272 ( .B1(n14344), .B2(n19621), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14345) );
  OAI21_X1 U16273 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n19622) );
  NOR2_X2 U16274 ( .A1(n19532), .A2(n19594), .ZN(n19582) );
  NAND2_X1 U16275 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19219), .ZN(n19354) );
  AOI22_X1 U16276 ( .A1(n19622), .A2(n19582), .B1(n19621), .B2(n19573), .ZN(
        n14348) );
  OAI211_X1 U16277 ( .C1(n19626), .C2(n14562), .A(n14349), .B(n14348), .ZN(
        P2_U3145) );
  INV_X1 U16278 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15852) );
  AOI22_X1 U16279 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19592), .ZN(n19276) );
  INV_X1 U16280 ( .A(n19276), .ZN(n19264) );
  INV_X1 U16281 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n22153) );
  INV_X1 U16282 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20599) );
  OAI22_X1 U16283 ( .A1(n22153), .A2(n19602), .B1(n20599), .B2(n19600), .ZN(
        n19272) );
  AOI22_X1 U16284 ( .A1(n19630), .A2(n19264), .B1(n19623), .B2(n19272), .ZN(
        n14351) );
  NOR2_X2 U16285 ( .A1(n19230), .A2(n19594), .ZN(n19273) );
  AND2_X1 U16286 ( .A1(n11873), .A2(n19596), .ZN(n19271) );
  AOI22_X1 U16287 ( .A1(n19622), .A2(n19273), .B1(n19621), .B2(n19271), .ZN(
        n14350) );
  OAI211_X1 U16288 ( .C1(n19626), .C2(n15852), .A(n14351), .B(n14350), .ZN(
        P2_U3150) );
  XNOR2_X1 U16289 ( .A(n14353), .B(n14352), .ZN(n14370) );
  XNOR2_X1 U16290 ( .A(n14382), .B(n14365), .ZN(n14384) );
  XNOR2_X1 U16291 ( .A(n14384), .B(n14354), .ZN(n14362) );
  NAND2_X1 U16292 ( .A1(n14362), .A2(n17032), .ZN(n14361) );
  INV_X1 U16293 ( .A(n15814), .ZN(n14355) );
  INV_X1 U16294 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15826) );
  OAI22_X1 U16295 ( .A1(n17018), .A2(n15826), .B1(n14356), .B2(n18475), .ZN(
        n14359) );
  OAI21_X1 U16296 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14357), .A(
        n14395), .ZN(n18062) );
  NOR2_X1 U16297 ( .A1(n17042), .A2(n18062), .ZN(n14358) );
  AOI211_X1 U16298 ( .C1(n17021), .C2(n14355), .A(n14359), .B(n14358), .ZN(
        n14360) );
  OAI211_X1 U16299 ( .C1(n14370), .C2(n17024), .A(n14361), .B(n14360), .ZN(
        P2_U3011) );
  NAND2_X1 U16300 ( .A1(n14362), .A2(n18501), .ZN(n14369) );
  NOR2_X1 U16301 ( .A1(n18489), .A2(n18486), .ZN(n14363) );
  OR2_X1 U16302 ( .A1(n14364), .A2(n14363), .ZN(n14615) );
  MUX2_X1 U16303 ( .A(n14615), .B(n14612), .S(n14365), .Z(n14367) );
  OAI22_X1 U16304 ( .A1(n17056), .A2(n18490), .B1(n14356), .B2(n18475), .ZN(
        n14366) );
  AOI211_X1 U16305 ( .C1(n18500), .C2(n14355), .A(n14367), .B(n14366), .ZN(
        n14368) );
  OAI211_X1 U16306 ( .C1(n14370), .C2(n18494), .A(n14369), .B(n14368), .ZN(
        P2_U3043) );
  INV_X1 U16307 ( .A(n21411), .ZN(n14381) );
  NAND2_X1 U16308 ( .A1(n16959), .A2(n21428), .ZN(n14380) );
  INV_X1 U16309 ( .A(n21553), .ZN(n21609) );
  INV_X1 U16310 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14374) );
  NAND2_X1 U16311 ( .A1(n21605), .A2(n21233), .ZN(n14373) );
  INV_X1 U16312 ( .A(n16957), .ZN(n14371) );
  AOI22_X1 U16313 ( .A1(n21586), .A2(n14371), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n15407), .ZN(n14372) );
  OAI211_X1 U16314 ( .C1(n21609), .C2(n14374), .A(n14373), .B(n14372), .ZN(
        n14378) );
  NAND2_X1 U16315 ( .A1(n21231), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U16316 ( .A1(n21597), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14375) );
  OAI21_X1 U16317 ( .B1(n14376), .B2(n21544), .A(n14375), .ZN(n14377) );
  NOR2_X1 U16318 ( .A1(n14378), .A2(n14377), .ZN(n14379) );
  OAI211_X1 U16319 ( .C1(n14381), .C2(n21850), .A(n14380), .B(n14379), .ZN(
        P1_U2838) );
  AOI22_X1 U16320 ( .A1(n14384), .A2(n14383), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14382), .ZN(n14386) );
  XNOR2_X1 U16321 ( .A(n18056), .B(n14544), .ZN(n14385) );
  XNOR2_X1 U16322 ( .A(n14386), .B(n14385), .ZN(n14402) );
  OAI21_X1 U16323 ( .B1(n14388), .B2(n14544), .A(n14387), .ZN(n14400) );
  NAND2_X1 U16324 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14612), .ZN(
        n14543) );
  NOR2_X1 U16325 ( .A1(n18422), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14389) );
  NOR2_X1 U16326 ( .A1(n14615), .A2(n14389), .ZN(n14549) );
  NAND2_X1 U16327 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16539), .ZN(n14390) );
  OAI221_X1 U16328 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14543), .C1(
        n14544), .C2(n14549), .A(n14390), .ZN(n14393) );
  INV_X1 U16329 ( .A(n18500), .ZN(n16567) );
  OAI22_X1 U16330 ( .A1(n18068), .A2(n16567), .B1(n18490), .B2(n14391), .ZN(
        n14392) );
  AOI211_X1 U16331 ( .C1(n14400), .C2(n18481), .A(n14393), .B(n14392), .ZN(
        n14394) );
  OAI21_X1 U16332 ( .B1(n14402), .B2(n18450), .A(n14394), .ZN(P2_U3042) );
  AOI21_X1 U16333 ( .B1(n14396), .B2(n14395), .A(n16967), .ZN(n18074) );
  OAI22_X1 U16334 ( .A1(n14396), .A2(n17018), .B1(n12673), .B2(n18240), .ZN(
        n14397) );
  AOI21_X1 U16335 ( .B1(n17005), .B2(n18074), .A(n14397), .ZN(n14398) );
  OAI21_X1 U16336 ( .B1(n17038), .B2(n18068), .A(n14398), .ZN(n14399) );
  AOI21_X1 U16337 ( .B1(n14400), .B2(n17035), .A(n14399), .ZN(n14401) );
  OAI21_X1 U16338 ( .B1(n14402), .B2(n17014), .A(n14401), .ZN(P2_U3010) );
  XNOR2_X1 U16339 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n14403), .ZN(
        n15185) );
  AOI22_X1 U16340 ( .A1(n15161), .A2(n15185), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14404) );
  OAI21_X1 U16341 ( .B1(n15087), .B2(n19799), .A(n14404), .ZN(n14405) );
  INV_X1 U16342 ( .A(n14405), .ZN(n14419) );
  AOI22_X1 U16343 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U16344 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U16345 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16346 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14407) );
  NAND4_X1 U16347 ( .A1(n14410), .A2(n14409), .A3(n14408), .A4(n14407), .ZN(
        n14417) );
  AOI22_X1 U16348 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U16349 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U16350 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U16351 ( .A1(n15145), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14412) );
  NAND4_X1 U16352 ( .A1(n14415), .A2(n14414), .A3(n14413), .A4(n14412), .ZN(
        n14416) );
  OAI21_X1 U16353 ( .B1(n14417), .B2(n14416), .A(n14656), .ZN(n14418) );
  AOI21_X1 U16354 ( .B1(n14423), .B2(n14422), .A(n11236), .ZN(n15187) );
  INV_X1 U16355 ( .A(n15509), .ZN(n19889) );
  OR2_X1 U16356 ( .A1(n14425), .A2(n14424), .ZN(n14426) );
  NAND2_X1 U16357 ( .A1(n14462), .A2(n14426), .ZN(n21286) );
  OAI22_X1 U16358 ( .A1(n21286), .A2(n15497), .B1(n14427), .B2(n19892), .ZN(
        n14428) );
  AOI21_X1 U16359 ( .B1(n15187), .B2(n19889), .A(n14428), .ZN(n14429) );
  INV_X1 U16360 ( .A(n14429), .ZN(P1_U2864) );
  NAND2_X1 U16361 ( .A1(n14431), .A2(n14430), .ZN(n14432) );
  AND2_X1 U16362 ( .A1(n14496), .A2(n14432), .ZN(n18186) );
  INV_X1 U16363 ( .A(n18186), .ZN(n14441) );
  NOR2_X1 U16364 ( .A1(n14435), .A2(n14433), .ZN(n14438) );
  INV_X1 U16365 ( .A(n14498), .ZN(n14436) );
  OAI211_X1 U16366 ( .C1(n14438), .C2(n14437), .A(n14436), .B(n16082), .ZN(
        n14440) );
  NAND2_X1 U16367 ( .A1(n16046), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14439) );
  OAI211_X1 U16368 ( .C1(n14441), .C2(n16046), .A(n14440), .B(n14439), .ZN(
        P2_U2873) );
  INV_X1 U16369 ( .A(n15187), .ZN(n14473) );
  OAI222_X1 U16370 ( .A1(n15585), .A2(n15541), .B1(n19799), .B2(n15553), .C1(
        n14473), .C2(n15587), .ZN(P1_U2896) );
  XOR2_X1 U16371 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n14442), .Z(n21468) );
  INV_X1 U16372 ( .A(n21468), .ZN(n15177) );
  INV_X1 U16373 ( .A(n14656), .ZN(n14862) );
  AOI22_X1 U16374 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15100), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U16375 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10981), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U16376 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U16377 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14443) );
  NAND4_X1 U16378 ( .A1(n14446), .A2(n14445), .A3(n14444), .A4(n14443), .ZN(
        n14452) );
  AOI22_X1 U16379 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U16380 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n13007), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U16381 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10966), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16382 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14447) );
  NAND4_X1 U16383 ( .A1(n14450), .A2(n14449), .A3(n14448), .A4(n14447), .ZN(
        n14451) );
  NOR2_X1 U16384 ( .A1(n14452), .A2(n14451), .ZN(n14455) );
  NAND2_X1 U16385 ( .A1(n15165), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n14454) );
  NAND2_X1 U16386 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14453) );
  OAI211_X1 U16387 ( .C1(n14862), .C2(n14455), .A(n14454), .B(n14453), .ZN(
        n14456) );
  AOI21_X1 U16388 ( .B1(n15177), .B2(n15161), .A(n14456), .ZN(n14459) );
  AOI21_X1 U16389 ( .B1(n14459), .B2(n14458), .A(n14492), .ZN(n15179) );
  INV_X1 U16390 ( .A(n15179), .ZN(n21466) );
  INV_X1 U16391 ( .A(n14798), .ZN(n14460) );
  AOI21_X1 U16392 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n21464) );
  AOI22_X1 U16393 ( .A1(n21464), .A2(n19888), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15507), .ZN(n14463) );
  OAI21_X1 U16394 ( .B1(n21466), .B2(n15509), .A(n14463), .ZN(P1_U2863) );
  NAND4_X1 U16395 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n21420)
         );
  INV_X1 U16396 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21432) );
  NOR2_X1 U16397 ( .A1(n21420), .A2(n21432), .ZN(n21433) );
  NAND2_X1 U16398 ( .A1(n21433), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n21445) );
  INV_X1 U16399 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21453) );
  NOR2_X1 U16400 ( .A1(n21445), .A2(n21453), .ZN(n14470) );
  NAND2_X1 U16401 ( .A1(n14470), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n21461) );
  AND2_X1 U16402 ( .A1(n21461), .A2(n21436), .ZN(n14471) );
  INV_X1 U16403 ( .A(n15185), .ZN(n14465) );
  NAND2_X1 U16404 ( .A1(n14709), .A2(n14464), .ZN(n21529) );
  AOI21_X1 U16405 ( .B1(n21586), .B2(n14465), .A(n21519), .ZN(n14466) );
  OAI21_X1 U16406 ( .B1(n21286), .B2(n21592), .A(n14466), .ZN(n14469) );
  INV_X1 U16407 ( .A(n14709), .ZN(n21435) );
  AOI21_X1 U16408 ( .B1(n21436), .B2(n21461), .A(n21435), .ZN(n21471) );
  INV_X1 U16409 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21285) );
  AOI22_X1 U16410 ( .A1(n21597), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n21553), .ZN(n14467) );
  OAI21_X1 U16411 ( .B1(n21471), .B2(n21285), .A(n14467), .ZN(n14468) );
  AOI211_X1 U16412 ( .C1(n14471), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        n14472) );
  OAI21_X1 U16413 ( .B1(n14473), .B2(n21602), .A(n14472), .ZN(P1_U2832) );
  OAI222_X1 U16414 ( .A1(n15585), .A2(n15537), .B1(n19801), .B2(n15553), .C1(
        n21466), .C2(n15587), .ZN(P1_U2895) );
  XNOR2_X1 U16415 ( .A(n14475), .B(n14474), .ZN(n15708) );
  NAND2_X1 U16416 ( .A1(n15708), .A2(n15161), .ZN(n14491) );
  AOI22_X1 U16417 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U16418 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U16419 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16420 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14476) );
  NAND4_X1 U16421 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14485) );
  AOI22_X1 U16422 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U16423 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U16424 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U16425 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14480) );
  NAND4_X1 U16426 ( .A1(n14483), .A2(n14482), .A3(n14481), .A4(n14480), .ZN(
        n14484) );
  NOR2_X1 U16427 ( .A1(n14485), .A2(n14484), .ZN(n14488) );
  NAND2_X1 U16428 ( .A1(n15165), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U16429 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14486) );
  OAI211_X1 U16430 ( .C1(n14862), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14489) );
  INV_X1 U16431 ( .A(n14489), .ZN(n14490) );
  NAND2_X1 U16432 ( .A1(n14491), .A2(n14490), .ZN(n14493) );
  OAI21_X1 U16433 ( .B1(n14492), .B2(n14493), .A(n14678), .ZN(n15706) );
  XNOR2_X1 U16434 ( .A(n14798), .B(n14795), .ZN(n21305) );
  AOI22_X1 U16435 ( .A1(n21305), .A2(n19888), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n15507), .ZN(n14494) );
  OAI21_X1 U16436 ( .B1(n15706), .B2(n15509), .A(n14494), .ZN(P1_U2862) );
  NAND2_X1 U16437 ( .A1(n14496), .A2(n14495), .ZN(n14497) );
  AND2_X1 U16438 ( .A1(n14535), .A2(n14497), .ZN(n18197) );
  INV_X1 U16439 ( .A(n18197), .ZN(n14503) );
  INV_X1 U16440 ( .A(n14521), .ZN(n14499) );
  OAI211_X1 U16441 ( .C1(n14498), .C2(n14500), .A(n14499), .B(n16082), .ZN(
        n14502) );
  NAND2_X1 U16442 ( .A1(n16046), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14501) );
  OAI211_X1 U16443 ( .C1(n14503), .C2(n16046), .A(n14502), .B(n14501), .ZN(
        P2_U2872) );
  AOI22_X1 U16444 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16445 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U16446 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14504) );
  NAND3_X1 U16447 ( .A1(n14506), .A2(n14505), .A3(n14504), .ZN(n14520) );
  NAND2_X1 U16448 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14508) );
  NAND2_X1 U16449 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14507) );
  OAI211_X1 U16450 ( .C1(n15874), .C2(n14509), .A(n14508), .B(n14507), .ZN(
        n14514) );
  INV_X1 U16451 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U16452 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14511) );
  NAND2_X1 U16453 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14510) );
  OAI211_X1 U16454 ( .C1(n12015), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14513) );
  NOR2_X1 U16455 ( .A1(n14514), .A2(n14513), .ZN(n14518) );
  AOI22_X1 U16456 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U16457 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14516) );
  NAND2_X1 U16458 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14515) );
  NAND4_X1 U16459 ( .A1(n14518), .A2(n14517), .A3(n14516), .A4(n14515), .ZN(
        n14519) );
  OR2_X1 U16460 ( .A1(n14520), .A2(n14519), .ZN(n14522) );
  OAI21_X1 U16461 ( .B1(n14521), .B2(n14522), .A(n14767), .ZN(n14539) );
  XNOR2_X1 U16462 ( .A(n10984), .B(n14523), .ZN(n18209) );
  INV_X1 U16463 ( .A(n18209), .ZN(n14532) );
  INV_X1 U16464 ( .A(n14529), .ZN(n14525) );
  NOR2_X1 U16465 ( .A1(n14525), .A2(n14524), .ZN(n16211) );
  INV_X1 U16466 ( .A(n16211), .ZN(n19462) );
  OAI22_X1 U16467 ( .A1(n19462), .A2(n19595), .B1(n19278), .B2(n13855), .ZN(
        n14531) );
  AND2_X1 U16468 ( .A1(n11873), .A2(n14526), .ZN(n14527) );
  INV_X1 U16469 ( .A(n18996), .ZN(n19463) );
  INV_X1 U16470 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18892) );
  AND2_X1 U16471 ( .A1(n11873), .A2(n16187), .ZN(n14528) );
  NAND2_X1 U16472 ( .A1(n14529), .A2(n14528), .ZN(n19474) );
  OAI22_X1 U16473 ( .A1(n19463), .A2(n21727), .B1(n18892), .B2(n19474), .ZN(
        n14530) );
  AOI211_X1 U16474 ( .C1(n14532), .C2(n19345), .A(n14531), .B(n14530), .ZN(
        n14533) );
  OAI21_X1 U16475 ( .B1(n19468), .B2(n14539), .A(n14533), .ZN(P2_U2903) );
  OAI222_X1 U16476 ( .A1(n15585), .A2(n15532), .B1(n19804), .B2(n15553), .C1(
        n15706), .C2(n15587), .ZN(P1_U2894) );
  AND2_X1 U16477 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  OR2_X1 U16478 ( .A1(n14536), .A2(n14582), .ZN(n18210) );
  NOR2_X1 U16479 ( .A1(n16046), .A2(n18210), .ZN(n14537) );
  AOI21_X1 U16480 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16046), .A(n14537), .ZN(
        n14538) );
  OAI21_X1 U16481 ( .B1(n14539), .B2(n16115), .A(n14538), .ZN(P2_U2871) );
  XNOR2_X1 U16482 ( .A(n14540), .B(n14548), .ZN(n16969) );
  XNOR2_X1 U16483 ( .A(n14541), .B(n14542), .ZN(n16968) );
  INV_X1 U16484 ( .A(n16968), .ZN(n14555) );
  AOI221_X1 U16485 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n14544), .C2(n14548), .A(
        n14543), .ZN(n14554) );
  OAI21_X1 U16486 ( .B1(n14207), .B2(n14546), .A(n14545), .ZN(n19286) );
  INV_X1 U16487 ( .A(n19286), .ZN(n14551) );
  INV_X1 U16488 ( .A(n18490), .ZN(n18466) );
  OAI22_X1 U16489 ( .A1(n14549), .A2(n14548), .B1(n18240), .B2(n14547), .ZN(
        n14550) );
  AOI21_X1 U16490 ( .B1(n14551), .B2(n18466), .A(n14550), .ZN(n14552) );
  OAI21_X1 U16491 ( .B1(n16567), .B2(n18076), .A(n14552), .ZN(n14553) );
  AOI211_X1 U16492 ( .C1(n14555), .C2(n18501), .A(n14554), .B(n14553), .ZN(
        n14556) );
  OAI21_X1 U16493 ( .B1(n18494), .B2(n16969), .A(n14556), .ZN(P2_U3041) );
  INV_X1 U16494 ( .A(n14767), .ZN(n14579) );
  AOI22_X1 U16495 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14559) );
  AOI22_X1 U16496 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U16497 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14557) );
  NAND3_X1 U16498 ( .A1(n14559), .A2(n14558), .A3(n14557), .ZN(n14577) );
  NAND2_X1 U16499 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14561) );
  NAND2_X1 U16500 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14560) );
  OAI211_X1 U16501 ( .C1(n15874), .C2(n14562), .A(n14561), .B(n14560), .ZN(
        n14567) );
  NAND2_X1 U16502 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14564) );
  NAND2_X1 U16503 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14563) );
  OAI211_X1 U16504 ( .C1(n12015), .C2(n14565), .A(n14564), .B(n14563), .ZN(
        n14566) );
  NOR2_X1 U16505 ( .A1(n14567), .A2(n14566), .ZN(n14575) );
  AOI22_X1 U16506 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14574) );
  OAI22_X1 U16507 ( .A1(n14571), .A2(n14570), .B1(n14569), .B2(n14568), .ZN(
        n14572) );
  INV_X1 U16508 ( .A(n14572), .ZN(n14573) );
  NAND3_X1 U16509 ( .A1(n14575), .A2(n14574), .A3(n14573), .ZN(n14576) );
  NOR2_X1 U16510 ( .A1(n14577), .A2(n14576), .ZN(n14764) );
  INV_X1 U16511 ( .A(n14764), .ZN(n14578) );
  OAI21_X1 U16512 ( .B1(n14579), .B2(n14578), .A(n14602), .ZN(n16214) );
  OAI21_X1 U16513 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n16382) );
  NOR2_X1 U16514 ( .A1(n16382), .A2(n16046), .ZN(n14583) );
  AOI21_X1 U16515 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16046), .A(n14583), .ZN(
        n14584) );
  OAI21_X1 U16516 ( .B1(n16214), .B2(n16115), .A(n14584), .ZN(P2_U2870) );
  AOI22_X1 U16517 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U16518 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14586) );
  AOI22_X1 U16519 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14585) );
  NAND3_X1 U16520 ( .A1(n14587), .A2(n14586), .A3(n14585), .ZN(n14601) );
  INV_X1 U16521 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U16522 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14589) );
  NAND2_X1 U16523 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14588) );
  OAI211_X1 U16524 ( .C1(n15874), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14595) );
  INV_X1 U16525 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U16526 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14592) );
  NAND2_X1 U16527 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14591) );
  OAI211_X1 U16528 ( .C1(n12015), .C2(n14593), .A(n14592), .B(n14591), .ZN(
        n14594) );
  NOR2_X1 U16529 ( .A1(n14595), .A2(n14594), .ZN(n14599) );
  AOI22_X1 U16530 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14598) );
  NAND2_X1 U16531 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14597) );
  NAND2_X1 U16532 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14596) );
  NAND4_X1 U16533 ( .A1(n14599), .A2(n14598), .A3(n14597), .A4(n14596), .ZN(
        n14600) );
  NOR2_X1 U16534 ( .A1(n14601), .A2(n14600), .ZN(n14763) );
  NAND2_X1 U16535 ( .A1(n14602), .A2(n14763), .ZN(n14603) );
  NAND2_X1 U16536 ( .A1(n14805), .A2(n14603), .ZN(n19469) );
  NAND2_X1 U16537 ( .A1(n16046), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14607) );
  NAND2_X1 U16538 ( .A1(n14580), .A2(n14604), .ZN(n14605) );
  AND2_X1 U16539 ( .A1(n11029), .A2(n14605), .ZN(n18235) );
  NAND2_X1 U16540 ( .A1(n18235), .A2(n16112), .ZN(n14606) );
  OAI211_X1 U16541 ( .C1(n19469), .C2(n16115), .A(n14607), .B(n14606), .ZN(
        P2_U2869) );
  XNOR2_X1 U16542 ( .A(n14609), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14629) );
  XOR2_X1 U16543 ( .A(n14610), .B(n14611), .Z(n14627) );
  INV_X1 U16544 ( .A(n14612), .ZN(n14614) );
  NAND3_X1 U16545 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14613) );
  NOR2_X1 U16546 ( .A1(n14614), .A2(n14613), .ZN(n14734) );
  AOI21_X1 U16547 ( .B1(n18460), .B2(n14616), .A(n14615), .ZN(n18485) );
  INV_X1 U16548 ( .A(n18485), .ZN(n14618) );
  NOR2_X1 U16549 ( .A1(n12682), .A2(n18240), .ZN(n14617) );
  AOI221_X1 U16550 ( .B1(n14734), .B2(n12221), .C1(n14618), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n14617), .ZN(n14620) );
  NAND2_X1 U16551 ( .A1(n18089), .A2(n18500), .ZN(n14619) );
  OAI211_X1 U16552 ( .C1(n18490), .C2(n18093), .A(n14620), .B(n14619), .ZN(
        n14621) );
  AOI21_X1 U16553 ( .B1(n14627), .B2(n18501), .A(n14621), .ZN(n14622) );
  OAI21_X1 U16554 ( .B1(n14629), .B2(n18494), .A(n14622), .ZN(P2_U3040) );
  AOI21_X1 U16555 ( .B1(n18083), .B2(n16966), .A(n14729), .ZN(n18099) );
  OAI22_X1 U16556 ( .A1(n18083), .A2(n17018), .B1(n12682), .B2(n18240), .ZN(
        n14623) );
  AOI21_X1 U16557 ( .B1(n17005), .B2(n18099), .A(n14623), .ZN(n14624) );
  OAI21_X1 U16558 ( .B1(n14625), .B2(n17038), .A(n14624), .ZN(n14626) );
  AOI21_X1 U16559 ( .B1(n14627), .B2(n17032), .A(n14626), .ZN(n14628) );
  OAI21_X1 U16560 ( .B1(n14629), .B2(n17024), .A(n14628), .ZN(P2_U3008) );
  OAI21_X1 U16561 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14631), .A(
        n14630), .ZN(n21480) );
  AOI22_X1 U16562 ( .A1(n15161), .A2(n21480), .B1(n15164), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14632) );
  OAI21_X1 U16563 ( .B1(n15087), .B2(n19806), .A(n14632), .ZN(n14633) );
  NAND2_X1 U16564 ( .A1(n14678), .A2(n11239), .ZN(n14634) );
  NAND2_X1 U16565 ( .A1(n14680), .A2(n14634), .ZN(n14713) );
  AOI22_X1 U16566 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U16567 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U16568 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U16569 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14635) );
  NAND4_X1 U16570 ( .A1(n14638), .A2(n14637), .A3(n14636), .A4(n14635), .ZN(
        n14644) );
  AOI22_X1 U16571 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14651), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14642) );
  AOI22_X1 U16572 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14641) );
  AOI22_X1 U16573 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16574 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14639) );
  NAND4_X1 U16575 ( .A1(n14642), .A2(n14641), .A3(n14640), .A4(n14639), .ZN(
        n14643) );
  OR2_X1 U16576 ( .A1(n14644), .A2(n14643), .ZN(n14645) );
  NAND2_X1 U16577 ( .A1(n14656), .A2(n14645), .ZN(n14714) );
  OAI21_X1 U16578 ( .B1(n14713), .B2(n14714), .A(n14680), .ZN(n14716) );
  XOR2_X1 U16579 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n14646), .Z(
        n21490) );
  AOI22_X1 U16580 ( .A1(n15165), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n15164), 
        .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U16581 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14650) );
  AOI22_X1 U16582 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U16583 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U16584 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14647) );
  NAND4_X1 U16585 ( .A1(n14650), .A2(n14649), .A3(n14648), .A4(n14647), .ZN(
        n14658) );
  AOI22_X1 U16586 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14651), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U16587 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U16588 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U16589 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14652) );
  NAND4_X1 U16590 ( .A1(n14655), .A2(n14654), .A3(n14653), .A4(n14652), .ZN(
        n14657) );
  OAI21_X1 U16591 ( .B1(n14658), .B2(n14657), .A(n14656), .ZN(n14659) );
  OAI211_X1 U16592 ( .C1(n21490), .C2(n14136), .A(n14660), .B(n14659), .ZN(
        n14715) );
  NAND2_X1 U16593 ( .A1(n14716), .A2(n14715), .ZN(n14718) );
  XOR2_X1 U16594 ( .A(n14662), .B(n14661), .Z(n14705) );
  AOI22_X1 U16595 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U16596 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U16597 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U16598 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14663) );
  NAND4_X1 U16599 ( .A1(n14666), .A2(n14665), .A3(n14664), .A4(n14663), .ZN(
        n14672) );
  AOI22_X1 U16600 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14670) );
  AOI22_X1 U16601 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15000), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14669) );
  AOI22_X1 U16602 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14668) );
  AOI22_X1 U16603 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14667) );
  NAND4_X1 U16604 ( .A1(n14670), .A2(n14669), .A3(n14668), .A4(n14667), .ZN(
        n14671) );
  NOR2_X1 U16605 ( .A1(n14672), .A2(n14671), .ZN(n14675) );
  NAND2_X1 U16606 ( .A1(n15165), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n14674) );
  NAND2_X1 U16607 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14673) );
  OAI211_X1 U16608 ( .C1(n14862), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14676) );
  INV_X1 U16609 ( .A(n14676), .ZN(n14677) );
  OAI21_X1 U16610 ( .B1(n14705), .B2(n14136), .A(n14677), .ZN(n14679) );
  INV_X1 U16611 ( .A(n14679), .ZN(n14681) );
  AOI21_X1 U16612 ( .B1(n14718), .B2(n14681), .A(n14704), .ZN(n15702) );
  INV_X1 U16613 ( .A(n15702), .ZN(n14721) );
  INV_X1 U16614 ( .A(n14799), .ZN(n14683) );
  AOI21_X1 U16615 ( .B1(n14683), .B2(n14719), .A(n14682), .ZN(n14684) );
  NOR2_X1 U16616 ( .A1(n14684), .A2(n14791), .ZN(n21212) );
  AOI22_X1 U16617 ( .A1(n21212), .A2(n19888), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15507), .ZN(n14685) );
  OAI21_X1 U16618 ( .B1(n14721), .B2(n15509), .A(n14685), .ZN(P1_U2859) );
  XNOR2_X1 U16619 ( .A(n14686), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15687) );
  NAND2_X1 U16620 ( .A1(n15687), .A2(n15161), .ZN(n14702) );
  AOI22_X1 U16621 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14690) );
  AOI22_X1 U16622 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U16623 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U16624 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14687) );
  NAND4_X1 U16625 ( .A1(n14690), .A2(n14689), .A3(n14688), .A4(n14687), .ZN(
        n14696) );
  AOI22_X1 U16626 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14694) );
  AOI22_X1 U16627 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U16628 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U16629 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14691) );
  NAND4_X1 U16630 ( .A1(n14694), .A2(n14693), .A3(n14692), .A4(n14691), .ZN(
        n14695) );
  NOR2_X1 U16631 ( .A1(n14696), .A2(n14695), .ZN(n14699) );
  NAND2_X1 U16632 ( .A1(n15165), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U16633 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14697) );
  OAI211_X1 U16634 ( .C1(n14862), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14700) );
  INV_X1 U16635 ( .A(n14700), .ZN(n14701) );
  NAND2_X1 U16636 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  OAI21_X1 U16637 ( .B1(n14704), .B2(n14703), .A(n14846), .ZN(n15398) );
  OAI222_X1 U16638 ( .A1(n15587), .A2(n15398), .B1(n15585), .B2(n15513), .C1(
        n19812), .C2(n15553), .ZN(P1_U2890) );
  INV_X1 U16639 ( .A(n14705), .ZN(n15700) );
  AOI21_X1 U16640 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21519), .ZN(n14707) );
  NAND2_X1 U16641 ( .A1(n21597), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14706) );
  OAI211_X1 U16642 ( .C1(n21600), .C2(n15700), .A(n14707), .B(n14706), .ZN(
        n14708) );
  AOI21_X1 U16643 ( .B1(n21212), .B2(n21605), .A(n14708), .ZN(n14712) );
  INV_X1 U16644 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21470) );
  NOR2_X1 U16645 ( .A1(n21461), .A2(n21470), .ZN(n15400) );
  NAND2_X1 U16646 ( .A1(n15400), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15367) );
  NOR2_X1 U16647 ( .A1(n21544), .A2(n15367), .ZN(n21486) );
  NAND3_X1 U16648 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(n21486), .ZN(n21494) );
  INV_X1 U16649 ( .A(n21494), .ZN(n15369) );
  NAND2_X1 U16650 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15369), .ZN(n15393) );
  NAND2_X1 U16651 ( .A1(n21544), .A2(n14709), .ZN(n21507) );
  INV_X1 U16652 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21207) );
  OAI21_X1 U16653 ( .B1(n21596), .B2(n21207), .A(n21494), .ZN(n14710) );
  NAND2_X1 U16654 ( .A1(n15393), .A2(n14710), .ZN(n14711) );
  OAI211_X1 U16655 ( .C1(n14721), .C2(n21602), .A(n14712), .B(n14711), .ZN(
        P1_U2827) );
  XOR2_X1 U16656 ( .A(n14714), .B(n14713), .Z(n21477) );
  INV_X1 U16657 ( .A(n21477), .ZN(n14801) );
  OAI222_X1 U16658 ( .A1(n14801), .A2(n15587), .B1(n19806), .B2(n15553), .C1(
        n15527), .C2(n15585), .ZN(P1_U2893) );
  OR2_X1 U16659 ( .A1(n14716), .A2(n14715), .ZN(n14717) );
  XNOR2_X1 U16660 ( .A(n14799), .B(n14719), .ZN(n21484) );
  AOI22_X1 U16661 ( .A1(n21484), .A2(n19888), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n15507), .ZN(n14720) );
  OAI21_X1 U16662 ( .B1(n21493), .B2(n15509), .A(n14720), .ZN(P1_U2860) );
  OAI222_X1 U16663 ( .A1(n15587), .A2(n14721), .B1(n15585), .B2(n15518), .C1(
        n19810), .C2(n15553), .ZN(P1_U2891) );
  XNOR2_X1 U16664 ( .A(n14723), .B(n14722), .ZN(n14741) );
  INV_X1 U16665 ( .A(n14724), .ZN(n14726) );
  NOR2_X1 U16666 ( .A1(n14726), .A2(n14725), .ZN(n14728) );
  XOR2_X1 U16667 ( .A(n14728), .B(n14727), .Z(n14739) );
  OAI21_X1 U16668 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14729), .A(
        n16975), .ZN(n18110) );
  OAI22_X1 U16669 ( .A1(n11177), .A2(n17018), .B1(n17042), .B2(n18110), .ZN(
        n14730) );
  AOI21_X1 U16670 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n16539), .A(n14730), .ZN(
        n14731) );
  OAI21_X1 U16671 ( .B1(n18105), .B2(n17038), .A(n14731), .ZN(n14732) );
  AOI21_X1 U16672 ( .B1(n14739), .B2(n17032), .A(n14732), .ZN(n14733) );
  OAI21_X1 U16673 ( .B1(n14741), .B2(n17024), .A(n14733), .ZN(P2_U3007) );
  NAND2_X1 U16674 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14734), .ZN(
        n18473) );
  NAND2_X1 U16675 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n16539), .ZN(n14735) );
  OAI221_X1 U16676 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18473), .C1(
        n18474), .C2(n18485), .A(n14735), .ZN(n14736) );
  AOI21_X1 U16677 ( .B1(n18101), .B2(n18466), .A(n14736), .ZN(n14737) );
  OAI21_X1 U16678 ( .B1(n16567), .B2(n18105), .A(n14737), .ZN(n14738) );
  AOI21_X1 U16679 ( .B1(n14739), .B2(n18501), .A(n14738), .ZN(n14740) );
  OAI21_X1 U16680 ( .B1(n14741), .B2(n18494), .A(n14740), .ZN(P2_U3039) );
  OAI222_X1 U16681 ( .A1(n21493), .A2(n15587), .B1(n19808), .B2(n15553), .C1(
        n15585), .C2(n15523), .ZN(P1_U2892) );
  NOR2_X1 U16682 ( .A1(n14743), .A2(n14744), .ZN(n14745) );
  OR2_X1 U16683 ( .A1(n14742), .A2(n14745), .ZN(n18269) );
  AOI22_X1 U16684 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14748) );
  AOI22_X1 U16685 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U16686 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14746) );
  NAND3_X1 U16687 ( .A1(n14748), .A2(n14747), .A3(n14746), .ZN(n14762) );
  NAND2_X1 U16688 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14750) );
  NAND2_X1 U16689 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14749) );
  OAI211_X1 U16690 ( .C1(n15874), .C2(n14751), .A(n14750), .B(n14749), .ZN(
        n14756) );
  INV_X1 U16691 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U16692 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14753) );
  NAND2_X1 U16693 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14752) );
  OAI211_X1 U16694 ( .C1(n12015), .C2(n14754), .A(n14753), .B(n14752), .ZN(
        n14755) );
  NOR2_X1 U16695 ( .A1(n14756), .A2(n14755), .ZN(n14760) );
  AOI22_X1 U16696 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14759) );
  NAND2_X1 U16697 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14758) );
  NAND2_X1 U16698 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14757) );
  NAND4_X1 U16699 ( .A1(n14760), .A2(n14759), .A3(n14758), .A4(n14757), .ZN(
        n14761) );
  NOR2_X1 U16700 ( .A1(n14762), .A2(n14761), .ZN(n14806) );
  OR2_X1 U16701 ( .A1(n14806), .A2(n14763), .ZN(n14765) );
  OR2_X1 U16702 ( .A1(n14765), .A2(n14764), .ZN(n14766) );
  AOI22_X1 U16703 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14770) );
  AOI22_X1 U16704 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14769) );
  AOI22_X1 U16705 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14768) );
  NAND3_X1 U16706 ( .A1(n14770), .A2(n14769), .A3(n14768), .ZN(n14784) );
  INV_X1 U16707 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14773) );
  NAND2_X1 U16708 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14772) );
  NAND2_X1 U16709 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14771) );
  OAI211_X1 U16710 ( .C1(n15874), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14778) );
  INV_X1 U16711 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U16712 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14775) );
  NAND2_X1 U16713 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14774) );
  OAI211_X1 U16714 ( .C1(n12015), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14777) );
  NOR2_X1 U16715 ( .A1(n14778), .A2(n14777), .ZN(n14782) );
  AOI22_X1 U16716 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14781) );
  NAND2_X1 U16717 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14780) );
  NAND2_X1 U16718 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14779) );
  NAND4_X1 U16719 ( .A1(n14782), .A2(n14781), .A3(n14780), .A4(n14779), .ZN(
        n14783) );
  OR2_X1 U16720 ( .A1(n14784), .A2(n14783), .ZN(n14785) );
  OR2_X1 U16721 ( .A1(n14786), .A2(n14785), .ZN(n14787) );
  AND2_X1 U16722 ( .A1(n14787), .A2(n14827), .ZN(n19347) );
  NAND2_X1 U16723 ( .A1(n19347), .A2(n16082), .ZN(n14789) );
  NAND2_X1 U16724 ( .A1(n16046), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14788) );
  OAI211_X1 U16725 ( .C1(n18269), .C2(n16046), .A(n14789), .B(n14788), .ZN(
        P2_U2867) );
  INV_X1 U16726 ( .A(n15398), .ZN(n15689) );
  OR2_X1 U16727 ( .A1(n14791), .A2(n14790), .ZN(n14792) );
  NAND2_X1 U16728 ( .A1(n15504), .A2(n14792), .ZN(n21227) );
  OAI22_X1 U16729 ( .A1(n21227), .A2(n15497), .B1(n15392), .B2(n19892), .ZN(
        n14793) );
  AOI21_X1 U16730 ( .B1(n15689), .B2(n19889), .A(n14793), .ZN(n14794) );
  INV_X1 U16731 ( .A(n14794), .ZN(P1_U2858) );
  INV_X1 U16732 ( .A(n14795), .ZN(n14797) );
  OAI21_X1 U16733 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14800) );
  NAND2_X1 U16734 ( .A1(n14800), .A2(n14799), .ZN(n21475) );
  INV_X1 U16735 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14802) );
  OAI222_X1 U16736 ( .A1(n21475), .A2(n15497), .B1(n14802), .B2(n19892), .C1(
        n14801), .C2(n15509), .ZN(P1_U2861) );
  AND2_X1 U16737 ( .A1(n11029), .A2(n14803), .ZN(n14804) );
  OR2_X1 U16738 ( .A1(n14804), .A2(n14743), .ZN(n16357) );
  AOI21_X1 U16739 ( .B1(n14806), .B2(n14805), .A(n14786), .ZN(n16196) );
  NAND2_X1 U16740 ( .A1(n16196), .A2(n16082), .ZN(n14808) );
  NAND2_X1 U16741 ( .A1(n16046), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14807) );
  OAI211_X1 U16742 ( .C1(n16357), .C2(n16046), .A(n14808), .B(n14807), .ZN(
        P2_U2868) );
  INV_X1 U16743 ( .A(n14827), .ZN(n14829) );
  AOI22_X1 U16744 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U16745 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16746 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14810) );
  NAND3_X1 U16747 ( .A1(n14812), .A2(n14811), .A3(n14810), .ZN(n14826) );
  NAND2_X1 U16748 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14814) );
  NAND2_X1 U16749 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14813) );
  OAI211_X1 U16750 ( .C1(n15874), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14820) );
  NAND2_X1 U16751 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14817) );
  NAND2_X1 U16752 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14816) );
  OAI211_X1 U16753 ( .C1(n12015), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        n14819) );
  NOR2_X1 U16754 ( .A1(n14820), .A2(n14819), .ZN(n14824) );
  AOI22_X1 U16755 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U16756 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14822) );
  NAND2_X1 U16757 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14821) );
  NAND4_X1 U16758 ( .A1(n14824), .A2(n14823), .A3(n14822), .A4(n14821), .ZN(
        n14825) );
  OR2_X1 U16759 ( .A1(n14826), .A2(n14825), .ZN(n14828) );
  INV_X1 U16760 ( .A(n15864), .ZN(n16106) );
  OAI21_X1 U16761 ( .B1(n14829), .B2(n14828), .A(n16106), .ZN(n16195) );
  NAND2_X1 U16762 ( .A1(n16046), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14836) );
  INV_X1 U16763 ( .A(n14742), .ZN(n14833) );
  INV_X1 U16764 ( .A(n14831), .ZN(n14832) );
  NAND2_X1 U16765 ( .A1(n14833), .A2(n14832), .ZN(n14834) );
  AND2_X1 U16766 ( .A1(n14830), .A2(n14834), .ZN(n18273) );
  NAND2_X1 U16767 ( .A1(n18273), .A2(n16112), .ZN(n14835) );
  OAI211_X1 U16768 ( .C1(n16195), .C2(n16115), .A(n14836), .B(n14835), .ZN(
        P2_U2866) );
  NAND2_X1 U16769 ( .A1(n16697), .A2(n21139), .ZN(n14837) );
  NAND2_X1 U16770 ( .A1(n20713), .A2(n14837), .ZN(n21138) );
  NOR2_X1 U16771 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20757) );
  INV_X1 U16772 ( .A(n20757), .ZN(n20730) );
  NOR2_X1 U16773 ( .A1(n21138), .A2(n20730), .ZN(n14845) );
  OR2_X1 U16774 ( .A1(n20085), .A2(n14838), .ZN(n16705) );
  INV_X1 U16775 ( .A(n14839), .ZN(n21127) );
  INV_X1 U16776 ( .A(n14840), .ZN(n14841) );
  NOR2_X2 U16777 ( .A1(n14841), .A2(n20029), .ZN(n20524) );
  AOI211_X1 U16778 ( .C1(n21127), .C2(n17133), .A(n20524), .B(n14842), .ZN(
        n14843) );
  OAI21_X1 U16779 ( .B1(n20029), .B2(n16705), .A(n14843), .ZN(n21141) );
  INV_X1 U16780 ( .A(n21141), .ZN(n21151) );
  NAND2_X1 U16781 ( .A1(n20082), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18566) );
  NOR2_X1 U16782 ( .A1(n20082), .A2(n17523), .ZN(n16703) );
  NAND2_X1 U16783 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n16703), .ZN(n14844) );
  OAI211_X1 U16784 ( .C1(n21188), .C2(n21151), .A(n18566), .B(n14844), .ZN(
        n20759) );
  INV_X1 U16785 ( .A(n20759), .ZN(n20762) );
  MUX2_X1 U16786 ( .A(n14845), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20762), .Z(P3_U3284) );
  XOR2_X1 U16787 ( .A(n14848), .B(n14847), .Z(n21501) );
  INV_X1 U16788 ( .A(n21501), .ZN(n14864) );
  AOI22_X1 U16789 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14852) );
  AOI22_X1 U16790 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14851) );
  AOI22_X1 U16791 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16792 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14849) );
  NAND4_X1 U16793 ( .A1(n14852), .A2(n14851), .A3(n14850), .A4(n14849), .ZN(
        n14858) );
  AOI22_X1 U16794 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14856) );
  AOI22_X1 U16795 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U16796 ( .A1(n15145), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16797 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14853) );
  NAND4_X1 U16798 ( .A1(n14856), .A2(n14855), .A3(n14854), .A4(n14853), .ZN(
        n14857) );
  NOR2_X1 U16799 ( .A1(n14858), .A2(n14857), .ZN(n14861) );
  NAND2_X1 U16800 ( .A1(n15165), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U16801 ( .A1(n15164), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14859) );
  OAI211_X1 U16802 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        n14863) );
  AOI21_X1 U16803 ( .B1(n14864), .B2(n15161), .A(n14863), .ZN(n15502) );
  NAND2_X2 U16804 ( .A1(n10970), .A2(n14865), .ZN(n15500) );
  INV_X1 U16805 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15675) );
  XNOR2_X1 U16806 ( .A(n14866), .B(n15675), .ZN(n21512) );
  NAND2_X1 U16807 ( .A1(n21512), .A2(n15161), .ZN(n14881) );
  AOI22_X1 U16808 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U16809 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U16810 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U16811 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14867) );
  NAND4_X1 U16812 ( .A1(n14870), .A2(n14869), .A3(n14868), .A4(n14867), .ZN(
        n14876) );
  AOI22_X1 U16813 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U16814 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14873) );
  AOI22_X1 U16815 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U16816 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14871) );
  NAND4_X1 U16817 ( .A1(n14874), .A2(n14873), .A3(n14872), .A4(n14871), .ZN(
        n14875) );
  NOR2_X1 U16818 ( .A1(n14876), .A2(n14875), .ZN(n14879) );
  AOI21_X1 U16819 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15675), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14877) );
  AOI21_X1 U16820 ( .B1(n15165), .B2(P1_EAX_REG_16__SCAN_IN), .A(n14877), .ZN(
        n14878) );
  OAI21_X1 U16821 ( .B1(n15158), .B2(n14879), .A(n14878), .ZN(n14880) );
  NAND2_X1 U16822 ( .A1(n14881), .A2(n14880), .ZN(n15491) );
  NOR2_X4 U16823 ( .A1(n15500), .A2(n15491), .ZN(n15492) );
  XOR2_X1 U16824 ( .A(n15383), .B(n14882), .Z(n19945) );
  AOI22_X1 U16825 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15005), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U16826 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n15000), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14885) );
  AOI22_X1 U16827 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10983), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U16828 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14883) );
  NAND4_X1 U16829 ( .A1(n14886), .A2(n14885), .A3(n14884), .A4(n14883), .ZN(
        n14892) );
  AOI22_X1 U16830 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16831 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10981), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14889) );
  AOI22_X1 U16832 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14888) );
  AOI22_X1 U16833 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n15095), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14887) );
  NAND4_X1 U16834 ( .A1(n14890), .A2(n14889), .A3(n14888), .A4(n14887), .ZN(
        n14891) );
  OR2_X1 U16835 ( .A1(n14892), .A2(n14891), .ZN(n14895) );
  INV_X1 U16836 ( .A(n15164), .ZN(n14893) );
  OAI22_X1 U16837 ( .A1(n15087), .A2(n14120), .B1(n14893), .B2(n15383), .ZN(
        n14894) );
  AOI21_X1 U16838 ( .B1(n15127), .B2(n14895), .A(n14894), .ZN(n14896) );
  OAI21_X1 U16839 ( .B1(n19945), .B2(n14136), .A(n14896), .ZN(n15378) );
  XNOR2_X1 U16840 ( .A(n14897), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21523) );
  NAND2_X1 U16841 ( .A1(n21523), .A2(n15161), .ZN(n14913) );
  AOI22_X1 U16842 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14901) );
  AOI22_X1 U16843 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U16844 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16845 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14898) );
  NAND4_X1 U16846 ( .A1(n14901), .A2(n14900), .A3(n14899), .A4(n14898), .ZN(
        n14907) );
  AOI22_X1 U16847 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U16848 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14904) );
  AOI22_X1 U16849 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14903) );
  AOI22_X1 U16850 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14902) );
  NAND4_X1 U16851 ( .A1(n14905), .A2(n14904), .A3(n14903), .A4(n14902), .ZN(
        n14906) );
  NOR2_X1 U16852 ( .A1(n14907), .A2(n14906), .ZN(n14910) );
  NAND2_X1 U16853 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14909) );
  NAND2_X1 U16854 ( .A1(n15165), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U16855 ( .C1(n15158), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n14911) );
  NAND2_X1 U16856 ( .A1(n14911), .A2(n14136), .ZN(n14912) );
  NAND2_X1 U16857 ( .A1(n14913), .A2(n14912), .ZN(n15482) );
  AOI22_X1 U16858 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U16859 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U16860 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U16861 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14914) );
  NAND4_X1 U16862 ( .A1(n14917), .A2(n14916), .A3(n14915), .A4(n14914), .ZN(
        n14923) );
  AOI22_X1 U16863 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U16864 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U16865 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14919) );
  AOI22_X1 U16866 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14918) );
  NAND4_X1 U16867 ( .A1(n14921), .A2(n14920), .A3(n14919), .A4(n14918), .ZN(
        n14922) );
  NOR2_X1 U16868 ( .A1(n14923), .A2(n14922), .ZN(n14927) );
  NAND2_X1 U16869 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14924) );
  OAI211_X1 U16870 ( .C1(n15087), .C2(n14322), .A(n14136), .B(n14924), .ZN(
        n14925) );
  INV_X1 U16871 ( .A(n14925), .ZN(n14926) );
  OAI21_X1 U16872 ( .B1(n15158), .B2(n14927), .A(n14926), .ZN(n14930) );
  OAI21_X1 U16873 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n14928), .A(
        n14944), .ZN(n21536) );
  OR2_X1 U16874 ( .A1(n14136), .A2(n21536), .ZN(n14929) );
  NAND2_X1 U16875 ( .A1(n14930), .A2(n14929), .ZN(n15473) );
  AOI22_X1 U16876 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14934) );
  AOI22_X1 U16877 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U16878 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U16879 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14931) );
  NAND4_X1 U16880 ( .A1(n14934), .A2(n14933), .A3(n14932), .A4(n14931), .ZN(
        n14940) );
  AOI22_X1 U16881 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14938) );
  AOI22_X1 U16882 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14937) );
  AOI22_X1 U16883 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14936) );
  AOI22_X1 U16884 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14935) );
  NAND4_X1 U16885 ( .A1(n14938), .A2(n14937), .A3(n14936), .A4(n14935), .ZN(
        n14939) );
  NOR2_X1 U16886 ( .A1(n14940), .A2(n14939), .ZN(n14943) );
  OAI21_X1 U16887 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15656), .A(n14136), 
        .ZN(n14941) );
  AOI21_X1 U16888 ( .B1(n15165), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14941), .ZN(
        n14942) );
  OAI21_X1 U16889 ( .B1(n15158), .B2(n14943), .A(n14942), .ZN(n14946) );
  XNOR2_X1 U16890 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n14944), .ZN(
        n15658) );
  NAND2_X1 U16891 ( .A1(n15161), .A2(n15658), .ZN(n14945) );
  AOI22_X1 U16892 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16893 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14949) );
  AOI22_X1 U16894 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14948) );
  AOI22_X1 U16895 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14947) );
  NAND4_X1 U16896 ( .A1(n14950), .A2(n14949), .A3(n14948), .A4(n14947), .ZN(
        n14956) );
  AOI22_X1 U16897 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14954) );
  AOI22_X1 U16898 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U16899 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U16900 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14951) );
  NAND4_X1 U16901 ( .A1(n14954), .A2(n14953), .A3(n14952), .A4(n14951), .ZN(
        n14955) );
  NOR2_X1 U16902 ( .A1(n14956), .A2(n14955), .ZN(n14960) );
  NAND2_X1 U16903 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14957) );
  OAI211_X1 U16904 ( .C1(n15087), .C2(n14320), .A(n14136), .B(n14957), .ZN(
        n14958) );
  INV_X1 U16905 ( .A(n14958), .ZN(n14959) );
  OAI21_X1 U16906 ( .B1(n15158), .B2(n14960), .A(n14959), .ZN(n14963) );
  OAI21_X1 U16907 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n14961), .A(
        n14977), .ZN(n21552) );
  OR2_X1 U16908 ( .A1(n21552), .A2(n14136), .ZN(n14962) );
  NAND2_X1 U16909 ( .A1(n14963), .A2(n14962), .ZN(n15462) );
  AOI22_X1 U16910 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16911 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U16912 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U16913 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14964) );
  NAND4_X1 U16914 ( .A1(n14967), .A2(n14966), .A3(n14965), .A4(n14964), .ZN(
        n14973) );
  AOI22_X1 U16915 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14971) );
  AOI22_X1 U16916 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U16917 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U16918 ( .A1(n15145), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14968) );
  NAND4_X1 U16919 ( .A1(n14971), .A2(n14970), .A3(n14969), .A4(n14968), .ZN(
        n14972) );
  NOR2_X1 U16920 ( .A1(n14973), .A2(n14972), .ZN(n14976) );
  INV_X1 U16921 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15649) );
  AOI21_X1 U16922 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15649), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14974) );
  AOI21_X1 U16923 ( .B1(n15165), .B2(P1_EAX_REG_22__SCAN_IN), .A(n14974), .ZN(
        n14975) );
  OAI21_X1 U16924 ( .B1(n15158), .B2(n14976), .A(n14975), .ZN(n14979) );
  XNOR2_X1 U16925 ( .A(n14977), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21558) );
  NAND2_X1 U16926 ( .A1(n21558), .A2(n15161), .ZN(n14978) );
  AOI22_X1 U16927 ( .A1(n15144), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14983) );
  AOI22_X1 U16928 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10966), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U16929 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10963), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14981) );
  AOI22_X1 U16930 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n15005), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14980) );
  NAND4_X1 U16931 ( .A1(n14983), .A2(n14982), .A3(n14981), .A4(n14980), .ZN(
        n14989) );
  AOI22_X1 U16932 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U16933 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15139), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U16934 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14985) );
  AOI22_X1 U16935 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n15095), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14984) );
  NAND4_X1 U16936 ( .A1(n14987), .A2(n14986), .A3(n14985), .A4(n14984), .ZN(
        n14988) );
  NOR2_X1 U16937 ( .A1(n14989), .A2(n14988), .ZN(n15032) );
  AOI22_X1 U16938 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U16939 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16940 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U16941 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14990) );
  NAND4_X1 U16942 ( .A1(n14993), .A2(n14992), .A3(n14991), .A4(n14990), .ZN(
        n14999) );
  AOI22_X1 U16943 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14997) );
  AOI22_X1 U16944 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U16945 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U16946 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14994) );
  NAND4_X1 U16947 ( .A1(n14997), .A2(n14996), .A3(n14995), .A4(n14994), .ZN(
        n14998) );
  OR2_X1 U16948 ( .A1(n14999), .A2(n14998), .ZN(n15039) );
  AOI22_X1 U16949 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15004) );
  AOI22_X1 U16950 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U16951 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U16952 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15001) );
  NAND4_X1 U16953 ( .A1(n15004), .A2(n15003), .A3(n15002), .A4(n15001), .ZN(
        n15011) );
  AOI22_X1 U16954 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U16955 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16956 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U16957 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15006) );
  NAND4_X1 U16958 ( .A1(n15009), .A2(n15008), .A3(n15007), .A4(n15006), .ZN(
        n15010) );
  OR2_X1 U16959 ( .A1(n15011), .A2(n15010), .ZN(n15040) );
  NAND2_X1 U16960 ( .A1(n15039), .A2(n15040), .ZN(n15031) );
  NOR2_X1 U16961 ( .A1(n15032), .A2(n15031), .ZN(n15064) );
  AOI22_X1 U16962 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15015) );
  AOI22_X1 U16963 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15014) );
  AOI22_X1 U16964 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15013) );
  AOI22_X1 U16965 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15012) );
  NAND4_X1 U16966 ( .A1(n15015), .A2(n15014), .A3(n15013), .A4(n15012), .ZN(
        n15021) );
  AOI22_X1 U16967 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15019) );
  AOI22_X1 U16968 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15018) );
  AOI22_X1 U16969 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15017) );
  AOI22_X1 U16970 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15016) );
  NAND4_X1 U16971 ( .A1(n15019), .A2(n15018), .A3(n15017), .A4(n15016), .ZN(
        n15020) );
  OR2_X1 U16972 ( .A1(n15021), .A2(n15020), .ZN(n15063) );
  INV_X1 U16973 ( .A(n15063), .ZN(n15022) );
  XNOR2_X1 U16974 ( .A(n15064), .B(n15022), .ZN(n15025) );
  NAND2_X1 U16975 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15023) );
  OAI211_X1 U16976 ( .C1(n15087), .C2(n14314), .A(n14136), .B(n15023), .ZN(
        n15024) );
  AOI21_X1 U16977 ( .B1(n15025), .B2(n15127), .A(n15024), .ZN(n15030) );
  NAND2_X1 U16978 ( .A1(n15027), .A2(n15026), .ZN(n15028) );
  NAND2_X1 U16979 ( .A1(n15069), .A2(n15028), .ZN(n21601) );
  NOR2_X1 U16980 ( .A1(n21601), .A2(n14136), .ZN(n15029) );
  INV_X1 U16981 ( .A(n15434), .ZN(n15051) );
  XOR2_X1 U16982 ( .A(n15032), .B(n15031), .Z(n15033) );
  NAND2_X1 U16983 ( .A1(n15033), .A2(n15127), .ZN(n15038) );
  NAND2_X1 U16984 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15034) );
  OAI211_X1 U16985 ( .C1(n15087), .C2(n14306), .A(n14136), .B(n15034), .ZN(
        n15035) );
  INV_X1 U16986 ( .A(n15035), .ZN(n15037) );
  XNOR2_X1 U16987 ( .A(n15048), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n21587) );
  AND2_X1 U16988 ( .A1(n21587), .A2(n15161), .ZN(n15036) );
  AOI21_X1 U16989 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15442) );
  XNOR2_X1 U16990 ( .A(n15040), .B(n15039), .ZN(n15044) );
  NAND2_X1 U16991 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15041) );
  OAI211_X1 U16992 ( .C1(n15087), .C2(n14297), .A(n14136), .B(n15041), .ZN(
        n15042) );
  INV_X1 U16993 ( .A(n15042), .ZN(n15043) );
  OAI21_X1 U16994 ( .B1(n15158), .B2(n15044), .A(n15043), .ZN(n15050) );
  INV_X1 U16995 ( .A(n15045), .ZN(n15046) );
  INV_X1 U16996 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15642) );
  NAND2_X1 U16997 ( .A1(n15046), .A2(n15642), .ZN(n15047) );
  AND2_X1 U16998 ( .A1(n15048), .A2(n15047), .ZN(n21571) );
  NAND2_X1 U16999 ( .A1(n21571), .A2(n15161), .ZN(n15049) );
  AOI22_X1 U17000 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15056) );
  AOI22_X1 U17001 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15055) );
  AOI22_X1 U17002 ( .A1(n15139), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15054) );
  AOI22_X1 U17003 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15053) );
  NAND4_X1 U17004 ( .A1(n15056), .A2(n15055), .A3(n15054), .A4(n15053), .ZN(
        n15062) );
  AOI22_X1 U17005 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15060) );
  AOI22_X1 U17006 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U17007 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U17008 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15057) );
  NAND4_X1 U17009 ( .A1(n15060), .A2(n15059), .A3(n15058), .A4(n15057), .ZN(
        n15061) );
  NOR2_X1 U17010 ( .A1(n15062), .A2(n15061), .ZN(n15073) );
  NAND2_X1 U17011 ( .A1(n15064), .A2(n15063), .ZN(n15072) );
  XOR2_X1 U17012 ( .A(n15073), .B(n15072), .Z(n15067) );
  NAND2_X1 U17013 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15065) );
  OAI211_X1 U17014 ( .C1(n15087), .C2(n14318), .A(n14136), .B(n15065), .ZN(
        n15066) );
  AOI21_X1 U17015 ( .B1(n15067), .B2(n15127), .A(n15066), .ZN(n15068) );
  INV_X1 U17016 ( .A(n15068), .ZN(n15071) );
  XNOR2_X1 U17017 ( .A(n15069), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15620) );
  NAND2_X1 U17018 ( .A1(n15620), .A2(n15161), .ZN(n15070) );
  NAND2_X1 U17019 ( .A1(n15071), .A2(n15070), .ZN(n15353) );
  NOR2_X1 U17020 ( .A1(n15073), .A2(n15072), .ZN(n15108) );
  AOI22_X1 U17021 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10966), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15077) );
  AOI22_X1 U17022 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U17023 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U17024 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15074) );
  NAND4_X1 U17025 ( .A1(n15077), .A2(n15076), .A3(n15075), .A4(n15074), .ZN(
        n15083) );
  AOI22_X1 U17026 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15081) );
  AOI22_X1 U17027 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15080) );
  AOI22_X1 U17028 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U17029 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15078) );
  NAND4_X1 U17030 ( .A1(n15081), .A2(n15080), .A3(n15079), .A4(n15078), .ZN(
        n15082) );
  OR2_X1 U17031 ( .A1(n15083), .A2(n15082), .ZN(n15107) );
  INV_X1 U17032 ( .A(n15107), .ZN(n15084) );
  XNOR2_X1 U17033 ( .A(n15108), .B(n15084), .ZN(n15085) );
  NAND2_X1 U17034 ( .A1(n15085), .A2(n15127), .ZN(n15094) );
  NAND2_X1 U17035 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15086) );
  OAI211_X1 U17036 ( .C1(n15087), .C2(n14310), .A(n14136), .B(n15086), .ZN(
        n15088) );
  INV_X1 U17037 ( .A(n15088), .ZN(n15093) );
  NAND2_X1 U17038 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  NAND2_X1 U17039 ( .A1(n15111), .A2(n15091), .ZN(n15615) );
  NOR2_X1 U17040 ( .A1(n15615), .A2(n14136), .ZN(n15092) );
  AOI21_X1 U17041 ( .B1(n15094), .B2(n15093), .A(n15092), .ZN(n15340) );
  AOI22_X1 U17042 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U17043 ( .A1(n10981), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15098) );
  AOI22_X1 U17044 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15147), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U17045 ( .A1(n15095), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13046), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15096) );
  NAND4_X1 U17046 ( .A1(n15099), .A2(n15098), .A3(n15097), .A4(n15096), .ZN(
        n15106) );
  AOI22_X1 U17047 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15104) );
  AOI22_X1 U17048 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10963), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15103) );
  AOI22_X1 U17049 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U17050 ( .A1(n10966), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15101) );
  NAND4_X1 U17051 ( .A1(n15104), .A2(n15103), .A3(n15102), .A4(n15101), .ZN(
        n15105) );
  NOR2_X1 U17052 ( .A1(n15106), .A2(n15105), .ZN(n15116) );
  NAND2_X1 U17053 ( .A1(n15108), .A2(n15107), .ZN(n15115) );
  XOR2_X1 U17054 ( .A(n15116), .B(n15115), .Z(n15109) );
  NAND2_X1 U17055 ( .A1(n15109), .A2(n15127), .ZN(n15114) );
  INV_X1 U17056 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15606) );
  AOI21_X1 U17057 ( .B1(n15606), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15110) );
  AOI21_X1 U17058 ( .B1(n15165), .B2(P1_EAX_REG_28__SCAN_IN), .A(n15110), .ZN(
        n15113) );
  XNOR2_X1 U17059 ( .A(n15111), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15610) );
  AOI21_X1 U17060 ( .B1(n15114), .B2(n15113), .A(n15112), .ZN(n15328) );
  NOR2_X1 U17061 ( .A1(n15116), .A2(n15115), .ZN(n15129) );
  AOI22_X1 U17062 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U17063 ( .A1(n13007), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U17064 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U17065 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12946), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15117) );
  NAND4_X1 U17066 ( .A1(n15120), .A2(n15119), .A3(n15118), .A4(n15117), .ZN(
        n15126) );
  AOI22_X1 U17067 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12901), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U17068 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15123) );
  AOI22_X1 U17069 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15122) );
  AOI22_X1 U17070 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12951), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15121) );
  NAND4_X1 U17071 ( .A1(n15124), .A2(n15123), .A3(n15122), .A4(n15121), .ZN(
        n15125) );
  OR2_X1 U17072 ( .A1(n15126), .A2(n15125), .ZN(n15128) );
  NAND2_X1 U17073 ( .A1(n15129), .A2(n15128), .ZN(n15155) );
  OAI211_X1 U17074 ( .C1(n15129), .C2(n15128), .A(n15155), .B(n15127), .ZN(
        n15132) );
  NAND2_X1 U17075 ( .A1(n15165), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n15131) );
  NAND2_X1 U17076 ( .A1(n21898), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15130) );
  NAND4_X1 U17077 ( .A1(n15132), .A2(n14136), .A3(n15131), .A4(n15130), .ZN(
        n15137) );
  NAND2_X1 U17078 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  NAND2_X1 U17079 ( .A1(n15160), .A2(n15135), .ZN(n15595) );
  NAND2_X1 U17080 ( .A1(n15137), .A2(n15136), .ZN(n15315) );
  AOI22_X1 U17081 ( .A1(n15000), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12941), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15143) );
  AOI22_X1 U17082 ( .A1(n10983), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U17083 ( .A1(n10963), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15138), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U17084 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15139), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15140) );
  NAND4_X1 U17085 ( .A1(n15143), .A2(n15142), .A3(n15141), .A4(n15140), .ZN(
        n15153) );
  AOI22_X1 U17086 ( .A1(n15100), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15144), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U17087 ( .A1(n15005), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15145), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U17088 ( .A1(n13046), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15146), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U17089 ( .A1(n15147), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15095), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15148) );
  NAND4_X1 U17090 ( .A1(n15151), .A2(n15150), .A3(n15149), .A4(n15148), .ZN(
        n15152) );
  NOR2_X1 U17091 ( .A1(n15153), .A2(n15152), .ZN(n15154) );
  XNOR2_X1 U17092 ( .A(n15155), .B(n15154), .ZN(n15159) );
  AOI21_X1 U17093 ( .B1(n15260), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n15156) );
  AOI21_X1 U17094 ( .B1(n15165), .B2(P1_EAX_REG_30__SCAN_IN), .A(n15156), .ZN(
        n15157) );
  OAI21_X1 U17095 ( .B1(n15159), .B2(n15158), .A(n15157), .ZN(n15163) );
  XNOR2_X1 U17096 ( .A(n15160), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15308) );
  NAND2_X1 U17097 ( .A1(n15308), .A2(n15161), .ZN(n15162) );
  NAND2_X1 U17098 ( .A1(n15163), .A2(n15162), .ZN(n15257) );
  AOI22_X1 U17099 ( .A1(n15165), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15164), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15166) );
  AOI21_X1 U17100 ( .B1(n19955), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15167), .ZN(n15168) );
  OAI21_X1 U17101 ( .B1(n19964), .B2(n15169), .A(n15168), .ZN(n15170) );
  AOI21_X1 U17102 ( .B1(n15295), .B2(n19952), .A(n15170), .ZN(n15171) );
  OAI21_X1 U17103 ( .B1(n15172), .B2(n21610), .A(n15171), .ZN(P1_U2968) );
  OAI21_X1 U17104 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n21295) );
  AOI22_X1 U17105 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n15176) );
  OAI21_X1 U17106 ( .B1(n19964), .B2(n15177), .A(n15176), .ZN(n15178) );
  AOI21_X1 U17107 ( .B1(n15179), .B2(n19952), .A(n15178), .ZN(n15180) );
  OAI21_X1 U17108 ( .B1(n21295), .B2(n21610), .A(n15180), .ZN(P1_U2990) );
  OAI21_X1 U17109 ( .B1(n15183), .B2(n15182), .A(n15181), .ZN(n21282) );
  AOI22_X1 U17110 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U17111 ( .B1(n19964), .B2(n15185), .A(n15184), .ZN(n15186) );
  AOI21_X1 U17112 ( .B1(n15187), .B2(n19952), .A(n15186), .ZN(n15188) );
  OAI21_X1 U17113 ( .B1(n21282), .B2(n21610), .A(n15188), .ZN(P1_U2991) );
  INV_X1 U17114 ( .A(n15189), .ZN(n15191) );
  NAND2_X1 U17115 ( .A1(n15191), .A2(n15190), .ZN(n15192) );
  NAND2_X1 U17116 ( .A1(n15204), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15200) );
  XOR2_X1 U17117 ( .A(n15200), .B(n15201), .Z(n18355) );
  OAI21_X1 U17118 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16243), .ZN(n15193) );
  INV_X1 U17119 ( .A(n16243), .ZN(n15194) );
  INV_X1 U17120 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16474) );
  NAND2_X1 U17121 ( .A1(n15194), .A2(n16474), .ZN(n15195) );
  NAND2_X1 U17122 ( .A1(n15196), .A2(n15195), .ZN(n15199) );
  INV_X1 U17123 ( .A(n15197), .ZN(n15198) );
  AND2_X1 U17124 ( .A1(n15204), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15202) );
  XOR2_X1 U17125 ( .A(n15202), .B(n15203), .Z(n18365) );
  NAND2_X1 U17126 ( .A1(n18365), .A2(n11337), .ZN(n15207) );
  INV_X1 U17127 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16458) );
  NAND2_X1 U17128 ( .A1(n15207), .A2(n16458), .ZN(n16229) );
  NAND2_X1 U17129 ( .A1(n16231), .A2(n16229), .ZN(n16215) );
  NAND2_X1 U17130 ( .A1(n15204), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15205) );
  XNOR2_X1 U17131 ( .A(n15209), .B(n15205), .ZN(n18379) );
  AOI21_X1 U17132 ( .B1(n18379), .B2(n11337), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16218) );
  INV_X1 U17133 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16441) );
  NOR2_X1 U17134 ( .A1(n15212), .A2(n16441), .ZN(n15206) );
  NAND2_X1 U17135 ( .A1(n18379), .A2(n15206), .ZN(n16216) );
  INV_X1 U17136 ( .A(n15207), .ZN(n15208) );
  NAND2_X1 U17137 ( .A1(n15208), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16230) );
  OAI21_X2 U17138 ( .B1(n16215), .B2(n16218), .A(n11391), .ZN(n15215) );
  INV_X1 U17139 ( .A(n15210), .ZN(n15211) );
  NOR2_X1 U17140 ( .A1(n18395), .A2(n15212), .ZN(n15213) );
  XOR2_X1 U17141 ( .A(n15213), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n15214) );
  XNOR2_X1 U17142 ( .A(n15215), .B(n15214), .ZN(n15280) );
  NAND2_X1 U17143 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15271) );
  INV_X1 U17144 ( .A(n15279), .ZN(n15235) );
  INV_X1 U17145 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16249) );
  NAND2_X1 U17146 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15218) );
  AOI22_X1 U17147 ( .A1(n15224), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n15217) );
  OAI211_X1 U17148 ( .C1(n15227), .C2(n16249), .A(n15218), .B(n15217), .ZN(
        n16064) );
  INV_X1 U17149 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17123) );
  NAND2_X1 U17150 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15220) );
  AOI22_X1 U17151 ( .A1(n15224), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n15219) );
  OAI211_X1 U17152 ( .C1(n15227), .C2(n17123), .A(n15220), .B(n15219), .ZN(
        n16056) );
  INV_X1 U17153 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n16222) );
  NAND2_X1 U17154 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15222) );
  AOI22_X1 U17155 ( .A1(n15224), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n15221) );
  OAI211_X1 U17156 ( .C1(n15227), .C2(n16222), .A(n15222), .B(n15221), .ZN(
        n16047) );
  NAND2_X1 U17157 ( .A1(n16058), .A2(n16047), .ZN(n15229) );
  INV_X1 U17158 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18397) );
  NAND2_X1 U17159 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15226) );
  AOI22_X1 U17160 ( .A1(n15224), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n15225) );
  OAI211_X1 U17161 ( .C1(n15227), .C2(n18397), .A(n15226), .B(n15225), .ZN(
        n15228) );
  INV_X1 U17162 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18163) );
  INV_X1 U17163 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18140) );
  INV_X1 U17164 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16403) );
  INV_X1 U17165 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16359) );
  INV_X1 U17166 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16334) );
  INV_X1 U17167 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18295) );
  INV_X1 U17168 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16286) );
  INV_X1 U17169 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16272) );
  INV_X1 U17170 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16235) );
  NOR2_X1 U17171 ( .A1(n18475), .A2(n18397), .ZN(n15273) );
  AOI21_X1 U17172 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15273), .ZN(n15230) );
  OAI21_X1 U17173 ( .B1(n15811), .B2(n17042), .A(n15230), .ZN(n15231) );
  INV_X1 U17174 ( .A(n15231), .ZN(n15232) );
  NAND2_X1 U17175 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  AOI21_X1 U17176 ( .B1(n15235), .B2(n17035), .A(n15234), .ZN(n15236) );
  OAI21_X1 U17177 ( .B1(n15280), .B2(n17014), .A(n15236), .ZN(P2_U2983) );
  NOR2_X1 U17178 ( .A1(n15239), .A2(n12967), .ZN(n15238) );
  NAND2_X1 U17179 ( .A1(n15238), .A2(n15237), .ZN(n15510) );
  INV_X1 U17180 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n22201) );
  NAND3_X1 U17181 ( .A1(n15295), .A2(n22202), .A3(n15553), .ZN(n15241) );
  AOI22_X1 U17182 ( .A1(n15581), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15239), .ZN(n15240) );
  OAI211_X1 U17183 ( .C1(n15510), .C2(n22201), .A(n15241), .B(n15240), .ZN(
        P1_U2873) );
  NAND2_X1 U17184 ( .A1(n15724), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15242) );
  OAI21_X1 U17185 ( .B1(n15612), .B2(n11387), .A(n15243), .ZN(n15245) );
  XNOR2_X1 U17186 ( .A(n15246), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15263) );
  INV_X1 U17187 ( .A(n15247), .ZN(n15248) );
  OAI22_X1 U17188 ( .A1(n15318), .A2(n13342), .B1(n15248), .B2(n15333), .ZN(
        n15250) );
  XNOR2_X1 U17189 ( .A(n15250), .B(n15249), .ZN(n15425) );
  NAND2_X1 U17190 ( .A1(n13790), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15258) );
  NAND3_X1 U17191 ( .A1(n15713), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15252), .ZN(n15251) );
  OAI211_X1 U17192 ( .C1(n15253), .C2(n15252), .A(n15258), .B(n15251), .ZN(
        n15254) );
  AOI21_X1 U17193 ( .B1(n15425), .B2(n21382), .A(n15254), .ZN(n15255) );
  OAI21_X1 U17194 ( .B1(n15263), .B2(n21353), .A(n15255), .ZN(P1_U3001) );
  NAND2_X1 U17195 ( .A1(n19946), .A2(n15308), .ZN(n15259) );
  OAI211_X1 U17196 ( .C1(n19923), .C2(n15260), .A(n15259), .B(n15258), .ZN(
        n15261) );
  AOI21_X1 U17197 ( .B1(n15304), .B2(n19952), .A(n15261), .ZN(n15262) );
  OAI21_X1 U17198 ( .B1(n15263), .B2(n21610), .A(n15262), .ZN(P1_U2969) );
  AOI22_X1 U17199 ( .A1(n12595), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15264) );
  OAI21_X1 U17200 ( .B1(n15269), .B2(n16249), .A(n15264), .ZN(n16133) );
  AOI22_X1 U17201 ( .A1(n12595), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15266) );
  OAI21_X1 U17202 ( .B1(n15269), .B2(n17123), .A(n15266), .ZN(n16126) );
  AOI22_X1 U17203 ( .A1(n12595), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15267) );
  OAI21_X1 U17204 ( .B1(n15269), .B2(n16222), .A(n15267), .ZN(n16116) );
  NAND2_X1 U17205 ( .A1(n11338), .A2(n16116), .ZN(n16119) );
  AOI22_X1 U17206 ( .A1(n12595), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12467), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15268) );
  OAI21_X1 U17207 ( .B1(n15269), .B2(n18397), .A(n15268), .ZN(n15270) );
  NOR2_X1 U17208 ( .A1(n15271), .A2(n15190), .ZN(n16439) );
  NAND2_X1 U17209 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16439), .ZN(
        n15272) );
  NOR3_X1 U17210 ( .A1(n16457), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15272), .ZN(n15277) );
  AOI21_X1 U17211 ( .B1(n15272), .B2(n18460), .A(n16455), .ZN(n16442) );
  OR2_X1 U17212 ( .A1(n16442), .A2(n15216), .ZN(n15275) );
  NAND2_X1 U17213 ( .A1(n15275), .A2(n15274), .ZN(n15276) );
  OAI21_X1 U17214 ( .B1(n15280), .B2(n18450), .A(n11010), .ZN(P2_U3015) );
  INV_X1 U17215 ( .A(n13325), .ZN(n15281) );
  OAI22_X1 U17216 ( .A1(n21623), .A2(n15281), .B1(n15288), .B2(n15287), .ZN(
        n15286) );
  NAND2_X1 U17217 ( .A1(n21623), .A2(n15282), .ZN(n15283) );
  OAI21_X1 U17218 ( .B1(n21623), .B2(n15284), .A(n15283), .ZN(n15285) );
  OR2_X1 U17219 ( .A1(n15286), .A2(n15285), .ZN(n16748) );
  INV_X1 U17220 ( .A(n21623), .ZN(n15292) );
  INV_X1 U17221 ( .A(n15287), .ZN(n15289) );
  AOI21_X1 U17222 ( .B1(n15289), .B2(n15288), .A(n13325), .ZN(n15290) );
  AOI21_X1 U17223 ( .B1(n15292), .B2(n15291), .A(n15290), .ZN(n19966) );
  OAI21_X1 U17224 ( .B1(n15294), .B2(n15293), .A(n21660), .ZN(n21194) );
  NAND2_X1 U17225 ( .A1(n19966), .A2(n21194), .ZN(n16752) );
  AND2_X1 U17226 ( .A1(n16752), .A2(n19965), .ZN(n21612) );
  MUX2_X1 U17227 ( .A(P1_MORE_REG_SCAN_IN), .B(n16748), .S(n21612), .Z(
        P1_U3484) );
  NAND2_X1 U17228 ( .A1(n15295), .A2(n21588), .ZN(n15303) );
  INV_X1 U17229 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16860) );
  INV_X1 U17230 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21595) );
  INV_X1 U17231 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21569) );
  NAND3_X1 U17232 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .ZN(n21495) );
  INV_X1 U17233 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15296) );
  INV_X1 U17234 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n19832) );
  NOR3_X1 U17235 ( .A1(n21495), .A2(n15296), .A3(n19832), .ZN(n15370) );
  INV_X1 U17236 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21537) );
  INV_X1 U17237 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21535) );
  NOR3_X1 U17238 ( .A1(n15655), .A2(n21537), .A3(n21535), .ZN(n21563) );
  NAND4_X1 U17239 ( .A1(n15370), .A2(n21563), .A3(P1_REIP_REG_11__SCAN_IN), 
        .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n15366) );
  NOR2_X1 U17240 ( .A1(n15366), .A2(n15367), .ZN(n21545) );
  NAND4_X1 U17241 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n21436), .A3(n21545), 
        .A4(P1_REIP_REG_22__SCAN_IN), .ZN(n21568) );
  NOR2_X1 U17242 ( .A1(n21569), .A2(n21568), .ZN(n21583) );
  NAND2_X1 U17243 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n21583), .ZN(n21594) );
  NOR2_X1 U17244 ( .A1(n21595), .A2(n21594), .ZN(n15356) );
  INV_X1 U17245 ( .A(n15356), .ZN(n21599) );
  NOR2_X1 U17246 ( .A1(n16860), .A2(n21599), .ZN(n15358) );
  NAND2_X1 U17247 ( .A1(n15351), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15338) );
  INV_X1 U17248 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n16933) );
  OR2_X1 U17249 ( .A1(n15338), .A2(n16933), .ZN(n15305) );
  INV_X1 U17250 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15297) );
  NOR2_X1 U17251 ( .A1(n15305), .A2(n15297), .ZN(n15298) );
  NOR2_X1 U17252 ( .A1(n15298), .A2(n21596), .ZN(n15306) );
  INV_X1 U17253 ( .A(n15298), .ZN(n15300) );
  AOI22_X1 U17254 ( .A1(n21597), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21553), .ZN(n15299) );
  OAI21_X1 U17255 ( .B1(n15300), .B2(P1_REIP_REG_31__SCAN_IN), .A(n15299), 
        .ZN(n15301) );
  AOI21_X1 U17256 ( .B1(n15306), .B2(P1_REIP_REG_31__SCAN_IN), .A(n15301), 
        .ZN(n15302) );
  OAI211_X1 U17257 ( .C1(n15424), .C2(n21592), .A(n15303), .B(n15302), .ZN(
        P1_U2809) );
  INV_X1 U17258 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15311) );
  INV_X1 U17259 ( .A(n15305), .ZN(n15307) );
  OAI21_X1 U17260 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n15307), .A(n15306), 
        .ZN(n15310) );
  AOI22_X1 U17261 ( .A1(n15308), .A2(n21586), .B1(n21553), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15309) );
  OAI211_X1 U17262 ( .C1(n21580), .C2(n15311), .A(n15310), .B(n15309), .ZN(
        n15312) );
  AOI21_X1 U17263 ( .B1(n15425), .B2(n21605), .A(n15312), .ZN(n15313) );
  OAI21_X1 U17264 ( .B1(n15517), .B2(n21602), .A(n15313), .ZN(P1_U2810) );
  NAND2_X1 U17265 ( .A1(n15314), .A2(n15315), .ZN(n15316) );
  AOI21_X1 U17266 ( .B1(n15319), .B2(n15333), .A(n15318), .ZN(n15719) );
  INV_X1 U17267 ( .A(n15595), .ZN(n15320) );
  AOI22_X1 U17268 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21553), .B1(
        n21586), .B2(n15320), .ZN(n15321) );
  OAI21_X1 U17269 ( .B1(n21580), .B2(n15322), .A(n15321), .ZN(n15325) );
  NAND3_X1 U17270 ( .A1(n15338), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n21507), 
        .ZN(n15323) );
  OAI21_X1 U17271 ( .B1(n15338), .B2(P1_REIP_REG_29__SCAN_IN), .A(n15323), 
        .ZN(n15324) );
  AOI211_X1 U17272 ( .C1(n15719), .C2(n21605), .A(n15325), .B(n15324), .ZN(
        n15326) );
  OAI21_X1 U17273 ( .B1(n15522), .B2(n21602), .A(n15326), .ZN(P1_U2811) );
  INV_X1 U17274 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15330) );
  INV_X1 U17275 ( .A(n15351), .ZN(n15329) );
  OAI21_X1 U17276 ( .B1(n21596), .B2(n15330), .A(n15329), .ZN(n15337) );
  OR2_X1 U17277 ( .A1(n15344), .A2(n15331), .ZN(n15332) );
  NAND2_X1 U17278 ( .A1(n15333), .A2(n15332), .ZN(n15722) );
  AOI22_X1 U17279 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n21553), .B1(
        n21586), .B2(n15610), .ZN(n15335) );
  NAND2_X1 U17280 ( .A1(n21597), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n15334) );
  OAI211_X1 U17281 ( .C1(n15722), .C2(n21592), .A(n15335), .B(n15334), .ZN(
        n15336) );
  AOI21_X1 U17282 ( .B1(n15338), .B2(n15337), .A(n15336), .ZN(n15339) );
  OAI21_X1 U17283 ( .B1(n15607), .B2(n21602), .A(n15339), .ZN(P1_U2812) );
  AOI21_X1 U17284 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n21507), .A(n15358), 
        .ZN(n15350) );
  INV_X1 U17285 ( .A(n15340), .ZN(n15343) );
  INV_X1 U17286 ( .A(n15341), .ZN(n15342) );
  AOI21_X1 U17287 ( .B1(n15343), .B2(n15342), .A(n15327), .ZN(n15617) );
  NAND2_X1 U17288 ( .A1(n15617), .A2(n21588), .ZN(n15349) );
  OAI22_X1 U17289 ( .A1(n15089), .A2(n21609), .B1(n21600), .B2(n15615), .ZN(
        n15347) );
  AOI21_X1 U17290 ( .B1(n15345), .B2(n15354), .A(n15344), .ZN(n15740) );
  INV_X1 U17291 ( .A(n15740), .ZN(n15429) );
  NOR2_X1 U17292 ( .A1(n15429), .A2(n21592), .ZN(n15346) );
  AOI211_X1 U17293 ( .C1(n21597), .C2(P1_EBX_REG_27__SCAN_IN), .A(n15347), .B(
        n15346), .ZN(n15348) );
  OAI211_X1 U17294 ( .C1(n15351), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        P1_U2813) );
  AOI21_X1 U17295 ( .B1(n15353), .B2(n15436), .A(n15341), .ZN(n15624) );
  INV_X1 U17296 ( .A(n15624), .ZN(n15536) );
  AOI21_X1 U17297 ( .B1(n15355), .B2(n15437), .A(n11202), .ZN(n15749) );
  AOI21_X1 U17298 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n21507), .A(n15356), 
        .ZN(n15357) );
  NOR2_X1 U17299 ( .A1(n15358), .A2(n15357), .ZN(n15362) );
  AOI22_X1 U17300 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21553), .B1(
        n21586), .B2(n15620), .ZN(n15359) );
  OAI21_X1 U17301 ( .B1(n21580), .B2(n15360), .A(n15359), .ZN(n15361) );
  AOI211_X1 U17302 ( .C1(n15749), .C2(n21605), .A(n15362), .B(n15361), .ZN(
        n15363) );
  OAI21_X1 U17303 ( .B1(n15536), .B2(n21602), .A(n15363), .ZN(P1_U2814) );
  OAI21_X1 U17304 ( .B1(n15364), .B2(n11385), .A(n15461), .ZN(n15661) );
  INV_X1 U17305 ( .A(n15366), .ZN(n15368) );
  NOR2_X1 U17306 ( .A1(n21435), .A2(n15367), .ZN(n21485) );
  AOI21_X1 U17307 ( .B1(n15368), .B2(n21485), .A(n21596), .ZN(n21559) );
  AND2_X1 U17308 ( .A1(n15370), .A2(n15369), .ZN(n21562) );
  NAND2_X1 U17309 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n21562), .ZN(n21531) );
  OAI21_X1 U17310 ( .B1(n21537), .B2(n21531), .A(n15655), .ZN(n15376) );
  AOI22_X1 U17311 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21553), .B1(
        n21586), .B2(n15658), .ZN(n15371) );
  OAI21_X1 U17312 ( .B1(n21580), .B2(n15469), .A(n15371), .ZN(n15375) );
  NOR2_X1 U17313 ( .A1(n15477), .A2(n15372), .ZN(n15373) );
  OR2_X1 U17314 ( .A1(n15463), .A2(n15373), .ZN(n21372) );
  NOR2_X1 U17315 ( .A1(n21372), .A2(n21592), .ZN(n15374) );
  AOI211_X1 U17316 ( .C1(n21559), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        n15377) );
  OAI21_X1 U17317 ( .B1(n15661), .B2(n21602), .A(n15377), .ZN(P1_U2820) );
  INV_X1 U17318 ( .A(n15378), .ZN(n15381) );
  INV_X1 U17319 ( .A(n15492), .ZN(n15380) );
  AOI21_X1 U17320 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n19947) );
  AOI22_X1 U17321 ( .A1(n21597), .A2(P1_EBX_REG_17__SCAN_IN), .B1(n21586), 
        .B2(n19945), .ZN(n15382) );
  OAI21_X1 U17322 ( .B1(n15383), .B2(n21609), .A(n15382), .ZN(n15388) );
  INV_X1 U17323 ( .A(n15484), .ZN(n15384) );
  AOI21_X1 U17324 ( .B1(n15385), .B2(n11189), .A(n15384), .ZN(n21348) );
  INV_X1 U17325 ( .A(n21348), .ZN(n15490) );
  NOR3_X1 U17326 ( .A1(n21495), .A2(n19832), .A3(n21494), .ZN(n21510) );
  NOR2_X1 U17327 ( .A1(n21596), .A2(n21562), .ZN(n21534) );
  OAI21_X1 U17328 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21510), .A(n21534), 
        .ZN(n15386) );
  OAI211_X1 U17329 ( .C1(n21592), .C2(n15490), .A(n15386), .B(n21529), .ZN(
        n15387) );
  AOI211_X1 U17330 ( .C1(n19947), .C2(n21588), .A(n15388), .B(n15387), .ZN(
        n15389) );
  INV_X1 U17331 ( .A(n15389), .ZN(P1_U2823) );
  INV_X1 U17332 ( .A(n21227), .ZN(n15396) );
  NOR2_X1 U17333 ( .A1(n21600), .A2(n15687), .ZN(n15390) );
  AOI211_X1 U17334 ( .C1(n21553), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21519), .B(n15390), .ZN(n15391) );
  OAI21_X1 U17335 ( .B1(n15392), .B2(n21580), .A(n15391), .ZN(n15395) );
  INV_X1 U17336 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21218) );
  NOR2_X1 U17337 ( .A1(n21218), .A2(n15393), .ZN(n21496) );
  AOI211_X1 U17338 ( .C1(n21218), .C2(n15393), .A(n21496), .B(n21596), .ZN(
        n15394) );
  AOI211_X1 U17339 ( .C1(n15396), .C2(n21605), .A(n15395), .B(n15394), .ZN(
        n15397) );
  OAI21_X1 U17340 ( .B1(n15398), .B2(n21602), .A(n15397), .ZN(P1_U2826) );
  NOR2_X1 U17341 ( .A1(n21596), .A2(n21485), .ZN(n21473) );
  AOI21_X1 U17342 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21519), .ZN(n15399) );
  OAI21_X1 U17343 ( .B1(n15708), .B2(n21600), .A(n15399), .ZN(n15404) );
  NAND2_X1 U17344 ( .A1(n21436), .A2(n15400), .ZN(n15402) );
  AOI22_X1 U17345 ( .A1(n21305), .A2(n21605), .B1(n21597), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15401) );
  OAI21_X1 U17346 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15402), .A(n15401), 
        .ZN(n15403) );
  AOI211_X1 U17347 ( .C1(n21473), .C2(P1_REIP_REG_10__SCAN_IN), .A(n15404), 
        .B(n15403), .ZN(n15405) );
  OAI21_X1 U17348 ( .B1(n15706), .B2(n21602), .A(n15405), .ZN(P1_U2830) );
  INV_X1 U17349 ( .A(n21805), .ZN(n21884) );
  MUX2_X1 U17350 ( .A(n21586), .B(n21553), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15406) );
  AOI21_X1 U17351 ( .B1(n21597), .B2(P1_EBX_REG_1__SCAN_IN), .A(n15406), .ZN(
        n15409) );
  OAI21_X1 U17352 ( .B1(n21436), .B2(P1_REIP_REG_1__SCAN_IN), .A(n15407), .ZN(
        n15408) );
  OAI211_X1 U17353 ( .C1(n15410), .C2(n21592), .A(n15409), .B(n15408), .ZN(
        n15411) );
  AOI21_X1 U17354 ( .B1(n21884), .B2(n21411), .A(n15411), .ZN(n15412) );
  OAI21_X1 U17355 ( .B1(n15414), .B2(n15413), .A(n15412), .ZN(P1_U2839) );
  INV_X1 U17356 ( .A(n15415), .ZN(n15416) );
  NAND2_X1 U17357 ( .A1(n15416), .A2(n21428), .ZN(n15422) );
  OR2_X1 U17358 ( .A1(n21553), .A2(n21586), .ZN(n15417) );
  AOI22_X1 U17359 ( .A1(n15417), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n21748), .B2(n21411), .ZN(n15421) );
  AOI22_X1 U17360 ( .A1(n21605), .A2(n15418), .B1(n21597), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n15420) );
  NAND2_X1 U17361 ( .A1(n21507), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15419) );
  NAND4_X1 U17362 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        P1_U2840) );
  INV_X1 U17363 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15423) );
  OAI22_X1 U17364 ( .A1(n15424), .A2(n15497), .B1(n19892), .B2(n15423), .ZN(
        P1_U2841) );
  AOI22_X1 U17365 ( .A1(n15425), .A2(n19888), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15507), .ZN(n15426) );
  OAI21_X1 U17366 ( .B1(n15517), .B2(n15509), .A(n15426), .ZN(P1_U2842) );
  AOI22_X1 U17367 ( .A1(n15719), .A2(n19888), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15507), .ZN(n15427) );
  OAI21_X1 U17368 ( .B1(n15522), .B2(n15509), .A(n15427), .ZN(P1_U2843) );
  INV_X1 U17369 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15428) );
  OAI222_X1 U17370 ( .A1(n15509), .A2(n15607), .B1(n15428), .B2(n19892), .C1(
        n15722), .C2(n15497), .ZN(P1_U2844) );
  INV_X1 U17371 ( .A(n15617), .ZN(n15531) );
  INV_X1 U17372 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15430) );
  OAI222_X1 U17373 ( .A1(n15509), .A2(n15531), .B1(n15430), .B2(n19892), .C1(
        n15429), .C2(n15497), .ZN(P1_U2845) );
  AOI22_X1 U17374 ( .A1(n15749), .A2(n19888), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n15507), .ZN(n15431) );
  OAI21_X1 U17375 ( .B1(n15536), .B2(n15509), .A(n15431), .ZN(P1_U2846) );
  NAND2_X1 U17376 ( .A1(n15432), .A2(n15433), .ZN(n15441) );
  NAND2_X1 U17377 ( .A1(n15441), .A2(n15434), .ZN(n15435) );
  NAND2_X1 U17378 ( .A1(n15436), .A2(n15435), .ZN(n21603) );
  INV_X1 U17379 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15440) );
  INV_X1 U17380 ( .A(n15445), .ZN(n15438) );
  AOI21_X1 U17381 ( .B1(n15439), .B2(n15438), .A(n11197), .ZN(n21606) );
  INV_X1 U17382 ( .A(n21606), .ZN(n15760) );
  OAI222_X1 U17383 ( .A1(n15509), .A2(n21603), .B1(n15440), .B2(n19892), .C1(
        n15760), .C2(n15497), .ZN(P1_U2847) );
  NOR2_X1 U17384 ( .A1(n15451), .A2(n15443), .ZN(n15444) );
  OR2_X1 U17385 ( .A1(n15445), .A2(n15444), .ZN(n21593) );
  OAI22_X1 U17386 ( .A1(n21593), .A2(n15497), .B1(n21579), .B2(n19892), .ZN(
        n15446) );
  INV_X1 U17387 ( .A(n15446), .ZN(n15447) );
  OAI21_X1 U17388 ( .B1(n21585), .B2(n15509), .A(n15447), .ZN(P1_U2848) );
  INV_X1 U17389 ( .A(n15448), .ZN(n15449) );
  OAI21_X1 U17390 ( .B1(n15450), .B2(n15432), .A(n15449), .ZN(n21573) );
  AOI21_X1 U17391 ( .B1(n15452), .B2(n15459), .A(n15451), .ZN(n21575) );
  AOI22_X1 U17392 ( .A1(n21575), .A2(n19888), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15507), .ZN(n15453) );
  OAI21_X1 U17393 ( .B1(n21573), .B2(n15509), .A(n15453), .ZN(P1_U2849) );
  INV_X1 U17394 ( .A(n15432), .ZN(n15455) );
  OAI21_X1 U17395 ( .B1(n15456), .B2(n15454), .A(n15455), .ZN(n21556) );
  NAND2_X1 U17396 ( .A1(n15464), .A2(n15457), .ZN(n15458) );
  AND2_X1 U17397 ( .A1(n15459), .A2(n15458), .ZN(n21554) );
  AOI22_X1 U17398 ( .A1(n21554), .A2(n19888), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15507), .ZN(n15460) );
  OAI21_X1 U17399 ( .B1(n21556), .B2(n15509), .A(n15460), .ZN(P1_U2850) );
  AOI21_X1 U17400 ( .B1(n15462), .B2(n15461), .A(n15454), .ZN(n19960) );
  INV_X1 U17401 ( .A(n19960), .ZN(n21548) );
  INV_X1 U17402 ( .A(n15463), .ZN(n15466) );
  INV_X1 U17403 ( .A(n15464), .ZN(n15465) );
  AOI21_X1 U17404 ( .B1(n15467), .B2(n15466), .A(n15465), .ZN(n21550) );
  AOI22_X1 U17405 ( .A1(n21550), .A2(n19888), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15507), .ZN(n15468) );
  OAI21_X1 U17406 ( .B1(n21548), .B2(n15509), .A(n15468), .ZN(P1_U2851) );
  OAI22_X1 U17407 ( .A1(n21372), .A2(n15497), .B1(n15469), .B2(n19892), .ZN(
        n15470) );
  INV_X1 U17408 ( .A(n15470), .ZN(n15471) );
  OAI21_X1 U17409 ( .B1(n15661), .B2(n15509), .A(n15471), .ZN(P1_U2852) );
  NAND2_X1 U17410 ( .A1(n15472), .A2(n15473), .ZN(n15474) );
  AND2_X1 U17411 ( .A1(n15475), .A2(n15474), .ZN(n21540) );
  AND2_X1 U17412 ( .A1(n15486), .A2(n15476), .ZN(n15478) );
  OR2_X1 U17413 ( .A1(n15478), .A2(n15477), .ZN(n21543) );
  INV_X1 U17414 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15479) );
  OAI22_X1 U17415 ( .A1(n21543), .A2(n15497), .B1(n15479), .B2(n19892), .ZN(
        n15480) );
  AOI21_X1 U17416 ( .B1(n21540), .B2(n19889), .A(n15480), .ZN(n15481) );
  INV_X1 U17417 ( .A(n15481), .ZN(P1_U2853) );
  OAI21_X1 U17418 ( .B1(n15379), .B2(n15482), .A(n15472), .ZN(n15571) );
  INV_X1 U17419 ( .A(n15571), .ZN(n21525) );
  NAND2_X1 U17420 ( .A1(n15484), .A2(n15483), .ZN(n15485) );
  NAND2_X1 U17421 ( .A1(n15486), .A2(n15485), .ZN(n21528) );
  OAI22_X1 U17422 ( .A1(n21528), .A2(n15497), .B1(n21521), .B2(n19892), .ZN(
        n15487) );
  AOI21_X1 U17423 ( .B1(n21525), .B2(n19889), .A(n15487), .ZN(n15488) );
  INV_X1 U17424 ( .A(n15488), .ZN(P1_U2854) );
  INV_X1 U17425 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15489) );
  INV_X1 U17426 ( .A(n19947), .ZN(n15576) );
  OAI222_X1 U17427 ( .A1(n15490), .A2(n15497), .B1(n15489), .B2(n19892), .C1(
        n15576), .C2(n15509), .ZN(P1_U2855) );
  AND2_X1 U17428 ( .A1(n15500), .A2(n15491), .ZN(n15493) );
  OR2_X1 U17429 ( .A1(n15493), .A2(n15492), .ZN(n21514) );
  AND2_X1 U17430 ( .A1(n15506), .A2(n15494), .ZN(n15496) );
  OR2_X1 U17431 ( .A1(n15496), .A2(n15495), .ZN(n21518) );
  OAI22_X1 U17432 ( .A1(n21518), .A2(n15497), .B1(n21508), .B2(n19892), .ZN(
        n15498) );
  INV_X1 U17433 ( .A(n15498), .ZN(n15499) );
  OAI21_X1 U17434 ( .B1(n21514), .B2(n15509), .A(n15499), .ZN(P1_U2856) );
  INV_X1 U17435 ( .A(n15500), .ZN(n15501) );
  AOI21_X1 U17436 ( .B1(n15502), .B2(n14846), .A(n15501), .ZN(n21502) );
  INV_X1 U17437 ( .A(n21502), .ZN(n15586) );
  NAND2_X1 U17438 ( .A1(n15504), .A2(n15503), .ZN(n15505) );
  AND2_X1 U17439 ( .A1(n15506), .A2(n15505), .ZN(n21500) );
  AOI22_X1 U17440 ( .A1(n21500), .A2(n19888), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n15507), .ZN(n15508) );
  OAI21_X1 U17441 ( .B1(n15586), .B2(n15509), .A(n15508), .ZN(P1_U2857) );
  AND2_X1 U17442 ( .A1(n22104), .A2(n15511), .ZN(n15512) );
  NAND2_X1 U17443 ( .A1(n15553), .A2(n15512), .ZN(n15578) );
  OAI22_X1 U17444 ( .A1(n15578), .A2(n15513), .B1(n15553), .B2(n14316), .ZN(
        n15514) );
  AOI21_X1 U17445 ( .B1(n15580), .B2(BUF1_REG_30__SCAN_IN), .A(n15514), .ZN(
        n15516) );
  NAND2_X1 U17446 ( .A1(n15581), .A2(DATAI_30_), .ZN(n15515) );
  OAI211_X1 U17447 ( .C1(n15517), .C2(n15587), .A(n15516), .B(n15515), .ZN(
        P1_U2874) );
  OAI22_X1 U17448 ( .A1(n15578), .A2(n15518), .B1(n15553), .B2(n14324), .ZN(
        n15519) );
  AOI21_X1 U17449 ( .B1(n15580), .B2(BUF1_REG_29__SCAN_IN), .A(n15519), .ZN(
        n15521) );
  NAND2_X1 U17450 ( .A1(n15581), .A2(DATAI_29_), .ZN(n15520) );
  OAI211_X1 U17451 ( .C1(n15522), .C2(n15587), .A(n15521), .B(n15520), .ZN(
        P1_U2875) );
  OAI22_X1 U17452 ( .A1(n15578), .A2(n15523), .B1(n15553), .B2(n14312), .ZN(
        n15524) );
  AOI21_X1 U17453 ( .B1(n15580), .B2(BUF1_REG_28__SCAN_IN), .A(n15524), .ZN(
        n15526) );
  NAND2_X1 U17454 ( .A1(n15581), .A2(DATAI_28_), .ZN(n15525) );
  OAI211_X1 U17455 ( .C1(n15607), .C2(n15587), .A(n15526), .B(n15525), .ZN(
        P1_U2876) );
  OAI22_X1 U17456 ( .A1(n15578), .A2(n15527), .B1(n15553), .B2(n14310), .ZN(
        n15528) );
  AOI21_X1 U17457 ( .B1(n15580), .B2(BUF1_REG_27__SCAN_IN), .A(n15528), .ZN(
        n15530) );
  NAND2_X1 U17458 ( .A1(n15581), .A2(DATAI_27_), .ZN(n15529) );
  OAI211_X1 U17459 ( .C1(n15531), .C2(n15587), .A(n15530), .B(n15529), .ZN(
        P1_U2877) );
  OAI22_X1 U17460 ( .A1(n15578), .A2(n15532), .B1(n15553), .B2(n14318), .ZN(
        n15533) );
  AOI21_X1 U17461 ( .B1(n15580), .B2(BUF1_REG_26__SCAN_IN), .A(n15533), .ZN(
        n15535) );
  NAND2_X1 U17462 ( .A1(n15581), .A2(DATAI_26_), .ZN(n15534) );
  OAI211_X1 U17463 ( .C1(n15536), .C2(n15587), .A(n15535), .B(n15534), .ZN(
        P1_U2878) );
  OAI22_X1 U17464 ( .A1(n15578), .A2(n15537), .B1(n15553), .B2(n14314), .ZN(
        n15538) );
  AOI21_X1 U17465 ( .B1(n15580), .B2(BUF1_REG_25__SCAN_IN), .A(n15538), .ZN(
        n15540) );
  NAND2_X1 U17466 ( .A1(n15581), .A2(DATAI_25_), .ZN(n15539) );
  OAI211_X1 U17467 ( .C1(n21603), .C2(n15587), .A(n15540), .B(n15539), .ZN(
        P1_U2879) );
  OAI22_X1 U17468 ( .A1(n15578), .A2(n15541), .B1(n15553), .B2(n14306), .ZN(
        n15542) );
  AOI21_X1 U17469 ( .B1(n15580), .B2(BUF1_REG_24__SCAN_IN), .A(n15542), .ZN(
        n15544) );
  NAND2_X1 U17470 ( .A1(n15581), .A2(DATAI_24_), .ZN(n15543) );
  OAI211_X1 U17471 ( .C1(n21585), .C2(n15587), .A(n15544), .B(n15543), .ZN(
        P1_U2880) );
  OAI22_X1 U17472 ( .A1(n15578), .A2(n15545), .B1(n15553), .B2(n14297), .ZN(
        n15546) );
  AOI21_X1 U17473 ( .B1(n15580), .B2(BUF1_REG_23__SCAN_IN), .A(n15546), .ZN(
        n15548) );
  NAND2_X1 U17474 ( .A1(n15581), .A2(DATAI_23_), .ZN(n15547) );
  OAI211_X1 U17475 ( .C1(n21573), .C2(n15587), .A(n15548), .B(n15547), .ZN(
        P1_U2881) );
  OAI22_X1 U17476 ( .A1(n15578), .A2(n15549), .B1(n15553), .B2(n14308), .ZN(
        n15550) );
  AOI21_X1 U17477 ( .B1(n15580), .B2(BUF1_REG_22__SCAN_IN), .A(n15550), .ZN(
        n15552) );
  NAND2_X1 U17478 ( .A1(n15581), .A2(DATAI_22_), .ZN(n15551) );
  OAI211_X1 U17479 ( .C1(n21556), .C2(n15587), .A(n15552), .B(n15551), .ZN(
        P1_U2882) );
  OAI22_X1 U17480 ( .A1(n15578), .A2(n15554), .B1(n15553), .B2(n14320), .ZN(
        n15555) );
  AOI21_X1 U17481 ( .B1(n15580), .B2(BUF1_REG_21__SCAN_IN), .A(n15555), .ZN(
        n15557) );
  NAND2_X1 U17482 ( .A1(n15581), .A2(DATAI_21_), .ZN(n15556) );
  OAI211_X1 U17483 ( .C1(n21548), .C2(n15587), .A(n15557), .B(n15556), .ZN(
        P1_U2883) );
  OAI22_X1 U17484 ( .A1(n15578), .A2(n15558), .B1(n15553), .B2(n14327), .ZN(
        n15559) );
  AOI21_X1 U17485 ( .B1(n15580), .B2(BUF1_REG_20__SCAN_IN), .A(n15559), .ZN(
        n15561) );
  NAND2_X1 U17486 ( .A1(n15581), .A2(DATAI_20_), .ZN(n15560) );
  OAI211_X1 U17487 ( .C1(n15661), .C2(n15587), .A(n15561), .B(n15560), .ZN(
        P1_U2884) );
  INV_X1 U17488 ( .A(n21540), .ZN(n15566) );
  OAI22_X1 U17489 ( .A1(n15578), .A2(n15562), .B1(n15553), .B2(n14322), .ZN(
        n15563) );
  AOI21_X1 U17490 ( .B1(n15580), .B2(BUF1_REG_19__SCAN_IN), .A(n15563), .ZN(
        n15565) );
  NAND2_X1 U17491 ( .A1(n15581), .A2(DATAI_19_), .ZN(n15564) );
  OAI211_X1 U17492 ( .C1(n15566), .C2(n15587), .A(n15565), .B(n15564), .ZN(
        P1_U2885) );
  OAI22_X1 U17493 ( .A1(n15578), .A2(n15567), .B1(n15553), .B2(n14122), .ZN(
        n15568) );
  AOI21_X1 U17494 ( .B1(n15580), .B2(BUF1_REG_18__SCAN_IN), .A(n15568), .ZN(
        n15570) );
  NAND2_X1 U17495 ( .A1(n15581), .A2(DATAI_18_), .ZN(n15569) );
  OAI211_X1 U17496 ( .C1(n15571), .C2(n15587), .A(n15570), .B(n15569), .ZN(
        P1_U2886) );
  OAI22_X1 U17497 ( .A1(n15578), .A2(n15572), .B1(n15553), .B2(n14120), .ZN(
        n15573) );
  AOI21_X1 U17498 ( .B1(n15580), .B2(BUF1_REG_17__SCAN_IN), .A(n15573), .ZN(
        n15575) );
  NAND2_X1 U17499 ( .A1(n15581), .A2(DATAI_17_), .ZN(n15574) );
  OAI211_X1 U17500 ( .C1(n15576), .C2(n15587), .A(n15575), .B(n15574), .ZN(
        P1_U2887) );
  OAI22_X1 U17501 ( .A1(n15578), .A2(n15577), .B1(n15553), .B2(n14295), .ZN(
        n15579) );
  AOI21_X1 U17502 ( .B1(n15580), .B2(BUF1_REG_16__SCAN_IN), .A(n15579), .ZN(
        n15583) );
  NAND2_X1 U17503 ( .A1(n15581), .A2(DATAI_16_), .ZN(n15582) );
  OAI211_X1 U17504 ( .C1(n21514), .C2(n15587), .A(n15583), .B(n15582), .ZN(
        P1_U2888) );
  OAI222_X1 U17505 ( .A1(n15587), .A2(n15586), .B1(n15553), .B2(n19816), .C1(
        n15585), .C2(n15584), .ZN(P1_U2889) );
  INV_X1 U17506 ( .A(n15588), .ZN(n15593) );
  OAI21_X1 U17507 ( .B1(n15592), .B2(n15590), .A(n15589), .ZN(n15591) );
  NOR2_X1 U17508 ( .A1(n21373), .A2(n16933), .ZN(n15714) );
  AOI21_X1 U17509 ( .B1(n19955), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15714), .ZN(n15594) );
  OAI21_X1 U17510 ( .B1(n19964), .B2(n15595), .A(n15594), .ZN(n15596) );
  AOI21_X1 U17511 ( .B1(n15597), .B2(n19952), .A(n15596), .ZN(n15598) );
  OAI21_X1 U17512 ( .B1(n15721), .B2(n21610), .A(n15598), .ZN(P1_U2970) );
  NAND3_X1 U17513 ( .A1(n15599), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15600), .ZN(n15604) );
  OR3_X1 U17514 ( .A1(n15599), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15601), .ZN(n15603) );
  MUX2_X1 U17515 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n15747), .S(
        n13221), .Z(n15602) );
  AOI21_X1 U17516 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15605) );
  XNOR2_X1 U17517 ( .A(n15605), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15733) );
  NAND2_X1 U17518 ( .A1(n13790), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15727) );
  OAI21_X1 U17519 ( .B1(n19923), .B2(n15606), .A(n15727), .ZN(n15609) );
  NOR2_X1 U17520 ( .A1(n15607), .A2(n15679), .ZN(n15608) );
  OAI21_X1 U17521 ( .B1(n15733), .B2(n21610), .A(n15611), .ZN(P1_U2971) );
  XNOR2_X1 U17522 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15613) );
  XNOR2_X1 U17523 ( .A(n15612), .B(n15613), .ZN(n15742) );
  NAND2_X1 U17524 ( .A1(n13790), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15736) );
  NAND2_X1 U17525 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15614) );
  OAI211_X1 U17526 ( .C1(n19964), .C2(n15615), .A(n15736), .B(n15614), .ZN(
        n15616) );
  AOI21_X1 U17527 ( .B1(n15617), .B2(n19952), .A(n15616), .ZN(n15618) );
  OAI21_X1 U17528 ( .B1(n15742), .B2(n21610), .A(n15618), .ZN(P1_U2972) );
  XNOR2_X1 U17529 ( .A(n15619), .B(n15747), .ZN(n15751) );
  INV_X1 U17530 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15622) );
  NAND2_X1 U17531 ( .A1(n19946), .A2(n15620), .ZN(n15621) );
  NAND2_X1 U17532 ( .A1(n13790), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15745) );
  OAI211_X1 U17533 ( .C1(n19923), .C2(n15622), .A(n15621), .B(n15745), .ZN(
        n15623) );
  AOI21_X1 U17534 ( .B1(n15624), .B2(n19952), .A(n15623), .ZN(n15625) );
  OAI21_X1 U17535 ( .B1(n15751), .B2(n21610), .A(n15625), .ZN(P1_U2973) );
  OAI21_X1 U17536 ( .B1(n15599), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15626), .ZN(n15628) );
  NAND2_X1 U17537 ( .A1(n13212), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15639) );
  NAND3_X1 U17538 ( .A1(n15628), .A2(n15627), .A3(n15639), .ZN(n15629) );
  XNOR2_X1 U17539 ( .A(n15629), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15752) );
  NAND2_X1 U17540 ( .A1(n15752), .A2(n19961), .ZN(n15632) );
  NOR2_X1 U17541 ( .A1(n21373), .A2(n21595), .ZN(n15755) );
  NOR2_X1 U17542 ( .A1(n19964), .A2(n21601), .ZN(n15630) );
  AOI211_X1 U17543 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15755), .B(n15630), .ZN(n15631) );
  OAI211_X1 U17544 ( .C1(n15679), .C2(n21603), .A(n15632), .B(n15631), .ZN(
        P1_U2974) );
  NAND2_X1 U17545 ( .A1(n15599), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15634) );
  INV_X1 U17546 ( .A(n15599), .ZN(n15641) );
  NAND2_X1 U17547 ( .A1(n15641), .A2(n15763), .ZN(n15633) );
  MUX2_X1 U17548 ( .A(n15634), .B(n15633), .S(n13212), .Z(n15635) );
  XNOR2_X1 U17549 ( .A(n15635), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15761) );
  NAND2_X1 U17550 ( .A1(n15761), .A2(n19961), .ZN(n15638) );
  INV_X1 U17551 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21582) );
  NOR2_X1 U17552 ( .A1(n21373), .A2(n21582), .ZN(n15765) );
  INV_X1 U17553 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21578) );
  NOR2_X1 U17554 ( .A1(n19923), .A2(n21578), .ZN(n15636) );
  AOI211_X1 U17555 ( .C1(n19946), .C2(n21587), .A(n15765), .B(n15636), .ZN(
        n15637) );
  OAI211_X1 U17556 ( .C1(n15679), .C2(n21585), .A(n15638), .B(n15637), .ZN(
        P1_U2975) );
  OAI21_X1 U17557 ( .B1(n13212), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15639), .ZN(n15640) );
  XNOR2_X1 U17558 ( .A(n15641), .B(n15640), .ZN(n15774) );
  NAND2_X1 U17559 ( .A1(n13790), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15769) );
  OAI21_X1 U17560 ( .B1(n19923), .B2(n15642), .A(n15769), .ZN(n15644) );
  NOR2_X1 U17561 ( .A1(n21573), .A2(n15679), .ZN(n15643) );
  AOI211_X1 U17562 ( .C1(n19946), .C2(n21571), .A(n15644), .B(n15643), .ZN(
        n15645) );
  OAI21_X1 U17563 ( .B1(n15774), .B2(n21610), .A(n15645), .ZN(P1_U2976) );
  NAND2_X1 U17564 ( .A1(n15647), .A2(n15646), .ZN(n15648) );
  XNOR2_X1 U17565 ( .A(n15648), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15775) );
  NAND2_X1 U17566 ( .A1(n15775), .A2(n19961), .ZN(n15652) );
  INV_X1 U17567 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21561) );
  NOR2_X1 U17568 ( .A1(n21373), .A2(n21561), .ZN(n15783) );
  NOR2_X1 U17569 ( .A1(n19923), .A2(n15649), .ZN(n15650) );
  AOI211_X1 U17570 ( .C1(n19946), .C2(n21558), .A(n15783), .B(n15650), .ZN(
        n15651) );
  OAI211_X1 U17571 ( .C1(n15679), .C2(n21556), .A(n15652), .B(n15651), .ZN(
        P1_U2977) );
  MUX2_X1 U17572 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n13388), .S(
        n13221), .Z(n15662) );
  NOR2_X1 U17573 ( .A1(n15653), .A2(n15662), .ZN(n15663) );
  AOI21_X1 U17574 ( .B1(n13212), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15663), .ZN(n19951) );
  OAI22_X1 U17575 ( .A1(n19951), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13212), .B2(n15663), .ZN(n19956) );
  AOI21_X1 U17576 ( .B1(n13212), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n19956), .ZN(n15654) );
  XNOR2_X1 U17577 ( .A(n15654), .B(n19958), .ZN(n21368) );
  NAND2_X1 U17578 ( .A1(n21368), .A2(n19961), .ZN(n15660) );
  INV_X1 U17579 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15655) );
  OAI22_X1 U17580 ( .A1(n19923), .A2(n15656), .B1(n21373), .B2(n15655), .ZN(
        n15657) );
  AOI21_X1 U17581 ( .B1(n19946), .B2(n15658), .A(n15657), .ZN(n15659) );
  OAI211_X1 U17582 ( .C1(n15679), .C2(n15661), .A(n15660), .B(n15659), .ZN(
        P1_U2979) );
  INV_X1 U17583 ( .A(n15662), .ZN(n15665) );
  INV_X1 U17584 ( .A(n15663), .ZN(n15664) );
  OAI21_X1 U17585 ( .B1(n15665), .B2(n13224), .A(n15664), .ZN(n21343) );
  AOI22_X1 U17586 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15666) );
  OAI21_X1 U17587 ( .B1(n19964), .B2(n21523), .A(n15666), .ZN(n15667) );
  AOI21_X1 U17588 ( .B1(n21525), .B2(n19952), .A(n15667), .ZN(n15668) );
  OAI21_X1 U17589 ( .B1(n21343), .B2(n21610), .A(n15668), .ZN(P1_U2981) );
  OAI21_X1 U17590 ( .B1(n15681), .B2(n15670), .A(n15669), .ZN(n19937) );
  INV_X1 U17591 ( .A(n15671), .ZN(n15672) );
  NOR3_X1 U17592 ( .A1(n19937), .A2(n19933), .A3(n15672), .ZN(n19935) );
  NOR2_X1 U17593 ( .A1(n19935), .A2(n19933), .ZN(n15674) );
  XNOR2_X1 U17594 ( .A(n15674), .B(n15673), .ZN(n21359) );
  NAND2_X1 U17595 ( .A1(n21359), .A2(n19961), .ZN(n15678) );
  OAI22_X1 U17596 ( .A1(n19923), .A2(n15675), .B1(n21373), .B2(n19832), .ZN(
        n15676) );
  AOI21_X1 U17597 ( .B1(n21512), .B2(n19946), .A(n15676), .ZN(n15677) );
  OAI211_X1 U17598 ( .C1(n15679), .C2(n21514), .A(n15678), .B(n15677), .ZN(
        P1_U2983) );
  NAND2_X1 U17599 ( .A1(n15681), .A2(n15680), .ZN(n15683) );
  AOI22_X1 U17600 ( .A1(n15683), .A2(n15682), .B1(n13212), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15685) );
  MUX2_X1 U17601 ( .A(n13377), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n13221), .Z(n15684) );
  XNOR2_X1 U17602 ( .A(n15685), .B(n15684), .ZN(n21224) );
  INV_X1 U17603 ( .A(n21224), .ZN(n15691) );
  AOI22_X1 U17604 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15686) );
  OAI21_X1 U17605 ( .B1(n19964), .B2(n15687), .A(n15686), .ZN(n15688) );
  AOI21_X1 U17606 ( .B1(n15689), .B2(n19952), .A(n15688), .ZN(n15690) );
  OAI21_X1 U17607 ( .B1(n15691), .B2(n21610), .A(n15690), .ZN(P1_U2985) );
  INV_X1 U17608 ( .A(n15693), .ZN(n15694) );
  AOI21_X1 U17609 ( .B1(n15692), .B2(n15695), .A(n15694), .ZN(n19924) );
  NAND3_X1 U17610 ( .A1(n19924), .A2(n19925), .A3(n15696), .ZN(n19926) );
  NAND2_X1 U17611 ( .A1(n19926), .A2(n19925), .ZN(n15697) );
  XOR2_X1 U17612 ( .A(n15698), .B(n15697), .Z(n21211) );
  AOI22_X1 U17613 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15699) );
  OAI21_X1 U17614 ( .B1(n19964), .B2(n15700), .A(n15699), .ZN(n15701) );
  AOI21_X1 U17615 ( .B1(n15702), .B2(n19952), .A(n15701), .ZN(n15703) );
  OAI21_X1 U17616 ( .B1(n21211), .B2(n21610), .A(n15703), .ZN(P1_U2986) );
  MUX2_X1 U17617 ( .A(n15173), .B(n15692), .S(n13212), .Z(n15704) );
  NOR2_X1 U17618 ( .A1(n15704), .A2(n15705), .ZN(n19917) );
  AOI21_X1 U17619 ( .B1(n15705), .B2(n15704), .A(n19917), .ZN(n21306) );
  INV_X1 U17620 ( .A(n21306), .ZN(n15712) );
  INV_X1 U17621 ( .A(n15706), .ZN(n15710) );
  AOI22_X1 U17622 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15707) );
  OAI21_X1 U17623 ( .B1(n19964), .B2(n15708), .A(n15707), .ZN(n15709) );
  AOI21_X1 U17624 ( .B1(n15710), .B2(n19952), .A(n15709), .ZN(n15711) );
  OAI21_X1 U17625 ( .B1(n15712), .B2(n21610), .A(n15711), .ZN(P1_U2989) );
  INV_X1 U17626 ( .A(n15713), .ZN(n15717) );
  AOI21_X1 U17627 ( .B1(n15715), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15714), .ZN(n15716) );
  OAI21_X1 U17628 ( .B1(n15717), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15716), .ZN(n15718) );
  AOI21_X1 U17629 ( .B1(n15719), .B2(n21382), .A(n15718), .ZN(n15720) );
  OAI21_X1 U17630 ( .B1(n15721), .B2(n21353), .A(n15720), .ZN(P1_U3002) );
  INV_X1 U17631 ( .A(n15722), .ZN(n15731) );
  NOR3_X1 U17632 ( .A1(n15738), .A2(n15724), .A3(n15723), .ZN(n15730) );
  INV_X1 U17633 ( .A(n15725), .ZN(n15735) );
  INV_X1 U17634 ( .A(n15726), .ZN(n15734) );
  NAND3_X1 U17635 ( .A1(n15735), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15734), .ZN(n15728) );
  NAND2_X1 U17636 ( .A1(n15728), .A2(n15727), .ZN(n15729) );
  AOI211_X1 U17637 ( .C1(n15731), .C2(n21382), .A(n15730), .B(n15729), .ZN(
        n15732) );
  OAI21_X1 U17638 ( .B1(n15733), .B2(n21353), .A(n15732), .ZN(P1_U3003) );
  NAND3_X1 U17639 ( .A1(n15735), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15734), .ZN(n15737) );
  OAI211_X1 U17640 ( .C1(n15738), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15737), .B(n15736), .ZN(n15739) );
  AOI21_X1 U17641 ( .B1(n15740), .B2(n21382), .A(n15739), .ZN(n15741) );
  OAI21_X1 U17642 ( .B1(n15742), .B2(n21353), .A(n15741), .ZN(P1_U3004) );
  INV_X1 U17643 ( .A(n15743), .ZN(n15753) );
  XNOR2_X1 U17644 ( .A(n15756), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15744) );
  NAND2_X1 U17645 ( .A1(n15757), .A2(n15744), .ZN(n15746) );
  OAI211_X1 U17646 ( .C1(n15753), .C2(n15747), .A(n15746), .B(n15745), .ZN(
        n15748) );
  AOI21_X1 U17647 ( .B1(n15749), .B2(n21382), .A(n15748), .ZN(n15750) );
  OAI21_X1 U17648 ( .B1(n15751), .B2(n21353), .A(n15750), .ZN(P1_U3005) );
  NAND2_X1 U17649 ( .A1(n15752), .A2(n21393), .ZN(n15759) );
  NOR2_X1 U17650 ( .A1(n15753), .A2(n15756), .ZN(n15754) );
  AOI211_X1 U17651 ( .C1(n15757), .C2(n15756), .A(n15755), .B(n15754), .ZN(
        n15758) );
  OAI211_X1 U17652 ( .C1(n21399), .C2(n15760), .A(n15759), .B(n15758), .ZN(
        P1_U3006) );
  NAND2_X1 U17653 ( .A1(n15761), .A2(n21393), .ZN(n15767) );
  NOR3_X1 U17654 ( .A1(n15771), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15763), .ZN(n15764) );
  AOI211_X1 U17655 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15768), .A(
        n15765), .B(n15764), .ZN(n15766) );
  OAI211_X1 U17656 ( .C1(n21399), .C2(n21593), .A(n15767), .B(n15766), .ZN(
        P1_U3007) );
  NAND2_X1 U17657 ( .A1(n15768), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15770) );
  OAI211_X1 U17658 ( .C1(n15771), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15770), .B(n15769), .ZN(n15772) );
  AOI21_X1 U17659 ( .B1(n21575), .B2(n21382), .A(n15772), .ZN(n15773) );
  OAI21_X1 U17660 ( .B1(n15774), .B2(n21353), .A(n15773), .ZN(P1_U3008) );
  INV_X1 U17661 ( .A(n15775), .ZN(n15789) );
  NAND2_X1 U17662 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21203) );
  NAND2_X1 U17663 ( .A1(n21314), .A2(n15776), .ZN(n21222) );
  NAND2_X1 U17664 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21206), .ZN(
        n15777) );
  OAI22_X1 U17665 ( .A1(n21203), .A2(n21222), .B1(n21205), .B2(n15777), .ZN(
        n21208) );
  NAND2_X1 U17666 ( .A1(n15778), .A2(n21208), .ZN(n21366) );
  NAND2_X1 U17667 ( .A1(n15779), .A2(n21366), .ZN(n21364) );
  INV_X1 U17668 ( .A(n21364), .ZN(n21379) );
  INV_X1 U17669 ( .A(n15780), .ZN(n15781) );
  NOR3_X1 U17670 ( .A1(n21379), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15781), .ZN(n15782) );
  AOI211_X1 U17671 ( .C1(n21554), .C2(n21382), .A(n15783), .B(n15782), .ZN(
        n15788) );
  INV_X1 U17672 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21378) );
  NOR4_X1 U17673 ( .A1(n21379), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n19958), .A4(n21378), .ZN(n21383) );
  AOI21_X1 U17674 ( .B1(n21314), .B2(n15785), .A(n15784), .ZN(n21377) );
  NOR2_X1 U17675 ( .A1(n21378), .A2(n19958), .ZN(n15786) );
  AOI22_X1 U17676 ( .A1(n21377), .A2(n15786), .B1(n21389), .B2(n21300), .ZN(
        n21381) );
  OAI21_X1 U17677 ( .B1(n21383), .B2(n21381), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15787) );
  OAI211_X1 U17678 ( .C1(n15789), .C2(n21353), .A(n15788), .B(n15787), .ZN(
        P1_U3009) );
  OAI211_X1 U17679 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n14068), .A(n21838), 
        .B(n21908), .ZN(n15790) );
  OAI21_X1 U17680 ( .B1(n15791), .B2(n21805), .A(n15790), .ZN(n15792) );
  MUX2_X1 U17681 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15792), .S(
        n16768), .Z(P1_U3477) );
  NOR2_X1 U17682 ( .A1(n14063), .A2(n13698), .ZN(n15800) );
  AOI22_X1 U17683 ( .A1(n15794), .A2(n12821), .B1(n15800), .B2(n15793), .ZN(
        n15795) );
  OAI21_X1 U17684 ( .B1(n21805), .B2(n15796), .A(n15795), .ZN(n16738) );
  INV_X1 U17685 ( .A(n16738), .ZN(n15803) );
  INV_X1 U17686 ( .A(n15797), .ZN(n15807) );
  AOI22_X1 U17687 ( .A1(n15801), .A2(n15800), .B1(n15799), .B2(n15798), .ZN(
        n15802) );
  OAI21_X1 U17688 ( .B1(n15803), .B2(n15807), .A(n15802), .ZN(n15804) );
  MUX2_X1 U17689 ( .A(n15804), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15809), .Z(P1_U3473) );
  OAI22_X1 U17690 ( .A1(n15808), .A2(n15807), .B1(n15806), .B2(n15805), .ZN(
        n15810) );
  MUX2_X1 U17691 ( .A(n15810), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15809), .Z(P1_U3469) );
  INV_X1 U17692 ( .A(n18049), .ZN(n18053) );
  AOI22_X1 U17693 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18022), .ZN(n15812) );
  INV_X1 U17694 ( .A(n15812), .ZN(n18039) );
  OAI22_X1 U17695 ( .A1(n18022), .A2(n18435), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n16680) );
  OR2_X1 U17696 ( .A1(n18039), .A2(n16680), .ZN(n15834) );
  NOR2_X1 U17697 ( .A1(n15835), .A2(n15834), .ZN(n18063) );
  NOR2_X1 U17698 ( .A1(n18246), .A2(n18063), .ZN(n15813) );
  XNOR2_X1 U17699 ( .A(n15813), .B(n18062), .ZN(n15832) );
  NAND4_X1 U17700 ( .A1(n18022), .A2(n19164), .A3(n21639), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n18516) );
  INV_X1 U17701 ( .A(n18516), .ZN(n18386) );
  NOR2_X1 U17702 ( .A1(n15814), .A2(n18283), .ZN(n15831) );
  NAND2_X1 U17703 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19164), .ZN(n18518) );
  NOR3_X1 U17704 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19183), .A3(n18518), 
        .ZN(n18521) );
  NOR4_X4 U17705 ( .A1(n16539), .A2(n18371), .A3(n16965), .A4(n18521), .ZN(
        n18378) );
  INV_X1 U17706 ( .A(n18527), .ZN(n21665) );
  OAI21_X1 U17707 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n21665), .A(
        P2_EBX_REG_31__SCAN_IN), .ZN(n15816) );
  INV_X1 U17708 ( .A(n15816), .ZN(n15817) );
  AND2_X1 U17709 ( .A1(n16011), .A2(n15817), .ZN(n15818) );
  OAI22_X1 U17710 ( .A1(n14356), .A2(n18396), .B1(n15819), .B2(n18394), .ZN(
        n15828) );
  OR2_X1 U17711 ( .A1(n15821), .A2(n15820), .ZN(n18398) );
  INV_X1 U17712 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n18399) );
  OAI21_X1 U17713 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n21665), .A(n18399), 
        .ZN(n15822) );
  INV_X1 U17714 ( .A(n15822), .ZN(n15823) );
  NAND2_X1 U17715 ( .A1(n15824), .A2(n15823), .ZN(n15825) );
  NAND2_X1 U17716 ( .A1(n18398), .A2(n15825), .ZN(n18381) );
  INV_X1 U17717 ( .A(n18381), .ZN(n18344) );
  OAI22_X1 U17718 ( .A1(n18344), .A2(n12148), .B1(n15826), .B2(n18340), .ZN(
        n15827) );
  NOR2_X1 U17719 ( .A1(n15828), .A2(n15827), .ZN(n15829) );
  OAI21_X1 U17720 ( .B1(n17056), .B2(n18354), .A(n15829), .ZN(n15830) );
  AOI211_X1 U17721 ( .C1(n15832), .C2(n18371), .A(n15831), .B(n15830), .ZN(
        n15833) );
  OAI21_X1 U17722 ( .B1(n19198), .B2(n18053), .A(n15833), .ZN(P2_U2852) );
  NAND2_X1 U17723 ( .A1(n18385), .A2(n15834), .ZN(n16679) );
  XNOR2_X1 U17724 ( .A(n15835), .B(n16679), .ZN(n15844) );
  NOR2_X1 U17725 ( .A1(n19142), .A2(n18053), .ZN(n15843) );
  OAI22_X1 U17726 ( .A1(n18491), .A2(n18354), .B1(n15836), .B2(n18340), .ZN(
        n15837) );
  INV_X1 U17727 ( .A(n15837), .ZN(n15841) );
  OAI22_X1 U17728 ( .A1(n11889), .A2(n18396), .B1(n15838), .B2(n18394), .ZN(
        n15839) );
  AOI21_X1 U17729 ( .B1(n18381), .B2(P2_EBX_REG_2__SCAN_IN), .A(n15839), .ZN(
        n15840) );
  OAI211_X1 U17730 ( .C1(n18283), .C2(n11138), .A(n15841), .B(n15840), .ZN(
        n15842) );
  AOI211_X1 U17731 ( .C1(n15844), .C2(n18371), .A(n15843), .B(n15842), .ZN(
        n15845) );
  INV_X1 U17732 ( .A(n15845), .ZN(P2_U2853) );
  NAND2_X1 U17733 ( .A1(n18403), .A2(n16112), .ZN(n15846) );
  OAI21_X1 U17734 ( .B1(n16112), .B2(n18399), .A(n15846), .ZN(P2_U2856) );
  AOI22_X1 U17735 ( .A1(n12126), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U17736 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15848) );
  AOI22_X1 U17737 ( .A1(n12092), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15847) );
  NAND3_X1 U17738 ( .A1(n15849), .A2(n15848), .A3(n15847), .ZN(n15863) );
  NAND2_X1 U17739 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n15851) );
  NAND2_X1 U17740 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15850) );
  OAI211_X1 U17741 ( .C1(n15874), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        n15857) );
  NAND2_X1 U17742 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n15854) );
  NAND2_X1 U17743 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n15853) );
  OAI211_X1 U17744 ( .C1(n12015), .C2(n15855), .A(n15854), .B(n15853), .ZN(
        n15856) );
  NOR2_X1 U17745 ( .A1(n15857), .A2(n15856), .ZN(n15861) );
  AOI22_X1 U17746 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15860) );
  NAND2_X1 U17747 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n15859) );
  NAND2_X1 U17748 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n15858) );
  NAND4_X1 U17749 ( .A1(n15861), .A2(n15860), .A3(n15859), .A4(n15858), .ZN(
        n15862) );
  OR2_X1 U17750 ( .A1(n15863), .A2(n15862), .ZN(n16108) );
  AOI22_X1 U17751 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12126), .B1(
        n14809), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15869) );
  AOI22_X1 U17752 ( .A1(n11998), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15865), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15868) );
  AOI22_X1 U17753 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12092), .B1(
        n15866), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15867) );
  NAND3_X1 U17754 ( .A1(n15869), .A2(n15868), .A3(n15867), .ZN(n15890) );
  NAND2_X1 U17755 ( .A1(n15870), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n15873) );
  NAND2_X1 U17756 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15872) );
  OAI211_X1 U17757 ( .C1(n15874), .C2(n19060), .A(n15873), .B(n15872), .ZN(
        n15881) );
  INV_X1 U17758 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15879) );
  NAND2_X1 U17759 ( .A1(n15875), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n15878) );
  NAND2_X1 U17760 ( .A1(n15876), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n15877) );
  OAI211_X1 U17761 ( .C1(n12015), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        n15880) );
  NOR2_X1 U17762 ( .A1(n15881), .A2(n15880), .ZN(n15888) );
  AOI22_X1 U17763 ( .A1(n12003), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15882), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15887) );
  NAND2_X1 U17764 ( .A1(n15883), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n15886) );
  NAND2_X1 U17765 ( .A1(n15884), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n15885) );
  NAND4_X1 U17766 ( .A1(n15888), .A2(n15887), .A3(n15886), .A4(n15885), .ZN(
        n15889) );
  OR2_X1 U17767 ( .A1(n15890), .A2(n15889), .ZN(n15912) );
  NAND2_X1 U17768 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15894) );
  AND2_X1 U17769 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15892) );
  OR2_X1 U17770 ( .A1(n15892), .A2(n15891), .ZN(n16037) );
  NAND2_X1 U17771 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n15893) );
  AND3_X1 U17772 ( .A1(n15894), .A2(n16037), .A3(n15893), .ZN(n15901) );
  AOI22_X1 U17773 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15900) );
  AOI22_X1 U17774 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U17775 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15898) );
  NAND4_X1 U17776 ( .A1(n15901), .A2(n15900), .A3(n15899), .A4(n15898), .ZN(
        n15909) );
  NAND2_X1 U17777 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15903) );
  INV_X1 U17778 ( .A(n16037), .ZN(n16001) );
  NAND2_X1 U17779 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15902) );
  AND3_X1 U17780 ( .A1(n15903), .A2(n16001), .A3(n15902), .ZN(n15907) );
  AOI22_X1 U17781 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15906) );
  AOI22_X1 U17782 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15905) );
  AOI22_X1 U17783 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15904) );
  NAND4_X1 U17784 ( .A1(n15907), .A2(n15906), .A3(n15905), .A4(n15904), .ZN(
        n15908) );
  NAND2_X1 U17785 ( .A1(n15909), .A2(n15908), .ZN(n15910) );
  XNOR2_X1 U17786 ( .A(n15912), .B(n15910), .ZN(n16099) );
  INV_X1 U17787 ( .A(n15910), .ZN(n15911) );
  AND2_X1 U17788 ( .A1(n15912), .A2(n15911), .ZN(n15914) );
  NAND2_X1 U17789 ( .A1(n15914), .A2(n15968), .ZN(n15913) );
  INV_X1 U17790 ( .A(n15914), .ZN(n15930) );
  NAND2_X1 U17791 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15916) );
  NAND2_X1 U17792 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n15915) );
  AND3_X1 U17793 ( .A1(n15916), .A2(n16037), .A3(n15915), .ZN(n15920) );
  AOI22_X1 U17794 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15919) );
  AOI22_X1 U17795 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15918) );
  AOI22_X1 U17796 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15917) );
  NAND4_X1 U17797 ( .A1(n15920), .A2(n15919), .A3(n15918), .A4(n15917), .ZN(
        n15928) );
  NAND2_X1 U17798 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15922) );
  NAND2_X1 U17799 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15921) );
  AND3_X1 U17800 ( .A1(n15922), .A2(n16001), .A3(n15921), .ZN(n15926) );
  AOI22_X1 U17801 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15925) );
  AOI22_X1 U17802 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15924) );
  AOI22_X1 U17803 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15923) );
  NAND4_X1 U17804 ( .A1(n15926), .A2(n15925), .A3(n15924), .A4(n15923), .ZN(
        n15927) );
  NAND2_X1 U17805 ( .A1(n15928), .A2(n15927), .ZN(n15929) );
  NOR2_X1 U17806 ( .A1(n15930), .A2(n15929), .ZN(n15948) );
  NAND2_X1 U17807 ( .A1(n15948), .A2(n16011), .ZN(n15933) );
  OAI21_X1 U17808 ( .B1(n15931), .B2(n15930), .A(n15929), .ZN(n15932) );
  AND2_X1 U17809 ( .A1(n15933), .A2(n15932), .ZN(n16092) );
  NAND2_X1 U17810 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15935) );
  NAND2_X1 U17811 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n15934) );
  AND3_X1 U17812 ( .A1(n15935), .A2(n16037), .A3(n15934), .ZN(n15939) );
  AOI22_X1 U17813 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U17814 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15937) );
  AOI22_X1 U17815 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15936) );
  NAND4_X1 U17816 ( .A1(n15939), .A2(n15938), .A3(n15937), .A4(n15936), .ZN(
        n15947) );
  NAND2_X1 U17817 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n15941) );
  NAND2_X1 U17818 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15940) );
  AND3_X1 U17819 ( .A1(n15941), .A2(n16001), .A3(n15940), .ZN(n15945) );
  AOI22_X1 U17820 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15944) );
  AOI22_X1 U17821 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15943) );
  AOI22_X1 U17822 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15942) );
  NAND4_X1 U17823 ( .A1(n15945), .A2(n15944), .A3(n15943), .A4(n15942), .ZN(
        n15946) );
  AND2_X1 U17824 ( .A1(n15947), .A2(n15946), .ZN(n15950) );
  NAND2_X1 U17825 ( .A1(n15948), .A2(n15950), .ZN(n15988) );
  OAI211_X1 U17826 ( .C1(n15948), .C2(n15950), .A(n15988), .B(n15990), .ZN(
        n15952) );
  INV_X1 U17827 ( .A(n15950), .ZN(n15951) );
  NOR2_X1 U17828 ( .A1(n16011), .A2(n15951), .ZN(n16086) );
  NAND2_X1 U17829 ( .A1(n16087), .A2(n16086), .ZN(n16085) );
  NAND2_X1 U17830 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15954) );
  NAND2_X1 U17831 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n15953) );
  AND3_X1 U17832 ( .A1(n15954), .A2(n16037), .A3(n15953), .ZN(n15958) );
  INV_X1 U17833 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n19443) );
  AOI22_X1 U17834 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15957) );
  AOI22_X1 U17835 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15956) );
  AOI22_X1 U17836 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15955) );
  NAND4_X1 U17837 ( .A1(n15958), .A2(n15957), .A3(n15956), .A4(n15955), .ZN(
        n15966) );
  NAND2_X1 U17838 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15960) );
  NAND2_X1 U17839 ( .A1(n16036), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n15959) );
  AND3_X1 U17840 ( .A1(n15960), .A2(n16001), .A3(n15959), .ZN(n15964) );
  AOI22_X1 U17841 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15963) );
  AOI22_X1 U17842 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U17843 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15961) );
  NAND4_X1 U17844 ( .A1(n15964), .A2(n15963), .A3(n15962), .A4(n15961), .ZN(
        n15965) );
  AND2_X1 U17845 ( .A1(n15966), .A2(n15965), .ZN(n15986) );
  XNOR2_X1 U17846 ( .A(n15988), .B(n15986), .ZN(n15967) );
  NAND2_X1 U17847 ( .A1(n15968), .A2(n15986), .ZN(n16080) );
  NOR2_X2 U17848 ( .A1(n16081), .A2(n16080), .ZN(n16079) );
  NOR2_X2 U17849 ( .A1(n16079), .A2(n15970), .ZN(n16010) );
  NAND2_X1 U17850 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15972) );
  NAND2_X1 U17851 ( .A1(n16036), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n15971) );
  AND3_X1 U17852 ( .A1(n15972), .A2(n16037), .A3(n15971), .ZN(n15977) );
  INV_X1 U17853 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19388) );
  AOI22_X1 U17854 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15976) );
  AOI22_X1 U17855 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15975) );
  AOI22_X1 U17856 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15973), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15974) );
  NAND4_X1 U17857 ( .A1(n15977), .A2(n15976), .A3(n15975), .A4(n15974), .ZN(
        n15985) );
  AOI22_X1 U17858 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U17859 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15979) );
  NAND2_X1 U17860 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15978) );
  AND3_X1 U17861 ( .A1(n16001), .A2(n15979), .A3(n15978), .ZN(n15982) );
  AOI22_X1 U17862 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15981) );
  AOI22_X1 U17863 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15980) );
  NAND4_X1 U17864 ( .A1(n15983), .A2(n15982), .A3(n15981), .A4(n15980), .ZN(
        n15984) );
  NAND2_X1 U17865 ( .A1(n15985), .A2(n15984), .ZN(n15993) );
  INV_X1 U17866 ( .A(n15993), .ZN(n15992) );
  INV_X1 U17867 ( .A(n15986), .ZN(n15987) );
  OR2_X1 U17868 ( .A1(n15988), .A2(n15987), .ZN(n15989) );
  INV_X1 U17869 ( .A(n15989), .ZN(n15991) );
  OR2_X1 U17870 ( .A1(n15989), .A2(n15993), .ZN(n16061) );
  OAI211_X1 U17871 ( .C1(n15992), .C2(n15991), .A(n15990), .B(n16061), .ZN(
        n16009) );
  NOR2_X1 U17872 ( .A1(n16011), .A2(n15993), .ZN(n16071) );
  NAND2_X1 U17873 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15995) );
  NAND2_X1 U17874 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n15994) );
  AND3_X1 U17875 ( .A1(n15995), .A2(n16037), .A3(n15994), .ZN(n15999) );
  AOI22_X1 U17876 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15998) );
  AOI22_X1 U17877 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U17878 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15996) );
  NAND4_X1 U17879 ( .A1(n15999), .A2(n15998), .A3(n15997), .A4(n15996), .ZN(
        n16008) );
  NAND2_X1 U17880 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n16002) );
  NAND2_X1 U17881 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n16000) );
  AND3_X1 U17882 ( .A1(n16002), .A2(n16001), .A3(n16000), .ZN(n16006) );
  AOI22_X1 U17883 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U17884 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16004) );
  AOI22_X1 U17885 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16003) );
  NAND4_X1 U17886 ( .A1(n16006), .A2(n16005), .A3(n16004), .A4(n16003), .ZN(
        n16007) );
  AND2_X1 U17887 ( .A1(n16008), .A2(n16007), .ZN(n16062) );
  INV_X1 U17888 ( .A(n16061), .ZN(n16012) );
  NAND3_X1 U17889 ( .A1(n16012), .A2(n16062), .A3(n16011), .ZN(n16053) );
  AOI22_X1 U17890 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U17891 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16013) );
  NAND2_X1 U17892 ( .A1(n16014), .A2(n16013), .ZN(n16028) );
  AOI21_X1 U17893 ( .B1(n10973), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n16037), .ZN(n16016) );
  AOI22_X1 U17894 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16015) );
  OAI211_X1 U17895 ( .C1(n11758), .C2(n16017), .A(n16016), .B(n16015), .ZN(
        n16027) );
  AOI22_X1 U17896 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U17897 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16020) );
  NAND2_X1 U17898 ( .A1(n16021), .A2(n16020), .ZN(n16026) );
  AOI22_X1 U17899 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16024) );
  NAND2_X1 U17900 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n16023) );
  NAND2_X1 U17901 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n16022) );
  NAND4_X1 U17902 ( .A1(n16024), .A2(n16037), .A3(n16023), .A4(n16022), .ZN(
        n16025) );
  OAI22_X1 U17903 ( .A1(n16028), .A2(n16027), .B1(n16026), .B2(n16025), .ZN(
        n16052) );
  AOI22_X1 U17904 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U17905 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16029) );
  NAND2_X1 U17906 ( .A1(n16030), .A2(n16029), .ZN(n16044) );
  INV_X1 U17907 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19033) );
  AOI21_X1 U17908 ( .B1(n10973), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n16037), .ZN(n16032) );
  AOI22_X1 U17909 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16031) );
  OAI211_X1 U17910 ( .C1(n10949), .C2(n19033), .A(n16032), .B(n16031), .ZN(
        n16043) );
  AOI22_X1 U17911 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16018), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16035) );
  AOI22_X1 U17912 ( .A1(n16019), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10950), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16034) );
  NAND2_X1 U17913 ( .A1(n16035), .A2(n16034), .ZN(n16042) );
  AOI22_X1 U17914 ( .A1(n15973), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16036), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U17915 ( .A1(n10973), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n16039) );
  NAND2_X1 U17916 ( .A1(n11825), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n16038) );
  NAND4_X1 U17917 ( .A1(n16040), .A2(n16039), .A3(n16038), .A4(n16037), .ZN(
        n16041) );
  OAI22_X1 U17918 ( .A1(n16044), .A2(n16043), .B1(n16042), .B2(n16041), .ZN(
        n16045) );
  NAND2_X1 U17919 ( .A1(n16046), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16050) );
  INV_X1 U17920 ( .A(n16047), .ZN(n16048) );
  NAND2_X1 U17921 ( .A1(n18383), .A2(n16112), .ZN(n16049) );
  OAI211_X1 U17922 ( .C1(n16124), .C2(n16115), .A(n16050), .B(n16049), .ZN(
        P2_U2857) );
  XNOR2_X1 U17923 ( .A(n16053), .B(n16052), .ZN(n16054) );
  XNOR2_X1 U17924 ( .A(n16051), .B(n16054), .ZN(n16132) );
  NOR2_X1 U17925 ( .A1(n16055), .A2(n16056), .ZN(n16057) );
  NOR2_X1 U17926 ( .A1(n16233), .A2(n16046), .ZN(n16059) );
  AOI21_X1 U17927 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16046), .A(n16059), .ZN(
        n16060) );
  OAI21_X1 U17928 ( .B1(n16132), .B2(n16115), .A(n16060), .ZN(P2_U2858) );
  NAND2_X1 U17929 ( .A1(n11004), .A2(n16061), .ZN(n16063) );
  XNOR2_X1 U17930 ( .A(n16063), .B(n16062), .ZN(n16140) );
  NOR2_X1 U17931 ( .A1(n16065), .A2(n16064), .ZN(n16066) );
  NOR2_X1 U17932 ( .A1(n16248), .A2(n16046), .ZN(n16067) );
  AOI21_X1 U17933 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16046), .A(n16067), .ZN(
        n16068) );
  OAI21_X1 U17934 ( .B1(n16140), .B2(n16115), .A(n16068), .ZN(P2_U2859) );
  NAND2_X1 U17935 ( .A1(n11004), .A2(n16069), .ZN(n16070) );
  XOR2_X1 U17936 ( .A(n16071), .B(n16070), .Z(n16146) );
  NOR2_X1 U17937 ( .A1(n16072), .A2(n16046), .ZN(n16073) );
  AOI21_X1 U17938 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16046), .A(n16073), .ZN(
        n16074) );
  OAI21_X1 U17939 ( .B1(n16146), .B2(n16115), .A(n16074), .ZN(P2_U2860) );
  NAND2_X1 U17940 ( .A1(n16075), .A2(n16076), .ZN(n16077) );
  NAND2_X1 U17941 ( .A1(n16078), .A2(n16077), .ZN(n18329) );
  AOI21_X1 U17942 ( .B1(n16081), .B2(n16080), .A(n16079), .ZN(n16153) );
  NAND2_X1 U17943 ( .A1(n16153), .A2(n16082), .ZN(n16084) );
  NAND2_X1 U17944 ( .A1(n16046), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16083) );
  OAI211_X1 U17945 ( .C1(n18329), .C2(n16046), .A(n16084), .B(n16083), .ZN(
        P2_U2861) );
  OAI21_X1 U17946 ( .B1(n16087), .B2(n16086), .A(n16085), .ZN(n16163) );
  INV_X1 U17947 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16089) );
  OAI21_X1 U17948 ( .B1(n16094), .B2(n16088), .A(n16075), .ZN(n16490) );
  MUX2_X1 U17949 ( .A(n16089), .B(n16490), .S(n16112), .Z(n16090) );
  OAI21_X1 U17950 ( .B1(n16163), .B2(n16115), .A(n16090), .ZN(P2_U2862) );
  OAI21_X1 U17951 ( .B1(n16093), .B2(n16092), .A(n16091), .ZN(n16172) );
  AOI21_X1 U17952 ( .B1(n16095), .B2(n16103), .A(n16094), .ZN(n18309) );
  INV_X1 U17953 ( .A(n18309), .ZN(n16508) );
  NOR2_X1 U17954 ( .A1(n16508), .A2(n16046), .ZN(n16096) );
  AOI21_X1 U17955 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16046), .A(n16096), .ZN(
        n16097) );
  OAI21_X1 U17956 ( .B1(n16172), .B2(n16115), .A(n16097), .ZN(P2_U2863) );
  XNOR2_X1 U17957 ( .A(n16098), .B(n16099), .ZN(n16178) );
  INV_X1 U17958 ( .A(n16100), .ZN(n16111) );
  NAND2_X1 U17959 ( .A1(n16111), .A2(n16101), .ZN(n16102) );
  NAND2_X1 U17960 ( .A1(n16103), .A2(n16102), .ZN(n18293) );
  NOR2_X1 U17961 ( .A1(n18293), .A2(n16046), .ZN(n16104) );
  AOI21_X1 U17962 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16046), .A(n16104), .ZN(
        n16105) );
  OAI21_X1 U17963 ( .B1(n16178), .B2(n16115), .A(n16105), .ZN(P2_U2864) );
  INV_X1 U17964 ( .A(n16098), .ZN(n16107) );
  OAI21_X1 U17965 ( .B1(n15864), .B2(n16108), .A(n16107), .ZN(n16185) );
  INV_X1 U17966 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16113) );
  NAND2_X1 U17967 ( .A1(n14830), .A2(n16109), .ZN(n16110) );
  NAND2_X1 U17968 ( .A1(n16111), .A2(n16110), .ZN(n18284) );
  MUX2_X1 U17969 ( .A(n16113), .B(n18284), .S(n16112), .Z(n16114) );
  OAI21_X1 U17970 ( .B1(n16185), .B2(n16115), .A(n16114), .ZN(P2_U2865) );
  INV_X1 U17971 ( .A(n19002), .ZN(n16122) );
  INV_X1 U17972 ( .A(n16116), .ZN(n16117) );
  NAND2_X1 U17973 ( .A1(n16125), .A2(n16117), .ZN(n16118) );
  NAND2_X1 U17974 ( .A1(n16119), .A2(n16118), .ZN(n16438) );
  OAI22_X1 U17975 ( .A1(n16438), .A2(n19467), .B1(n19278), .B2(n13906), .ZN(
        n16121) );
  INV_X1 U17976 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n22151) );
  INV_X1 U17977 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18647) );
  OAI22_X1 U17978 ( .A1(n19463), .A2(n22151), .B1(n19474), .B2(n18647), .ZN(
        n16120) );
  OAI21_X1 U17979 ( .B1(n16124), .B2(n19468), .A(n16123), .ZN(P2_U2889) );
  INV_X1 U17980 ( .A(n19005), .ZN(n16129) );
  OAI21_X1 U17981 ( .B1(n16134), .B2(n16126), .A(n16125), .ZN(n18366) );
  OAI22_X1 U17982 ( .A1(n19467), .A2(n18366), .B1(n19278), .B2(n16127), .ZN(
        n16128) );
  AOI21_X1 U17983 ( .B1(n16211), .B2(n16129), .A(n16128), .ZN(n16131) );
  AOI22_X1 U17984 ( .A1(n18995), .A2(BUF2_REG_29__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16130) );
  OAI211_X1 U17985 ( .C1(n16132), .C2(n19468), .A(n16131), .B(n16130), .ZN(
        P2_U2890) );
  INV_X1 U17986 ( .A(n19008), .ZN(n16137) );
  INV_X1 U17987 ( .A(n15265), .ZN(n16135) );
  AOI21_X1 U17988 ( .B1(n11343), .B2(n16135), .A(n16134), .ZN(n18356) );
  INV_X1 U17989 ( .A(n18356), .ZN(n16471) );
  OAI22_X1 U17990 ( .A1(n19467), .A2(n16471), .B1(n19278), .B2(n13886), .ZN(
        n16136) );
  AOI21_X1 U17991 ( .B1(n16211), .B2(n16137), .A(n16136), .ZN(n16139) );
  AOI22_X1 U17992 ( .A1(n18995), .A2(BUF2_REG_28__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16138) );
  OAI211_X1 U17993 ( .C1(n16140), .C2(n19468), .A(n16139), .B(n16138), .ZN(
        P2_U2891) );
  INV_X1 U17994 ( .A(n19011), .ZN(n16143) );
  OAI22_X1 U17995 ( .A1(n19467), .A2(n18353), .B1(n19278), .B2(n16141), .ZN(
        n16142) );
  AOI21_X1 U17996 ( .B1(n16211), .B2(n16143), .A(n16142), .ZN(n16145) );
  AOI22_X1 U17997 ( .A1(n18995), .A2(BUF2_REG_27__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16144) );
  OAI211_X1 U17998 ( .C1(n16146), .C2(n19468), .A(n16145), .B(n16144), .ZN(
        P2_U2892) );
  AOI22_X1 U17999 ( .A1(n18995), .A2(BUF2_REG_26__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16151) );
  AND2_X1 U18000 ( .A1(n16155), .A2(n16147), .ZN(n16148) );
  NOR2_X1 U18001 ( .A1(n16149), .A2(n16148), .ZN(n18330) );
  AOI22_X1 U18002 ( .A1(n19345), .A2(n18330), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19465), .ZN(n16150) );
  OAI211_X1 U18003 ( .C1(n19014), .C2(n19462), .A(n16151), .B(n16150), .ZN(
        n16152) );
  AOI21_X1 U18004 ( .B1(n16153), .B2(n19346), .A(n16152), .ZN(n16154) );
  INV_X1 U18005 ( .A(n16154), .ZN(P2_U2893) );
  INV_X1 U18006 ( .A(n19017), .ZN(n16160) );
  INV_X1 U18007 ( .A(n16167), .ZN(n16157) );
  OAI21_X1 U18008 ( .B1(n16157), .B2(n16156), .A(n16155), .ZN(n16491) );
  OAI22_X1 U18009 ( .A1(n16491), .A2(n19467), .B1(n19278), .B2(n16158), .ZN(
        n16159) );
  AOI21_X1 U18010 ( .B1(n16211), .B2(n16160), .A(n16159), .ZN(n16162) );
  AOI22_X1 U18011 ( .A1(n18995), .A2(BUF2_REG_25__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16161) );
  OAI211_X1 U18012 ( .C1(n16163), .C2(n19468), .A(n16162), .B(n16161), .ZN(
        P2_U2894) );
  INV_X1 U18013 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n19601) );
  NOR2_X1 U18014 ( .A1(n19474), .A2(n19601), .ZN(n16170) );
  NAND2_X1 U18015 ( .A1(n16164), .A2(n16165), .ZN(n16166) );
  AND2_X1 U18016 ( .A1(n16167), .A2(n16166), .ZN(n18308) );
  AOI22_X1 U18017 ( .A1(n19345), .A2(n18308), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19465), .ZN(n16168) );
  OAI21_X1 U18018 ( .B1(n19462), .B2(n19020), .A(n16168), .ZN(n16169) );
  AOI211_X1 U18019 ( .C1(n18996), .C2(BUF1_REG_24__SCAN_IN), .A(n16170), .B(
        n16169), .ZN(n16171) );
  OAI21_X1 U18020 ( .B1(n16172), .B2(n19468), .A(n16171), .ZN(P2_U2895) );
  INV_X1 U18021 ( .A(n19029), .ZN(n16175) );
  OAI21_X1 U18022 ( .B1(n16173), .B2(n10991), .A(n16164), .ZN(n18306) );
  OAI22_X1 U18023 ( .A1(n18306), .A2(n19467), .B1(n19278), .B2(n13899), .ZN(
        n16174) );
  AOI21_X1 U18024 ( .B1(n16211), .B2(n16175), .A(n16174), .ZN(n16177) );
  AOI22_X1 U18025 ( .A1(n18995), .A2(BUF2_REG_23__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16176) );
  OAI211_X1 U18026 ( .C1(n16178), .C2(n19468), .A(n16177), .B(n16176), .ZN(
        P2_U2896) );
  INV_X1 U18027 ( .A(n19230), .ZN(n16182) );
  XNOR2_X1 U18028 ( .A(n16180), .B(n16179), .ZN(n18282) );
  OAI22_X1 U18029 ( .A1(n18282), .A2(n19467), .B1(n19278), .B2(n13888), .ZN(
        n16181) );
  AOI21_X1 U18030 ( .B1(n16211), .B2(n16182), .A(n16181), .ZN(n16184) );
  AOI22_X1 U18031 ( .A1(n18995), .A2(BUF2_REG_22__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16183) );
  OAI211_X1 U18032 ( .C1(n16185), .C2(n19468), .A(n16184), .B(n16183), .ZN(
        P2_U2897) );
  INV_X1 U18033 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16186) );
  OR2_X1 U18034 ( .A1(n16187), .A2(n16186), .ZN(n16189) );
  NAND2_X1 U18035 ( .A1(n16187), .A2(BUF2_REG_5__SCAN_IN), .ZN(n16188) );
  AND2_X1 U18036 ( .A1(n16189), .A2(n16188), .ZN(n19290) );
  INV_X1 U18037 ( .A(n19290), .ZN(n16192) );
  OAI21_X1 U18038 ( .B1(n16562), .B2(n16190), .A(n16179), .ZN(n18271) );
  OAI22_X1 U18039 ( .A1(n18271), .A2(n19467), .B1(n19278), .B2(n13891), .ZN(
        n16191) );
  AOI21_X1 U18040 ( .B1(n16211), .B2(n16192), .A(n16191), .ZN(n16194) );
  AOI22_X1 U18041 ( .A1(n18995), .A2(BUF2_REG_21__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16193) );
  OAI211_X1 U18042 ( .C1(n16195), .C2(n19468), .A(n16194), .B(n16193), .ZN(
        P2_U2898) );
  INV_X1 U18043 ( .A(n16196), .ZN(n16204) );
  INV_X1 U18044 ( .A(n16585), .ZN(n16199) );
  INV_X1 U18045 ( .A(n16197), .ZN(n16198) );
  OAI21_X1 U18046 ( .B1(n16199), .B2(n16198), .A(n16560), .ZN(n18252) );
  OAI22_X1 U18047 ( .A1(n18252), .A2(n19467), .B1(n19278), .B2(n13903), .ZN(
        n16200) );
  AOI21_X1 U18048 ( .B1(n16211), .B2(n16201), .A(n16200), .ZN(n16203) );
  AOI22_X1 U18049 ( .A1(n18995), .A2(BUF2_REG_19__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16202) );
  OAI211_X1 U18050 ( .C1(n16204), .C2(n19468), .A(n16203), .B(n16202), .ZN(
        P2_U2900) );
  INV_X1 U18051 ( .A(n16205), .ZN(n16206) );
  OAI21_X1 U18052 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n18229) );
  OAI22_X1 U18053 ( .A1(n18229), .A2(n19467), .B1(n19278), .B2(n13719), .ZN(
        n16209) );
  AOI21_X1 U18054 ( .B1(n16211), .B2(n16210), .A(n16209), .ZN(n16213) );
  AOI22_X1 U18055 ( .A1(n18995), .A2(BUF2_REG_17__SCAN_IN), .B1(n18996), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16212) );
  OAI211_X1 U18056 ( .C1(n16214), .C2(n19468), .A(n16213), .B(n16212), .ZN(
        P2_U2902) );
  NAND2_X1 U18057 ( .A1(n16215), .A2(n16230), .ZN(n16220) );
  INV_X1 U18058 ( .A(n16216), .ZN(n16217) );
  NOR2_X1 U18059 ( .A1(n16218), .A2(n16217), .ZN(n16219) );
  XNOR2_X1 U18060 ( .A(n16220), .B(n16219), .ZN(n16454) );
  XOR2_X1 U18061 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n16238), .Z(
        n16452) );
  XNOR2_X1 U18062 ( .A(n16221), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18387) );
  NOR2_X1 U18063 ( .A1(n18240), .A2(n16222), .ZN(n16443) );
  AOI21_X1 U18064 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16443), .ZN(n16223) );
  OAI21_X1 U18065 ( .B1(n18387), .B2(n17042), .A(n16223), .ZN(n16224) );
  INV_X1 U18066 ( .A(n16224), .ZN(n16225) );
  AOI21_X1 U18067 ( .B1(n16452), .B2(n17035), .A(n16227), .ZN(n16228) );
  OAI21_X1 U18068 ( .B1(n16454), .B2(n17014), .A(n16228), .ZN(P2_U2984) );
  NAND2_X1 U18069 ( .A1(n16230), .A2(n16229), .ZN(n16232) );
  XOR2_X1 U18070 ( .A(n16232), .B(n16231), .Z(n16467) );
  AOI21_X1 U18071 ( .B1(n16235), .B2(n16247), .A(n16221), .ZN(n18370) );
  NAND2_X1 U18072 ( .A1(n18368), .A2(n17021), .ZN(n16234) );
  NAND2_X1 U18073 ( .A1(n18072), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16461) );
  OAI211_X1 U18074 ( .C1(n17018), .C2(n16235), .A(n16234), .B(n16461), .ZN(
        n16236) );
  AOI21_X1 U18075 ( .B1(n17005), .B2(n18370), .A(n16236), .ZN(n16241) );
  AOI21_X1 U18076 ( .B1(n16237), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16239) );
  NOR2_X1 U18077 ( .A1(n16239), .A2(n16238), .ZN(n16464) );
  NAND2_X1 U18078 ( .A1(n16464), .A2(n17035), .ZN(n16240) );
  OAI211_X1 U18079 ( .C1(n16467), .C2(n17014), .A(n16241), .B(n16240), .ZN(
        P2_U2985) );
  XNOR2_X1 U18080 ( .A(n16243), .B(n16474), .ZN(n16244) );
  XNOR2_X1 U18081 ( .A(n16245), .B(n16244), .ZN(n16479) );
  XNOR2_X1 U18082 ( .A(n16246), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16477) );
  OAI21_X1 U18083 ( .B1(n16255), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16247), .ZN(n18359) );
  NAND2_X1 U18084 ( .A1(n18357), .A2(n17021), .ZN(n16251) );
  NOR2_X1 U18085 ( .A1(n18240), .A2(n16249), .ZN(n16468) );
  AOI21_X1 U18086 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16468), .ZN(n16250) );
  OAI211_X1 U18087 ( .C1(n18359), .C2(n17042), .A(n16251), .B(n16250), .ZN(
        n16252) );
  AOI21_X1 U18088 ( .B1(n16477), .B2(n17035), .A(n16252), .ZN(n16253) );
  OAI21_X1 U18089 ( .B1(n16479), .B2(n17014), .A(n16253), .ZN(P2_U2986) );
  NOR2_X1 U18090 ( .A1(n16273), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16254) );
  OR2_X1 U18091 ( .A1(n16255), .A2(n16254), .ZN(n18349) );
  INV_X1 U18092 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18341) );
  NOR2_X1 U18093 ( .A1(n17018), .A2(n18341), .ZN(n16256) );
  AOI211_X1 U18094 ( .C1(n18347), .C2(n17021), .A(n16257), .B(n16256), .ZN(
        n16258) );
  OAI21_X1 U18095 ( .B1(n17042), .B2(n18349), .A(n16258), .ZN(n16259) );
  AOI21_X1 U18096 ( .B1(n16260), .B2(n17035), .A(n16259), .ZN(n16261) );
  OAI21_X1 U18097 ( .B1(n16262), .B2(n17014), .A(n16261), .ZN(P2_U2987) );
  INV_X1 U18098 ( .A(n16263), .ZN(n16268) );
  AOI21_X1 U18099 ( .B1(n16264), .B2(n16280), .A(n16282), .ZN(n16266) );
  MUX2_X1 U18100 ( .A(n16280), .B(n16266), .S(n16265), .Z(n16267) );
  NAND2_X1 U18101 ( .A1(n16268), .A2(n16267), .ZN(n16489) );
  AOI21_X1 U18102 ( .B1(n10968), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16271) );
  INV_X1 U18103 ( .A(n16269), .ZN(n16270) );
  NOR2_X1 U18104 ( .A1(n16271), .A2(n16270), .ZN(n16487) );
  AND2_X1 U18105 ( .A1(n16284), .A2(n16272), .ZN(n16274) );
  OR2_X1 U18106 ( .A1(n16274), .A2(n16273), .ZN(n18333) );
  NOR2_X1 U18107 ( .A1(n18475), .A2(n16275), .ZN(n16483) );
  NOR2_X1 U18108 ( .A1(n18329), .A2(n17038), .ZN(n16276) );
  AOI211_X1 U18109 ( .C1(n17031), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16483), .B(n16276), .ZN(n16277) );
  OAI21_X1 U18110 ( .B1(n17042), .B2(n18333), .A(n16277), .ZN(n16278) );
  AOI21_X1 U18111 ( .B1(n16487), .B2(n17035), .A(n16278), .ZN(n16279) );
  OAI21_X1 U18112 ( .B1(n16489), .B2(n17014), .A(n16279), .ZN(P2_U2988) );
  XNOR2_X1 U18113 ( .A(n10968), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16502) );
  INV_X1 U18114 ( .A(n16280), .ZN(n16281) );
  NOR2_X1 U18115 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  XNOR2_X1 U18116 ( .A(n16264), .B(n16283), .ZN(n16500) );
  INV_X1 U18117 ( .A(n16284), .ZN(n16285) );
  AOI21_X1 U18118 ( .B1(n16286), .B2(n16295), .A(n16285), .ZN(n18321) );
  NAND2_X1 U18119 ( .A1(n18321), .A2(n17005), .ZN(n16288) );
  NOR2_X1 U18120 ( .A1(n18240), .A2(n17120), .ZN(n16494) );
  AOI21_X1 U18121 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16494), .ZN(n16287) );
  OAI211_X1 U18122 ( .C1(n17038), .C2(n16490), .A(n16288), .B(n16287), .ZN(
        n16289) );
  AOI21_X1 U18123 ( .B1(n16500), .B2(n17032), .A(n16289), .ZN(n16290) );
  OAI21_X1 U18124 ( .B1(n17024), .B2(n16502), .A(n16290), .ZN(P2_U2989) );
  XNOR2_X1 U18125 ( .A(n16292), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16293) );
  XNOR2_X1 U18126 ( .A(n16291), .B(n16293), .ZN(n16512) );
  INV_X1 U18127 ( .A(n16306), .ZN(n16294) );
  AOI21_X1 U18128 ( .B1(n11228), .B2(n16294), .A(n10968), .ZN(n16510) );
  OAI21_X1 U18129 ( .B1(n11039), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16295), .ZN(n18311) );
  NAND2_X1 U18130 ( .A1(n18309), .A2(n17021), .ZN(n16297) );
  NOR2_X1 U18131 ( .A1(n18240), .A2(n17119), .ZN(n16503) );
  AOI21_X1 U18132 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16503), .ZN(n16296) );
  OAI211_X1 U18133 ( .C1(n18311), .C2(n17042), .A(n16297), .B(n16296), .ZN(
        n16298) );
  AOI21_X1 U18134 ( .B1(n16510), .B2(n17035), .A(n16298), .ZN(n16299) );
  OAI21_X1 U18135 ( .B1(n16512), .B2(n17014), .A(n16299), .ZN(P2_U2990) );
  INV_X1 U18136 ( .A(n16301), .ZN(n16303) );
  NAND2_X1 U18137 ( .A1(n16303), .A2(n16302), .ZN(n16304) );
  XNOR2_X1 U18138 ( .A(n16300), .B(n16304), .ZN(n16523) );
  AOI21_X1 U18139 ( .B1(n16515), .B2(n16305), .A(n16306), .ZN(n16513) );
  NAND2_X1 U18140 ( .A1(n16513), .A2(n17035), .ZN(n16310) );
  AOI21_X1 U18141 ( .B1(n17029), .B2(n18295), .A(n11039), .ZN(n18302) );
  NOR2_X1 U18142 ( .A1(n18240), .A2(n18294), .ZN(n16517) );
  AOI21_X1 U18143 ( .B1(n17031), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16517), .ZN(n16307) );
  OAI21_X1 U18144 ( .B1(n18293), .B2(n17038), .A(n16307), .ZN(n16308) );
  AOI21_X1 U18145 ( .B1(n17005), .B2(n18302), .A(n16308), .ZN(n16309) );
  OAI211_X1 U18146 ( .C1(n17014), .C2(n16523), .A(n16310), .B(n16309), .ZN(
        P2_U2991) );
  AND2_X1 U18147 ( .A1(n16986), .A2(n16989), .ZN(n16424) );
  AND2_X1 U18148 ( .A1(n16424), .A2(n16420), .ZN(n16312) );
  INV_X1 U18149 ( .A(n16998), .ZN(n16313) );
  INV_X1 U18150 ( .A(n16314), .ZN(n16315) );
  NAND2_X1 U18151 ( .A1(n16317), .A2(n16316), .ZN(n16395) );
  INV_X1 U18152 ( .A(n16377), .ZN(n16319) );
  NAND2_X1 U18153 ( .A1(n16321), .A2(n16349), .ZN(n16323) );
  NOR2_X1 U18154 ( .A1(n16324), .A2(n16325), .ZN(n16327) );
  XNOR2_X1 U18155 ( .A(n16325), .B(n16324), .ZN(n16341) );
  NOR2_X1 U18156 ( .A1(n16341), .A2(n16558), .ZN(n16326) );
  NOR2_X1 U18157 ( .A1(n16329), .A2(n16328), .ZN(n16330) );
  XOR2_X1 U18158 ( .A(n16331), .B(n16330), .Z(n16547) );
  NAND2_X1 U18159 ( .A1(n16432), .A2(n16536), .ZN(n16340) );
  NAND2_X1 U18160 ( .A1(n16340), .A2(n16537), .ZN(n16332) );
  NAND2_X1 U18161 ( .A1(n16332), .A2(n16532), .ZN(n16542) );
  OAI22_X1 U18162 ( .A1(n16334), .A2(n17018), .B1(n17118), .B2(n18475), .ZN(
        n16333) );
  AOI21_X1 U18163 ( .B1(n18273), .B2(n17021), .A(n16333), .ZN(n16336) );
  AOI21_X1 U18164 ( .B1(n16334), .B2(n16344), .A(n17030), .ZN(n18274) );
  NAND2_X1 U18165 ( .A1(n18274), .A2(n17005), .ZN(n16335) );
  OAI211_X1 U18166 ( .C1(n16542), .C2(n17024), .A(n16336), .B(n16335), .ZN(
        n16337) );
  INV_X1 U18167 ( .A(n16337), .ZN(n16338) );
  OAI21_X1 U18168 ( .B1(n16547), .B2(n17014), .A(n16338), .ZN(P2_U2993) );
  NOR2_X2 U18169 ( .A1(n16380), .A2(n16563), .ZN(n16355) );
  OAI21_X1 U18170 ( .B1(n16355), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16340), .ZN(n16572) );
  XNOR2_X1 U18171 ( .A(n16341), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16570) );
  NOR2_X1 U18172 ( .A1(n18240), .A2(n16342), .ZN(n16565) );
  OR2_X1 U18173 ( .A1(n11041), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16343) );
  NAND2_X1 U18174 ( .A1(n16344), .A2(n16343), .ZN(n18253) );
  NOR2_X1 U18175 ( .A1(n17042), .A2(n18253), .ZN(n16345) );
  AOI211_X1 U18176 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n17031), .A(
        n16565), .B(n16345), .ZN(n16346) );
  OAI21_X1 U18177 ( .B1(n17038), .B2(n18269), .A(n16346), .ZN(n16347) );
  AOI21_X1 U18178 ( .B1(n16570), .B2(n17032), .A(n16347), .ZN(n16348) );
  OAI21_X1 U18179 ( .B1(n16572), .B2(n17024), .A(n16348), .ZN(P2_U2994) );
  OAI21_X1 U18180 ( .B1(n16351), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16352), .ZN(n16364) );
  OR2_X1 U18181 ( .A1(n16364), .A2(n16363), .ZN(n16366) );
  NAND2_X1 U18182 ( .A1(n16366), .A2(n16352), .ZN(n16353) );
  INV_X1 U18183 ( .A(n16380), .ZN(n16354) );
  AOI21_X1 U18184 ( .B1(n16354), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16356) );
  NOR2_X2 U18185 ( .A1(n16356), .A2(n16355), .ZN(n16573) );
  NAND2_X1 U18186 ( .A1(n16573), .A2(n17035), .ZN(n16362) );
  AOI21_X1 U18187 ( .B1(n16359), .B2(n16367), .A(n11041), .ZN(n18254) );
  NAND2_X1 U18188 ( .A1(n17005), .A2(n18254), .ZN(n16358) );
  NAND2_X1 U18189 ( .A1(n18072), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16575) );
  OAI211_X1 U18190 ( .C1(n16359), .C2(n17018), .A(n16358), .B(n16575), .ZN(
        n16360) );
  AOI21_X1 U18191 ( .B1(n18249), .B2(n17021), .A(n16360), .ZN(n16361) );
  NAND2_X1 U18192 ( .A1(n16364), .A2(n16363), .ZN(n16365) );
  NAND2_X1 U18193 ( .A1(n16366), .A2(n16365), .ZN(n16594) );
  XNOR2_X1 U18194 ( .A(n16380), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16582) );
  NAND2_X1 U18195 ( .A1(n16582), .A2(n17035), .ZN(n16373) );
  INV_X1 U18196 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16370) );
  OAI21_X1 U18197 ( .B1(n16385), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16367), .ZN(n16368) );
  INV_X1 U18198 ( .A(n16368), .ZN(n18245) );
  NAND2_X1 U18199 ( .A1(n17005), .A2(n18245), .ZN(n16369) );
  OR2_X1 U18200 ( .A1(n18240), .A2(n17117), .ZN(n16586) );
  OAI211_X1 U18201 ( .C1(n16370), .C2(n17018), .A(n16369), .B(n16586), .ZN(
        n16371) );
  AOI21_X1 U18202 ( .B1(n17021), .B2(n18235), .A(n16371), .ZN(n16372) );
  OAI211_X1 U18203 ( .C1(n16594), .C2(n17014), .A(n16373), .B(n16372), .ZN(
        P2_U2996) );
  NAND2_X1 U18204 ( .A1(n16374), .A2(n16375), .ZN(n16379) );
  NAND2_X1 U18205 ( .A1(n16377), .A2(n16376), .ZN(n16378) );
  XNOR2_X1 U18206 ( .A(n16379), .B(n16378), .ZN(n16606) );
  INV_X1 U18207 ( .A(n16606), .ZN(n16390) );
  INV_X1 U18208 ( .A(n16598), .ZN(n16381) );
  OAI211_X1 U18209 ( .C1(n16381), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17035), .B(n16380), .ZN(n16389) );
  INV_X1 U18210 ( .A(n16382), .ZN(n18222) );
  NOR2_X1 U18211 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16383), .ZN(
        n16384) );
  NOR2_X1 U18212 ( .A1(n16385), .A2(n16384), .ZN(n18216) );
  INV_X1 U18213 ( .A(n18216), .ZN(n18225) );
  NAND2_X1 U18214 ( .A1(n18072), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16599) );
  NAND2_X1 U18215 ( .A1(n17031), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16386) );
  OAI211_X1 U18216 ( .C1(n17042), .C2(n18225), .A(n16599), .B(n16386), .ZN(
        n16387) );
  AOI21_X1 U18217 ( .B1(n17021), .B2(n18222), .A(n16387), .ZN(n16388) );
  OAI211_X1 U18218 ( .C1(n16390), .C2(n17014), .A(n16389), .B(n16388), .ZN(
        P2_U2997) );
  OAI211_X1 U18219 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16400), .A(
        n16598), .B(n17035), .ZN(n16398) );
  INV_X1 U18220 ( .A(n18210), .ZN(n16616) );
  OAI21_X1 U18221 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16401), .A(
        n16391), .ZN(n18205) );
  AOI22_X1 U18222 ( .A1(n17031), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n16539), .ZN(n16392) );
  OAI21_X1 U18223 ( .B1(n17042), .B2(n18205), .A(n16392), .ZN(n16393) );
  AOI21_X1 U18224 ( .B1(n17021), .B2(n16616), .A(n16393), .ZN(n16397) );
  OR2_X1 U18225 ( .A1(n16395), .A2(n16394), .ZN(n16614) );
  NAND3_X1 U18226 ( .A1(n16614), .A2(n17032), .A3(n16374), .ZN(n16396) );
  NAND3_X1 U18227 ( .A1(n16398), .A2(n16397), .A3(n16396), .ZN(P2_U2998) );
  INV_X1 U18228 ( .A(n16400), .ZN(n16612) );
  OAI21_X1 U18229 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16399), .A(
        n16612), .ZN(n16636) );
  AOI21_X1 U18230 ( .B1(n17019), .B2(n16403), .A(n16401), .ZN(n18192) );
  NAND2_X1 U18231 ( .A1(n17005), .A2(n18192), .ZN(n16402) );
  OR2_X1 U18232 ( .A1(n18240), .A2(n18191), .ZN(n16624) );
  OAI211_X1 U18233 ( .C1(n16403), .C2(n17018), .A(n16402), .B(n16624), .ZN(
        n16414) );
  NAND2_X1 U18234 ( .A1(n16405), .A2(n16404), .ZN(n16412) );
  NAND2_X1 U18235 ( .A1(n16406), .A2(n16999), .ZN(n17012) );
  AND2_X1 U18236 ( .A1(n16638), .A2(n16407), .ZN(n17011) );
  NAND2_X1 U18237 ( .A1(n17012), .A2(n17011), .ZN(n17010) );
  NAND2_X1 U18238 ( .A1(n16409), .A2(n16408), .ZN(n16639) );
  AOI21_X1 U18239 ( .B1(n17010), .B2(n16638), .A(n16639), .ZN(n16641) );
  INV_X1 U18240 ( .A(n16409), .ZN(n16410) );
  NOR2_X1 U18241 ( .A1(n16641), .A2(n16410), .ZN(n16411) );
  XOR2_X1 U18242 ( .A(n16412), .B(n16411), .Z(n16631) );
  NOR2_X1 U18243 ( .A1(n16631), .A2(n17014), .ZN(n16413) );
  AOI211_X1 U18244 ( .C1(n17021), .C2(n18197), .A(n16414), .B(n16413), .ZN(
        n16415) );
  OAI21_X1 U18245 ( .B1(n17024), .B2(n16636), .A(n16415), .ZN(P2_U2999) );
  INV_X1 U18246 ( .A(n16416), .ZN(n16993) );
  OAI21_X1 U18247 ( .B1(n16993), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17007), .ZN(n16663) );
  NOR2_X1 U18248 ( .A1(n18475), .A2(n16417), .ZN(n16656) );
  AOI21_X1 U18249 ( .B1(n18140), .B2(n16984), .A(n11023), .ZN(n16418) );
  INV_X1 U18250 ( .A(n16418), .ZN(n18154) );
  OAI22_X1 U18251 ( .A1(n18140), .A2(n17018), .B1(n17042), .B2(n18154), .ZN(
        n16419) );
  AOI211_X1 U18252 ( .C1(n11379), .C2(n17021), .A(n16656), .B(n16419), .ZN(
        n16428) );
  INV_X1 U18253 ( .A(n16420), .ZN(n16421) );
  NOR2_X1 U18254 ( .A1(n16422), .A2(n16421), .ZN(n16426) );
  NAND2_X1 U18255 ( .A1(n16423), .A2(n16424), .ZN(n16425) );
  XOR2_X1 U18256 ( .A(n16426), .B(n16425), .Z(n16661) );
  NAND2_X1 U18257 ( .A1(n16661), .A2(n17032), .ZN(n16427) );
  OAI211_X1 U18258 ( .C1(n16663), .C2(n17024), .A(n16428), .B(n16427), .ZN(
        P2_U3003) );
  NAND2_X1 U18259 ( .A1(n16989), .A2(n16429), .ZN(n16431) );
  XOR2_X1 U18260 ( .A(n16431), .B(n16430), .Z(n16674) );
  INV_X1 U18261 ( .A(n16432), .ZN(n16601) );
  NAND2_X1 U18262 ( .A1(n16601), .A2(n16668), .ZN(n16664) );
  NAND3_X1 U18263 ( .A1(n16664), .A2(n17035), .A3(n16994), .ZN(n16437) );
  OAI21_X1 U18264 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16974), .A(
        n16433), .ZN(n18132) );
  OAI22_X1 U18265 ( .A1(n11174), .A2(n17018), .B1(n17042), .B2(n18132), .ZN(
        n16435) );
  NOR2_X1 U18266 ( .A1(n18124), .A2(n17038), .ZN(n16434) );
  AOI211_X1 U18267 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n16539), .A(n16435), .B(
        n16434), .ZN(n16436) );
  OAI211_X1 U18268 ( .C1(n17014), .C2(n16674), .A(n16437), .B(n16436), .ZN(
        P2_U3005) );
  NAND2_X1 U18269 ( .A1(n18383), .A2(n18500), .ZN(n16450) );
  INV_X1 U18270 ( .A(n16438), .ZN(n18382) );
  INV_X1 U18271 ( .A(n16439), .ZN(n16440) );
  NOR3_X1 U18272 ( .A1(n16457), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16440), .ZN(n16447) );
  OR2_X1 U18273 ( .A1(n16442), .A2(n16441), .ZN(n16445) );
  INV_X1 U18274 ( .A(n16443), .ZN(n16444) );
  NAND2_X1 U18275 ( .A1(n16445), .A2(n16444), .ZN(n16446) );
  AOI21_X1 U18276 ( .B1(n16452), .B2(n18481), .A(n16451), .ZN(n16453) );
  OAI21_X1 U18277 ( .B1(n16454), .B2(n18450), .A(n16453), .ZN(P2_U3016) );
  AOI21_X1 U18278 ( .B1(n15190), .B2(n18460), .A(n16455), .ZN(n16475) );
  NAND2_X1 U18279 ( .A1(n16474), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16456) );
  OR2_X1 U18280 ( .A1(n16457), .A2(n16456), .ZN(n16469) );
  AOI21_X1 U18281 ( .B1(n16475), .B2(n16469), .A(n16458), .ZN(n16463) );
  INV_X1 U18282 ( .A(n16457), .ZN(n16459) );
  NAND4_X1 U18283 ( .A1(n16459), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n16458), .ZN(n16460) );
  OAI211_X1 U18284 ( .C1(n18490), .C2(n18366), .A(n16461), .B(n16460), .ZN(
        n16462) );
  AOI211_X1 U18285 ( .C1(n18368), .C2(n18500), .A(n16463), .B(n16462), .ZN(
        n16466) );
  NAND2_X1 U18286 ( .A1(n16464), .A2(n18481), .ZN(n16465) );
  OAI211_X1 U18287 ( .C1(n16467), .C2(n18450), .A(n16466), .B(n16465), .ZN(
        P2_U3017) );
  INV_X1 U18288 ( .A(n16468), .ZN(n16470) );
  OAI211_X1 U18289 ( .C1(n18490), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        n16472) );
  AOI21_X1 U18290 ( .B1(n18357), .B2(n18500), .A(n16472), .ZN(n16473) );
  OAI21_X1 U18291 ( .B1(n16475), .B2(n16474), .A(n16473), .ZN(n16476) );
  AOI21_X1 U18292 ( .B1(n16477), .B2(n18481), .A(n16476), .ZN(n16478) );
  OAI21_X1 U18293 ( .B1(n16479), .B2(n18450), .A(n16478), .ZN(P2_U3018) );
  INV_X1 U18294 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16480) );
  NOR2_X1 U18295 ( .A1(n16498), .A2(n16480), .ZN(n16486) );
  XNOR2_X1 U18296 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16481) );
  NOR2_X1 U18297 ( .A1(n16492), .A2(n16481), .ZN(n16482) );
  AOI211_X1 U18298 ( .C1(n18466), .C2(n18330), .A(n16483), .B(n16482), .ZN(
        n16484) );
  OAI21_X1 U18299 ( .B1(n18329), .B2(n16567), .A(n16484), .ZN(n16485) );
  AOI211_X1 U18300 ( .C1(n16487), .C2(n18481), .A(n16486), .B(n16485), .ZN(
        n16488) );
  OAI21_X1 U18301 ( .B1(n16489), .B2(n18450), .A(n16488), .ZN(P2_U3020) );
  INV_X1 U18302 ( .A(n16490), .ZN(n18319) );
  NAND2_X1 U18303 ( .A1(n18319), .A2(n18500), .ZN(n16496) );
  INV_X1 U18304 ( .A(n16491), .ZN(n18318) );
  NOR2_X1 U18305 ( .A1(n16492), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16493) );
  AOI211_X1 U18306 ( .C1(n18466), .C2(n18318), .A(n16494), .B(n16493), .ZN(
        n16495) );
  OAI211_X1 U18307 ( .C1(n16498), .C2(n16497), .A(n16496), .B(n16495), .ZN(
        n16499) );
  AOI21_X1 U18308 ( .B1(n16500), .B2(n18501), .A(n16499), .ZN(n16501) );
  OAI21_X1 U18309 ( .B1(n18494), .B2(n16502), .A(n16501), .ZN(P2_U3021) );
  AOI21_X1 U18310 ( .B1(n18466), .B2(n18308), .A(n16503), .ZN(n16507) );
  OAI21_X1 U18311 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16505), .A(
        n16504), .ZN(n16506) );
  OAI211_X1 U18312 ( .C1(n16508), .C2(n16567), .A(n16507), .B(n16506), .ZN(
        n16509) );
  AOI21_X1 U18313 ( .B1(n16510), .B2(n18481), .A(n16509), .ZN(n16511) );
  OAI21_X1 U18314 ( .B1(n16512), .B2(n18450), .A(n16511), .ZN(P2_U3022) );
  NAND2_X1 U18315 ( .A1(n16513), .A2(n18481), .ZN(n16522) );
  INV_X1 U18316 ( .A(n16514), .ZN(n16545) );
  XNOR2_X1 U18317 ( .A(n16515), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16518) );
  NOR2_X1 U18318 ( .A1(n18490), .A2(n18306), .ZN(n16516) );
  AOI211_X1 U18319 ( .C1(n16529), .C2(n16518), .A(n16517), .B(n16516), .ZN(
        n16519) );
  OAI21_X1 U18320 ( .B1(n18293), .B2(n16567), .A(n16519), .ZN(n16520) );
  AOI21_X1 U18321 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16545), .A(
        n16520), .ZN(n16521) );
  OAI211_X1 U18322 ( .C1(n16523), .C2(n18450), .A(n16522), .B(n16521), .ZN(
        P2_U3023) );
  XNOR2_X1 U18323 ( .A(n16525), .B(n11355), .ZN(n16526) );
  XNOR2_X1 U18324 ( .A(n16524), .B(n16526), .ZN(n17033) );
  INV_X1 U18325 ( .A(n17033), .ZN(n16535) );
  NOR2_X1 U18326 ( .A1(n12737), .A2(n18240), .ZN(n16528) );
  NOR2_X1 U18327 ( .A1(n18490), .A2(n18282), .ZN(n16527) );
  AOI211_X1 U18328 ( .C1(n16529), .C2(n11355), .A(n16528), .B(n16527), .ZN(
        n16530) );
  OAI21_X1 U18329 ( .B1(n18284), .B2(n16567), .A(n16530), .ZN(n16531) );
  AOI21_X1 U18330 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16545), .A(
        n16531), .ZN(n16534) );
  NAND2_X1 U18331 ( .A1(n16532), .A2(n11355), .ZN(n17034) );
  NAND3_X1 U18332 ( .A1(n16305), .A2(n18481), .A3(n17034), .ZN(n16533) );
  OAI211_X1 U18333 ( .C1(n16535), .C2(n18450), .A(n16534), .B(n16533), .ZN(
        P2_U3024) );
  NAND2_X1 U18334 ( .A1(n18273), .A2(n18500), .ZN(n16541) );
  INV_X1 U18335 ( .A(n16651), .ZN(n16666) );
  AND2_X1 U18336 ( .A1(n16536), .A2(n16666), .ZN(n16538) );
  AOI22_X1 U18337 ( .A1(n16539), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n16538), 
        .B2(n16537), .ZN(n16540) );
  OAI211_X1 U18338 ( .C1(n18490), .C2(n18271), .A(n16541), .B(n16540), .ZN(
        n16544) );
  NOR2_X1 U18339 ( .A1(n16542), .A2(n18494), .ZN(n16543) );
  AOI211_X1 U18340 ( .C1(n16545), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16544), .B(n16543), .ZN(n16546) );
  OAI21_X1 U18341 ( .B1(n16547), .B2(n18450), .A(n16546), .ZN(P2_U3025) );
  NAND2_X1 U18342 ( .A1(n16588), .A2(n16666), .ZN(n16554) );
  NAND2_X1 U18343 ( .A1(n16548), .A2(n16626), .ZN(n16595) );
  INV_X1 U18344 ( .A(n16549), .ZN(n16550) );
  NAND2_X1 U18345 ( .A1(n16550), .A2(n16556), .ZN(n16552) );
  NAND4_X1 U18346 ( .A1(n18489), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16551) );
  NAND3_X1 U18347 ( .A1(n18460), .A2(n16552), .A3(n16551), .ZN(n16553) );
  AND4_X1 U18348 ( .A1(n16555), .A2(n16554), .A3(n16595), .A4(n16553), .ZN(
        n16587) );
  NAND2_X1 U18349 ( .A1(n16556), .A2(n16666), .ZN(n16589) );
  INV_X1 U18350 ( .A(n16589), .ZN(n16557) );
  NAND3_X1 U18351 ( .A1(n16576), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16557), .ZN(n16574) );
  AOI21_X1 U18352 ( .B1(n16587), .B2(n16574), .A(n16558), .ZN(n16569) );
  AND2_X1 U18353 ( .A1(n16560), .A2(n16559), .ZN(n16561) );
  NOR2_X1 U18354 ( .A1(n16562), .A2(n16561), .ZN(n19344) );
  NOR3_X1 U18355 ( .A1(n16563), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16589), .ZN(n16564) );
  AOI211_X1 U18356 ( .C1(n18466), .C2(n19344), .A(n16565), .B(n16564), .ZN(
        n16566) );
  OAI21_X1 U18357 ( .B1(n18269), .B2(n16567), .A(n16566), .ZN(n16568) );
  AOI211_X1 U18358 ( .C1(n16570), .C2(n18501), .A(n16569), .B(n16568), .ZN(
        n16571) );
  OAI21_X1 U18359 ( .B1(n18494), .B2(n16572), .A(n16571), .ZN(P2_U3026) );
  NAND2_X1 U18360 ( .A1(n16573), .A2(n18481), .ZN(n16580) );
  OAI211_X1 U18361 ( .C1(n18490), .C2(n18252), .A(n16575), .B(n16574), .ZN(
        n16578) );
  NOR2_X1 U18362 ( .A1(n16587), .A2(n16576), .ZN(n16577) );
  AOI211_X1 U18363 ( .C1(n18249), .C2(n18500), .A(n16578), .B(n16577), .ZN(
        n16579) );
  OAI211_X1 U18364 ( .C1(n16581), .C2(n18450), .A(n16580), .B(n16579), .ZN(
        P2_U3027) );
  NAND2_X1 U18365 ( .A1(n16582), .A2(n18481), .ZN(n16593) );
  OR2_X1 U18366 ( .A1(n16205), .A2(n16583), .ZN(n16584) );
  AND2_X1 U18367 ( .A1(n16585), .A2(n16584), .ZN(n18234) );
  INV_X1 U18368 ( .A(n18234), .ZN(n19466) );
  OAI21_X1 U18369 ( .B1(n18490), .B2(n19466), .A(n16586), .ZN(n16591) );
  AOI21_X1 U18370 ( .B1(n16589), .B2(n16588), .A(n16587), .ZN(n16590) );
  AOI211_X1 U18371 ( .C1(n18500), .C2(n18235), .A(n16591), .B(n16590), .ZN(
        n16592) );
  OAI211_X1 U18372 ( .C1(n18450), .C2(n16594), .A(n16593), .B(n16592), .ZN(
        P2_U3028) );
  NAND2_X1 U18373 ( .A1(n18494), .A2(n18495), .ZN(n16611) );
  OAI21_X1 U18374 ( .B1(n16602), .B2(n18489), .A(n16595), .ZN(n16596) );
  NOR2_X1 U18375 ( .A1(n18459), .A2(n16596), .ZN(n16630) );
  OAI21_X1 U18376 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18422), .A(
        n16630), .ZN(n16597) );
  AOI21_X1 U18377 ( .B1(n16598), .B2(n16611), .A(n16597), .ZN(n16609) );
  NAND2_X1 U18378 ( .A1(n18222), .A2(n18500), .ZN(n16600) );
  OAI211_X1 U18379 ( .C1(n18490), .C2(n18229), .A(n16600), .B(n16599), .ZN(
        n16605) );
  OAI21_X1 U18380 ( .B1(n16601), .B2(n18494), .A(n16651), .ZN(n16603) );
  NAND2_X1 U18381 ( .A1(n16603), .A2(n16602), .ZN(n16613) );
  NOR3_X1 U18382 ( .A1(n16613), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16622), .ZN(n16604) );
  AOI211_X1 U18383 ( .C1(n16606), .C2(n18501), .A(n16605), .B(n16604), .ZN(
        n16607) );
  OAI21_X1 U18384 ( .B1(n16609), .B2(n16608), .A(n16607), .ZN(P2_U3029) );
  INV_X1 U18385 ( .A(n16630), .ZN(n16610) );
  AOI21_X1 U18386 ( .B1(n16612), .B2(n16611), .A(n16610), .ZN(n16623) );
  INV_X1 U18387 ( .A(n16613), .ZN(n16620) );
  NAND3_X1 U18388 ( .A1(n16614), .A2(n18501), .A3(n16374), .ZN(n16618) );
  NOR2_X1 U18389 ( .A1(n18475), .A2(n12721), .ZN(n16615) );
  AOI21_X1 U18390 ( .B1(n18500), .B2(n16616), .A(n16615), .ZN(n16617) );
  OAI211_X1 U18391 ( .C1(n18209), .C2(n18490), .A(n16618), .B(n16617), .ZN(
        n16619) );
  AOI21_X1 U18392 ( .B1(n16620), .B2(n16622), .A(n16619), .ZN(n16621) );
  OAI21_X1 U18393 ( .B1(n16623), .B2(n16622), .A(n16621), .ZN(P2_U3030) );
  INV_X1 U18394 ( .A(n18204), .ZN(n16634) );
  INV_X1 U18395 ( .A(n16624), .ZN(n16625) );
  AOI21_X1 U18396 ( .B1(n18500), .B2(n18197), .A(n16625), .ZN(n16628) );
  OR3_X1 U18397 ( .A1(n16651), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16626), .ZN(n16627) );
  OAI211_X1 U18398 ( .C1(n16630), .C2(n16629), .A(n16628), .B(n16627), .ZN(
        n16633) );
  NOR2_X1 U18399 ( .A1(n16631), .A2(n18450), .ZN(n16632) );
  AOI211_X1 U18400 ( .C1(n18466), .C2(n16634), .A(n16633), .B(n16632), .ZN(
        n16635) );
  OAI21_X1 U18401 ( .B1(n18494), .B2(n16636), .A(n16635), .ZN(P2_U3031) );
  NOR2_X1 U18402 ( .A1(n17006), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16637) );
  OR2_X1 U18403 ( .A1(n16399), .A2(n16637), .ZN(n17025) );
  AND3_X1 U18404 ( .A1(n17010), .A2(n16639), .A3(n16638), .ZN(n16640) );
  OR2_X1 U18405 ( .A1(n16641), .A2(n16640), .ZN(n17022) );
  NOR4_X1 U18406 ( .A1(n16651), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18461), .A4(n16642), .ZN(n16647) );
  INV_X1 U18407 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16645) );
  NOR3_X1 U18408 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18461), .A3(
        n16651), .ZN(n18464) );
  AOI211_X1 U18409 ( .C1(n18461), .C2(n18460), .A(n18464), .B(n18459), .ZN(
        n18458) );
  NOR2_X1 U18410 ( .A1(n18461), .A2(n16651), .ZN(n16643) );
  NAND2_X1 U18411 ( .A1(n16643), .A2(n18457), .ZN(n18447) );
  NAND2_X1 U18412 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n16539), .ZN(n16644) );
  OAI221_X1 U18413 ( .B1(n16645), .B2(n18458), .C1(n16645), .C2(n18447), .A(
        n16644), .ZN(n16646) );
  AOI211_X1 U18414 ( .C1(n18186), .C2(n18500), .A(n16647), .B(n16646), .ZN(
        n16648) );
  OAI21_X1 U18415 ( .B1(n18490), .B2(n18184), .A(n16648), .ZN(n16649) );
  AOI21_X1 U18416 ( .B1(n17022), .B2(n18501), .A(n16649), .ZN(n16650) );
  OAI21_X1 U18417 ( .B1(n17025), .B2(n18494), .A(n16650), .ZN(P2_U3032) );
  OR2_X1 U18418 ( .A1(n18459), .A2(n16668), .ZN(n16652) );
  NOR3_X1 U18419 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16668), .A3(
        n16651), .ZN(n18436) );
  AOI21_X1 U18420 ( .B1(n16653), .B2(n16652), .A(n18436), .ZN(n18446) );
  NAND2_X1 U18421 ( .A1(n11379), .A2(n18500), .ZN(n16658) );
  INV_X1 U18422 ( .A(n16654), .ZN(n18142) );
  AND4_X1 U18423 ( .A1(n16659), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A4(n16666), .ZN(n16655) );
  AOI211_X1 U18424 ( .C1(n18466), .C2(n18142), .A(n16656), .B(n16655), .ZN(
        n16657) );
  OAI211_X1 U18425 ( .C1(n18446), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        n16660) );
  AOI21_X1 U18426 ( .B1(n16661), .B2(n18501), .A(n16660), .ZN(n16662) );
  OAI21_X1 U18427 ( .B1(n16663), .B2(n18494), .A(n16662), .ZN(P2_U3035) );
  NAND3_X1 U18428 ( .A1(n16664), .A2(n18481), .A3(n16994), .ZN(n16673) );
  INV_X1 U18429 ( .A(n18459), .ZN(n16669) );
  OAI22_X1 U18430 ( .A1(n18490), .A2(n18123), .B1(n12694), .B2(n18475), .ZN(
        n16665) );
  AOI21_X1 U18431 ( .B1(n16666), .B2(n16668), .A(n16665), .ZN(n16667) );
  OAI21_X1 U18432 ( .B1(n16669), .B2(n16668), .A(n16667), .ZN(n16670) );
  AOI21_X1 U18433 ( .B1(n16671), .B2(n18500), .A(n16670), .ZN(n16672) );
  OAI211_X1 U18434 ( .C1(n16674), .C2(n18450), .A(n16673), .B(n16672), .ZN(
        P2_U3037) );
  INV_X1 U18435 ( .A(n16694), .ZN(n18525) );
  AOI22_X1 U18436 ( .A1(n18246), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18039), .B2(n18257), .ZN(n16678) );
  AOI222_X1 U18437 ( .A1(n16675), .A2(n16687), .B1(n18038), .B2(n18525), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n16678), .ZN(n16677) );
  NAND2_X1 U18438 ( .A1(n16690), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16676) );
  OAI21_X1 U18439 ( .B1(n16677), .B2(n16690), .A(n16676), .ZN(P2_U3601) );
  NOR2_X1 U18440 ( .A1(n16678), .A2(n16714), .ZN(n16685) );
  AOI21_X1 U18441 ( .B1(n18039), .B2(n16680), .A(n16679), .ZN(n18050) );
  AOI21_X1 U18442 ( .B1(n18246), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18050), .ZN(n16684) );
  AOI222_X1 U18443 ( .A1(n16681), .A2(n16687), .B1(n16685), .B2(n16684), .C1(
        n19035), .C2(n18525), .ZN(n16683) );
  NAND2_X1 U18444 ( .A1(n16690), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16682) );
  OAI21_X1 U18445 ( .B1(n16683), .B2(n16690), .A(n16682), .ZN(P2_U3600) );
  INV_X1 U18446 ( .A(n16684), .ZN(n16686) );
  AOI222_X1 U18447 ( .A1(n16688), .A2(n16687), .B1(n18525), .B2(n19085), .C1(
        n16686), .C2(n16685), .ZN(n16691) );
  NAND2_X1 U18448 ( .A1(n16690), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16689) );
  OAI21_X1 U18449 ( .B1(n16691), .B2(n16690), .A(n16689), .ZN(P2_U3599) );
  INV_X1 U18450 ( .A(n16692), .ZN(n16693) );
  OAI22_X1 U18451 ( .A1(n19198), .A2(n16694), .B1(n16693), .B2(n18511), .ZN(
        n16696) );
  MUX2_X1 U18452 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16696), .S(
        n16695), .Z(P2_U3596) );
  NAND2_X1 U18453 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18590) );
  NAND2_X1 U18454 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17829) );
  INV_X1 U18455 ( .A(n17829), .ZN(n17876) );
  NOR2_X1 U18456 ( .A1(n17876), .A2(n20018), .ZN(n16699) );
  NOR2_X1 U18457 ( .A1(n21176), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17525) );
  INV_X1 U18458 ( .A(n17525), .ZN(n18568) );
  NAND3_X1 U18459 ( .A1(n11377), .A2(n16697), .A3(n21139), .ZN(n17524) );
  NOR2_X1 U18460 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17524), .ZN(n16698) );
  INV_X1 U18461 ( .A(n16703), .ZN(n21174) );
  OAI21_X1 U18462 ( .B1(n16698), .B2(n21174), .A(n18765), .ZN(n17527) );
  NAND2_X1 U18463 ( .A1(n18568), .A2(n17527), .ZN(n17928) );
  AOI221_X1 U18464 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18590), .C1(n16699), 
        .C2(n18590), .A(n17928), .ZN(n17926) );
  NOR2_X1 U18465 ( .A1(n21176), .A2(n21144), .ZN(n18581) );
  OAI21_X1 U18466 ( .B1(n16699), .B2(n18581), .A(n17527), .ZN(n17930) );
  INV_X1 U18467 ( .A(n17930), .ZN(n16700) );
  INV_X1 U18468 ( .A(n18609), .ZN(n17927) );
  AOI22_X1 U18469 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16700), .B1(
        n17927), .B2(n17527), .ZN(n17925) );
  AOI22_X1 U18470 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17926), .B1(
        n17925), .B2(n21153), .ZN(P3_U2865) );
  INV_X1 U18471 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16701) );
  INV_X1 U18472 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21690) );
  AOI221_X1 U18473 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n21690), .C1(
        P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18006), 
        .ZN(n21647) );
  INV_X1 U18474 ( .A(BS16), .ZN(n16861) );
  NAND2_X1 U18475 ( .A1(n21698), .A2(n21690), .ZN(n21648) );
  AOI21_X1 U18476 ( .B1(n16861), .B2(n21648), .A(n16702), .ZN(n21643) );
  AOI21_X1 U18477 ( .B1(n16701), .B2(n16702), .A(n21643), .ZN(P3_U3280) );
  AND2_X1 U18478 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16702), .ZN(P3_U3028) );
  AND2_X1 U18479 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16702), .ZN(P3_U3027) );
  AND2_X1 U18480 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16702), .ZN(P3_U3026) );
  AND2_X1 U18481 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16702), .ZN(P3_U3025) );
  AND2_X1 U18482 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16702), .ZN(P3_U3024) );
  AND2_X1 U18483 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16702), .ZN(P3_U3023) );
  AND2_X1 U18484 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16702), .ZN(P3_U3022) );
  AND2_X1 U18485 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16702), .ZN(P3_U3021) );
  AND2_X1 U18486 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16702), .ZN(
        P3_U3020) );
  AND2_X1 U18487 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16702), .ZN(
        P3_U3019) );
  AND2_X1 U18488 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16702), .ZN(
        P3_U3018) );
  AND2_X1 U18489 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16702), .ZN(
        P3_U3017) );
  AND2_X1 U18490 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16702), .ZN(
        P3_U3016) );
  AND2_X1 U18491 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16702), .ZN(
        P3_U3015) );
  AND2_X1 U18492 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16702), .ZN(
        P3_U3014) );
  AND2_X1 U18493 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16702), .ZN(
        P3_U3013) );
  AND2_X1 U18494 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16702), .ZN(
        P3_U3012) );
  AND2_X1 U18495 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16702), .ZN(
        P3_U3011) );
  AND2_X1 U18496 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16702), .ZN(
        P3_U3010) );
  AND2_X1 U18497 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16702), .ZN(
        P3_U3009) );
  AND2_X1 U18498 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16702), .ZN(
        P3_U3008) );
  AND2_X1 U18499 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16702), .ZN(
        P3_U3007) );
  AND2_X1 U18500 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16702), .ZN(
        P3_U3006) );
  AND2_X1 U18501 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16702), .ZN(
        P3_U3005) );
  AND2_X1 U18502 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16702), .ZN(
        P3_U3004) );
  AND2_X1 U18503 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16702), .ZN(
        P3_U3003) );
  AND2_X1 U18504 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16702), .ZN(
        P3_U3002) );
  AND2_X1 U18505 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16702), .ZN(
        P3_U3001) );
  AND2_X1 U18506 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16702), .ZN(
        P3_U3000) );
  AND2_X1 U18507 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16702), .ZN(
        P3_U2999) );
  AOI21_X1 U18508 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16704)
         );
  NOR4_X1 U18509 ( .A1(n17919), .A2(n20082), .A3(n21649), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21124) );
  AOI211_X1 U18510 ( .C1(n17829), .C2(n16704), .A(n16703), .B(n21124), .ZN(
        P3_U2998) );
  INV_X1 U18511 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21157) );
  NOR2_X1 U18512 ( .A1(n21157), .A2(n17527), .ZN(P3_U2867) );
  NOR2_X1 U18513 ( .A1(n17919), .A2(n17917), .ZN(n21177) );
  NAND2_X1 U18514 ( .A1(n21164), .A2(n21130), .ZN(n20027) );
  AND2_X1 U18515 ( .A1(n17982), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U18516 ( .A(n20016), .ZN(n20090) );
  OAI21_X1 U18517 ( .B1(n17520), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n20090), 
        .ZN(n16706) );
  OAI21_X1 U18518 ( .B1(n20090), .B2(n16707), .A(n16706), .ZN(P3_U3298) );
  NOR2_X1 U18519 ( .A1(n17520), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n16708)
         );
  OAI21_X1 U18520 ( .B1(n20016), .B2(n16708), .A(n20088), .ZN(P3_U3299) );
  INV_X1 U18521 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21677) );
  NOR2_X1 U18522 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21677), .ZN(n21671) );
  AOI21_X1 U18523 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21671), .A(n16709), 
        .ZN(n16711) );
  INV_X1 U18524 ( .A(n16711), .ZN(n21642) );
  INV_X1 U18525 ( .A(n21642), .ZN(n16712) );
  INV_X1 U18526 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16728) );
  NAND2_X1 U18527 ( .A1(n21682), .A2(n21677), .ZN(n16710) );
  AOI21_X1 U18528 ( .B1(n16861), .B2(n16710), .A(n16712), .ZN(n21638) );
  AOI21_X1 U18529 ( .B1(n16712), .B2(n16728), .A(n21638), .ZN(P2_U3591) );
  AND2_X1 U18530 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n16712), .ZN(P2_U3208) );
  AND2_X1 U18531 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n16712), .ZN(P2_U3207) );
  AND2_X1 U18532 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n16712), .ZN(P2_U3206) );
  AND2_X1 U18533 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n16712), .ZN(P2_U3205) );
  AND2_X1 U18534 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n16712), .ZN(P2_U3204) );
  AND2_X1 U18535 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n16712), .ZN(P2_U3203) );
  AND2_X1 U18536 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n16712), .ZN(P2_U3202) );
  AND2_X1 U18537 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n16712), .ZN(P2_U3201) );
  AND2_X1 U18538 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16712), .ZN(
        P2_U3200) );
  AND2_X1 U18539 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16712), .ZN(
        P2_U3199) );
  AND2_X1 U18540 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16712), .ZN(
        P2_U3198) );
  AND2_X1 U18541 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16712), .ZN(
        P2_U3197) );
  AND2_X1 U18542 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16712), .ZN(
        P2_U3196) );
  AND2_X1 U18543 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16712), .ZN(
        P2_U3195) );
  AND2_X1 U18544 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16711), .ZN(
        P2_U3194) );
  AND2_X1 U18545 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n16711), .ZN(
        P2_U3193) );
  AND2_X1 U18546 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n16711), .ZN(
        P2_U3192) );
  AND2_X1 U18547 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n16711), .ZN(
        P2_U3191) );
  AND2_X1 U18548 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n16711), .ZN(
        P2_U3190) );
  AND2_X1 U18549 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n16711), .ZN(
        P2_U3189) );
  AND2_X1 U18550 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n16711), .ZN(
        P2_U3188) );
  AND2_X1 U18551 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n16711), .ZN(
        P2_U3187) );
  AND2_X1 U18552 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n16711), .ZN(
        P2_U3186) );
  AND2_X1 U18553 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n16711), .ZN(
        P2_U3185) );
  AND2_X1 U18554 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n16711), .ZN(
        P2_U3184) );
  AND2_X1 U18555 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n16711), .ZN(
        P2_U3183) );
  AND2_X1 U18556 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n16712), .ZN(
        P2_U3182) );
  AND2_X1 U18557 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n16712), .ZN(
        P2_U3181) );
  AND2_X1 U18558 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n16712), .ZN(
        P2_U3180) );
  AND2_X1 U18559 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n16712), .ZN(
        P2_U3179) );
  NAND2_X1 U18560 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18527), .ZN(n18512) );
  AOI21_X1 U18561 ( .B1(n16713), .B2(n18022), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16715) );
  AOI221_X1 U18562 ( .B1(n18512), .B2(n16715), .C1(n16714), .C2(n16715), .A(
        n16716), .ZN(P2_U3178) );
  AOI221_X1 U18563 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16716), .C1(n18520), .C2(
        n16716), .A(n19219), .ZN(n17064) );
  INV_X1 U18564 ( .A(n17064), .ZN(n17062) );
  NOR2_X1 U18565 ( .A1(n16717), .A2(n17062), .ZN(P2_U3047) );
  AND2_X1 U18566 ( .A1(n17095), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18567 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16721) );
  NOR4_X1 U18568 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16720) );
  NOR4_X1 U18569 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16719) );
  NOR4_X1 U18570 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16718) );
  NAND4_X1 U18571 ( .A1(n16721), .A2(n16720), .A3(n16719), .A4(n16718), .ZN(
        n16727) );
  NOR4_X1 U18572 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16725) );
  AOI211_X1 U18573 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16724) );
  NOR4_X1 U18574 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16723) );
  NOR4_X1 U18575 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16722) );
  NAND4_X1 U18576 ( .A1(n16725), .A2(n16724), .A3(n16723), .A4(n16722), .ZN(
        n16726) );
  NOR2_X1 U18577 ( .A1(n16727), .A2(n16726), .ZN(n17072) );
  INV_X1 U18578 ( .A(n17072), .ZN(n17070) );
  NOR2_X1 U18579 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17070), .ZN(n17065) );
  INV_X1 U18580 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21641) );
  NAND3_X1 U18581 ( .A1(n11137), .A2(n21641), .A3(n16728), .ZN(n17069) );
  INV_X1 U18582 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16729) );
  AOI22_X1 U18583 ( .A1(n17065), .A2(n17069), .B1(n17070), .B2(n16729), .ZN(
        P2_U2821) );
  INV_X1 U18584 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n16730) );
  AOI22_X1 U18585 ( .A1(n17065), .A2(n11137), .B1(n17070), .B2(n16730), .ZN(
        P2_U2820) );
  INV_X1 U18586 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16731) );
  INV_X1 U18587 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21659) );
  NOR2_X1 U18588 ( .A1(n21659), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21656) );
  OAI21_X1 U18589 ( .B1(n21656), .B2(n13264), .A(n11057), .ZN(n16732) );
  INV_X1 U18590 ( .A(n16732), .ZN(n21634) );
  OAI221_X1 U18591 ( .B1(n21659), .B2(BS16), .C1(n12962), .C2(BS16), .A(n21634), .ZN(n21633) );
  INV_X1 U18592 ( .A(n21633), .ZN(n21635) );
  AOI21_X1 U18593 ( .B1(n16731), .B2(n21636), .A(n21635), .ZN(P1_U3464) );
  AND2_X1 U18594 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21636), .ZN(P1_U3193) );
  AND2_X1 U18595 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n16732), .ZN(P1_U3192) );
  AND2_X1 U18596 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21636), .ZN(P1_U3191) );
  AND2_X1 U18597 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21636), .ZN(P1_U3190) );
  AND2_X1 U18598 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21636), .ZN(P1_U3189) );
  AND2_X1 U18599 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21636), .ZN(P1_U3188) );
  AND2_X1 U18600 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21636), .ZN(P1_U3187) );
  AND2_X1 U18601 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21636), .ZN(P1_U3186) );
  AND2_X1 U18602 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21636), .ZN(
        P1_U3185) );
  AND2_X1 U18603 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21636), .ZN(
        P1_U3184) );
  AND2_X1 U18604 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21636), .ZN(
        P1_U3183) );
  AND2_X1 U18605 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21636), .ZN(
        P1_U3182) );
  AND2_X1 U18606 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21636), .ZN(
        P1_U3181) );
  AND2_X1 U18607 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21636), .ZN(
        P1_U3180) );
  AND2_X1 U18608 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21636), .ZN(
        P1_U3179) );
  AND2_X1 U18609 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21636), .ZN(
        P1_U3178) );
  AND2_X1 U18610 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n16732), .ZN(
        P1_U3177) );
  AND2_X1 U18611 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21636), .ZN(
        P1_U3176) );
  AND2_X1 U18612 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21636), .ZN(
        P1_U3175) );
  AND2_X1 U18613 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21636), .ZN(
        P1_U3174) );
  AND2_X1 U18614 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21636), .ZN(
        P1_U3173) );
  AND2_X1 U18615 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21636), .ZN(
        P1_U3172) );
  AND2_X1 U18616 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n16732), .ZN(
        P1_U3171) );
  AND2_X1 U18617 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21636), .ZN(
        P1_U3170) );
  AND2_X1 U18618 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21636), .ZN(
        P1_U3169) );
  AND2_X1 U18619 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21636), .ZN(
        P1_U3168) );
  AND2_X1 U18620 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21636), .ZN(
        P1_U3167) );
  AND2_X1 U18621 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21636), .ZN(
        P1_U3166) );
  AND2_X1 U18622 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21636), .ZN(
        P1_U3165) );
  AND2_X1 U18623 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21636), .ZN(
        P1_U3164) );
  NAND2_X1 U18624 ( .A1(n16747), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16744) );
  NAND2_X1 U18625 ( .A1(n16733), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16734) );
  OR2_X1 U18626 ( .A1(n16735), .A2(n16734), .ZN(n16739) );
  INV_X1 U18627 ( .A(n16739), .ZN(n16742) );
  NAND2_X1 U18628 ( .A1(n16745), .A2(n21853), .ZN(n16741) );
  INV_X1 U18629 ( .A(n16736), .ZN(n16737) );
  OAI211_X1 U18630 ( .C1(n21827), .C2(n16739), .A(n16738), .B(n16737), .ZN(
        n16740) );
  OAI211_X1 U18631 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16742), .A(
        n16741), .B(n16740), .ZN(n16743) );
  OAI211_X1 U18632 ( .C1(n16745), .C2(n21853), .A(n16744), .B(n16743), .ZN(
        n16746) );
  OAI21_X1 U18633 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16747), .A(
        n16746), .ZN(n16755) );
  NOR2_X1 U18634 ( .A1(P1_MORE_REG_SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(
        n16751) );
  INV_X1 U18635 ( .A(n16748), .ZN(n16750) );
  OAI211_X1 U18636 ( .C1(n16752), .C2(n16751), .A(n16750), .B(n16749), .ZN(
        n16754) );
  AOI211_X1 U18637 ( .C1(n16769), .C2(n16755), .A(n16754), .B(n16753), .ZN(
        n21632) );
  OR2_X1 U18638 ( .A1(n21660), .A2(n16756), .ZN(n16763) );
  INV_X1 U18639 ( .A(n16757), .ZN(n16758) );
  NOR4_X1 U18640 ( .A1(n16760), .A2(n16759), .A3(n21657), .A4(n16758), .ZN(
        n16761) );
  AOI21_X1 U18641 ( .B1(n16763), .B2(n16762), .A(n16761), .ZN(n21626) );
  AND2_X1 U18642 ( .A1(n21632), .A2(n21626), .ZN(n21613) );
  OAI21_X1 U18643 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21660), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n16764) );
  NOR3_X1 U18644 ( .A1(n21622), .A2(n21613), .A3(n16764), .ZN(n21625) );
  NOR2_X1 U18645 ( .A1(n16765), .A2(n16764), .ZN(n21617) );
  AOI21_X1 U18646 ( .B1(n21627), .B2(n14136), .A(n21617), .ZN(n16766) );
  OAI22_X1 U18647 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21625), .B1(n21626), 
        .B2(n16766), .ZN(n16767) );
  INV_X1 U18648 ( .A(n16767), .ZN(P1_U3162) );
  NOR2_X1 U18649 ( .A1(n16769), .A2(n16768), .ZN(P1_U3032) );
  AND2_X1 U18650 ( .A1(n19802), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18651 ( .A1(n21656), .A2(n13264), .ZN(n16770) );
  INV_X1 U18652 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n16909) );
  AOI21_X1 U18653 ( .B1(n16770), .B2(n16909), .A(n22319), .ZN(P1_U2802) );
  OAI22_X1 U18654 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_63), .B1(
        keyinput_61), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16771) );
  AOI221_X1 U18655 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_63), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_61), .A(n16771), .ZN(n16857) );
  INV_X1 U18656 ( .A(keyinput_56), .ZN(n16850) );
  INV_X1 U18657 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16942) );
  INV_X1 U18658 ( .A(keyinput_55), .ZN(n16848) );
  INV_X1 U18659 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19868) );
  INV_X1 U18660 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19875) );
  OAI22_X1 U18661 ( .A1(n19868), .A2(keyinput_50), .B1(n19875), .B2(
        keyinput_49), .ZN(n16772) );
  AOI221_X1 U18662 ( .B1(n19868), .B2(keyinput_50), .C1(keyinput_49), .C2(
        n19875), .A(n16772), .ZN(n16846) );
  INV_X1 U18663 ( .A(keyinput_48), .ZN(n16838) );
  INV_X1 U18664 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n16930) );
  INV_X1 U18665 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n16924) );
  OAI22_X1 U18666 ( .A1(n16924), .A2(keyinput_45), .B1(P1_FLUSH_REG_SCAN_IN), 
        .B2(keyinput_46), .ZN(n16773) );
  AOI221_X1 U18667 ( .B1(n16924), .B2(keyinput_45), .C1(keyinput_46), .C2(
        P1_FLUSH_REG_SCAN_IN), .A(n16773), .ZN(n16835) );
  XOR2_X1 U18668 ( .A(n16861), .B(keyinput_35), .Z(n16827) );
  OAI22_X1 U18669 ( .A1(DATAI_0_), .A2(keyinput_32), .B1(keyinput_33), .B2(
        HOLD), .ZN(n16774) );
  AOI221_X1 U18670 ( .B1(DATAI_0_), .B2(keyinput_32), .C1(HOLD), .C2(
        keyinput_33), .A(n16774), .ZN(n16819) );
  INV_X1 U18671 ( .A(DATAI_10_), .ZN(n16892) );
  INV_X1 U18672 ( .A(keyinput_22), .ZN(n16804) );
  INV_X1 U18673 ( .A(DATAI_17_), .ZN(n21916) );
  INV_X1 U18674 ( .A(DATAI_19_), .ZN(n22010) );
  AOI22_X1 U18675 ( .A1(DATAI_18_), .A2(keyinput_14), .B1(n22010), .B2(
        keyinput_13), .ZN(n16775) );
  OAI221_X1 U18676 ( .B1(DATAI_18_), .B2(keyinput_14), .C1(n22010), .C2(
        keyinput_13), .A(n16775), .ZN(n16792) );
  INV_X1 U18677 ( .A(DATAI_23_), .ZN(n22206) );
  XOR2_X1 U18678 ( .A(n22206), .B(keyinput_9), .Z(n16790) );
  INV_X1 U18679 ( .A(DATAI_20_), .ZN(n22057) );
  AOI22_X1 U18680 ( .A1(DATAI_22_), .A2(keyinput_10), .B1(n22057), .B2(
        keyinput_12), .ZN(n16776) );
  OAI221_X1 U18681 ( .B1(DATAI_22_), .B2(keyinput_10), .C1(n22057), .C2(
        keyinput_12), .A(n16776), .ZN(n16789) );
  AOI22_X1 U18682 ( .A1(DATAI_26_), .A2(keyinput_6), .B1(DATAI_27_), .B2(
        keyinput_5), .ZN(n16777) );
  OAI221_X1 U18683 ( .B1(DATAI_26_), .B2(keyinput_6), .C1(DATAI_27_), .C2(
        keyinput_5), .A(n16777), .ZN(n16784) );
  INV_X1 U18684 ( .A(DATAI_28_), .ZN(n22055) );
  OAI22_X1 U18685 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(keyinput_2), .B2(
        DATAI_30_), .ZN(n16778) );
  AOI221_X1 U18686 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(DATAI_30_), .C2(
        keyinput_2), .A(n16778), .ZN(n16781) );
  OAI22_X1 U18687 ( .A1(DATAI_29_), .A2(keyinput_3), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .ZN(n16779) );
  AOI221_X1 U18688 ( .B1(DATAI_29_), .B2(keyinput_3), .C1(keyinput_0), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n16779), .ZN(n16780) );
  AOI22_X1 U18689 ( .A1(n16781), .A2(n16780), .B1(keyinput_4), .B2(n22055), 
        .ZN(n16782) );
  OAI21_X1 U18690 ( .B1(keyinput_4), .B2(n22055), .A(n16782), .ZN(n16783) );
  OAI22_X1 U18691 ( .A1(n16784), .A2(n16783), .B1(keyinput_7), .B2(DATAI_25_), 
        .ZN(n16785) );
  AOI21_X1 U18692 ( .B1(keyinput_7), .B2(DATAI_25_), .A(n16785), .ZN(n16788)
         );
  AOI22_X1 U18693 ( .A1(DATAI_21_), .A2(keyinput_11), .B1(DATAI_24_), .B2(
        keyinput_8), .ZN(n16786) );
  OAI221_X1 U18694 ( .B1(DATAI_21_), .B2(keyinput_11), .C1(DATAI_24_), .C2(
        keyinput_8), .A(n16786), .ZN(n16787) );
  NOR4_X1 U18695 ( .A1(n16790), .A2(n16789), .A3(n16788), .A4(n16787), .ZN(
        n16791) );
  OAI22_X1 U18696 ( .A1(n16792), .A2(n16791), .B1(n21916), .B2(keyinput_15), 
        .ZN(n16793) );
  AOI21_X1 U18697 ( .B1(n21916), .B2(keyinput_15), .A(n16793), .ZN(n16802) );
  OAI22_X1 U18698 ( .A1(n13667), .A2(keyinput_17), .B1(keyinput_16), .B2(
        DATAI_16_), .ZN(n16794) );
  AOI221_X1 U18699 ( .B1(n13667), .B2(keyinput_17), .C1(DATAI_16_), .C2(
        keyinput_16), .A(n16794), .ZN(n16801) );
  AOI22_X1 U18700 ( .A1(n16797), .A2(keyinput_19), .B1(n16796), .B2(
        keyinput_18), .ZN(n16795) );
  OAI221_X1 U18701 ( .B1(n16797), .B2(keyinput_19), .C1(n16796), .C2(
        keyinput_18), .A(n16795), .ZN(n16800) );
  AOI22_X1 U18702 ( .A1(DATAI_11_), .A2(keyinput_21), .B1(DATAI_12_), .B2(
        keyinput_20), .ZN(n16798) );
  OAI221_X1 U18703 ( .B1(DATAI_11_), .B2(keyinput_21), .C1(DATAI_12_), .C2(
        keyinput_20), .A(n16798), .ZN(n16799) );
  AOI211_X1 U18704 ( .C1(n16802), .C2(n16801), .A(n16800), .B(n16799), .ZN(
        n16803) );
  AOI221_X1 U18705 ( .B1(DATAI_10_), .B2(keyinput_22), .C1(n16892), .C2(n16804), .A(n16803), .ZN(n16813) );
  AOI22_X1 U18706 ( .A1(DATAI_4_), .A2(keyinput_28), .B1(DATAI_6_), .B2(
        keyinput_26), .ZN(n16805) );
  OAI221_X1 U18707 ( .B1(DATAI_4_), .B2(keyinput_28), .C1(DATAI_6_), .C2(
        keyinput_26), .A(n16805), .ZN(n16812) );
  INV_X1 U18708 ( .A(DATAI_9_), .ZN(n16807) );
  AOI22_X1 U18709 ( .A1(DATAI_7_), .A2(keyinput_25), .B1(n16807), .B2(
        keyinput_23), .ZN(n16806) );
  OAI221_X1 U18710 ( .B1(DATAI_7_), .B2(keyinput_25), .C1(n16807), .C2(
        keyinput_23), .A(n16806), .ZN(n16811) );
  INV_X1 U18711 ( .A(DATAI_8_), .ZN(n16809) );
  AOI22_X1 U18712 ( .A1(n13590), .A2(keyinput_27), .B1(n16809), .B2(
        keyinput_24), .ZN(n16808) );
  OAI221_X1 U18713 ( .B1(n13590), .B2(keyinput_27), .C1(n16809), .C2(
        keyinput_24), .A(n16808), .ZN(n16810) );
  NOR4_X1 U18714 ( .A1(n16813), .A2(n16812), .A3(n16811), .A4(n16810), .ZN(
        n16816) );
  AOI22_X1 U18715 ( .A1(DATAI_3_), .A2(keyinput_29), .B1(n13618), .B2(
        keyinput_31), .ZN(n16814) );
  OAI221_X1 U18716 ( .B1(DATAI_3_), .B2(keyinput_29), .C1(n13618), .C2(
        keyinput_31), .A(n16814), .ZN(n16815) );
  AOI211_X1 U18717 ( .C1(n13607), .C2(keyinput_30), .A(n16816), .B(n16815), 
        .ZN(n16817) );
  OAI21_X1 U18718 ( .B1(n13607), .B2(keyinput_30), .A(n16817), .ZN(n16818) );
  AOI22_X1 U18719 ( .A1(n16819), .A2(n16818), .B1(keyinput_34), .B2(NA), .ZN(
        n16820) );
  OAI21_X1 U18720 ( .B1(keyinput_34), .B2(NA), .A(n16820), .ZN(n16826) );
  INV_X1 U18721 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n16822) );
  AOI22_X1 U18722 ( .A1(keyinput_36), .A2(READY1), .B1(n16822), .B2(
        keyinput_38), .ZN(n16821) );
  OAI221_X1 U18723 ( .B1(keyinput_36), .B2(READY1), .C1(n16822), .C2(
        keyinput_38), .A(n16821), .ZN(n16825) );
  AOI22_X1 U18724 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_39), .B1(READY2), 
        .B2(keyinput_37), .ZN(n16823) );
  OAI221_X1 U18725 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_39), .C1(READY2), 
        .C2(keyinput_37), .A(n16823), .ZN(n16824) );
  AOI211_X1 U18726 ( .C1(n16827), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        n16833) );
  INV_X1 U18727 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n19968) );
  AOI22_X1 U18728 ( .A1(keyinput_41), .A2(P1_M_IO_N_REG_SCAN_IN), .B1(n19968), 
        .B2(keyinput_40), .ZN(n16828) );
  OAI221_X1 U18729 ( .B1(keyinput_41), .B2(P1_M_IO_N_REG_SCAN_IN), .C1(n19968), 
        .C2(keyinput_40), .A(n16828), .ZN(n16832) );
  OAI22_X1 U18730 ( .A1(n21881), .A2(keyinput_44), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(keyinput_42), .ZN(n16829) );
  AOI221_X1 U18731 ( .B1(n21881), .B2(keyinput_44), .C1(keyinput_42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n16829), .ZN(n16831) );
  XNOR2_X1 U18732 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .ZN(
        n16830) );
  OAI211_X1 U18733 ( .C1(n16833), .C2(n16832), .A(n16831), .B(n16830), .ZN(
        n16834) );
  AOI22_X1 U18734 ( .A1(n16835), .A2(n16834), .B1(keyinput_47), .B2(
        P1_W_R_N_REG_SCAN_IN), .ZN(n16836) );
  OAI21_X1 U18735 ( .B1(keyinput_47), .B2(P1_W_R_N_REG_SCAN_IN), .A(n16836), 
        .ZN(n16837) );
  OAI221_X1 U18736 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n16838), .C1(
        n16930), .C2(keyinput_48), .A(n16837), .ZN(n16845) );
  INV_X1 U18737 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U18738 ( .A1(n16841), .A2(keyinput_52), .B1(keyinput_51), .B2(
        n16840), .ZN(n16839) );
  OAI221_X1 U18739 ( .B1(n16841), .B2(keyinput_52), .C1(n16840), .C2(
        keyinput_51), .A(n16839), .ZN(n16844) );
  AOI22_X1 U18740 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_53), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .ZN(n16842) );
  OAI221_X1 U18741 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_53), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_54), .A(n16842), .ZN(n16843) );
  AOI211_X1 U18742 ( .C1(n16846), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        n16847) );
  AOI221_X1 U18743 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .C1(
        n15330), .C2(n16848), .A(n16847), .ZN(n16849) );
  AOI221_X1 U18744 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n16850), .C1(n16942), 
        .C2(keyinput_56), .A(n16849), .ZN(n16855) );
  AOI22_X1 U18745 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_58), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .ZN(n16851) );
  OAI221_X1 U18746 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_57), .A(n16851), .ZN(n16854) );
  OAI22_X1 U18747 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_59), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .ZN(n16852) );
  AOI221_X1 U18748 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .C1(
        keyinput_60), .C2(P1_REIP_REG_23__SCAN_IN), .A(n16852), .ZN(n16853) );
  OAI21_X1 U18749 ( .B1(n16855), .B2(n16854), .A(n16853), .ZN(n16856) );
  OAI211_X1 U18750 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(keyinput_62), .A(n16857), .B(n16856), .ZN(n16858) );
  AOI21_X1 U18751 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .A(n16858), 
        .ZN(n16952) );
  OAI22_X1 U18752 ( .A1(n16860), .A2(keyinput_121), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_122), .ZN(n16859) );
  AOI221_X1 U18753 ( .B1(n16860), .B2(keyinput_121), .C1(keyinput_122), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n16859), .ZN(n16947) );
  INV_X1 U18754 ( .A(keyinput_120), .ZN(n16943) );
  INV_X1 U18755 ( .A(keyinput_119), .ZN(n16940) );
  INV_X1 U18756 ( .A(keyinput_112), .ZN(n16929) );
  XNOR2_X1 U18757 ( .A(n16861), .B(keyinput_99), .ZN(n16915) );
  OAI22_X1 U18758 ( .A1(n13623), .A2(keyinput_96), .B1(keyinput_97), .B2(HOLD), 
        .ZN(n16862) );
  AOI221_X1 U18759 ( .B1(n13623), .B2(keyinput_96), .C1(HOLD), .C2(keyinput_97), .A(n16862), .ZN(n16905) );
  INV_X1 U18760 ( .A(keyinput_86), .ZN(n16891) );
  INV_X1 U18761 ( .A(DATAI_16_), .ZN(n21726) );
  AOI22_X1 U18762 ( .A1(DATAI_18_), .A2(keyinput_78), .B1(DATAI_19_), .B2(
        keyinput_77), .ZN(n16863) );
  OAI221_X1 U18763 ( .B1(DATAI_18_), .B2(keyinput_78), .C1(DATAI_19_), .C2(
        keyinput_77), .A(n16863), .ZN(n16880) );
  XOR2_X1 U18764 ( .A(keyinput_72), .B(DATAI_24_), .Z(n16878) );
  INV_X1 U18765 ( .A(DATAI_21_), .ZN(n22105) );
  AOI22_X1 U18766 ( .A1(n22105), .A2(keyinput_75), .B1(keyinput_76), .B2(
        n22057), .ZN(n16864) );
  OAI221_X1 U18767 ( .B1(n22105), .B2(keyinput_75), .C1(n22057), .C2(
        keyinput_76), .A(n16864), .ZN(n16877) );
  INV_X1 U18768 ( .A(DATAI_27_), .ZN(n22008) );
  AOI22_X1 U18769 ( .A1(DATAI_28_), .A2(keyinput_68), .B1(n22008), .B2(
        keyinput_69), .ZN(n16865) );
  OAI221_X1 U18770 ( .B1(DATAI_28_), .B2(keyinput_68), .C1(n22008), .C2(
        keyinput_69), .A(n16865), .ZN(n16872) );
  INV_X1 U18771 ( .A(DATAI_26_), .ZN(n21960) );
  OAI22_X1 U18772 ( .A1(DATAI_30_), .A2(keyinput_66), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .ZN(n16866) );
  AOI221_X1 U18773 ( .B1(DATAI_30_), .B2(keyinput_66), .C1(keyinput_64), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n16866), .ZN(n16869) );
  OAI22_X1 U18774 ( .A1(DATAI_31_), .A2(keyinput_65), .B1(DATAI_29_), .B2(
        keyinput_67), .ZN(n16867) );
  AOI221_X1 U18775 ( .B1(DATAI_31_), .B2(keyinput_65), .C1(keyinput_67), .C2(
        DATAI_29_), .A(n16867), .ZN(n16868) );
  AOI22_X1 U18776 ( .A1(n16869), .A2(n16868), .B1(keyinput_70), .B2(n21960), 
        .ZN(n16870) );
  OAI21_X1 U18777 ( .B1(keyinput_70), .B2(n21960), .A(n16870), .ZN(n16871) );
  OAI22_X1 U18778 ( .A1(n16872), .A2(n16871), .B1(keyinput_71), .B2(DATAI_25_), 
        .ZN(n16873) );
  AOI21_X1 U18779 ( .B1(keyinput_71), .B2(DATAI_25_), .A(n16873), .ZN(n16876)
         );
  INV_X1 U18780 ( .A(DATAI_22_), .ZN(n22152) );
  AOI22_X1 U18781 ( .A1(n22206), .A2(keyinput_73), .B1(keyinput_74), .B2(
        n22152), .ZN(n16874) );
  OAI221_X1 U18782 ( .B1(n22206), .B2(keyinput_73), .C1(n22152), .C2(
        keyinput_74), .A(n16874), .ZN(n16875) );
  NOR4_X1 U18783 ( .A1(n16878), .A2(n16877), .A3(n16876), .A4(n16875), .ZN(
        n16879) );
  OAI22_X1 U18784 ( .A1(n16880), .A2(n16879), .B1(n21726), .B2(keyinput_80), 
        .ZN(n16881) );
  AOI21_X1 U18785 ( .B1(n21726), .B2(keyinput_80), .A(n16881), .ZN(n16889) );
  OAI22_X1 U18786 ( .A1(n13667), .A2(keyinput_81), .B1(DATAI_17_), .B2(
        keyinput_79), .ZN(n16882) );
  AOI221_X1 U18787 ( .B1(n13667), .B2(keyinput_81), .C1(keyinput_79), .C2(
        DATAI_17_), .A(n16882), .ZN(n16888) );
  INV_X1 U18788 ( .A(DATAI_11_), .ZN(n16884) );
  AOI22_X1 U18789 ( .A1(DATAI_13_), .A2(keyinput_83), .B1(n16884), .B2(
        keyinput_85), .ZN(n16883) );
  OAI221_X1 U18790 ( .B1(DATAI_13_), .B2(keyinput_83), .C1(n16884), .C2(
        keyinput_85), .A(n16883), .ZN(n16887) );
  AOI22_X1 U18791 ( .A1(DATAI_12_), .A2(keyinput_84), .B1(DATAI_14_), .B2(
        keyinput_82), .ZN(n16885) );
  OAI221_X1 U18792 ( .B1(DATAI_12_), .B2(keyinput_84), .C1(DATAI_14_), .C2(
        keyinput_82), .A(n16885), .ZN(n16886) );
  AOI211_X1 U18793 ( .C1(n16889), .C2(n16888), .A(n16887), .B(n16886), .ZN(
        n16890) );
  AOI221_X1 U18794 ( .B1(DATAI_10_), .B2(keyinput_86), .C1(n16892), .C2(n16891), .A(n16890), .ZN(n16899) );
  AOI22_X1 U18795 ( .A1(DATAI_8_), .A2(keyinput_88), .B1(n13568), .B2(
        keyinput_90), .ZN(n16893) );
  OAI221_X1 U18796 ( .B1(DATAI_8_), .B2(keyinput_88), .C1(n13568), .C2(
        keyinput_90), .A(n16893), .ZN(n16898) );
  AOI22_X1 U18797 ( .A1(DATAI_9_), .A2(keyinput_87), .B1(n13590), .B2(
        keyinput_91), .ZN(n16894) );
  OAI221_X1 U18798 ( .B1(DATAI_9_), .B2(keyinput_87), .C1(n13590), .C2(
        keyinput_91), .A(n16894), .ZN(n16897) );
  AOI22_X1 U18799 ( .A1(n13610), .A2(keyinput_92), .B1(n13580), .B2(
        keyinput_89), .ZN(n16895) );
  OAI221_X1 U18800 ( .B1(n13610), .B2(keyinput_92), .C1(n13580), .C2(
        keyinput_89), .A(n16895), .ZN(n16896) );
  NOR4_X1 U18801 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16902) );
  AOI22_X1 U18802 ( .A1(DATAI_2_), .A2(keyinput_94), .B1(n13618), .B2(
        keyinput_95), .ZN(n16900) );
  OAI221_X1 U18803 ( .B1(DATAI_2_), .B2(keyinput_94), .C1(n13618), .C2(
        keyinput_95), .A(n16900), .ZN(n16901) );
  AOI211_X1 U18804 ( .C1(n13613), .C2(keyinput_93), .A(n16902), .B(n16901), 
        .ZN(n16903) );
  OAI21_X1 U18805 ( .B1(n13613), .B2(keyinput_93), .A(n16903), .ZN(n16904) );
  AOI22_X1 U18806 ( .A1(n16905), .A2(n16904), .B1(keyinput_98), .B2(NA), .ZN(
        n16906) );
  OAI21_X1 U18807 ( .B1(keyinput_98), .B2(NA), .A(n16906), .ZN(n16914) );
  INV_X1 U18808 ( .A(READY1), .ZN(n16908) );
  AOI22_X1 U18809 ( .A1(n16909), .A2(keyinput_103), .B1(n16908), .B2(
        keyinput_100), .ZN(n16907) );
  OAI221_X1 U18810 ( .B1(n16909), .B2(keyinput_103), .C1(n16908), .C2(
        keyinput_100), .A(n16907), .ZN(n16913) );
  INV_X1 U18811 ( .A(READY2), .ZN(n16911) );
  AOI22_X1 U18812 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_102), .B1(
        n16911), .B2(keyinput_101), .ZN(n16910) );
  OAI221_X1 U18813 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_102), .C1(
        n16911), .C2(keyinput_101), .A(n16910), .ZN(n16912) );
  AOI211_X1 U18814 ( .C1(n16915), .C2(n16914), .A(n16913), .B(n16912), .ZN(
        n16922) );
  AOI22_X1 U18815 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_104), .B1(
        n16917), .B2(keyinput_105), .ZN(n16916) );
  OAI221_X1 U18816 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_104), .C1(
        n16917), .C2(keyinput_105), .A(n16916), .ZN(n16921) );
  OAI22_X1 U18817 ( .A1(n21881), .A2(keyinput_108), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(keyinput_106), .ZN(n16918) );
  AOI221_X1 U18818 ( .B1(n21881), .B2(keyinput_108), .C1(keyinput_106), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n16918), .ZN(n16920) );
  XNOR2_X1 U18819 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_107), .ZN(
        n16919) );
  OAI211_X1 U18820 ( .C1(n16922), .C2(n16921), .A(n16920), .B(n16919), .ZN(
        n16927) );
  OAI22_X1 U18821 ( .A1(n16924), .A2(keyinput_109), .B1(keyinput_110), .B2(
        P1_FLUSH_REG_SCAN_IN), .ZN(n16923) );
  AOI221_X1 U18822 ( .B1(n16924), .B2(keyinput_109), .C1(P1_FLUSH_REG_SCAN_IN), 
        .C2(keyinput_110), .A(n16923), .ZN(n16926) );
  NOR2_X1 U18823 ( .A1(n20015), .A2(keyinput_111), .ZN(n16925) );
  AOI221_X1 U18824 ( .B1(n16927), .B2(n16926), .C1(keyinput_111), .C2(n20015), 
        .A(n16925), .ZN(n16928) );
  AOI221_X1 U18825 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_112), 
        .C1(n16930), .C2(n16929), .A(n16928), .ZN(n16938) );
  AOI22_X1 U18826 ( .A1(n19875), .A2(keyinput_113), .B1(n19868), .B2(
        keyinput_114), .ZN(n16931) );
  OAI221_X1 U18827 ( .B1(n19875), .B2(keyinput_113), .C1(n19868), .C2(
        keyinput_114), .A(n16931), .ZN(n16937) );
  OAI22_X1 U18828 ( .A1(n16933), .A2(keyinput_118), .B1(n15297), .B2(
        keyinput_117), .ZN(n16932) );
  AOI221_X1 U18829 ( .B1(n16933), .B2(keyinput_118), .C1(keyinput_117), .C2(
        n15297), .A(n16932), .ZN(n16936) );
  OAI22_X1 U18830 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_116), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_115), .ZN(n16934) );
  AOI221_X1 U18831 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_116), .C1(
        keyinput_115), .C2(P1_BYTEENABLE_REG_3__SCAN_IN), .A(n16934), .ZN(
        n16935) );
  OAI211_X1 U18832 ( .C1(n16938), .C2(n16937), .A(n16936), .B(n16935), .ZN(
        n16939) );
  OAI221_X1 U18833 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n16940), .C1(n15330), 
        .C2(keyinput_119), .A(n16939), .ZN(n16941) );
  OAI221_X1 U18834 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n16943), .C1(n16942), 
        .C2(keyinput_120), .A(n16941), .ZN(n16946) );
  AOI22_X1 U18835 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_124), .B1(
        n21582), .B2(keyinput_123), .ZN(n16944) );
  OAI221_X1 U18836 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_124), .C1(
        n21582), .C2(keyinput_123), .A(n16944), .ZN(n16945) );
  AOI21_X1 U18837 ( .B1(n16947), .B2(n16946), .A(n16945), .ZN(n16951) );
  XOR2_X1 U18838 ( .A(n15655), .B(keyinput_127), .Z(n16950) );
  AOI22_X1 U18839 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_125), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_126), .ZN(n16948) );
  OAI221_X1 U18840 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_125), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_126), .A(n16948), .ZN(n16949)
         );
  NOR4_X1 U18841 ( .A1(n16952), .A2(n16951), .A3(n16950), .A4(n16949), .ZN(
        n16963) );
  AOI21_X1 U18842 ( .B1(n16953), .B2(n16955), .A(n16954), .ZN(n21234) );
  INV_X1 U18843 ( .A(n21234), .ZN(n16961) );
  AOI22_X1 U18844 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13790), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n16956) );
  OAI21_X1 U18845 ( .B1(n19964), .B2(n16957), .A(n16956), .ZN(n16958) );
  AOI21_X1 U18846 ( .B1(n16959), .B2(n19952), .A(n16958), .ZN(n16960) );
  OAI21_X1 U18847 ( .B1(n16961), .B2(n21610), .A(n16960), .ZN(n16962) );
  XOR2_X1 U18848 ( .A(n16963), .B(n16962), .Z(P1_U2997) );
  INV_X1 U18849 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n16964) );
  OAI22_X1 U18850 ( .A1(n16965), .A2(n16964), .B1(n18511), .B2(n18518), .ZN(
        P2_U2816) );
  OAI21_X1 U18851 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16967), .A(
        n16966), .ZN(n18086) );
  AOI22_X1 U18852 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17031), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n16539), .ZN(n16973) );
  OAI22_X1 U18853 ( .A1(n16969), .A2(n17024), .B1(n17014), .B2(n16968), .ZN(
        n16970) );
  AOI21_X1 U18854 ( .B1(n17021), .B2(n16971), .A(n16970), .ZN(n16972) );
  OAI211_X1 U18855 ( .C1(n17042), .C2(n18086), .A(n16973), .B(n16972), .ZN(
        P2_U3009) );
  AOI21_X1 U18856 ( .B1(n18107), .B2(n16975), .A(n16974), .ZN(n18119) );
  AOI22_X1 U18857 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16539), .B1(n17005), 
        .B2(n18119), .ZN(n16983) );
  XOR2_X1 U18858 ( .A(n16977), .B(n16976), .Z(n18482) );
  INV_X1 U18859 ( .A(n18117), .ZN(n18480) );
  NOR2_X1 U18860 ( .A1(n16980), .A2(n16979), .ZN(n16981) );
  XNOR2_X1 U18861 ( .A(n16978), .B(n16981), .ZN(n18479) );
  AOI222_X1 U18862 ( .A1(n18482), .A2(n17035), .B1(n17021), .B2(n18480), .C1(
        n17032), .C2(n18479), .ZN(n16982) );
  OAI211_X1 U18863 ( .C1(n18107), .C2(n17018), .A(n16983), .B(n16982), .ZN(
        P2_U3006) );
  OAI21_X1 U18864 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16985), .A(
        n16984), .ZN(n18147) );
  AOI22_X1 U18865 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17031), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16539), .ZN(n16997) );
  NAND2_X1 U18866 ( .A1(n16987), .A2(n16986), .ZN(n16992) );
  INV_X1 U18867 ( .A(n16989), .ZN(n16990) );
  NOR2_X1 U18868 ( .A1(n16988), .A2(n16990), .ZN(n16991) );
  XOR2_X1 U18869 ( .A(n16992), .B(n16991), .Z(n18442) );
  INV_X1 U18870 ( .A(n18139), .ZN(n18441) );
  AOI21_X1 U18871 ( .B1(n16995), .B2(n16994), .A(n16993), .ZN(n18440) );
  AOI222_X1 U18872 ( .A1(n18442), .A2(n17032), .B1(n17021), .B2(n18441), .C1(
        n17035), .C2(n18440), .ZN(n16996) );
  OAI211_X1 U18873 ( .C1(n17042), .C2(n18147), .A(n16997), .B(n16996), .ZN(
        P2_U3004) );
  OAI21_X1 U18874 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11023), .A(
        n17004), .ZN(n18169) );
  AOI22_X1 U18875 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17031), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n16539), .ZN(n17003) );
  NAND2_X1 U18876 ( .A1(n16999), .A2(n16998), .ZN(n17000) );
  XNOR2_X1 U18877 ( .A(n17001), .B(n17000), .ZN(n18469) );
  INV_X1 U18878 ( .A(n18162), .ZN(n18468) );
  XOR2_X1 U18879 ( .A(n12702), .B(n17007), .Z(n18467) );
  AOI222_X1 U18880 ( .A1(n18469), .A2(n17032), .B1(n17021), .B2(n18468), .C1(
        n18467), .C2(n17035), .ZN(n17002) );
  OAI211_X1 U18881 ( .C1(n17042), .C2(n18169), .A(n17003), .B(n17002), .ZN(
        P2_U3002) );
  AOI21_X1 U18882 ( .B1(n18163), .B2(n17004), .A(n17020), .ZN(n18172) );
  AOI22_X1 U18883 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16539), .B1(n17005), 
        .B2(n18172), .ZN(n17017) );
  INV_X1 U18884 ( .A(n17006), .ZN(n17009) );
  OAI21_X1 U18885 ( .B1(n17007), .B2(n12702), .A(n18457), .ZN(n17008) );
  NAND2_X1 U18886 ( .A1(n17009), .A2(n17008), .ZN(n18452) );
  OAI21_X1 U18887 ( .B1(n17012), .B2(n17011), .A(n17010), .ZN(n17013) );
  INV_X1 U18888 ( .A(n17013), .ZN(n18451) );
  OAI22_X1 U18889 ( .A1(n18452), .A2(n17024), .B1(n18451), .B2(n17014), .ZN(
        n17015) );
  AOI21_X1 U18890 ( .B1(n17021), .B2(n18454), .A(n17015), .ZN(n17016) );
  OAI211_X1 U18891 ( .C1(n18163), .C2(n17018), .A(n17017), .B(n17016), .ZN(
        P2_U3001) );
  OAI21_X1 U18892 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17020), .A(
        n17019), .ZN(n18178) );
  AOI22_X1 U18893 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17031), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16539), .ZN(n17028) );
  AOI22_X1 U18894 ( .A1(n17022), .A2(n17032), .B1(n17021), .B2(n18186), .ZN(
        n17023) );
  OAI21_X1 U18895 ( .B1(n17025), .B2(n17024), .A(n17023), .ZN(n17026) );
  INV_X1 U18896 ( .A(n17026), .ZN(n17027) );
  OAI211_X1 U18897 ( .C1(n17042), .C2(n18178), .A(n17028), .B(n17027), .ZN(
        P2_U3000) );
  OAI21_X1 U18898 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17030), .A(
        n17029), .ZN(n18287) );
  AOI22_X1 U18899 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17031), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n16539), .ZN(n17041) );
  NAND2_X1 U18900 ( .A1(n17033), .A2(n17032), .ZN(n17037) );
  NAND3_X1 U18901 ( .A1(n16305), .A2(n17035), .A3(n17034), .ZN(n17036) );
  OAI211_X1 U18902 ( .C1(n17038), .C2(n18284), .A(n17037), .B(n17036), .ZN(
        n17039) );
  INV_X1 U18903 ( .A(n17039), .ZN(n17040) );
  OAI211_X1 U18904 ( .C1(n17042), .C2(n18287), .A(n17041), .B(n17040), .ZN(
        P2_U2992) );
  INV_X1 U18905 ( .A(n17043), .ZN(n18019) );
  OAI22_X1 U18906 ( .A1(n19034), .A2(n18019), .B1(n19164), .B2(n17044), .ZN(
        n17045) );
  AOI21_X1 U18907 ( .B1(n19146), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17045), 
        .ZN(n17046) );
  OAI22_X1 U18908 ( .A1(n19146), .A2(n17062), .B1(n17064), .B2(n17046), .ZN(
        P2_U3605) );
  AND2_X1 U18909 ( .A1(n19035), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17047) );
  NAND2_X1 U18910 ( .A1(n19142), .A2(n17047), .ZN(n19169) );
  INV_X1 U18911 ( .A(n19169), .ZN(n17050) );
  INV_X1 U18912 ( .A(n17047), .ZN(n19107) );
  NAND2_X1 U18913 ( .A1(n19107), .A2(n19200), .ZN(n17052) );
  NAND2_X1 U18914 ( .A1(n18511), .A2(n17052), .ZN(n17061) );
  INV_X1 U18915 ( .A(n17061), .ZN(n17048) );
  OAI22_X1 U18916 ( .A1(n19142), .A2(n17048), .B1(n18491), .B2(n19183), .ZN(
        n17049) );
  AOI21_X1 U18917 ( .B1(n19200), .B2(n17050), .A(n17049), .ZN(n17051) );
  AOI22_X1 U18918 ( .A1(n17064), .A2(n19160), .B1(n17051), .B2(n17062), .ZN(
        P2_U3603) );
  AOI21_X1 U18919 ( .B1(n19049), .B2(n21639), .A(n17052), .ZN(n17054) );
  OAI22_X1 U18920 ( .A1(n19049), .A2(n18511), .B1(n18425), .B2(n19183), .ZN(
        n17053) );
  NOR2_X1 U18921 ( .A1(n17054), .A2(n17053), .ZN(n17055) );
  AOI22_X1 U18922 ( .A1(n17064), .A2(n19179), .B1(n17055), .B2(n17062), .ZN(
        P2_U3604) );
  NOR2_X1 U18923 ( .A1(n17056), .A2(n19183), .ZN(n17060) );
  INV_X1 U18924 ( .A(n19131), .ZN(n17057) );
  NAND2_X1 U18925 ( .A1(n17057), .A2(n19035), .ZN(n17058) );
  AOI211_X1 U18926 ( .C1(n17058), .C2(n19083), .A(n13500), .B(n21639), .ZN(
        n17059) );
  AOI211_X1 U18927 ( .C1(n17061), .C2(n19170), .A(n17060), .B(n17059), .ZN(
        n17063) );
  AOI22_X1 U18928 ( .A1(n17064), .A2(n19159), .B1(n17063), .B2(n17062), .ZN(
        P2_U3602) );
  NAND2_X1 U18929 ( .A1(n17065), .A2(n21641), .ZN(n17068) );
  OAI21_X1 U18930 ( .B1(n11901), .B2(n11137), .A(n17072), .ZN(n17066) );
  OAI21_X1 U18931 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17072), .A(n17066), 
        .ZN(n17067) );
  OAI221_X1 U18932 ( .B1(n17068), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17068), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17067), .ZN(P2_U2822) );
  INV_X1 U18933 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17071) );
  OAI221_X1 U18934 ( .B1(n17072), .B2(n17071), .C1(n17070), .C2(n17069), .A(
        n17068), .ZN(P2_U2823) );
  OAI22_X1 U18935 ( .A1(n21666), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17128), .ZN(n17073) );
  INV_X1 U18936 ( .A(n17073), .ZN(P2_U3611) );
  INV_X1 U18937 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17074) );
  AOI22_X1 U18938 ( .A1(n17128), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17074), 
        .B2(n21666), .ZN(P2_U3608) );
  AOI21_X1 U18939 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21642), .ZN(n17075) );
  INV_X1 U18940 ( .A(n17075), .ZN(P2_U2815) );
  AOI22_X1 U18941 ( .A1(n17108), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17077) );
  OAI21_X1 U18942 ( .B1(n13754), .B2(n17110), .A(n17077), .ZN(P2_U2951) );
  AOI22_X1 U18943 ( .A1(n17108), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17078) );
  OAI21_X1 U18944 ( .B1(n17079), .B2(n17110), .A(n17078), .ZN(P2_U2950) );
  INV_X1 U18945 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U18946 ( .A1(n17108), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17080) );
  OAI21_X1 U18947 ( .B1(n17081), .B2(n17110), .A(n17080), .ZN(P2_U2949) );
  INV_X1 U18948 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U18949 ( .A1(n17096), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17082) );
  OAI21_X1 U18950 ( .B1(n17083), .B2(n17110), .A(n17082), .ZN(P2_U2948) );
  INV_X1 U18951 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U18952 ( .A1(n17108), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17084) );
  OAI21_X1 U18953 ( .B1(n17085), .B2(n17110), .A(n17084), .ZN(P2_U2947) );
  INV_X1 U18954 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19277) );
  AOI22_X1 U18955 ( .A1(n17096), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17086) );
  OAI21_X1 U18956 ( .B1(n19277), .B2(n17110), .A(n17086), .ZN(P2_U2946) );
  AOI22_X1 U18957 ( .A1(n17096), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17087) );
  OAI21_X1 U18958 ( .B1(n17088), .B2(n17110), .A(n17087), .ZN(P2_U2945) );
  AOI22_X1 U18959 ( .A1(n17096), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17089) );
  OAI21_X1 U18960 ( .B1(n17090), .B2(n17110), .A(n17089), .ZN(P2_U2944) );
  AOI22_X1 U18961 ( .A1(n17096), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17091) );
  OAI21_X1 U18962 ( .B1(n17092), .B2(n17110), .A(n17091), .ZN(P2_U2943) );
  AOI22_X1 U18963 ( .A1(n17108), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17093) );
  OAI21_X1 U18964 ( .B1(n17094), .B2(n17110), .A(n17093), .ZN(P2_U2942) );
  AOI22_X1 U18965 ( .A1(n17096), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17095), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17097) );
  OAI21_X1 U18966 ( .B1(n17098), .B2(n17110), .A(n17097), .ZN(P2_U2941) );
  AOI22_X1 U18967 ( .A1(n17108), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17099) );
  OAI21_X1 U18968 ( .B1(n17100), .B2(n17110), .A(n17099), .ZN(P2_U2940) );
  AOI22_X1 U18969 ( .A1(n17108), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17101) );
  OAI21_X1 U18970 ( .B1(n17102), .B2(n17110), .A(n17101), .ZN(P2_U2939) );
  AOI22_X1 U18971 ( .A1(n17108), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17103) );
  OAI21_X1 U18972 ( .B1(n17104), .B2(n17110), .A(n17103), .ZN(P2_U2938) );
  AOI22_X1 U18973 ( .A1(n17108), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17105) );
  OAI21_X1 U18974 ( .B1(n17106), .B2(n17110), .A(n17105), .ZN(P2_U2937) );
  AOI22_X1 U18975 ( .A1(n17108), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17107), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17109) );
  OAI21_X1 U18976 ( .B1(n17111), .B2(n17110), .A(n17109), .ZN(P2_U2936) );
  AOI21_X1 U18977 ( .B1(n21682), .B2(n21685), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17112) );
  AOI22_X1 U18978 ( .A1(n17128), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n17112), 
        .B2(n21666), .ZN(P2_U2817) );
  OAI222_X1 U18979 ( .A1(n17125), .A2(n11889), .B1(n17113), .B2(n17128), .C1(
        n11901), .C2(n17124), .ZN(P2_U3212) );
  INV_X1 U18980 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17114) );
  OAI222_X1 U18981 ( .A1(n17125), .A2(n14356), .B1(n17114), .B2(n17128), .C1(
        n11889), .C2(n17124), .ZN(P2_U3213) );
  INV_X1 U18982 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19725) );
  OAI222_X1 U18983 ( .A1(n17125), .A2(n12673), .B1(n19725), .B2(n17128), .C1(
        n14356), .C2(n17124), .ZN(P2_U3214) );
  INV_X1 U18984 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n17115) );
  OAI222_X1 U18985 ( .A1(n17125), .A2(n14547), .B1(n17115), .B2(n17128), .C1(
        n12673), .C2(n17124), .ZN(P2_U3215) );
  INV_X1 U18986 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n17116) );
  OAI222_X1 U18987 ( .A1(n17125), .A2(n12682), .B1(n17116), .B2(n17128), .C1(
        n14547), .C2(n17124), .ZN(P2_U3216) );
  INV_X1 U18988 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19729) );
  OAI222_X1 U18989 ( .A1(n17125), .A2(n18096), .B1(n19729), .B2(n17128), .C1(
        n12682), .C2(n17124), .ZN(P2_U3217) );
  INV_X1 U18990 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19731) );
  OAI222_X1 U18991 ( .A1(n17125), .A2(n12688), .B1(n19731), .B2(n17128), .C1(
        n18096), .C2(n17124), .ZN(P2_U3218) );
  INV_X1 U18992 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19733) );
  OAI222_X1 U18993 ( .A1(n17125), .A2(n12694), .B1(n19733), .B2(n17128), .C1(
        n12688), .C2(n17124), .ZN(P2_U3219) );
  INV_X1 U18994 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19735) );
  OAI222_X1 U18995 ( .A1(n17124), .A2(n12694), .B1(n19735), .B2(n17128), .C1(
        n18437), .C2(n17125), .ZN(P2_U3220) );
  INV_X1 U18996 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19737) );
  OAI222_X1 U18997 ( .A1(n17124), .A2(n18437), .B1(n19737), .B2(n17128), .C1(
        n16417), .C2(n17125), .ZN(P2_U3221) );
  INV_X1 U18998 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19739) );
  INV_X1 U18999 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n18462) );
  OAI222_X1 U19000 ( .A1(n17124), .A2(n16417), .B1(n19739), .B2(n17128), .C1(
        n18462), .C2(n17125), .ZN(P2_U3222) );
  INV_X1 U19001 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19741) );
  OAI222_X1 U19002 ( .A1(n17124), .A2(n18462), .B1(n19741), .B2(n17128), .C1(
        n12706), .C2(n17125), .ZN(P2_U3223) );
  INV_X1 U19003 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19743) );
  OAI222_X1 U19004 ( .A1(n17124), .A2(n12706), .B1(n19743), .B2(n17128), .C1(
        n12714), .C2(n17125), .ZN(P2_U3224) );
  INV_X1 U19005 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19745) );
  OAI222_X1 U19006 ( .A1(n17124), .A2(n12714), .B1(n19745), .B2(n17128), .C1(
        n18191), .C2(n17125), .ZN(P2_U3225) );
  INV_X1 U19007 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19747) );
  OAI222_X1 U19008 ( .A1(n17124), .A2(n18191), .B1(n19747), .B2(n17128), .C1(
        n12721), .C2(n17125), .ZN(P2_U3226) );
  INV_X1 U19009 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19749) );
  OAI222_X1 U19010 ( .A1(n17124), .A2(n12721), .B1(n19749), .B2(n17128), .C1(
        n18219), .C2(n17125), .ZN(P2_U3227) );
  INV_X1 U19011 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19751) );
  OAI222_X1 U19012 ( .A1(n17124), .A2(n18219), .B1(n19751), .B2(n17128), .C1(
        n17117), .C2(n17125), .ZN(P2_U3228) );
  INV_X1 U19013 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19753) );
  OAI222_X1 U19014 ( .A1(n17125), .A2(n18242), .B1(n19753), .B2(n17128), .C1(
        n17117), .C2(n17124), .ZN(P2_U3229) );
  INV_X1 U19015 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19755) );
  OAI222_X1 U19016 ( .A1(n17124), .A2(n18242), .B1(n19755), .B2(n17128), .C1(
        n16342), .C2(n17125), .ZN(P2_U3230) );
  INV_X1 U19017 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19757) );
  OAI222_X1 U19018 ( .A1(n17125), .A2(n17118), .B1(n19757), .B2(n17128), .C1(
        n16342), .C2(n17124), .ZN(P2_U3231) );
  INV_X1 U19019 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19759) );
  OAI222_X1 U19020 ( .A1(n17125), .A2(n12737), .B1(n19759), .B2(n17128), .C1(
        n17118), .C2(n17124), .ZN(P2_U3232) );
  INV_X1 U19021 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19761) );
  OAI222_X1 U19022 ( .A1(n17125), .A2(n18294), .B1(n19761), .B2(n17128), .C1(
        n12737), .C2(n17124), .ZN(P2_U3233) );
  INV_X1 U19023 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19763) );
  OAI222_X1 U19024 ( .A1(n17125), .A2(n17119), .B1(n19763), .B2(n17128), .C1(
        n18294), .C2(n17124), .ZN(P2_U3234) );
  INV_X1 U19025 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19765) );
  OAI222_X1 U19026 ( .A1(n17125), .A2(n17120), .B1(n19765), .B2(n17128), .C1(
        n17119), .C2(n17124), .ZN(P2_U3235) );
  INV_X1 U19027 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19767) );
  OAI222_X1 U19028 ( .A1(n17124), .A2(n17120), .B1(n19767), .B2(n17128), .C1(
        n16275), .C2(n17125), .ZN(P2_U3236) );
  INV_X1 U19029 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19769) );
  OAI222_X1 U19030 ( .A1(n17125), .A2(n18339), .B1(n19769), .B2(n17128), .C1(
        n16275), .C2(n17124), .ZN(P2_U3237) );
  INV_X1 U19031 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19771) );
  OAI222_X1 U19032 ( .A1(n17124), .A2(n18339), .B1(n19771), .B2(n17128), .C1(
        n16249), .C2(n17125), .ZN(P2_U3238) );
  INV_X1 U19033 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n17121) );
  OAI222_X1 U19034 ( .A1(n17124), .A2(n16249), .B1(n17121), .B2(n17128), .C1(
        n17123), .C2(n17125), .ZN(P2_U3239) );
  INV_X1 U19035 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n17122) );
  OAI222_X1 U19036 ( .A1(n17124), .A2(n17123), .B1(n17122), .B2(n17128), .C1(
        n16222), .C2(n17125), .ZN(P2_U3240) );
  INV_X1 U19037 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19777) );
  OAI222_X1 U19038 ( .A1(n17125), .A2(n18397), .B1(n19777), .B2(n17128), .C1(
        n16222), .C2(n17124), .ZN(P2_U3241) );
  OAI22_X1 U19039 ( .A1(n21666), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17128), .ZN(n17126) );
  INV_X1 U19040 ( .A(n17126), .ZN(P2_U3588) );
  OAI22_X1 U19041 ( .A1(n21666), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17128), .ZN(n17127) );
  INV_X1 U19042 ( .A(n17127), .ZN(P2_U3587) );
  MUX2_X1 U19043 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n21666), .Z(P2_U3586) );
  OAI22_X1 U19044 ( .A1(n21666), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17128), .ZN(n17129) );
  INV_X1 U19045 ( .A(n17129), .ZN(P2_U3585) );
  INV_X1 U19046 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20112) );
  INV_X1 U19047 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20099) );
  INV_X1 U19048 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20098) );
  NOR2_X1 U19049 ( .A1(n20099), .A2(n20098), .ZN(n17511) );
  NOR4_X1 U19050 ( .A1(n20625), .A2(n17131), .A3(n17130), .A4(n20723), .ZN(
        n17132) );
  AOI21_X1 U19051 ( .B1(n17133), .B2(n21127), .A(n17132), .ZN(n20522) );
  NOR4_X2 U19052 ( .A1(n18898), .A2(n20084), .A3(n20522), .A4(n21188), .ZN(
        n17519) );
  NOR2_X1 U19053 ( .A1(n20625), .A2(n17506), .ZN(n17516) );
  NAND3_X1 U19054 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17511), .A3(n17516), .ZN(
        n17136) );
  NOR2_X1 U19055 ( .A1(n20112), .A2(n17136), .ZN(n17138) );
  NAND2_X1 U19056 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17138), .ZN(n17160) );
  INV_X1 U19057 ( .A(n17160), .ZN(n17163) );
  NOR2_X2 U19058 ( .A1(n17506), .A2(n20597), .ZN(n17517) );
  AOI21_X1 U19059 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17513), .A(n17138), .ZN(
        n17135) );
  INV_X1 U19060 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17134) );
  OAI22_X1 U19061 ( .A1(n17163), .A2(n17135), .B1(n17134), .B2(n17513), .ZN(
        P3_U2699) );
  INV_X1 U19062 ( .A(n17136), .ZN(n17139) );
  AOI21_X1 U19063 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17513), .A(n17139), .ZN(
        n17137) );
  OAI22_X1 U19064 ( .A1(n17138), .A2(n17137), .B1(n17342), .B2(n17513), .ZN(
        P3_U2700) );
  INV_X1 U19065 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17141) );
  AOI221_X1 U19066 ( .B1(n17511), .B2(n17519), .C1(n20625), .C2(n17519), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17140) );
  AOI211_X1 U19067 ( .C1(n17517), .C2(n17141), .A(n17140), .B(n17139), .ZN(
        P3_U2701) );
  AOI22_X1 U19068 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U19069 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U19070 ( .A1(n11578), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17142) );
  OAI21_X1 U19071 ( .B1(n17261), .B2(n17143), .A(n17142), .ZN(n17149) );
  AOI22_X1 U19072 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U19073 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U19074 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U19075 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17144) );
  NAND4_X1 U19076 ( .A1(n17147), .A2(n17146), .A3(n17145), .A4(n17144), .ZN(
        n17148) );
  AOI211_X1 U19077 ( .C1(n10955), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n17149), .B(n17148), .ZN(n17150) );
  NAND3_X1 U19078 ( .A1(n17152), .A2(n17151), .A3(n17150), .ZN(n20693) );
  INV_X1 U19079 ( .A(n20693), .ZN(n17155) );
  INV_X1 U19080 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20170) );
  AND3_X1 U19081 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .A3(n17511), .ZN(n17153) );
  NAND4_X1 U19082 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(P3_EBX_REG_4__SCAN_IN), .A4(n17153), .ZN(n17156) );
  NOR2_X1 U19083 ( .A1(n20170), .A2(n17156), .ZN(n17166) );
  AND2_X1 U19084 ( .A1(n17519), .A2(n17166), .ZN(n17159) );
  NAND3_X1 U19085 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17519), .A3(n17166), .ZN(
        n17258) );
  OAI21_X1 U19086 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17159), .A(n17258), .ZN(
        n17154) );
  AOI22_X1 U19087 ( .A1(n17517), .A2(n17155), .B1(n17154), .B2(n17513), .ZN(
        P3_U2695) );
  INV_X1 U19088 ( .A(n17516), .ZN(n17515) );
  NOR2_X1 U19089 ( .A1(n17156), .A2(n17515), .ZN(n17162) );
  OAI21_X1 U19090 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17162), .A(n17513), .ZN(
        n17158) );
  OAI22_X1 U19091 ( .A1(n17159), .A2(n17158), .B1(n17157), .B2(n17513), .ZN(
        P3_U2696) );
  INV_X1 U19092 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20146) );
  NOR2_X1 U19093 ( .A1(n20146), .A2(n17160), .ZN(n17165) );
  AOI21_X1 U19094 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17513), .A(n17165), .ZN(
        n17161) );
  INV_X1 U19095 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17206) );
  OAI22_X1 U19096 ( .A1(n17162), .A2(n17161), .B1(n17206), .B2(n17513), .ZN(
        P3_U2697) );
  AOI21_X1 U19097 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17513), .A(n17163), .ZN(
        n17164) );
  OAI22_X1 U19098 ( .A1(n17165), .A2(n17164), .B1(n17353), .B2(n17513), .ZN(
        P3_U2698) );
  INV_X1 U19099 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20283) );
  INV_X1 U19100 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20273) );
  INV_X1 U19101 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20260) );
  NOR3_X1 U19102 ( .A1(n20283), .A2(n20273), .A3(n20260), .ZN(n17275) );
  INV_X1 U19103 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20243) );
  INV_X1 U19104 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20227) );
  NAND4_X1 U19105 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17166), .ZN(n17277) );
  NOR3_X1 U19106 ( .A1(n20227), .A2(n17506), .A3(n17277), .ZN(n17219) );
  NAND2_X1 U19107 ( .A1(n20597), .A2(n17219), .ZN(n17233) );
  NOR2_X1 U19108 ( .A1(n20243), .A2(n17233), .ZN(n17204) );
  NAND2_X1 U19109 ( .A1(n17275), .A2(n17204), .ZN(n17188) );
  AOI22_X1 U19110 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U19111 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10952), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U19112 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U19113 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17167) );
  NAND4_X1 U19114 ( .A1(n17170), .A2(n17169), .A3(n17168), .A4(n17167), .ZN(
        n17176) );
  AOI22_X1 U19115 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U19116 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U19117 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U19118 ( .A1(n11578), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17171) );
  NAND4_X1 U19119 ( .A1(n17174), .A2(n17173), .A3(n17172), .A4(n17171), .ZN(
        n17175) );
  NOR2_X1 U19120 ( .A1(n17176), .A2(n17175), .ZN(n20678) );
  NAND3_X1 U19121 ( .A1(n17188), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17513), 
        .ZN(n17177) );
  OAI221_X1 U19122 ( .B1(n17188), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17513), 
        .C2(n20678), .A(n17177), .ZN(P3_U2687) );
  AOI22_X1 U19123 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U19124 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U19125 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U19126 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17178) );
  NAND4_X1 U19127 ( .A1(n17181), .A2(n17180), .A3(n17179), .A4(n17178), .ZN(
        n17187) );
  AOI22_X1 U19128 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U19129 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U19130 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U19131 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17182) );
  NAND4_X1 U19132 ( .A1(n17185), .A2(n17184), .A3(n17183), .A4(n17182), .ZN(
        n17186) );
  NOR2_X1 U19133 ( .A1(n17187), .A2(n17186), .ZN(n20692) );
  NAND2_X1 U19134 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17219), .ZN(n17191) );
  NOR3_X1 U19135 ( .A1(n20273), .A2(n20260), .A3(n17191), .ZN(n17189) );
  OAI211_X1 U19136 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17189), .A(n17188), .B(
        n17513), .ZN(n17190) );
  OAI21_X1 U19137 ( .B1(n20692), .B2(n17513), .A(n17190), .ZN(P3_U2688) );
  NAND3_X1 U19138 ( .A1(n17513), .A2(P3_EBX_REG_13__SCAN_IN), .A3(n17191), 
        .ZN(n17203) );
  AOI22_X1 U19139 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U19140 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U19141 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17192) );
  OAI21_X1 U19142 ( .B1(n17261), .B2(n17353), .A(n17192), .ZN(n17198) );
  AOI22_X1 U19143 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U19144 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U19145 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U19146 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17193) );
  NAND4_X1 U19147 ( .A1(n17196), .A2(n17195), .A3(n17194), .A4(n17193), .ZN(
        n17197) );
  AOI211_X1 U19148 ( .C1(n17491), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17198), .B(n17197), .ZN(n17199) );
  NAND3_X1 U19149 ( .A1(n17201), .A2(n17200), .A3(n17199), .ZN(n20529) );
  AOI22_X1 U19150 ( .A1(n17517), .A2(n20529), .B1(n17204), .B2(n20260), .ZN(
        n17202) );
  NAND2_X1 U19151 ( .A1(n17203), .A2(n17202), .ZN(P3_U2690) );
  NAND2_X1 U19152 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17204), .ZN(n17218) );
  AOI22_X1 U19153 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U19154 ( .A1(n17435), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U19155 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U19156 ( .B1(n17261), .B2(n17206), .A(n17205), .ZN(n17212) );
  AOI22_X1 U19157 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U19158 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U19159 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U19160 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17207) );
  NAND4_X1 U19161 ( .A1(n17210), .A2(n17209), .A3(n17208), .A4(n17207), .ZN(
        n17211) );
  AOI211_X1 U19162 ( .C1(n17262), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17212), .B(n17211), .ZN(n17213) );
  NAND3_X1 U19163 ( .A1(n17215), .A2(n17214), .A3(n17213), .ZN(n20680) );
  INV_X1 U19164 ( .A(n20680), .ZN(n17217) );
  NAND3_X1 U19165 ( .A1(n17218), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17513), 
        .ZN(n17216) );
  OAI221_X1 U19166 ( .B1(n17218), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17513), 
        .C2(n17217), .A(n17216), .ZN(P3_U2689) );
  NOR2_X1 U19167 ( .A1(n17517), .A2(n17219), .ZN(n17244) );
  AOI22_X1 U19168 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U19169 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U19170 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U19171 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17221) );
  NAND4_X1 U19172 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17230) );
  AOI22_X1 U19173 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U19174 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U19175 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U19176 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17225) );
  NAND4_X1 U19177 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17229) );
  NOR2_X1 U19178 ( .A1(n17230), .A2(n17229), .ZN(n20533) );
  INV_X1 U19179 ( .A(n20533), .ZN(n17231) );
  AOI22_X1 U19180 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17244), .B1(n17517), 
        .B2(n17231), .ZN(n17232) );
  OAI21_X1 U19181 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17233), .A(n17232), .ZN(
        P3_U2691) );
  AOI22_X1 U19182 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U19183 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U19184 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U19185 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17234) );
  NAND4_X1 U19186 ( .A1(n17237), .A2(n17236), .A3(n17235), .A4(n17234), .ZN(
        n17243) );
  AOI22_X1 U19187 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U19188 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U19189 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U19190 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17238) );
  NAND4_X1 U19191 ( .A1(n17241), .A2(n17240), .A3(n17239), .A4(n17238), .ZN(
        n17242) );
  NOR2_X1 U19192 ( .A1(n17243), .A2(n17242), .ZN(n20538) );
  NOR2_X1 U19193 ( .A1(n17506), .A2(n17277), .ZN(n17245) );
  OAI21_X1 U19194 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17245), .A(n17244), .ZN(
        n17246) );
  OAI21_X1 U19195 ( .B1(n20538), .B2(n17513), .A(n17246), .ZN(P3_U2692) );
  AOI22_X1 U19196 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U19197 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U19198 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U19199 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17247) );
  NAND4_X1 U19200 ( .A1(n17250), .A2(n17249), .A3(n17248), .A4(n17247), .ZN(
        n17256) );
  AOI22_X1 U19201 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U19202 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U19203 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U19204 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17251) );
  NAND4_X1 U19205 ( .A1(n17254), .A2(n17253), .A3(n17252), .A4(n17251), .ZN(
        n17255) );
  NOR2_X1 U19206 ( .A1(n17256), .A2(n17255), .ZN(n20545) );
  INV_X1 U19207 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20192) );
  NOR2_X1 U19208 ( .A1(n20192), .A2(n17258), .ZN(n17274) );
  OAI22_X1 U19209 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17274), .B1(n17277), 
        .B2(n17506), .ZN(n17257) );
  AOI22_X1 U19210 ( .A1(n17517), .A2(n20545), .B1(n17257), .B2(n17513), .ZN(
        P3_U2693) );
  INV_X1 U19211 ( .A(n17258), .ZN(n17259) );
  OAI21_X1 U19212 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17259), .A(n17513), .ZN(
        n17273) );
  AOI22_X1 U19213 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10960), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U19214 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U19215 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U19216 ( .B1(n17261), .B2(n17514), .A(n17260), .ZN(n17268) );
  AOI22_X1 U19217 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U19218 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n10953), .ZN(n17265) );
  AOI22_X1 U19219 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10948), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17457), .ZN(n17264) );
  AOI22_X1 U19220 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17492), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17475), .ZN(n17263) );
  NAND4_X1 U19221 ( .A1(n17266), .A2(n17265), .A3(n17264), .A4(n17263), .ZN(
        n17267) );
  AOI211_X1 U19222 ( .C1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .C2(n17300), .A(
        n17268), .B(n17267), .ZN(n17269) );
  NAND3_X1 U19223 ( .A1(n17271), .A2(n17270), .A3(n17269), .ZN(n20549) );
  INV_X1 U19224 ( .A(n20549), .ZN(n17272) );
  OAI22_X1 U19225 ( .A1(n17274), .A2(n17273), .B1(n17272), .B2(n17513), .ZN(
        P3_U2694) );
  INV_X1 U19226 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20471) );
  INV_X1 U19227 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20346) );
  NAND4_X1 U19228 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(n17275), .ZN(n17276) );
  NOR2_X1 U19229 ( .A1(n17277), .A2(n17276), .ZN(n17508) );
  NAND2_X1 U19230 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17508), .ZN(n17507) );
  NOR2_X1 U19231 ( .A1(n17506), .A2(n17507), .ZN(n17470) );
  NAND2_X1 U19232 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17470), .ZN(n17472) );
  NAND2_X1 U19233 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17490), .ZN(n17389) );
  AND2_X1 U19234 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .ZN(n17278) );
  AND4_X1 U19235 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n17391)
         );
  NAND4_X1 U19236 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17278), .A4(n17391), .ZN(n17395) );
  NOR3_X1 U19237 ( .A1(n20471), .A2(n17389), .A3(n17395), .ZN(n17376) );
  NAND2_X1 U19238 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17376), .ZN(n17375) );
  INV_X1 U19239 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20499) );
  INV_X1 U19240 ( .A(n17375), .ZN(n17279) );
  OAI33_X1 U19241 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20625), .A3(n17375), 
        .B1(n20499), .B2(n17517), .B3(n17279), .ZN(P3_U2672) );
  AOI22_X1 U19242 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U19243 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U19244 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U19245 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U19246 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17289) );
  AOI22_X1 U19247 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U19248 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U19249 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U19250 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U19251 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  NOR2_X1 U19252 ( .A1(n17289), .A2(n17288), .ZN(n17398) );
  AOI22_X1 U19253 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U19254 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U19255 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U19256 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17290) );
  NAND4_X1 U19257 ( .A1(n17293), .A2(n17292), .A3(n17291), .A4(n17290), .ZN(
        n17299) );
  AOI22_X1 U19258 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U19259 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10952), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U19260 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U19261 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17294) );
  NAND4_X1 U19262 ( .A1(n17297), .A2(n17296), .A3(n17295), .A4(n17294), .ZN(
        n17298) );
  NOR2_X1 U19263 ( .A1(n17299), .A2(n17298), .ZN(n17392) );
  AOI22_X1 U19264 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U19265 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17300), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U19266 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U19267 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17301) );
  NAND4_X1 U19268 ( .A1(n17304), .A2(n17303), .A3(n17302), .A4(n17301), .ZN(
        n17310) );
  AOI22_X1 U19269 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U19270 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U19271 ( .A1(n10956), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U19272 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17305) );
  NAND4_X1 U19273 ( .A1(n17308), .A2(n17307), .A3(n17306), .A4(n17305), .ZN(
        n17309) );
  NOR2_X1 U19274 ( .A1(n17310), .A2(n17309), .ZN(n17416) );
  AOI22_X1 U19275 ( .A1(n11578), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U19276 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U19277 ( .A1(n10948), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U19278 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17311) );
  NAND4_X1 U19279 ( .A1(n17314), .A2(n17313), .A3(n17312), .A4(n17311), .ZN(
        n17320) );
  AOI22_X1 U19280 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U19281 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U19282 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U19283 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17315) );
  NAND4_X1 U19284 ( .A1(n17318), .A2(n17317), .A3(n17316), .A4(n17315), .ZN(
        n17319) );
  NOR2_X1 U19285 ( .A1(n17320), .A2(n17319), .ZN(n17425) );
  AOI22_X1 U19286 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U19287 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U19288 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U19289 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17321) );
  NAND4_X1 U19290 ( .A1(n17324), .A2(n17323), .A3(n17322), .A4(n17321), .ZN(
        n17330) );
  AOI22_X1 U19291 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10965), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U19292 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U19293 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U19294 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17325) );
  NAND4_X1 U19295 ( .A1(n17328), .A2(n17327), .A3(n17326), .A4(n17325), .ZN(
        n17329) );
  NOR2_X1 U19296 ( .A1(n17330), .A2(n17329), .ZN(n17426) );
  NOR2_X1 U19297 ( .A1(n17425), .A2(n17426), .ZN(n17424) );
  AOI22_X1 U19298 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10976), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n11578), .ZN(n17340) );
  AOI22_X1 U19299 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17498), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n10953), .ZN(n17339) );
  AOI22_X1 U19300 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17491), .B1(
        n17499), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17331) );
  OAI21_X1 U19301 ( .B1(n17354), .B2(n17514), .A(n17331), .ZN(n17337) );
  AOI22_X1 U19302 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17444), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n10974), .ZN(n17335) );
  AOI22_X1 U19303 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10956), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U19304 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17457), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17474), .ZN(n17333) );
  AOI22_X1 U19305 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17492), .ZN(n17332) );
  NAND4_X1 U19306 ( .A1(n17335), .A2(n17334), .A3(n17333), .A4(n17332), .ZN(
        n17336) );
  AOI211_X1 U19307 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n17337), .B(n17336), .ZN(n17338) );
  NAND3_X1 U19308 ( .A1(n17340), .A2(n17339), .A3(n17338), .ZN(n17421) );
  NAND2_X1 U19309 ( .A1(n17424), .A2(n17421), .ZN(n17420) );
  NOR2_X1 U19310 ( .A1(n17416), .A2(n17420), .ZN(n17415) );
  AOI22_X1 U19311 ( .A1(n10974), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U19312 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U19313 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17341) );
  OAI21_X1 U19314 ( .B1(n17354), .B2(n17342), .A(n17341), .ZN(n17348) );
  AOI22_X1 U19315 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U19316 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U19317 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U19318 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17343) );
  NAND4_X1 U19319 ( .A1(n17346), .A2(n17345), .A3(n17344), .A4(n17343), .ZN(
        n17347) );
  AOI211_X1 U19320 ( .C1(n17491), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17348), .B(n17347), .ZN(n17349) );
  NAND3_X1 U19321 ( .A1(n17351), .A2(n17350), .A3(n17349), .ZN(n17411) );
  NAND2_X1 U19322 ( .A1(n17415), .A2(n17411), .ZN(n17410) );
  NOR2_X1 U19323 ( .A1(n17392), .A2(n17410), .ZN(n17404) );
  AOI22_X1 U19324 ( .A1(n11578), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U19325 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17463), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U19326 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17352) );
  OAI21_X1 U19327 ( .B1(n17354), .B2(n17353), .A(n17352), .ZN(n17360) );
  AOI22_X1 U19328 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U19329 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U19330 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U19331 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17355) );
  NAND4_X1 U19332 ( .A1(n17358), .A2(n17357), .A3(n17356), .A4(n17355), .ZN(
        n17359) );
  AOI211_X1 U19333 ( .C1(n10957), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17360), .B(n17359), .ZN(n17361) );
  NAND3_X1 U19334 ( .A1(n17363), .A2(n17362), .A3(n17361), .ZN(n17403) );
  NAND2_X1 U19335 ( .A1(n17404), .A2(n17403), .ZN(n17402) );
  NOR2_X1 U19336 ( .A1(n17398), .A2(n17402), .ZN(n17397) );
  AOI22_X1 U19337 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U19338 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U19339 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U19340 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17364) );
  NAND4_X1 U19341 ( .A1(n17367), .A2(n17366), .A3(n17365), .A4(n17364), .ZN(
        n17373) );
  AOI22_X1 U19342 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U19343 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U19344 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U19345 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17368) );
  NAND4_X1 U19346 ( .A1(n17371), .A2(n17370), .A3(n17369), .A4(n17368), .ZN(
        n17372) );
  NOR2_X1 U19347 ( .A1(n17373), .A2(n17372), .ZN(n17374) );
  XOR2_X1 U19348 ( .A(n17397), .B(n17374), .Z(n20641) );
  OAI211_X1 U19349 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17376), .A(n17375), .B(
        n17513), .ZN(n17377) );
  OAI21_X1 U19350 ( .B1(n20641), .B2(n17513), .A(n17377), .ZN(P3_U2673) );
  AOI22_X1 U19351 ( .A1(n17463), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U19352 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U19353 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17378), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U19354 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17379) );
  NAND4_X1 U19355 ( .A1(n17382), .A2(n17381), .A3(n17380), .A4(n17379), .ZN(
        n17388) );
  AOI22_X1 U19356 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U19357 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U19358 ( .A1(n10957), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U19359 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U19360 ( .A1(n17386), .A2(n17385), .A3(n17384), .A4(n17383), .ZN(
        n17387) );
  NOR2_X1 U19361 ( .A1(n17388), .A2(n17387), .ZN(n20588) );
  AND2_X1 U19362 ( .A1(n17513), .A2(n17389), .ZN(n17455) );
  NOR2_X1 U19363 ( .A1(n20625), .A2(n17389), .ZN(n17430) );
  INV_X1 U19364 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20372) );
  AOI22_X1 U19365 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17455), .B1(n17430), 
        .B2(n20372), .ZN(n17390) );
  OAI21_X1 U19366 ( .B1(n20588), .B2(n17513), .A(n17390), .ZN(P3_U2682) );
  NAND3_X1 U19367 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17430), .ZN(n17429) );
  NAND2_X1 U19368 ( .A1(n17443), .A2(n17391), .ZN(n17409) );
  AOI21_X1 U19369 ( .B1(n17392), .B2(n17410), .A(n17404), .ZN(n20658) );
  INV_X1 U19370 ( .A(n20658), .ZN(n17394) );
  NAND3_X1 U19371 ( .A1(n17409), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17513), 
        .ZN(n17393) );
  OAI221_X1 U19372 ( .B1(n17409), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17513), 
        .C2(n17394), .A(n17393), .ZN(P3_U2676) );
  INV_X1 U19373 ( .A(n17430), .ZN(n17396) );
  NOR2_X1 U19374 ( .A1(n17396), .A2(n17395), .ZN(n17399) );
  NOR2_X1 U19375 ( .A1(n17517), .A2(n17399), .ZN(n17407) );
  INV_X1 U19376 ( .A(n17407), .ZN(n17401) );
  AOI21_X1 U19377 ( .B1(n17398), .B2(n17402), .A(n17397), .ZN(n20646) );
  AOI22_X1 U19378 ( .A1(n17517), .A2(n20646), .B1(n17399), .B2(n20471), .ZN(
        n17400) );
  OAI21_X1 U19379 ( .B1(n20471), .B2(n17401), .A(n17400), .ZN(P3_U2674) );
  OAI21_X1 U19380 ( .B1(n17404), .B2(n17403), .A(n17402), .ZN(n20652) );
  INV_X1 U19381 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20449) );
  NOR2_X1 U19382 ( .A1(n20449), .A2(n17409), .ZN(n17406) );
  INV_X1 U19383 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U19384 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17407), .B1(n17406), 
        .B2(n17405), .ZN(n17408) );
  OAI21_X1 U19385 ( .B1(n20652), .B2(n17513), .A(n17408), .ZN(P3_U2675) );
  INV_X1 U19386 ( .A(n17409), .ZN(n17413) );
  INV_X1 U19387 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20417) );
  NAND3_X1 U19388 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n17443), .ZN(n17414) );
  NOR2_X1 U19389 ( .A1(n20417), .A2(n17414), .ZN(n17419) );
  AOI21_X1 U19390 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17513), .A(n17419), .ZN(
        n17412) );
  OAI21_X1 U19391 ( .B1(n17415), .B2(n17411), .A(n17410), .ZN(n20635) );
  OAI22_X1 U19392 ( .A1(n17413), .A2(n17412), .B1(n20635), .B2(n17513), .ZN(
        P3_U2677) );
  INV_X1 U19393 ( .A(n17414), .ZN(n17423) );
  AOI21_X1 U19394 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17513), .A(n17423), .ZN(
        n17418) );
  AOI21_X1 U19395 ( .B1(n17416), .B2(n17420), .A(n17415), .ZN(n20622) );
  INV_X1 U19396 ( .A(n20622), .ZN(n17417) );
  OAI22_X1 U19397 ( .A1(n17419), .A2(n17418), .B1(n17417), .B2(n17513), .ZN(
        P3_U2678) );
  AOI22_X1 U19398 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17513), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n17443), .ZN(n17422) );
  OAI21_X1 U19399 ( .B1(n17424), .B2(n17421), .A(n17420), .ZN(n20665) );
  OAI22_X1 U19400 ( .A1(n17423), .A2(n17422), .B1(n20665), .B2(n17513), .ZN(
        P3_U2679) );
  AOI21_X1 U19401 ( .B1(n17426), .B2(n17425), .A(n17424), .ZN(n20666) );
  INV_X1 U19402 ( .A(n20666), .ZN(n17428) );
  NAND3_X1 U19403 ( .A1(n17429), .A2(P3_EBX_REG_23__SCAN_IN), .A3(n17513), 
        .ZN(n17427) );
  OAI221_X1 U19404 ( .B1(n17429), .B2(P3_EBX_REG_23__SCAN_IN), .C1(n17513), 
        .C2(n17428), .A(n17427), .ZN(P3_U2680) );
  AOI22_X1 U19405 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17513), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17430), .ZN(n17442) );
  AOI22_X1 U19406 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U19407 ( .A1(n11578), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U19408 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U19409 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17431) );
  NAND4_X1 U19410 ( .A1(n17434), .A2(n17433), .A3(n17432), .A4(n17431), .ZN(
        n17441) );
  AOI22_X1 U19411 ( .A1(n10975), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U19412 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U19413 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U19414 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17435), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17436) );
  NAND4_X1 U19415 ( .A1(n17439), .A2(n17438), .A3(n17437), .A4(n17436), .ZN(
        n17440) );
  NOR2_X1 U19416 ( .A1(n17441), .A2(n17440), .ZN(n20600) );
  OAI22_X1 U19417 ( .A1(n17443), .A2(n17442), .B1(n20600), .B2(n17513), .ZN(
        P3_U2681) );
  AOI22_X1 U19418 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U19419 ( .A1(n10953), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U19420 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10948), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U19421 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17445) );
  NAND4_X1 U19422 ( .A1(n17448), .A2(n17447), .A3(n17446), .A4(n17445), .ZN(
        n17454) );
  AOI22_X1 U19423 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10955), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U19424 ( .A1(n17499), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19425 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U19426 ( .A1(n10976), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17449) );
  NAND4_X1 U19427 ( .A1(n17452), .A2(n17451), .A3(n17450), .A4(n17449), .ZN(
        n17453) );
  NOR2_X1 U19428 ( .A1(n17454), .A2(n17453), .ZN(n20595) );
  OAI21_X1 U19429 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17490), .A(n17455), .ZN(
        n17456) );
  OAI21_X1 U19430 ( .B1(n20595), .B2(n17513), .A(n17456), .ZN(P3_U2683) );
  AOI22_X1 U19431 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U19432 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10953), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U19433 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U19434 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17458) );
  NAND4_X1 U19435 ( .A1(n17461), .A2(n17460), .A3(n17459), .A4(n17458), .ZN(
        n17469) );
  AOI22_X1 U19436 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19437 ( .A1(n17435), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U19438 ( .A1(n11434), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U19439 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17464) );
  NAND4_X1 U19440 ( .A1(n17467), .A2(n17466), .A3(n17465), .A4(n17464), .ZN(
        n17468) );
  NOR2_X1 U19441 ( .A1(n17469), .A2(n17468), .ZN(n20615) );
  OAI21_X1 U19442 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17470), .A(n17472), .ZN(
        n17471) );
  AOI22_X1 U19443 ( .A1(n17517), .A2(n20615), .B1(n17471), .B2(n17513), .ZN(
        P3_U2685) );
  AOI21_X1 U19444 ( .B1(n20346), .B2(n17472), .A(n17517), .ZN(n17473) );
  INV_X1 U19445 ( .A(n17473), .ZN(n17489) );
  AOI22_X1 U19446 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U19447 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10957), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U19448 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U19449 ( .A1(n17475), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17492), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17476) );
  NAND4_X1 U19450 ( .A1(n17479), .A2(n17478), .A3(n17477), .A4(n17476), .ZN(
        n17488) );
  AOI22_X1 U19451 ( .A1(n17435), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10974), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U19452 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U19453 ( .A1(n17491), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U19454 ( .A1(n10952), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10976), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17483) );
  NAND4_X1 U19455 ( .A1(n17486), .A2(n17485), .A3(n17484), .A4(n17483), .ZN(
        n17487) );
  NOR2_X1 U19456 ( .A1(n17488), .A2(n17487), .ZN(n20611) );
  OAI22_X1 U19457 ( .A1(n17490), .A2(n17489), .B1(n20611), .B2(n17513), .ZN(
        P3_U2684) );
  AOI22_X1 U19458 ( .A1(n17262), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17444), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19459 ( .A1(n10965), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17491), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U19460 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17492), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17457), .ZN(n17494) );
  AOI22_X1 U19461 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17474), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17475), .ZN(n17493) );
  NAND4_X1 U19462 ( .A1(n17496), .A2(n17495), .A3(n17494), .A4(n17493), .ZN(
        n17505) );
  AOI22_X1 U19463 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17463), .ZN(n17503) );
  AOI22_X1 U19464 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11578), .ZN(n17502) );
  AOI22_X1 U19465 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10974), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17499), .ZN(n17501) );
  AOI22_X1 U19466 ( .A1(n10955), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10952), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17500) );
  NAND4_X1 U19467 ( .A1(n17503), .A2(n17502), .A3(n17501), .A4(n17500), .ZN(
        n17504) );
  NOR2_X1 U19468 ( .A1(n17505), .A2(n17504), .ZN(n20621) );
  NAND2_X1 U19469 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17506), .ZN(n17510) );
  OAI211_X1 U19470 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17508), .A(n17516), .B(
        n17507), .ZN(n17509) );
  OAI211_X1 U19471 ( .C1(n20621), .C2(n17513), .A(n17510), .B(n17509), .ZN(
        P3_U2686) );
  AOI21_X1 U19472 ( .B1(n20099), .B2(n20098), .A(n17511), .ZN(n17512) );
  INV_X1 U19473 ( .A(n17512), .ZN(n20091) );
  OAI222_X1 U19474 ( .A1(n17515), .A2(n20091), .B1(n20098), .B2(n17519), .C1(
        n17514), .C2(n17513), .ZN(P3_U2702) );
  AOI22_X1 U19475 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17517), .B1(
        n17516), .B2(n20099), .ZN(n17518) );
  OAI21_X1 U19476 ( .B1(n17519), .B2(n20099), .A(n17518), .ZN(P3_U2703) );
  INV_X1 U19477 ( .A(n17520), .ZN(n17522) );
  OAI21_X1 U19478 ( .B1(n21135), .B2(n20027), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17521) );
  OAI21_X1 U19479 ( .B1(n17522), .B2(n20082), .A(n17521), .ZN(P3_U2634) );
  INV_X1 U19480 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21192) );
  AOI21_X1 U19481 ( .B1(n21192), .B2(n17524), .A(n17523), .ZN(n21182) );
  OAI21_X1 U19482 ( .B1(n21182), .B2(n17525), .A(n17527), .ZN(n17526) );
  OAI221_X1 U19483 ( .B1(n21144), .B2(n20018), .C1(n21144), .C2(n17527), .A(
        n17526), .ZN(P3_U2863) );
  NAND2_X1 U19484 ( .A1(n17530), .A2(n21071), .ZN(n21077) );
  AOI21_X1 U19485 ( .B1(n17876), .B2(n17528), .A(n17875), .ZN(n17762) );
  OAI21_X1 U19486 ( .B1(n11026), .B2(n17917), .A(n17762), .ZN(n17542) );
  NOR3_X1 U19487 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17680), .A3(
        n17528), .ZN(n17543) );
  OAI21_X1 U19488 ( .B1(n11026), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17541), .ZN(n20328) );
  NAND2_X1 U19489 ( .A1(n10958), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n21075) );
  OAI21_X1 U19490 ( .B1(n17755), .B2(n20328), .A(n21075), .ZN(n17529) );
  AOI211_X1 U19491 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17542), .A(
        n17543), .B(n17529), .ZN(n17533) );
  AOI22_X1 U19492 ( .A1(n17908), .A2(n21061), .B1(n17836), .B2(n20920), .ZN(
        n17570) );
  OAI21_X1 U19493 ( .B1(n17530), .B2(n17753), .A(n17570), .ZN(n17760) );
  OAI21_X1 U19494 ( .B1(n17708), .B2(n21071), .A(n17619), .ZN(n17531) );
  XNOR2_X1 U19495 ( .A(n17531), .B(n17535), .ZN(n21074) );
  AOI22_X1 U19496 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17760), .B1(
        n17837), .B2(n21074), .ZN(n17532) );
  OAI211_X1 U19497 ( .C1(n17753), .C2(n21077), .A(n17533), .B(n17532), .ZN(
        P3_U2812) );
  NOR2_X2 U19498 ( .A1(n17821), .A2(n17534), .ZN(n17669) );
  INV_X1 U19499 ( .A(n17669), .ZN(n17549) );
  NAND3_X1 U19500 ( .A1(n17626), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21017), .ZN(n21039) );
  NAND3_X1 U19501 ( .A1(n17626), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21018), .ZN(n21038) );
  AOI22_X1 U19502 ( .A1(n17836), .A2(n21039), .B1(n17908), .B2(n21038), .ZN(
        n17628) );
  INV_X1 U19503 ( .A(n17619), .ZN(n17536) );
  NAND2_X1 U19504 ( .A1(n17536), .A2(n17535), .ZN(n17613) );
  NAND3_X1 U19505 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17537), .ZN(n17620) );
  NAND2_X1 U19506 ( .A1(n17613), .A2(n17620), .ZN(n17538) );
  XNOR2_X1 U19507 ( .A(n21048), .B(n17538), .ZN(n21044) );
  NOR3_X1 U19508 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17680), .A3(
        n17539), .ZN(n17547) );
  AOI21_X1 U19509 ( .B1(n17541), .B2(n20355), .A(n17540), .ZN(n20333) );
  INV_X1 U19510 ( .A(n20333), .ZN(n17545) );
  NAND2_X1 U19511 ( .A1(n10958), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21045) );
  OAI21_X1 U19512 ( .B1(n17543), .B2(n17542), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17544) );
  OAI211_X1 U19513 ( .C1(n17755), .C2(n17545), .A(n21045), .B(n17544), .ZN(
        n17546) );
  AOI211_X1 U19514 ( .C1(n17837), .C2(n21044), .A(n17547), .B(n17546), .ZN(
        n17548) );
  OAI221_X1 U19515 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17549), 
        .C1(n21048), .C2(n17628), .A(n17548), .ZN(P3_U2811) );
  NOR2_X1 U19516 ( .A1(n17550), .A2(n20096), .ZN(n17767) );
  NAND2_X1 U19517 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17767), .ZN(
        n17562) );
  OAI21_X1 U19518 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17767), .A(
        n17562), .ZN(n20286) );
  NOR2_X1 U19519 ( .A1(n17680), .A2(n17550), .ZN(n17565) );
  INV_X1 U19520 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17551) );
  AOI21_X1 U19521 ( .B1(n17876), .B2(n17550), .A(n17875), .ZN(n17772) );
  OAI21_X1 U19522 ( .B1(n17767), .B2(n17917), .A(n17772), .ZN(n17563) );
  INV_X1 U19523 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20297) );
  NOR2_X1 U19524 ( .A1(n21105), .A2(n20297), .ZN(n20923) );
  AOI221_X1 U19525 ( .B1(n17565), .B2(n17551), .C1(n17563), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n20923), .ZN(n17559) );
  INV_X1 U19526 ( .A(n17764), .ZN(n20921) );
  AOI21_X1 U19527 ( .B1(n20921), .B2(n20915), .A(n17570), .ZN(n17557) );
  NAND2_X1 U19528 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20890) );
  INV_X1 U19529 ( .A(n20880), .ZN(n20873) );
  NOR3_X1 U19530 ( .A1(n11516), .A2(n17708), .A3(n17552), .ZN(n17796) );
  NAND2_X1 U19531 ( .A1(n20873), .A2(n17796), .ZN(n17783) );
  NOR2_X1 U19532 ( .A1(n20890), .A2(n17783), .ZN(n17583) );
  NAND2_X1 U19533 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17583), .ZN(
        n17778) );
  NAND2_X1 U19534 ( .A1(n17553), .A2(n20858), .ZN(n17812) );
  INV_X1 U19535 ( .A(n17812), .ZN(n17577) );
  NAND2_X1 U19536 ( .A1(n17554), .A2(n17577), .ZN(n17779) );
  AOI22_X1 U19537 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17778), .B1(
        n17779), .B2(n20918), .ZN(n17555) );
  XOR2_X1 U19538 ( .A(n20915), .B(n17555), .Z(n20930) );
  NAND2_X1 U19539 ( .A1(n17776), .A2(n20915), .ZN(n20922) );
  OAI22_X1 U19540 ( .A1(n20930), .A2(n17810), .B1(n17923), .B2(n20922), .ZN(
        n17556) );
  NOR2_X1 U19541 ( .A1(n17557), .A2(n17556), .ZN(n17558) );
  OAI211_X1 U19542 ( .C1(n17755), .C2(n20286), .A(n17559), .B(n17558), .ZN(
        P3_U2815) );
  AOI22_X1 U19543 ( .A1(n17793), .A2(n21090), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17708), .ZN(n17560) );
  XOR2_X1 U19544 ( .A(n17561), .B(n17560), .Z(n21087) );
  INV_X1 U19545 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20298) );
  INV_X1 U19546 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20304) );
  AND2_X1 U19547 ( .A1(n17751), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20306) );
  AOI21_X1 U19548 ( .B1(n20304), .B2(n17562), .A(n20306), .ZN(n20296) );
  AOI22_X1 U19549 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17563), .B1(
        n17747), .B2(n20296), .ZN(n17567) );
  OAI211_X1 U19550 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17565), .B(n17564), .ZN(n17566) );
  OAI211_X1 U19551 ( .C1(n20298), .C2(n21105), .A(n17567), .B(n17566), .ZN(
        n17568) );
  AOI21_X1 U19552 ( .B1(n17837), .B2(n21087), .A(n17568), .ZN(n17569) );
  OAI221_X1 U19553 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17753), 
        .C1(n21090), .C2(n17570), .A(n17569), .ZN(P3_U2814) );
  INV_X1 U19554 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20244) );
  NAND2_X1 U19555 ( .A1(n17571), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17788) );
  NOR2_X1 U19556 ( .A1(n20244), .A2(n17788), .ZN(n17588) );
  AOI21_X1 U19557 ( .B1(n20244), .B2(n17788), .A(n17588), .ZN(n20241) );
  NOR2_X1 U19558 ( .A1(n20880), .A2(n20875), .ZN(n20868) );
  INV_X1 U19559 ( .A(n20868), .ZN(n20895) );
  NOR3_X1 U19560 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17821), .A3(
        n20895), .ZN(n17575) );
  NAND2_X1 U19561 ( .A1(n17571), .A2(n17683), .ZN(n17587) );
  OAI21_X1 U19562 ( .B1(n17571), .B2(n17829), .A(n17918), .ZN(n17572) );
  AOI21_X1 U19563 ( .B1(n17635), .B2(n17788), .A(n17572), .ZN(n17589) );
  NAND2_X1 U19564 ( .A1(n10958), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17573) );
  OAI221_X1 U19565 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17587), .C1(
        n20244), .C2(n17589), .A(n17573), .ZN(n17574) );
  AOI211_X1 U19566 ( .C1(n17747), .C2(n20241), .A(n17575), .B(n17574), .ZN(
        n17582) );
  AND2_X1 U19567 ( .A1(n20869), .A2(n20900), .ZN(n20894) );
  INV_X1 U19568 ( .A(n17786), .ZN(n21062) );
  INV_X1 U19569 ( .A(n20900), .ZN(n20891) );
  NOR2_X1 U19570 ( .A1(n21062), .A2(n20891), .ZN(n17576) );
  OAI22_X1 U19571 ( .A1(n20894), .A2(n17923), .B1(n17576), .B2(n17785), .ZN(
        n17592) );
  NOR2_X1 U19572 ( .A1(n17708), .A2(n20895), .ZN(n17579) );
  AOI22_X1 U19573 ( .A1(n17826), .A2(n17579), .B1(n17578), .B2(n17577), .ZN(
        n17580) );
  XOR2_X1 U19574 ( .A(n20899), .B(n17580), .Z(n20885) );
  AOI22_X1 U19575 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17592), .B1(
        n17837), .B2(n20885), .ZN(n17581) );
  NAND2_X1 U19576 ( .A1(n17582), .A2(n17581), .ZN(P3_U2818) );
  INV_X1 U19577 ( .A(n17583), .ZN(n17584) );
  OAI21_X1 U19578 ( .B1(n17812), .B2(n17585), .A(n17584), .ZN(n17586) );
  INV_X1 U19579 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20903) );
  XOR2_X1 U19580 ( .A(n17586), .B(n20903), .Z(n21099) );
  INV_X1 U19581 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17766) );
  AOI211_X1 U19582 ( .C1(n20244), .C2(n17766), .A(n17771), .B(n17587), .ZN(
        n17591) );
  INV_X1 U19583 ( .A(n17588), .ZN(n20252) );
  AOI22_X1 U19584 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20252), .B1(
        n17588), .B2(n17766), .ZN(n20258) );
  OAI22_X1 U19585 ( .A1(n17589), .A2(n17766), .B1(n17755), .B2(n20258), .ZN(
        n17590) );
  AOI211_X1 U19586 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n10958), .A(n17591), 
        .B(n17590), .ZN(n17594) );
  NOR2_X1 U19587 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20891), .ZN(
        n21092) );
  AOI22_X1 U19588 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17592), .B1(
        n21092), .B2(n17806), .ZN(n17593) );
  OAI211_X1 U19589 ( .C1(n21099), .C2(n17810), .A(n17594), .B(n17593), .ZN(
        P3_U2817) );
  NAND2_X1 U19590 ( .A1(n17596), .A2(n17669), .ZN(n17740) );
  NOR2_X1 U19591 ( .A1(n20920), .A2(n17595), .ZN(n17658) );
  INV_X1 U19592 ( .A(n17658), .ZN(n20766) );
  AOI22_X1 U19593 ( .A1(n17836), .A2(n20766), .B1(n17908), .B2(n20765), .ZN(
        n17617) );
  NAND2_X1 U19594 ( .A1(n17597), .A2(n17596), .ZN(n17599) );
  AOI21_X1 U19595 ( .B1(n17599), .B2(n17598), .A(n17618), .ZN(n17644) );
  XOR2_X1 U19596 ( .A(n17644), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n20939) );
  INV_X1 U19597 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20367) );
  NOR2_X1 U19598 ( .A1(n17622), .A2(n20367), .ZN(n17601) );
  OAI21_X1 U19599 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17601), .A(
        n17600), .ZN(n20382) );
  OAI21_X1 U19600 ( .B1(n17540), .B2(n17917), .A(n17918), .ZN(n17602) );
  AOI21_X1 U19601 ( .B1(n17876), .B2(n17603), .A(n17602), .ZN(n17625) );
  OAI21_X1 U19602 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17754), .A(
        n17625), .ZN(n17611) );
  AOI22_X1 U19603 ( .A1(n10958), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17611), .ZN(n17606) );
  NOR2_X1 U19604 ( .A1(n17680), .A2(n17603), .ZN(n17612) );
  OAI211_X1 U19605 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17612), .B(n17604), .ZN(n17605) );
  OAI211_X1 U19606 ( .C1(n17755), .C2(n20382), .A(n17606), .B(n17605), .ZN(
        n17607) );
  AOI21_X1 U19607 ( .B1(n17837), .B2(n20939), .A(n17607), .ZN(n17608) );
  OAI221_X1 U19608 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17740), 
        .C1(n20942), .C2(n17617), .A(n17608), .ZN(P3_U2808) );
  INV_X1 U19609 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20370) );
  INV_X1 U19610 ( .A(n17622), .ZN(n17609) );
  AOI22_X1 U19611 ( .A1(n17609), .A2(n20367), .B1(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17622), .ZN(n20363) );
  OAI22_X1 U19612 ( .A1(n21105), .A2(n20370), .B1(n17755), .B2(n20363), .ZN(
        n17610) );
  AOI221_X1 U19613 ( .B1(n17612), .B2(n20367), .C1(n17611), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17610), .ZN(n17616) );
  OAI22_X1 U19614 ( .A1(n20769), .A2(n17620), .B1(n21051), .B2(n17613), .ZN(
        n17614) );
  XOR2_X1 U19615 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17614), .Z(
        n20772) );
  NOR2_X1 U19616 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n20769), .ZN(
        n20771) );
  AOI22_X1 U19617 ( .A1(n17837), .A2(n20772), .B1(n17669), .B2(n20771), .ZN(
        n17615) );
  OAI211_X1 U19618 ( .C1(n17617), .C2(n20937), .A(n17616), .B(n17615), .ZN(
        P3_U2809) );
  AOI221_X1 U19619 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17620), 
        .C1(n21048), .C2(n17619), .A(n17618), .ZN(n17621) );
  XOR2_X1 U19620 ( .A(n21053), .B(n17621), .Z(n21057) );
  OAI21_X1 U19621 ( .B1(n17540), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17622), .ZN(n20357) );
  AOI21_X1 U19622 ( .B1(n17755), .B2(n17754), .A(n20357), .ZN(n17633) );
  AOI21_X1 U19623 ( .B1(n17623), .B2(n18894), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17624) );
  NAND2_X1 U19624 ( .A1(n10958), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21055) );
  OAI21_X1 U19625 ( .B1(n17625), .B2(n17624), .A(n21055), .ZN(n17632) );
  NAND2_X1 U19626 ( .A1(n17626), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17627) );
  NOR2_X1 U19627 ( .A1(n17753), .A2(n17627), .ZN(n17630) );
  INV_X1 U19628 ( .A(n17628), .ZN(n17629) );
  MUX2_X1 U19629 ( .A(n17630), .B(n17629), .S(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n17631) );
  NOR3_X1 U19630 ( .A1(n17633), .A2(n17632), .A3(n17631), .ZN(n17634) );
  OAI21_X1 U19631 ( .B1(n17810), .B2(n21057), .A(n17634), .ZN(P3_U2810) );
  AOI21_X1 U19632 ( .B1(n21019), .B2(n21018), .A(n17923), .ZN(n17643) );
  AOI21_X1 U19633 ( .B1(n21019), .B2(n21017), .A(n17785), .ZN(n17642) );
  AOI22_X1 U19634 ( .A1(n17651), .A2(n17643), .B1(n17658), .B2(n17642), .ZN(
        n17649) );
  AND2_X1 U19635 ( .A1(n17654), .A2(n18894), .ZN(n17640) );
  INV_X1 U19636 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18000) );
  NOR2_X1 U19637 ( .A1(n21105), .A2(n18000), .ZN(n21027) );
  AOI211_X1 U19638 ( .C1(n17635), .C2(n17670), .A(n17640), .B(n17875), .ZN(
        n17675) );
  AOI21_X1 U19639 ( .B1(n17637), .B2(n17636), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17638) );
  OAI21_X1 U19640 ( .B1(n17637), .B2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17670), .ZN(n20399) );
  OAI22_X1 U19641 ( .A1(n17675), .A2(n17638), .B1(n17755), .B2(n20399), .ZN(
        n17639) );
  AOI211_X1 U19642 ( .C1(n17641), .C2(n17640), .A(n21027), .B(n17639), .ZN(
        n17648) );
  OR2_X1 U19643 ( .A1(n17643), .A2(n17642), .ZN(n17677) );
  OAI221_X1 U19644 ( .B1(n17645), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n17645), .C2(n17793), .A(n17644), .ZN(n17646) );
  XOR2_X1 U19645 ( .A(n17650), .B(n17646), .Z(n21028) );
  AOI22_X1 U19646 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17677), .B1(
        n17837), .B2(n21028), .ZN(n17647) );
  OAI211_X1 U19647 ( .C1(n17649), .C2(n20942), .A(n17648), .B(n17647), .ZN(
        P3_U2807) );
  NOR2_X1 U19648 ( .A1(n17666), .A2(n17650), .ZN(n20948) );
  NAND3_X1 U19649 ( .A1(n20948), .A2(n17651), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17652) );
  XOR2_X1 U19650 ( .A(n17652), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n20952) );
  INV_X1 U19651 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17657) );
  NAND2_X1 U19652 ( .A1(n17671), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17653) );
  AOI21_X1 U19653 ( .B1(n17657), .B2(n17653), .A(n17713), .ZN(n20413) );
  NAND2_X1 U19654 ( .A1(n10958), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n20958) );
  NOR2_X1 U19655 ( .A1(n17680), .A2(n17654), .ZN(n17672) );
  OAI211_X1 U19656 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17672), .B(n17655), .ZN(n17656) );
  OAI211_X1 U19657 ( .C1(n17675), .C2(n17657), .A(n20958), .B(n17656), .ZN(
        n17663) );
  NAND3_X1 U19658 ( .A1(n20948), .A2(n17658), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17659) );
  XOR2_X1 U19659 ( .A(n17659), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n20950) );
  NAND2_X1 U19660 ( .A1(n17708), .A2(n17665), .ZN(n17707) );
  OAI21_X1 U19661 ( .B1(n17708), .B2(n17660), .A(n17707), .ZN(n17661) );
  XOR2_X1 U19662 ( .A(n17661), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n20954) );
  OAI22_X1 U19663 ( .A1(n17785), .A2(n20950), .B1(n17810), .B2(n20954), .ZN(
        n17662) );
  AOI211_X1 U19664 ( .C1(n17747), .C2(n20413), .A(n17663), .B(n17662), .ZN(
        n17664) );
  OAI21_X1 U19665 ( .B1(n17923), .B2(n20952), .A(n17664), .ZN(P3_U2805) );
  OAI21_X1 U19666 ( .B1(n17667), .B2(n17666), .A(n17665), .ZN(n21033) );
  NOR2_X1 U19667 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17668), .ZN(
        n21032) );
  AOI22_X1 U19668 ( .A1(n17837), .A2(n21033), .B1(n17669), .B2(n21032), .ZN(
        n17679) );
  INV_X1 U19669 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19670 ( .A1(n17671), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n17674), .B2(n17670), .ZN(n20402) );
  AOI22_X1 U19671 ( .A1(n20402), .A2(n17747), .B1(n17672), .B2(n17674), .ZN(
        n17673) );
  NAND2_X1 U19672 ( .A1(n10958), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n21034) );
  OAI211_X1 U19673 ( .C1(n17675), .C2(n17674), .A(n17673), .B(n21034), .ZN(
        n17676) );
  AOI21_X1 U19674 ( .B1(n17677), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17676), .ZN(n17678) );
  NAND2_X1 U19675 ( .A1(n17679), .A2(n17678), .ZN(P3_U2806) );
  NOR3_X1 U19676 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17680), .A3(
        n17682), .ZN(n17697) );
  OAI21_X1 U19677 ( .B1(n17713), .B2(n17917), .A(n17918), .ZN(n17681) );
  AOI21_X1 U19678 ( .B1(n17876), .B2(n17682), .A(n17681), .ZN(n17717) );
  OAI21_X1 U19679 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17754), .A(
        n17717), .ZN(n17700) );
  OAI21_X1 U19680 ( .B1(n11040), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17745), .ZN(n20458) );
  NAND2_X1 U19681 ( .A1(n10958), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17686) );
  NAND3_X1 U19682 ( .A1(n17684), .A2(n11096), .A3(n17683), .ZN(n17685) );
  OAI211_X1 U19683 ( .C1(n17755), .C2(n20458), .A(n17686), .B(n17685), .ZN(
        n17687) );
  AOI221_X1 U19684 ( .B1(n17697), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n17700), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17687), .ZN(
        n17696) );
  OR2_X1 U19685 ( .A1(n17688), .A2(n20765), .ZN(n20964) );
  AOI22_X1 U19686 ( .A1(n17908), .A2(n20964), .B1(n17836), .B2(n20976), .ZN(
        n17721) );
  NAND2_X1 U19687 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17721), .ZN(
        n17702) );
  OAI211_X1 U19688 ( .C1(n17836), .C2(n17908), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17702), .ZN(n17695) );
  INV_X1 U19689 ( .A(n17753), .ZN(n17729) );
  NAND3_X1 U19690 ( .A1(n17689), .A2(n17729), .A3(n20998), .ZN(n17694) );
  OAI211_X1 U19691 ( .C1(n17692), .C2(n17691), .A(n17837), .B(n17690), .ZN(
        n17693) );
  NAND4_X1 U19692 ( .A1(n17696), .A2(n17695), .A3(n17694), .A4(n17693), .ZN(
        P3_U2802) );
  AOI21_X1 U19693 ( .B1(n17712), .B2(n20446), .A(n11040), .ZN(n20443) );
  AOI21_X1 U19694 ( .B1(n17747), .B2(n20443), .A(n17697), .ZN(n17706) );
  OAI21_X1 U19695 ( .B1(n17793), .B2(n17699), .A(n17698), .ZN(n20985) );
  AOI22_X1 U19696 ( .A1(n17837), .A2(n20985), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17700), .ZN(n17705) );
  NOR2_X1 U19697 ( .A1(n17701), .A2(n17753), .ZN(n17703) );
  OAI21_X1 U19698 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17703), .A(
        n17702), .ZN(n17704) );
  NAND2_X1 U19699 ( .A1(n10958), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n20986) );
  NAND4_X1 U19700 ( .A1(n17706), .A2(n17705), .A3(n17704), .A4(n20986), .ZN(
        P3_U2803) );
  OAI221_X1 U19701 ( .B1(n17709), .B2(n17708), .C1(n17709), .C2(n20963), .A(
        n17707), .ZN(n17710) );
  XOR2_X1 U19702 ( .A(n20962), .B(n17710), .Z(n20960) );
  NOR4_X1 U19703 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n20942), .A3(
        n20968), .A4(n17740), .ZN(n17719) );
  AOI21_X1 U19704 ( .B1(n17711), .B2(n18894), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17716) );
  OAI21_X1 U19705 ( .B1(n17713), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17712), .ZN(n17714) );
  INV_X1 U19706 ( .A(n17714), .ZN(n20435) );
  OAI21_X1 U19707 ( .B1(n17747), .B2(n17636), .A(n20435), .ZN(n17715) );
  NAND2_X1 U19708 ( .A1(n10958), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n20972) );
  OAI211_X1 U19709 ( .C1(n17717), .C2(n17716), .A(n17715), .B(n20972), .ZN(
        n17718) );
  AOI211_X1 U19710 ( .C1(n17837), .C2(n20960), .A(n17719), .B(n17718), .ZN(
        n17720) );
  OAI21_X1 U19711 ( .B1(n17721), .B2(n20962), .A(n17720), .ZN(P3_U2804) );
  AOI22_X1 U19712 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17737), .B1(
        n17738), .B2(n21008), .ZN(n17722) );
  XOR2_X1 U19713 ( .A(n21007), .B(n17722), .Z(n21015) );
  NOR2_X1 U19714 ( .A1(n20988), .A2(n21008), .ZN(n20996) );
  NOR3_X1 U19715 ( .A1(n17728), .A2(n20976), .A3(n21008), .ZN(n20994) );
  OAI22_X1 U19716 ( .A1(n20996), .A2(n17923), .B1(n20994), .B2(n17785), .ZN(
        n17743) );
  INV_X1 U19717 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20485) );
  OAI21_X1 U19718 ( .B1(n17744), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17723), .ZN(n20494) );
  OAI22_X1 U19719 ( .A1(n17724), .A2(n20485), .B1(n17755), .B2(n20494), .ZN(
        n17727) );
  INV_X1 U19720 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20497) );
  OAI22_X1 U19721 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17725), .B1(
        n21105), .B2(n20497), .ZN(n17726) );
  AOI211_X1 U19722 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17743), .A(
        n17727), .B(n17726), .ZN(n17733) );
  NOR2_X1 U19723 ( .A1(n17728), .A2(n21008), .ZN(n17730) );
  NAND4_X1 U19724 ( .A1(n17731), .A2(n17730), .A3(n17729), .A4(n21007), .ZN(
        n17732) );
  OAI211_X1 U19725 ( .C1(n21015), .C2(n17810), .A(n17733), .B(n17732), .ZN(
        P3_U2800) );
  OAI21_X1 U19726 ( .B1(n17734), .B2(n18893), .A(n20481), .ZN(n17735) );
  AOI22_X1 U19727 ( .A1(n10958), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17736), 
        .B2(n17735), .ZN(n17750) );
  NAND2_X1 U19728 ( .A1(n17738), .A2(n17737), .ZN(n17739) );
  XOR2_X1 U19729 ( .A(n17739), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n20992) );
  OAI21_X1 U19730 ( .B1(n17741), .B2(n17740), .A(n21008), .ZN(n17742) );
  AOI22_X1 U19731 ( .A1(n17837), .A2(n20992), .B1(n17743), .B2(n17742), .ZN(
        n17749) );
  AOI21_X1 U19732 ( .B1(n17745), .B2(n20481), .A(n17744), .ZN(n20476) );
  OAI21_X1 U19733 ( .B1(n17747), .B2(n17746), .A(n20476), .ZN(n17748) );
  NAND3_X1 U19734 ( .A1(n17750), .A2(n17749), .A3(n17748), .ZN(P3_U2801) );
  AOI21_X1 U19735 ( .B1(n17751), .B2(n18894), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17763) );
  INV_X1 U19736 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17752) );
  OAI21_X1 U19737 ( .B1(n21090), .B2(n17753), .A(n17752), .ZN(n17759) );
  INV_X1 U19738 ( .A(n11026), .ZN(n20325) );
  OAI21_X1 U19739 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20306), .A(
        n20325), .ZN(n20308) );
  AOI21_X1 U19740 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17757), .A(
        n17756), .ZN(n21083) );
  OAI22_X1 U19741 ( .A1(n17895), .A2(n20308), .B1(n21083), .B2(n17810), .ZN(
        n17758) );
  AOI21_X1 U19742 ( .B1(n17760), .B2(n17759), .A(n17758), .ZN(n17761) );
  NAND2_X1 U19743 ( .A1(n10958), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21081) );
  OAI211_X1 U19744 ( .C1(n17763), .C2(n17762), .A(n17761), .B(n21081), .ZN(
        P3_U2813) );
  AOI21_X1 U19745 ( .B1(n20918), .B2(n17765), .A(n17764), .ZN(n20908) );
  INV_X1 U19746 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20271) );
  NOR2_X1 U19747 ( .A1(n21105), .A2(n20271), .ZN(n17775) );
  NOR2_X1 U19748 ( .A1(n17766), .A2(n20252), .ZN(n17769) );
  INV_X1 U19749 ( .A(n17767), .ZN(n17768) );
  OAI21_X1 U19750 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17769), .A(
        n17768), .ZN(n20266) );
  NOR3_X1 U19751 ( .A1(n17855), .A2(n20159), .A3(n18893), .ZN(n17842) );
  NAND2_X1 U19752 ( .A1(n17770), .A2(n17842), .ZN(n17802) );
  NOR2_X1 U19753 ( .A1(n20231), .A2(n17802), .ZN(n17787) );
  AOI21_X1 U19754 ( .B1(n17771), .B2(n17787), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17773) );
  OAI22_X1 U19755 ( .A1(n17895), .A2(n20266), .B1(n17773), .B2(n17772), .ZN(
        n17774) );
  AOI211_X1 U19756 ( .C1(n20908), .C2(n17836), .A(n17775), .B(n17774), .ZN(
        n17782) );
  AOI21_X1 U19757 ( .B1(n20918), .B2(n17777), .A(n17776), .ZN(n20909) );
  NAND2_X1 U19758 ( .A1(n17779), .A2(n17778), .ZN(n17780) );
  XOR2_X1 U19759 ( .A(n17780), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n20910) );
  AOI22_X1 U19760 ( .A1(n17908), .A2(n20909), .B1(n17837), .B2(n20910), .ZN(
        n17781) );
  NAND2_X1 U19761 ( .A1(n17782), .A2(n17781), .ZN(P3_U2816) );
  OAI21_X1 U19762 ( .B1(n17812), .B2(n17807), .A(n17783), .ZN(n17784) );
  XOR2_X1 U19763 ( .A(n17784), .B(n20875), .Z(n20884) );
  OAI22_X1 U19764 ( .A1(n17786), .A2(n17785), .B1(n17923), .B2(n20869), .ZN(
        n17811) );
  NOR2_X1 U19765 ( .A1(n17875), .A2(n17876), .ZN(n17915) );
  AOI211_X1 U19766 ( .C1(n17802), .C2(n20231), .A(n17915), .B(n17787), .ZN(
        n17790) );
  NOR2_X1 U19767 ( .A1(n20213), .A2(n20096), .ZN(n17800) );
  OAI21_X1 U19768 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17800), .A(
        n17788), .ZN(n20224) );
  INV_X1 U19769 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20235) );
  OAI22_X1 U19770 ( .A1(n17895), .A2(n20224), .B1(n21105), .B2(n20235), .ZN(
        n17789) );
  AOI211_X1 U19771 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n17811), .A(
        n17790), .B(n17789), .ZN(n17792) );
  OAI211_X1 U19772 ( .C1(n20873), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n20895), .B(n17806), .ZN(n17791) );
  OAI211_X1 U19773 ( .C1(n20884), .C2(n17810), .A(n17792), .B(n17791), .ZN(
        P3_U2819) );
  NOR2_X1 U19774 ( .A1(n17793), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17795) );
  OAI22_X1 U19775 ( .A1(n17796), .A2(n17795), .B1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17794), .ZN(n17798) );
  INV_X1 U19776 ( .A(n17796), .ZN(n17813) );
  OAI221_X1 U19777 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17812), .C1(
        n21115), .C2(n17813), .A(n20874), .ZN(n17797) );
  OAI21_X1 U19778 ( .B1(n20874), .B2(n17798), .A(n17797), .ZN(n21111) );
  INV_X1 U19779 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20222) );
  NOR2_X1 U19780 ( .A1(n21105), .A2(n20222), .ZN(n17805) );
  NAND3_X1 U19781 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n17842), .ZN(n17816) );
  NOR2_X1 U19782 ( .A1(n20201), .A2(n17816), .ZN(n17815) );
  INV_X1 U19783 ( .A(n17815), .ZN(n17799) );
  OAI21_X1 U19784 ( .B1(n20220), .B2(n17915), .A(n17799), .ZN(n17801) );
  NAND2_X1 U19785 ( .A1(n17830), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20175) );
  NOR2_X1 U19786 ( .A1(n20174), .A2(n20175), .ZN(n17843) );
  INV_X1 U19787 ( .A(n17843), .ZN(n17825) );
  NOR2_X1 U19788 ( .A1(n20185), .A2(n17825), .ZN(n17824) );
  NAND2_X1 U19789 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17824), .ZN(
        n20214) );
  AOI21_X1 U19790 ( .B1(n20220), .B2(n20214), .A(n17800), .ZN(n20217) );
  AOI22_X1 U19791 ( .A1(n17802), .A2(n17801), .B1(n17911), .B2(n20217), .ZN(
        n17803) );
  INV_X1 U19792 ( .A(n17803), .ZN(n17804) );
  AOI211_X1 U19793 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17811), .A(
        n17805), .B(n17804), .ZN(n17809) );
  NAND3_X1 U19794 ( .A1(n20880), .A2(n17807), .A3(n17806), .ZN(n17808) );
  OAI211_X1 U19795 ( .C1(n21111), .C2(n17810), .A(n17809), .B(n17808), .ZN(
        P3_U2820) );
  INV_X1 U19796 ( .A(n17811), .ZN(n17820) );
  NAND2_X1 U19797 ( .A1(n17813), .A2(n17812), .ZN(n17814) );
  XOR2_X1 U19798 ( .A(n17814), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21119) );
  AOI211_X1 U19799 ( .C1(n17816), .C2(n20201), .A(n17915), .B(n17815), .ZN(
        n17818) );
  OAI21_X1 U19800 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17824), .A(
        n20214), .ZN(n20195) );
  NAND2_X1 U19801 ( .A1(n10958), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n21121) );
  OAI21_X1 U19802 ( .B1(n17895), .B2(n20195), .A(n21121), .ZN(n17817) );
  AOI211_X1 U19803 ( .C1(n17837), .C2(n21119), .A(n17818), .B(n17817), .ZN(
        n17819) );
  OAI221_X1 U19804 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17821), .C1(
        n21115), .C2(n17820), .A(n17819), .ZN(P3_U2821) );
  OAI21_X1 U19805 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17823), .A(
        n17822), .ZN(n20866) );
  AOI21_X1 U19806 ( .B1(n20185), .B2(n17825), .A(n17824), .ZN(n20178) );
  AOI22_X1 U19807 ( .A1(n10958), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n20178), 
        .B2(n17911), .ZN(n17839) );
  AOI21_X1 U19808 ( .B1(n17828), .B2(n17827), .A(n17826), .ZN(n20862) );
  INV_X1 U19809 ( .A(n20862), .ZN(n17835) );
  NAND2_X1 U19810 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17842), .ZN(
        n17833) );
  NAND2_X1 U19811 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17831) );
  OAI21_X1 U19812 ( .B1(n17830), .B2(n17829), .A(n17918), .ZN(n17844) );
  AOI21_X1 U19813 ( .B1(n18894), .B2(n17831), .A(n17844), .ZN(n17832) );
  AOI21_X1 U19814 ( .B1(n20185), .B2(n17833), .A(n17832), .ZN(n17834) );
  AOI221_X1 U19815 ( .B1(n17837), .B2(n20862), .C1(n17836), .C2(n17835), .A(
        n17834), .ZN(n17838) );
  OAI211_X1 U19816 ( .C1(n17923), .C2(n20866), .A(n17839), .B(n17838), .ZN(
        P3_U2822) );
  AOI21_X1 U19817 ( .B1(n20850), .B2(n17841), .A(n17840), .ZN(n20846) );
  AOI22_X1 U19818 ( .A1(n17912), .A2(n20846), .B1(n17842), .B2(n20174), .ZN(
        n17851) );
  AOI21_X1 U19819 ( .B1(n20174), .B2(n20175), .A(n17843), .ZN(n20161) );
  AOI22_X1 U19820 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17844), .B1(
        n20161), .B2(n17911), .ZN(n17850) );
  AOI21_X1 U19821 ( .B1(n17847), .B2(n17846), .A(n17845), .ZN(n17848) );
  XOR2_X1 U19822 ( .A(n17848), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n20845) );
  NAND2_X1 U19823 ( .A1(n17908), .A2(n20845), .ZN(n17849) );
  NAND2_X1 U19824 ( .A1(n10958), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n20856) );
  NAND4_X1 U19825 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n20856), .ZN(
        P3_U2823) );
  INV_X1 U19826 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20834) );
  AOI21_X1 U19827 ( .B1(n11047), .B2(n17853), .A(n17852), .ZN(n20842) );
  NOR2_X1 U19828 ( .A1(n17855), .A2(n18893), .ZN(n17854) );
  AOI22_X1 U19829 ( .A1(n17912), .A2(n20842), .B1(n17854), .B2(n20159), .ZN(
        n17860) );
  NOR2_X1 U19830 ( .A1(n17915), .A2(n17854), .ZN(n17870) );
  NOR2_X1 U19831 ( .A1(n17855), .A2(n20096), .ZN(n17861) );
  OAI21_X1 U19832 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17861), .A(
        n20175), .ZN(n20153) );
  OAI21_X1 U19833 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17857), .A(
        n17856), .ZN(n20844) );
  OAI22_X1 U19834 ( .A1(n17895), .A2(n20153), .B1(n17923), .B2(n20844), .ZN(
        n17858) );
  AOI21_X1 U19835 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17870), .A(
        n17858), .ZN(n17859) );
  OAI211_X1 U19836 ( .C1(n21105), .C2(n20834), .A(n17860), .B(n17859), .ZN(
        P3_U2824) );
  INV_X1 U19837 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20150) );
  NAND2_X1 U19838 ( .A1(n20128), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17874) );
  AOI21_X1 U19839 ( .B1(n20150), .B2(n17874), .A(n17861), .ZN(n20142) );
  INV_X1 U19840 ( .A(n20142), .ZN(n17873) );
  OAI21_X1 U19841 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17862), .A(
        n20798), .ZN(n17867) );
  OAI211_X1 U19842 ( .C1(n17865), .C2(n17864), .A(n21125), .B(n17863), .ZN(
        n17866) );
  OAI21_X1 U19843 ( .B1(n17868), .B2(n17867), .A(n17866), .ZN(n20829) );
  AOI22_X1 U19844 ( .A1(n10958), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17869), 
        .B2(n20829), .ZN(n17872) );
  OAI221_X1 U19845 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20128), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17918), .A(n17870), .ZN(n17871) );
  OAI211_X1 U19846 ( .C1(n17895), .C2(n17873), .A(n17872), .B(n17871), .ZN(
        P3_U2825) );
  NOR2_X1 U19847 ( .A1(n17891), .A2(n20096), .ZN(n20127) );
  OAI21_X1 U19848 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20127), .A(
        n17874), .ZN(n20131) );
  NOR3_X1 U19849 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17891), .A3(
        n18893), .ZN(n17886) );
  AOI21_X1 U19850 ( .B1(n17876), .B2(n17891), .A(n17875), .ZN(n17899) );
  AOI21_X1 U19851 ( .B1(n20819), .B2(n17877), .A(n20995), .ZN(n17883) );
  AOI211_X1 U19852 ( .C1(n17880), .C2(n17879), .A(n17878), .B(n21132), .ZN(
        n17881) );
  AOI21_X1 U19853 ( .B1(n17883), .B2(n17882), .A(n17881), .ZN(n20822) );
  OAI22_X1 U19854 ( .A1(n17899), .A2(n17884), .B1(n20822), .B2(n21191), .ZN(
        n17885) );
  AOI211_X1 U19855 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n10958), .A(n17886), .B(
        n17885), .ZN(n17887) );
  OAI21_X1 U19856 ( .B1(n17895), .B2(n20131), .A(n17887), .ZN(P3_U2826) );
  INV_X1 U19857 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17898) );
  NAND2_X1 U19858 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17918), .ZN(
        n17903) );
  AOI21_X1 U19859 ( .B1(n17890), .B2(n17889), .A(n17888), .ZN(n20809) );
  INV_X1 U19860 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20116) );
  NOR2_X1 U19861 ( .A1(n21105), .A2(n20116), .ZN(n20808) );
  INV_X1 U19862 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20097) );
  NOR2_X1 U19863 ( .A1(n20097), .A2(n20096), .ZN(n20108) );
  OAI22_X1 U19864 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20108), .B1(
        n20096), .B2(n17891), .ZN(n20121) );
  OAI21_X1 U19865 ( .B1(n17894), .B2(n17893), .A(n17892), .ZN(n20817) );
  OAI22_X1 U19866 ( .A1(n17895), .A2(n20121), .B1(n17923), .B2(n20817), .ZN(
        n17896) );
  AOI211_X1 U19867 ( .C1(n17912), .C2(n20809), .A(n20808), .B(n17896), .ZN(
        n17897) );
  OAI221_X1 U19868 ( .B1(n17899), .B2(n17898), .C1(n17899), .C2(n17903), .A(
        n17897), .ZN(P3_U2827) );
  AOI21_X1 U19869 ( .B1(n17902), .B2(n17901), .A(n17900), .ZN(n20797) );
  AOI21_X1 U19870 ( .B1(n20097), .B2(n20096), .A(n20108), .ZN(n20103) );
  AOI22_X1 U19871 ( .A1(n17912), .A2(n20797), .B1(n20103), .B2(n17911), .ZN(
        n17906) );
  OAI21_X1 U19872 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18894), .A(
        n17903), .ZN(n17905) );
  NAND2_X1 U19873 ( .A1(n10958), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n20804) );
  OAI211_X1 U19874 ( .C1(n20794), .C2(n20793), .A(n17908), .B(n20792), .ZN(
        n17904) );
  NAND4_X1 U19875 ( .A1(n17906), .A2(n17905), .A3(n20804), .A4(n17904), .ZN(
        P3_U2828) );
  NOR2_X1 U19876 ( .A1(n20703), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17907) );
  XNOR2_X1 U19877 ( .A(n17907), .B(n17910), .ZN(n20783) );
  AOI22_X1 U19878 ( .A1(n10958), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17908), 
        .B2(n20783), .ZN(n17914) );
  AOI21_X1 U19879 ( .B1(n17916), .B2(n17910), .A(n17909), .ZN(n20787) );
  AOI22_X1 U19880 ( .A1(n17912), .A2(n20787), .B1(n20096), .B2(n17911), .ZN(
        n17913) );
  OAI211_X1 U19881 ( .C1(n17915), .C2(n20096), .A(n17914), .B(n17913), .ZN(
        P3_U2829) );
  OAI21_X1 U19882 ( .B1(n20703), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17916), .ZN(n20780) );
  INV_X1 U19883 ( .A(n20780), .ZN(n20779) );
  NAND3_X1 U19884 ( .A1(n17919), .A2(n17918), .A3(n17917), .ZN(n17920) );
  AOI22_X1 U19885 ( .A1(n10958), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17920), .ZN(n17921) );
  OAI221_X1 U19886 ( .B1(n20779), .B2(n17923), .C1(n20780), .C2(n17922), .A(
        n17921), .ZN(P3_U2830) );
  NAND2_X1 U19887 ( .A1(n21156), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18613) );
  INV_X1 U19888 ( .A(n18613), .ZN(n18614) );
  NAND2_X1 U19889 ( .A1(n21153), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18595) );
  INV_X1 U19890 ( .A(n18595), .ZN(n18596) );
  NOR2_X1 U19891 ( .A1(n18614), .A2(n18596), .ZN(n17924) );
  OAI22_X1 U19892 ( .A1(n17926), .A2(n21156), .B1(n17925), .B2(n17924), .ZN(
        P3_U2866) );
  OAI21_X1 U19893 ( .B1(n17928), .B2(n17927), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17929) );
  OAI21_X1 U19894 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17930), .A(
        n17929), .ZN(P3_U2864) );
  NOR4_X1 U19895 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17934) );
  NOR4_X1 U19896 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17933) );
  NOR4_X1 U19897 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17932) );
  NOR4_X1 U19898 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17931) );
  NAND4_X1 U19899 ( .A1(n17934), .A2(n17933), .A3(n17932), .A4(n17931), .ZN(
        n17940) );
  NOR4_X1 U19900 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17938) );
  AOI211_X1 U19901 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17937) );
  NOR4_X1 U19902 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17936) );
  NOR4_X1 U19903 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17935) );
  NAND4_X1 U19904 ( .A1(n17938), .A2(n17937), .A3(n17936), .A4(n17935), .ZN(
        n17939) );
  NOR2_X1 U19905 ( .A1(n17940), .A2(n17939), .ZN(n17952) );
  INV_X1 U19906 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17942) );
  OAI21_X1 U19907 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n17952), .ZN(n17941) );
  OAI21_X1 U19908 ( .B1(n17952), .B2(n17942), .A(n17941), .ZN(P3_U3293) );
  INV_X1 U19909 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n17945) );
  AOI21_X1 U19910 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n17943) );
  INV_X1 U19911 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n17995) );
  OAI221_X1 U19912 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17943), .C1(n17995), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n17952), .ZN(n17944) );
  OAI21_X1 U19913 ( .B1(n17952), .B2(n17945), .A(n17944), .ZN(P3_U3292) );
  INV_X1 U19914 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17947) );
  NOR3_X1 U19915 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17948) );
  OAI21_X1 U19916 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17948), .A(n17952), .ZN(
        n17946) );
  OAI21_X1 U19917 ( .B1(n17952), .B2(n17947), .A(n17946), .ZN(P3_U2638) );
  INV_X1 U19918 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21646) );
  AOI21_X1 U19919 ( .B1(n17995), .B2(n21646), .A(n17948), .ZN(n17951) );
  INV_X1 U19920 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17950) );
  INV_X1 U19921 ( .A(n17952), .ZN(n17949) );
  AOI22_X1 U19922 ( .A1(n17952), .A2(n17951), .B1(n17950), .B2(n17949), .ZN(
        P3_U2639) );
  OAI22_X1 U19923 ( .A1(n18012), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18006), .ZN(n17953) );
  INV_X1 U19924 ( .A(n17953), .ZN(P3_U3297) );
  INV_X1 U19925 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n17954) );
  AOI22_X1 U19926 ( .A1(n18006), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n17954), 
        .B2(n18012), .ZN(P3_U3294) );
  AOI21_X1 U19927 ( .B1(n21698), .B2(n21689), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17955) );
  AOI22_X1 U19928 ( .A1(n18006), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17955), 
        .B2(n18012), .ZN(P3_U2635) );
  INV_X1 U19929 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20708) );
  AOI22_X1 U19930 ( .A1(n21177), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17956) );
  OAI21_X1 U19931 ( .B1(n20708), .B2(n17972), .A(n17956), .ZN(P3_U2767) );
  INV_X1 U19932 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U19933 ( .A1(n21177), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17957) );
  OAI21_X1 U19934 ( .B1(n20057), .B2(n17972), .A(n17957), .ZN(P3_U2766) );
  INV_X1 U19935 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20576) );
  AOI22_X1 U19936 ( .A1(n21177), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17958) );
  OAI21_X1 U19937 ( .B1(n20576), .B2(n17972), .A(n17958), .ZN(P3_U2765) );
  INV_X1 U19938 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20547) );
  AOI22_X1 U19939 ( .A1(n21177), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17959) );
  OAI21_X1 U19940 ( .B1(n20547), .B2(n17972), .A(n17959), .ZN(P3_U2764) );
  INV_X1 U19941 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20525) );
  AOI22_X1 U19942 ( .A1(n21177), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17960) );
  OAI21_X1 U19943 ( .B1(n20525), .B2(n17972), .A(n17960), .ZN(P3_U2763) );
  INV_X1 U19944 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20548) );
  AOI22_X1 U19945 ( .A1(n21177), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17961) );
  OAI21_X1 U19946 ( .B1(n20548), .B2(n17972), .A(n17961), .ZN(P3_U2762) );
  INV_X1 U19947 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20526) );
  AOI22_X1 U19948 ( .A1(n21177), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17962) );
  OAI21_X1 U19949 ( .B1(n20526), .B2(n17972), .A(n17962), .ZN(P3_U2761) );
  INV_X1 U19950 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20064) );
  AOI22_X1 U19951 ( .A1(n17990), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17963) );
  OAI21_X1 U19952 ( .B1(n20064), .B2(n17972), .A(n17963), .ZN(P3_U2760) );
  INV_X1 U19953 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20066) );
  AOI22_X1 U19954 ( .A1(n17990), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17964) );
  OAI21_X1 U19955 ( .B1(n20066), .B2(n17972), .A(n17964), .ZN(P3_U2759) );
  INV_X1 U19956 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20068) );
  AOI22_X1 U19957 ( .A1(n17990), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17965) );
  OAI21_X1 U19958 ( .B1(n20068), .B2(n17972), .A(n17965), .ZN(P3_U2758) );
  INV_X1 U19959 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20580) );
  AOI22_X1 U19960 ( .A1(n17990), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17966) );
  OAI21_X1 U19961 ( .B1(n20580), .B2(n17972), .A(n17966), .ZN(P3_U2757) );
  INV_X1 U19962 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20536) );
  AOI22_X1 U19963 ( .A1(n17990), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17967) );
  OAI21_X1 U19964 ( .B1(n20536), .B2(n17972), .A(n17967), .ZN(P3_U2756) );
  INV_X1 U19965 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20582) );
  AOI22_X1 U19966 ( .A1(n17990), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17968) );
  OAI21_X1 U19967 ( .B1(n20582), .B2(n17972), .A(n17968), .ZN(P3_U2755) );
  INV_X1 U19968 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20074) );
  AOI22_X1 U19969 ( .A1(n17990), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17969) );
  OAI21_X1 U19970 ( .B1(n20074), .B2(n17972), .A(n17969), .ZN(P3_U2754) );
  INV_X1 U19971 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20683) );
  AOI22_X1 U19972 ( .A1(n17990), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17970) );
  OAI21_X1 U19973 ( .B1(n20683), .B2(n17972), .A(n17970), .ZN(P3_U2753) );
  INV_X1 U19974 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20687) );
  AOI22_X1 U19975 ( .A1(n17990), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17971) );
  OAI21_X1 U19976 ( .B1(n20687), .B2(n17972), .A(n17971), .ZN(P3_U2752) );
  INV_X1 U19977 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20032) );
  NAND2_X1 U19978 ( .A1(n17973), .A2(n20521), .ZN(n17992) );
  AOI22_X1 U19979 ( .A1(n17990), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17974) );
  OAI21_X1 U19980 ( .B1(n20032), .B2(n17992), .A(n17974), .ZN(P3_U2751) );
  INV_X1 U19981 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20584) );
  AOI22_X1 U19982 ( .A1(n17990), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17975) );
  OAI21_X1 U19983 ( .B1(n20584), .B2(n17992), .A(n17975), .ZN(P3_U2750) );
  INV_X1 U19984 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20035) );
  AOI22_X1 U19985 ( .A1(n17990), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17976) );
  OAI21_X1 U19986 ( .B1(n20035), .B2(n17992), .A(n17976), .ZN(P3_U2749) );
  INV_X1 U19987 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20607) );
  AOI22_X1 U19988 ( .A1(n17990), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17977) );
  OAI21_X1 U19989 ( .B1(n20607), .B2(n17992), .A(n17977), .ZN(P3_U2748) );
  INV_X1 U19990 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20038) );
  AOI22_X1 U19991 ( .A1(n17990), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17978) );
  OAI21_X1 U19992 ( .B1(n20038), .B2(n17992), .A(n17978), .ZN(P3_U2747) );
  INV_X1 U19993 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20591) );
  AOI22_X1 U19994 ( .A1(n17990), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17979) );
  OAI21_X1 U19995 ( .B1(n20591), .B2(n17992), .A(n17979), .ZN(P3_U2746) );
  INV_X1 U19996 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20041) );
  AOI22_X1 U19997 ( .A1(n17990), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17980) );
  OAI21_X1 U19998 ( .B1(n20041), .B2(n17992), .A(n17980), .ZN(P3_U2745) );
  INV_X1 U19999 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20043) );
  AOI22_X1 U20000 ( .A1(n17990), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17981) );
  OAI21_X1 U20001 ( .B1(n20043), .B2(n17992), .A(n17981), .ZN(P3_U2744) );
  INV_X1 U20002 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U20003 ( .A1(n17990), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17982), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17983) );
  OAI21_X1 U20004 ( .B1(n20045), .B2(n17992), .A(n17983), .ZN(P3_U2743) );
  INV_X1 U20005 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20626) );
  AOI22_X1 U20006 ( .A1(n17990), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17984) );
  OAI21_X1 U20007 ( .B1(n20626), .B2(n17992), .A(n17984), .ZN(P3_U2742) );
  INV_X1 U20008 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20048) );
  AOI22_X1 U20009 ( .A1(n17990), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17985) );
  OAI21_X1 U20010 ( .B1(n20048), .B2(n17992), .A(n17985), .ZN(P3_U2741) );
  INV_X1 U20011 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U20012 ( .A1(n17990), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17986) );
  OAI21_X1 U20013 ( .B1(n20655), .B2(n17992), .A(n17986), .ZN(P3_U2740) );
  INV_X1 U20014 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U20015 ( .A1(n17990), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17987) );
  OAI21_X1 U20016 ( .B1(n20051), .B2(n17992), .A(n17987), .ZN(P3_U2739) );
  INV_X1 U20017 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20643) );
  AOI22_X1 U20018 ( .A1(n17990), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17988) );
  OAI21_X1 U20019 ( .B1(n20643), .B2(n17992), .A(n17988), .ZN(P3_U2738) );
  INV_X1 U20020 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20054) );
  AOI22_X1 U20021 ( .A1(n17990), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17989), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17991) );
  OAI21_X1 U20022 ( .B1(n20054), .B2(n17992), .A(n17991), .ZN(P3_U2737) );
  AOI21_X1 U20023 ( .B1(n18012), .B2(P3_ADS_N_REG_SCAN_IN), .A(n21647), .ZN(
        n17993) );
  INV_X1 U20024 ( .A(n17993), .ZN(P3_U2633) );
  AND2_X1 U20025 ( .A1(n21698), .A2(n18006), .ZN(n18001) );
  AOI22_X1 U20026 ( .A1(n18001), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18012), .ZN(n17994) );
  OAI21_X1 U20027 ( .B1(n18005), .B2(n17995), .A(n17994), .ZN(P3_U3032) );
  AOI22_X1 U20028 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18003), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18012), .ZN(n17996) );
  OAI21_X1 U20029 ( .B1(n20116), .B2(n18008), .A(n17996), .ZN(P3_U3033) );
  INV_X1 U20030 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20825) );
  INV_X1 U20031 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19726) );
  OAI222_X1 U20032 ( .A1(n18008), .A2(n20825), .B1(n19726), .B2(n18006), .C1(
        n20116), .C2(n18005), .ZN(P3_U3034) );
  AOI22_X1 U20033 ( .A1(n18001), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n18012), .ZN(n17997) );
  OAI21_X1 U20034 ( .B1(n18005), .B2(n20825), .A(n17997), .ZN(P3_U3035) );
  AOI22_X1 U20035 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18003), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n18012), .ZN(n17998) );
  OAI21_X1 U20036 ( .B1(n20834), .B2(n18008), .A(n17998), .ZN(P3_U3036) );
  INV_X1 U20037 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20165) );
  INV_X1 U20038 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19730) );
  OAI222_X1 U20039 ( .A1(n18008), .A2(n20165), .B1(n19730), .B2(n18006), .C1(
        n20834), .C2(n18005), .ZN(P3_U3037) );
  INV_X1 U20040 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20182) );
  INV_X1 U20041 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19732) );
  OAI222_X1 U20042 ( .A1(n18008), .A2(n20182), .B1(n19732), .B2(n18006), .C1(
        n20165), .C2(n18005), .ZN(P3_U3038) );
  INV_X1 U20043 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20199) );
  INV_X1 U20044 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19734) );
  OAI222_X1 U20045 ( .A1(n18008), .A2(n20199), .B1(n19734), .B2(n18006), .C1(
        n20182), .C2(n18005), .ZN(P3_U3039) );
  INV_X1 U20046 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19736) );
  OAI222_X1 U20047 ( .A1(n18008), .A2(n20222), .B1(n19736), .B2(n18006), .C1(
        n20199), .C2(n18005), .ZN(P3_U3040) );
  INV_X1 U20048 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19738) );
  OAI222_X1 U20049 ( .A1(n18008), .A2(n20235), .B1(n19738), .B2(n18006), .C1(
        n20222), .C2(n18005), .ZN(P3_U3041) );
  INV_X1 U20050 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19740) );
  INV_X1 U20051 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20249) );
  OAI222_X1 U20052 ( .A1(n20235), .A2(n18005), .B1(n19740), .B2(n18006), .C1(
        n20249), .C2(n18008), .ZN(P3_U3042) );
  INV_X1 U20053 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20254) );
  INV_X1 U20054 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19742) );
  OAI222_X1 U20055 ( .A1(n18008), .A2(n20254), .B1(n19742), .B2(n18006), .C1(
        n20249), .C2(n18005), .ZN(P3_U3043) );
  INV_X1 U20056 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19744) );
  OAI222_X1 U20057 ( .A1(n18008), .A2(n20271), .B1(n19744), .B2(n18006), .C1(
        n20254), .C2(n18005), .ZN(P3_U3044) );
  INV_X1 U20058 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19746) );
  OAI222_X1 U20059 ( .A1(n20271), .A2(n18005), .B1(n19746), .B2(n18006), .C1(
        n20297), .C2(n18008), .ZN(P3_U3045) );
  INV_X1 U20060 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19748) );
  OAI222_X1 U20061 ( .A1(n18008), .A2(n20298), .B1(n19748), .B2(n18006), .C1(
        n20297), .C2(n18005), .ZN(P3_U3046) );
  INV_X1 U20062 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n17999) );
  INV_X1 U20063 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19750) );
  OAI222_X1 U20064 ( .A1(n18008), .A2(n17999), .B1(n19750), .B2(n18006), .C1(
        n20298), .C2(n18005), .ZN(P3_U3047) );
  INV_X1 U20065 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20337) );
  INV_X1 U20066 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19752) );
  OAI222_X1 U20067 ( .A1(n18008), .A2(n20337), .B1(n19752), .B2(n18006), .C1(
        n17999), .C2(n18005), .ZN(P3_U3048) );
  INV_X1 U20068 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20338) );
  INV_X1 U20069 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19754) );
  OAI222_X1 U20070 ( .A1(n18008), .A2(n20338), .B1(n19754), .B2(n18006), .C1(
        n20337), .C2(n18005), .ZN(P3_U3049) );
  INV_X1 U20071 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20349) );
  INV_X1 U20072 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19756) );
  OAI222_X1 U20073 ( .A1(n18008), .A2(n20349), .B1(n19756), .B2(n18006), .C1(
        n20338), .C2(n18005), .ZN(P3_U3050) );
  INV_X1 U20074 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19758) );
  OAI222_X1 U20075 ( .A1(n18008), .A2(n20370), .B1(n19758), .B2(n18006), .C1(
        n20349), .C2(n18005), .ZN(P3_U3051) );
  INV_X1 U20076 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20389) );
  INV_X1 U20077 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U20078 ( .A1(n18008), .A2(n20389), .B1(n19760), .B2(n18006), .C1(
        n20370), .C2(n18005), .ZN(P3_U3052) );
  INV_X1 U20079 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19762) );
  OAI222_X1 U20080 ( .A1(n18008), .A2(n18000), .B1(n19762), .B2(n18006), .C1(
        n20389), .C2(n18005), .ZN(P3_U3053) );
  INV_X1 U20081 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19764) );
  INV_X1 U20082 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20420) );
  OAI222_X1 U20083 ( .A1(n18000), .A2(n18005), .B1(n19764), .B2(n18006), .C1(
        n20420), .C2(n18008), .ZN(P3_U3054) );
  INV_X1 U20084 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20421) );
  INV_X1 U20085 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19766) );
  OAI222_X1 U20086 ( .A1(n18008), .A2(n20421), .B1(n19766), .B2(n18006), .C1(
        n20420), .C2(n18005), .ZN(P3_U3055) );
  INV_X1 U20087 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20428) );
  INV_X1 U20088 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19768) );
  OAI222_X1 U20089 ( .A1(n18008), .A2(n20428), .B1(n19768), .B2(n18006), .C1(
        n20421), .C2(n18005), .ZN(P3_U3056) );
  INV_X1 U20090 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20454) );
  INV_X1 U20091 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19770) );
  OAI222_X1 U20092 ( .A1(n18008), .A2(n20454), .B1(n19770), .B2(n18006), .C1(
        n20428), .C2(n18005), .ZN(P3_U3057) );
  INV_X1 U20093 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19772) );
  OAI222_X1 U20094 ( .A1(n18008), .A2(n20466), .B1(n19772), .B2(n18006), .C1(
        n20454), .C2(n18005), .ZN(P3_U3058) );
  AOI22_X1 U20095 ( .A1(n18001), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n18012), .ZN(n18002) );
  OAI21_X1 U20096 ( .B1(n18005), .B2(n20466), .A(n18002), .ZN(P3_U3059) );
  AOI22_X1 U20097 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18003), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n18012), .ZN(n18004) );
  OAI21_X1 U20098 ( .B1(n20497), .B2(n18008), .A(n18004), .ZN(P3_U3060) );
  INV_X1 U20099 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19778) );
  OAI222_X1 U20100 ( .A1(n18008), .A2(n18007), .B1(n19778), .B2(n18006), .C1(
        n20497), .C2(n18005), .ZN(P3_U3061) );
  OAI22_X1 U20101 ( .A1(n18012), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18006), .ZN(n18009) );
  INV_X1 U20102 ( .A(n18009), .ZN(P3_U3277) );
  OAI22_X1 U20103 ( .A1(n18012), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18006), .ZN(n18010) );
  INV_X1 U20104 ( .A(n18010), .ZN(P3_U3276) );
  OAI22_X1 U20105 ( .A1(n18012), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18006), .ZN(n18011) );
  INV_X1 U20106 ( .A(n18011), .ZN(P3_U3275) );
  OAI22_X1 U20107 ( .A1(n18012), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18006), .ZN(n18013) );
  INV_X1 U20108 ( .A(n18013), .ZN(P3_U3274) );
  NOR4_X1 U20109 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18016)
         );
  INV_X1 U20110 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18014) );
  NOR4_X1 U20111 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18014), .ZN(n18015) );
  NAND3_X1 U20112 ( .A1(n18016), .A2(n18015), .A3(U215), .ZN(U213) );
  NAND4_X1 U20113 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n18022), .A4(n18527), .ZN(n18017) );
  OAI211_X1 U20114 ( .C1(n18535), .C2(n18019), .A(n18018), .B(n18017), .ZN(
        n18028) );
  INV_X1 U20115 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21676) );
  NOR2_X1 U20116 ( .A1(n21665), .A2(n19164), .ZN(n18020) );
  NOR2_X1 U20117 ( .A1(n18020), .A2(n18528), .ZN(n18026) );
  AOI21_X1 U20118 ( .B1(n21669), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n18021), 
        .ZN(n18024) );
  NOR3_X1 U20119 ( .A1(n19597), .A2(n18022), .A3(n21669), .ZN(n18023) );
  MUX2_X1 U20120 ( .A(n18024), .B(n18023), .S(n16011), .Z(n18025) );
  OAI21_X1 U20121 ( .B1(n18026), .B2(n18025), .A(n18028), .ZN(n18027) );
  OAI21_X1 U20122 ( .B1(n18028), .B2(n21676), .A(n18027), .ZN(P2_U3610) );
  INV_X1 U20123 ( .A(n18410), .ZN(n18029) );
  NAND2_X1 U20124 ( .A1(n18405), .A2(n18029), .ZN(n18032) );
  NAND2_X1 U20125 ( .A1(n18380), .A2(n18030), .ZN(n18031) );
  OAI211_X1 U20126 ( .C1(n11137), .C2(n18396), .A(n18032), .B(n18031), .ZN(
        n18033) );
  INV_X1 U20127 ( .A(n18033), .ZN(n18035) );
  NAND2_X1 U20128 ( .A1(n18381), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18034) );
  OAI211_X1 U20129 ( .C1(n18283), .C2(n18036), .A(n18035), .B(n18034), .ZN(
        n18037) );
  INV_X1 U20130 ( .A(n18037), .ZN(n18042) );
  AOI22_X1 U20131 ( .A1(n18393), .A2(n18039), .B1(n18038), .B2(n18049), .ZN(
        n18041) );
  NAND2_X1 U20132 ( .A1(n18246), .A2(n18371), .ZN(n18193) );
  OAI21_X1 U20133 ( .B1(n18402), .B2(n18260), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18040) );
  NAND3_X1 U20134 ( .A1(n18042), .A2(n18041), .A3(n18040), .ZN(P2_U2855) );
  OAI22_X1 U20135 ( .A1(n18396), .A2(n11901), .B1(n18340), .B2(n13531), .ZN(
        n18045) );
  NOR2_X1 U20136 ( .A1(n18394), .A2(n18043), .ZN(n18044) );
  AOI211_X1 U20137 ( .C1(n18405), .C2(n18046), .A(n18045), .B(n18044), .ZN(
        n18047) );
  OAI21_X1 U20138 ( .B1(n18344), .B2(n12136), .A(n18047), .ZN(n18048) );
  AOI21_X1 U20139 ( .B1(n18427), .B2(n18404), .A(n18048), .ZN(n18052) );
  AOI22_X1 U20140 ( .A1(n18050), .A2(n18371), .B1(n18049), .B2(n19035), .ZN(
        n18051) );
  OAI211_X1 U20141 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18193), .A(
        n18052), .B(n18051), .ZN(P2_U2854) );
  AOI22_X1 U20142 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18381), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18402), .ZN(n18061) );
  OR2_X1 U20143 ( .A1(n19281), .A2(n18053), .ZN(n18060) );
  OAI21_X1 U20144 ( .B1(n12673), .B2(n18396), .A(n18475), .ZN(n18054) );
  AOI21_X1 U20145 ( .B1(n18405), .B2(n18055), .A(n18054), .ZN(n18059) );
  INV_X1 U20146 ( .A(n18056), .ZN(n18057) );
  NAND2_X1 U20147 ( .A1(n18380), .A2(n18057), .ZN(n18058) );
  AND4_X1 U20148 ( .A1(n18061), .A2(n18060), .A3(n18059), .A4(n18058), .ZN(
        n18067) );
  NAND2_X1 U20149 ( .A1(n18063), .A2(n18062), .ZN(n18073) );
  AND2_X1 U20150 ( .A1(n18385), .A2(n18073), .ZN(n18065) );
  AOI21_X1 U20151 ( .B1(n18074), .B2(n18065), .A(n18516), .ZN(n18064) );
  OAI21_X1 U20152 ( .B1(n18074), .B2(n18065), .A(n18064), .ZN(n18066) );
  OAI211_X1 U20153 ( .C1(n18068), .C2(n18283), .A(n18067), .B(n18066), .ZN(
        P2_U2851) );
  INV_X1 U20154 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18070) );
  OAI22_X1 U20155 ( .A1(n18070), .A2(n18340), .B1(n18069), .B2(n18394), .ZN(
        n18071) );
  AOI211_X1 U20156 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18378), .A(n18072), .B(
        n18071), .ZN(n18080) );
  NOR2_X1 U20157 ( .A1(n18074), .A2(n18073), .ZN(n18087) );
  NOR2_X1 U20158 ( .A1(n18246), .A2(n18087), .ZN(n18075) );
  XNOR2_X1 U20159 ( .A(n18086), .B(n18075), .ZN(n18078) );
  OAI22_X1 U20160 ( .A1(n18354), .A2(n19286), .B1(n18283), .B2(n18076), .ZN(
        n18077) );
  AOI21_X1 U20161 ( .B1(n18078), .B2(n18386), .A(n18077), .ZN(n18079) );
  OAI211_X1 U20162 ( .C1(n18344), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P2_U2850) );
  OAI21_X1 U20163 ( .B1(n12682), .B2(n18396), .A(n18475), .ZN(n18085) );
  OAI22_X1 U20164 ( .A1(n18083), .A2(n18340), .B1(n18082), .B2(n18394), .ZN(
        n18084) );
  AOI211_X1 U20165 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n18381), .A(n18085), .B(
        n18084), .ZN(n18092) );
  NAND2_X1 U20166 ( .A1(n18087), .A2(n18086), .ZN(n18098) );
  NAND2_X1 U20167 ( .A1(n18385), .A2(n18098), .ZN(n18088) );
  XNOR2_X1 U20168 ( .A(n18099), .B(n18088), .ZN(n18090) );
  AOI22_X1 U20169 ( .A1(n18371), .A2(n18090), .B1(n18404), .B2(n18089), .ZN(
        n18091) );
  OAI211_X1 U20170 ( .C1(n18354), .C2(n18093), .A(n18092), .B(n18091), .ZN(
        P2_U2849) );
  AOI22_X1 U20171 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n18381), .B1(n18094), .B2(
        n18380), .ZN(n18095) );
  OAI211_X1 U20172 ( .C1(n18096), .C2(n18396), .A(n18095), .B(n18475), .ZN(
        n18097) );
  AOI21_X1 U20173 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18402), .A(
        n18097), .ZN(n18104) );
  NOR2_X1 U20174 ( .A1(n18099), .A2(n18098), .ZN(n18111) );
  NOR2_X1 U20175 ( .A1(n18246), .A2(n18111), .ZN(n18100) );
  XNOR2_X1 U20176 ( .A(n18100), .B(n18110), .ZN(n18102) );
  AOI22_X1 U20177 ( .A1(n18371), .A2(n18102), .B1(n18405), .B2(n18101), .ZN(
        n18103) );
  OAI211_X1 U20178 ( .C1(n18283), .C2(n18105), .A(n18104), .B(n18103), .ZN(
        P2_U2848) );
  OAI21_X1 U20179 ( .B1(n12688), .B2(n18396), .A(n18475), .ZN(n18109) );
  OAI22_X1 U20180 ( .A1(n18107), .A2(n18340), .B1(n18106), .B2(n18394), .ZN(
        n18108) );
  AOI211_X1 U20181 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18381), .A(n18109), .B(
        n18108), .ZN(n18116) );
  NAND2_X1 U20182 ( .A1(n18111), .A2(n18110), .ZN(n18118) );
  NAND2_X1 U20183 ( .A1(n18257), .A2(n18118), .ZN(n18112) );
  XNOR2_X1 U20184 ( .A(n18119), .B(n18112), .ZN(n18114) );
  AOI22_X1 U20185 ( .A1(n18371), .A2(n18114), .B1(n18405), .B2(n18113), .ZN(
        n18115) );
  OAI211_X1 U20186 ( .C1(n18283), .C2(n18117), .A(n18116), .B(n18115), .ZN(
        P2_U2847) );
  NOR2_X1 U20187 ( .A1(n18119), .A2(n18118), .ZN(n18133) );
  NOR2_X1 U20188 ( .A1(n18246), .A2(n18133), .ZN(n18120) );
  XOR2_X1 U20189 ( .A(n18132), .B(n18120), .Z(n18128) );
  AOI22_X1 U20190 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18402), .B1(
        n18121), .B2(n18380), .ZN(n18122) );
  OAI211_X1 U20191 ( .C1(n12694), .C2(n18396), .A(n18122), .B(n18475), .ZN(
        n18126) );
  OAI22_X1 U20192 ( .A1(n18124), .A2(n18283), .B1(n18123), .B2(n18354), .ZN(
        n18125) );
  AOI211_X1 U20193 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18381), .A(n18126), .B(
        n18125), .ZN(n18127) );
  OAI21_X1 U20194 ( .B1(n18516), .B2(n18128), .A(n18127), .ZN(P2_U2846) );
  AOI22_X1 U20195 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18402), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n18381), .ZN(n18129) );
  OAI21_X1 U20196 ( .B1(n18130), .B2(n18394), .A(n18129), .ZN(n18131) );
  AOI211_X1 U20197 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18378), .A(n16539), 
        .B(n18131), .ZN(n18138) );
  NAND2_X1 U20198 ( .A1(n18133), .A2(n18132), .ZN(n18148) );
  NAND2_X1 U20199 ( .A1(n18385), .A2(n18148), .ZN(n18134) );
  XOR2_X1 U20200 ( .A(n18147), .B(n18134), .Z(n18135) );
  AOI22_X1 U20201 ( .A1(n18136), .A2(n18405), .B1(n18371), .B2(n18135), .ZN(
        n18137) );
  OAI211_X1 U20202 ( .C1(n18139), .C2(n18283), .A(n18138), .B(n18137), .ZN(
        P2_U2845) );
  OAI22_X1 U20203 ( .A1(n18344), .A2(n18141), .B1(n18140), .B2(n18340), .ZN(
        n18146) );
  AOI22_X1 U20204 ( .A1(n18143), .A2(n18380), .B1(n18142), .B2(n18405), .ZN(
        n18144) );
  OAI211_X1 U20205 ( .C1(n16417), .C2(n18396), .A(n18144), .B(n18240), .ZN(
        n18145) );
  AOI211_X1 U20206 ( .C1(n11379), .C2(n18404), .A(n18146), .B(n18145), .ZN(
        n18153) );
  INV_X1 U20207 ( .A(n18147), .ZN(n18149) );
  NOR2_X1 U20208 ( .A1(n18149), .A2(n18148), .ZN(n18151) );
  NAND2_X1 U20209 ( .A1(n18151), .A2(n18154), .ZN(n18170) );
  NAND2_X1 U20210 ( .A1(n18257), .A2(n18170), .ZN(n18158) );
  INV_X1 U20211 ( .A(n18158), .ZN(n18150) );
  OAI211_X1 U20212 ( .C1(n18151), .C2(n18154), .A(n18386), .B(n18150), .ZN(
        n18152) );
  OAI211_X1 U20213 ( .C1(n18193), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        P2_U2844) );
  AOI22_X1 U20214 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18402), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18381), .ZN(n18155) );
  OAI21_X1 U20215 ( .B1(n18156), .B2(n18394), .A(n18155), .ZN(n18157) );
  AOI211_X1 U20216 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18378), .A(n16539), 
        .B(n18157), .ZN(n18161) );
  XOR2_X1 U20217 ( .A(n18169), .B(n18158), .Z(n18159) );
  AOI22_X1 U20218 ( .A1(n18465), .A2(n18405), .B1(n18386), .B2(n18159), .ZN(
        n18160) );
  OAI211_X1 U20219 ( .C1(n18162), .C2(n18283), .A(n18161), .B(n18160), .ZN(
        P2_U2843) );
  OAI22_X1 U20220 ( .A1(n18344), .A2(n18164), .B1(n18163), .B2(n18340), .ZN(
        n18168) );
  AOI22_X1 U20221 ( .A1(n18165), .A2(n18380), .B1(n18172), .B2(n18260), .ZN(
        n18166) );
  OAI211_X1 U20222 ( .C1(n12706), .C2(n18396), .A(n18166), .B(n18240), .ZN(
        n18167) );
  AOI211_X1 U20223 ( .C1(n18454), .C2(n18404), .A(n18168), .B(n18167), .ZN(
        n18177) );
  INV_X1 U20224 ( .A(n18169), .ZN(n18171) );
  NOR2_X1 U20225 ( .A1(n18171), .A2(n18170), .ZN(n18175) );
  INV_X1 U20226 ( .A(n18172), .ZN(n18174) );
  NAND2_X1 U20227 ( .A1(n18175), .A2(n18174), .ZN(n18198) );
  NAND2_X1 U20228 ( .A1(n18393), .A2(n18198), .ZN(n18189) );
  INV_X1 U20229 ( .A(n18189), .ZN(n18173) );
  OAI21_X1 U20230 ( .B1(n18175), .B2(n18174), .A(n18173), .ZN(n18176) );
  OAI211_X1 U20231 ( .C1(n18354), .C2(n18448), .A(n18177), .B(n18176), .ZN(
        P2_U2842) );
  INV_X1 U20232 ( .A(n18178), .ZN(n18199) );
  AOI22_X1 U20233 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n18381), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18402), .ZN(n18181) );
  INV_X1 U20234 ( .A(n18198), .ZN(n18179) );
  OAI211_X1 U20235 ( .C1(n18246), .C2(n18179), .A(n18199), .B(n18371), .ZN(
        n18180) );
  OAI211_X1 U20236 ( .C1(n18394), .C2(n18182), .A(n18181), .B(n18180), .ZN(
        n18183) );
  AOI211_X1 U20237 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18378), .A(n16539), 
        .B(n18183), .ZN(n18188) );
  INV_X1 U20238 ( .A(n18184), .ZN(n18185) );
  AOI22_X1 U20239 ( .A1(n18186), .A2(n18404), .B1(n18185), .B2(n18405), .ZN(
        n18187) );
  OAI211_X1 U20240 ( .C1(n18199), .C2(n18189), .A(n18188), .B(n18187), .ZN(
        P2_U2841) );
  AOI22_X1 U20241 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18402), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n18381), .ZN(n18190) );
  OAI211_X1 U20242 ( .C1(n18191), .C2(n18396), .A(n18190), .B(n18240), .ZN(
        n18196) );
  INV_X1 U20243 ( .A(n18192), .ZN(n18200) );
  OAI22_X1 U20244 ( .A1(n18194), .A2(n18394), .B1(n18200), .B2(n18193), .ZN(
        n18195) );
  AOI211_X1 U20245 ( .C1(n18197), .C2(n18404), .A(n18196), .B(n18195), .ZN(
        n18203) );
  NOR2_X1 U20246 ( .A1(n18199), .A2(n18198), .ZN(n18201) );
  NAND2_X1 U20247 ( .A1(n18201), .A2(n18200), .ZN(n18223) );
  AND2_X1 U20248 ( .A1(n18257), .A2(n18223), .ZN(n18206) );
  OAI211_X1 U20249 ( .C1(n18201), .C2(n18200), .A(n18386), .B(n18206), .ZN(
        n18202) );
  OAI211_X1 U20250 ( .C1(n18354), .C2(n18204), .A(n18203), .B(n18202), .ZN(
        P2_U2840) );
  INV_X1 U20251 ( .A(n18205), .ZN(n18224) );
  XNOR2_X1 U20252 ( .A(n18206), .B(n18224), .ZN(n18214) );
  AOI22_X1 U20253 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18402), .B1(
        n18207), .B2(n18380), .ZN(n18208) );
  OAI211_X1 U20254 ( .C1(n12721), .C2(n18396), .A(n18208), .B(n18240), .ZN(
        n18212) );
  OAI22_X1 U20255 ( .A1(n18210), .A2(n18283), .B1(n18209), .B2(n18354), .ZN(
        n18211) );
  AOI211_X1 U20256 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18381), .A(n18212), .B(
        n18211), .ZN(n18213) );
  OAI21_X1 U20257 ( .B1(n18214), .B2(n18516), .A(n18213), .ZN(P2_U2839) );
  AOI22_X1 U20258 ( .A1(n18381), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18402), .ZN(n18215) );
  INV_X1 U20259 ( .A(n18215), .ZN(n18221) );
  AOI22_X1 U20260 ( .A1(n18217), .A2(n18380), .B1(n18216), .B2(n18260), .ZN(
        n18218) );
  OAI211_X1 U20261 ( .C1(n18219), .C2(n18396), .A(n18218), .B(n18240), .ZN(
        n18220) );
  AOI211_X1 U20262 ( .C1(n18222), .C2(n18404), .A(n18221), .B(n18220), .ZN(
        n18228) );
  NOR2_X1 U20263 ( .A1(n18224), .A2(n18223), .ZN(n18226) );
  NAND2_X1 U20264 ( .A1(n18226), .A2(n18225), .ZN(n18244) );
  OAI211_X1 U20265 ( .C1(n18226), .C2(n18225), .A(n18393), .B(n18244), .ZN(
        n18227) );
  OAI211_X1 U20266 ( .C1(n18354), .C2(n18229), .A(n18228), .B(n18227), .ZN(
        P2_U2838) );
  NAND2_X1 U20267 ( .A1(n18257), .A2(n18244), .ZN(n18230) );
  XOR2_X1 U20268 ( .A(n18245), .B(n18230), .Z(n18238) );
  AOI22_X1 U20269 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18402), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18381), .ZN(n18231) );
  OAI21_X1 U20270 ( .B1(n18232), .B2(n18394), .A(n18231), .ZN(n18233) );
  AOI211_X1 U20271 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18378), .A(n16539), 
        .B(n18233), .ZN(n18237) );
  AOI22_X1 U20272 ( .A1(n18235), .A2(n18404), .B1(n18234), .B2(n18405), .ZN(
        n18236) );
  OAI211_X1 U20273 ( .C1(n18516), .C2(n18238), .A(n18237), .B(n18236), .ZN(
        P2_U2837) );
  AOI22_X1 U20274 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n18381), .B1(n18239), 
        .B2(n18380), .ZN(n18241) );
  OAI211_X1 U20275 ( .C1(n18242), .C2(n18396), .A(n18241), .B(n18240), .ZN(
        n18243) );
  AOI21_X1 U20276 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18402), .A(
        n18243), .ZN(n18251) );
  NOR2_X1 U20277 ( .A1(n18245), .A2(n18244), .ZN(n18256) );
  NOR2_X1 U20278 ( .A1(n18246), .A2(n18256), .ZN(n18247) );
  XOR2_X1 U20279 ( .A(n18247), .B(n18254), .Z(n18248) );
  AOI22_X1 U20280 ( .A1(n18249), .A2(n18404), .B1(n18386), .B2(n18248), .ZN(
        n18250) );
  OAI211_X1 U20281 ( .C1(n18252), .C2(n18354), .A(n18251), .B(n18250), .ZN(
        P2_U2836) );
  INV_X1 U20282 ( .A(n18253), .ZN(n18261) );
  INV_X1 U20283 ( .A(n18254), .ZN(n18255) );
  NAND2_X1 U20284 ( .A1(n18256), .A2(n18255), .ZN(n18258) );
  OAI21_X1 U20285 ( .B1(n18261), .B2(n18258), .A(n18257), .ZN(n18276) );
  AOI21_X1 U20286 ( .B1(n18261), .B2(n18258), .A(n18276), .ZN(n18259) );
  AOI22_X1 U20287 ( .A1(n18261), .A2(n18260), .B1(n18371), .B2(n18259), .ZN(
        n18268) );
  INV_X1 U20288 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18263) );
  OAI22_X1 U20289 ( .A1(n18344), .A2(n18263), .B1(n18262), .B2(n18394), .ZN(
        n18266) );
  AOI22_X1 U20290 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18378), .ZN(n18264) );
  INV_X1 U20291 ( .A(n18264), .ZN(n18265) );
  AOI211_X1 U20292 ( .C1(n19344), .C2(n18405), .A(n18266), .B(n18265), .ZN(
        n18267) );
  OAI211_X1 U20293 ( .C1(n18269), .C2(n18283), .A(n18268), .B(n18267), .ZN(
        P2_U2835) );
  AOI22_X1 U20294 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18378), .ZN(n18280) );
  AOI22_X1 U20295 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18381), .B1(n18270), 
        .B2(n18380), .ZN(n18279) );
  INV_X1 U20296 ( .A(n18271), .ZN(n18272) );
  AOI22_X1 U20297 ( .A1(n18273), .A2(n18404), .B1(n18272), .B2(n18405), .ZN(
        n18278) );
  INV_X1 U20298 ( .A(n18274), .ZN(n18275) );
  NAND2_X1 U20299 ( .A1(n18275), .A2(n18276), .ZN(n18286) );
  OAI211_X1 U20300 ( .C1(n18276), .C2(n18275), .A(n18386), .B(n18286), .ZN(
        n18277) );
  NAND4_X1 U20301 ( .A1(n18280), .A2(n18279), .A3(n18278), .A4(n18277), .ZN(
        P2_U2834) );
  AOI22_X1 U20302 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18378), .ZN(n18292) );
  AOI22_X1 U20303 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18381), .B1(n18281), 
        .B2(n18380), .ZN(n18291) );
  OAI22_X1 U20304 ( .A1(n18284), .A2(n18283), .B1(n18282), .B2(n18354), .ZN(
        n18285) );
  INV_X1 U20305 ( .A(n18285), .ZN(n18290) );
  NAND2_X1 U20306 ( .A1(n18385), .A2(n18286), .ZN(n18288) );
  NAND2_X1 U20307 ( .A1(n18287), .A2(n18288), .ZN(n18301) );
  OAI211_X1 U20308 ( .C1(n18288), .C2(n18287), .A(n18386), .B(n18301), .ZN(
        n18289) );
  NAND4_X1 U20309 ( .A1(n18292), .A2(n18291), .A3(n18290), .A4(n18289), .ZN(
        P2_U2833) );
  INV_X1 U20310 ( .A(n18293), .ZN(n18300) );
  OAI22_X1 U20311 ( .A1(n18295), .A2(n18340), .B1(n18294), .B2(n18396), .ZN(
        n18299) );
  INV_X1 U20312 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n18297) );
  OAI22_X1 U20313 ( .A1(n18344), .A2(n18297), .B1(n18296), .B2(n18394), .ZN(
        n18298) );
  AOI211_X1 U20314 ( .C1(n18300), .C2(n18404), .A(n18299), .B(n18298), .ZN(
        n18305) );
  INV_X1 U20315 ( .A(n18302), .ZN(n18303) );
  OAI211_X1 U20316 ( .C1(n18354), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P2_U2832) );
  AOI22_X1 U20317 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18378), .ZN(n18316) );
  AOI22_X1 U20318 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18381), .B1(n18307), 
        .B2(n18380), .ZN(n18315) );
  AOI22_X1 U20319 ( .A1(n18309), .A2(n18404), .B1(n18308), .B2(n18405), .ZN(
        n18314) );
  NAND2_X1 U20320 ( .A1(n18385), .A2(n18310), .ZN(n18312) );
  NAND2_X1 U20321 ( .A1(n18311), .A2(n18312), .ZN(n18320) );
  OAI211_X1 U20322 ( .C1(n18312), .C2(n18311), .A(n18386), .B(n18320), .ZN(
        n18313) );
  NAND4_X1 U20323 ( .A1(n18316), .A2(n18315), .A3(n18314), .A4(n18313), .ZN(
        P2_U2831) );
  AOI22_X1 U20324 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18378), .ZN(n18327) );
  AOI22_X1 U20325 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18381), .B1(n18317), 
        .B2(n18380), .ZN(n18326) );
  AOI22_X1 U20326 ( .A1(n18319), .A2(n18404), .B1(n18318), .B2(n18405), .ZN(
        n18325) );
  NAND2_X1 U20327 ( .A1(n18385), .A2(n18320), .ZN(n18323) );
  INV_X1 U20328 ( .A(n18321), .ZN(n18322) );
  NAND2_X1 U20329 ( .A1(n18322), .A2(n18323), .ZN(n18332) );
  OAI211_X1 U20330 ( .C1(n18323), .C2(n18322), .A(n18371), .B(n18332), .ZN(
        n18324) );
  NAND4_X1 U20331 ( .A1(n18327), .A2(n18326), .A3(n18325), .A4(n18324), .ZN(
        P2_U2830) );
  AOI22_X1 U20332 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18378), .ZN(n18338) );
  AOI22_X1 U20333 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18381), .B1(n18328), 
        .B2(n18380), .ZN(n18337) );
  INV_X1 U20334 ( .A(n18329), .ZN(n18331) );
  AOI22_X1 U20335 ( .A1(n18331), .A2(n18404), .B1(n18330), .B2(n18405), .ZN(
        n18336) );
  OAI211_X1 U20336 ( .C1(n18334), .C2(n18333), .A(n18371), .B(n18348), .ZN(
        n18335) );
  NAND4_X1 U20337 ( .A1(n18338), .A2(n18337), .A3(n18336), .A4(n18335), .ZN(
        P2_U2829) );
  OAI22_X1 U20338 ( .A1(n18341), .A2(n18340), .B1(n18339), .B2(n18396), .ZN(
        n18346) );
  INV_X1 U20339 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n18343) );
  OAI22_X1 U20340 ( .A1(n18344), .A2(n18343), .B1(n18342), .B2(n18394), .ZN(
        n18345) );
  AOI211_X1 U20341 ( .C1(n18347), .C2(n18404), .A(n18346), .B(n18345), .ZN(
        n18352) );
  NAND2_X1 U20342 ( .A1(n18385), .A2(n18348), .ZN(n18350) );
  NAND2_X1 U20343 ( .A1(n18349), .A2(n18350), .ZN(n18358) );
  OAI211_X1 U20344 ( .C1(n18350), .C2(n18349), .A(n18371), .B(n18358), .ZN(
        n18351) );
  OAI211_X1 U20345 ( .C1(n18354), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        P2_U2828) );
  AOI22_X1 U20346 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18378), .ZN(n18364) );
  AOI22_X1 U20347 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18381), .B1(n18355), 
        .B2(n18380), .ZN(n18363) );
  AOI22_X1 U20348 ( .A1(n18357), .A2(n18404), .B1(n18356), .B2(n18405), .ZN(
        n18362) );
  OAI211_X1 U20349 ( .C1(n18360), .C2(n18359), .A(n18371), .B(n18369), .ZN(
        n18361) );
  NAND4_X1 U20350 ( .A1(n18364), .A2(n18363), .A3(n18362), .A4(n18361), .ZN(
        P2_U2827) );
  AOI22_X1 U20351 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18378), .ZN(n18377) );
  AOI22_X1 U20352 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18381), .B1(n18365), 
        .B2(n18380), .ZN(n18376) );
  INV_X1 U20353 ( .A(n18366), .ZN(n18367) );
  AOI22_X1 U20354 ( .A1(n18368), .A2(n18404), .B1(n18367), .B2(n18405), .ZN(
        n18375) );
  NAND2_X1 U20355 ( .A1(n18257), .A2(n18369), .ZN(n18373) );
  INV_X1 U20356 ( .A(n18370), .ZN(n18372) );
  NAND2_X1 U20357 ( .A1(n18372), .A2(n18373), .ZN(n18384) );
  OAI211_X1 U20358 ( .C1(n18373), .C2(n18372), .A(n18371), .B(n18384), .ZN(
        n18374) );
  NAND4_X1 U20359 ( .A1(n18377), .A2(n18376), .A3(n18375), .A4(n18374), .ZN(
        P2_U2826) );
  AOI22_X1 U20360 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18402), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18378), .ZN(n18392) );
  AOI22_X1 U20361 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18381), .B1(n18380), 
        .B2(n18379), .ZN(n18391) );
  AOI22_X1 U20362 ( .A1(n18383), .A2(n18404), .B1(n18382), .B2(n18405), .ZN(
        n18390) );
  NAND2_X1 U20363 ( .A1(n18385), .A2(n18384), .ZN(n18388) );
  NAND2_X1 U20364 ( .A1(n18387), .A2(n18388), .ZN(n18409) );
  OAI211_X1 U20365 ( .C1(n18388), .C2(n18387), .A(n18386), .B(n18409), .ZN(
        n18389) );
  NAND4_X1 U20366 ( .A1(n18392), .A2(n18391), .A3(n18390), .A4(n18389), .ZN(
        P2_U2825) );
  INV_X1 U20367 ( .A(n18393), .ZN(n18408) );
  NOR2_X1 U20368 ( .A1(n18395), .A2(n18394), .ZN(n18401) );
  OAI22_X1 U20369 ( .A1(n18399), .A2(n18398), .B1(n18397), .B2(n18396), .ZN(
        n18400) );
  AOI211_X1 U20370 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n18402), .A(
        n18401), .B(n18400), .ZN(n18407) );
  AOI22_X1 U20371 ( .A1(n18405), .A2(n18994), .B1(n18404), .B2(n18403), .ZN(
        n18406) );
  OAI211_X1 U20372 ( .C1(n18409), .C2(n18408), .A(n18407), .B(n18406), .ZN(
        P2_U2824) );
  OAI22_X1 U20373 ( .A1(n18411), .A2(n18450), .B1(n18490), .B2(n18410), .ZN(
        n18412) );
  INV_X1 U20374 ( .A(n18412), .ZN(n18421) );
  AOI21_X1 U20375 ( .B1(n18481), .B2(n18414), .A(n18413), .ZN(n18417) );
  NAND2_X1 U20376 ( .A1(n18500), .A2(n18415), .ZN(n18416) );
  OAI211_X1 U20377 ( .C1(n18418), .C2(n18509), .A(n18417), .B(n18416), .ZN(
        n18419) );
  INV_X1 U20378 ( .A(n18419), .ZN(n18420) );
  OAI211_X1 U20379 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18422), .A(
        n18421), .B(n18420), .ZN(P2_U3046) );
  OR2_X1 U20380 ( .A1(n18423), .A2(n18450), .ZN(n18432) );
  OAI22_X1 U20381 ( .A1(n18425), .A2(n18490), .B1(n18494), .B2(n18424), .ZN(
        n18426) );
  INV_X1 U20382 ( .A(n18426), .ZN(n18431) );
  NAND2_X1 U20383 ( .A1(n18500), .A2(n18427), .ZN(n18430) );
  OAI211_X1 U20384 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n18460), .B(n18428), .ZN(n18429) );
  AND4_X1 U20385 ( .A1(n18432), .A2(n18431), .A3(n18430), .A4(n18429), .ZN(
        n18434) );
  OAI211_X1 U20386 ( .C1(n18509), .C2(n18435), .A(n18434), .B(n18433), .ZN(
        P2_U3045) );
  NOR2_X1 U20387 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18436), .ZN(
        n18445) );
  OAI22_X1 U20388 ( .A1(n18490), .A2(n18438), .B1(n18475), .B2(n18437), .ZN(
        n18439) );
  INV_X1 U20389 ( .A(n18439), .ZN(n18444) );
  AOI222_X1 U20390 ( .A1(n18442), .A2(n18501), .B1(n18500), .B2(n18441), .C1(
        n18481), .C2(n18440), .ZN(n18443) );
  OAI211_X1 U20391 ( .C1(n18446), .C2(n18445), .A(n18444), .B(n18443), .ZN(
        P2_U3036) );
  OAI22_X1 U20392 ( .A1(n18448), .A2(n18490), .B1(n12702), .B2(n18447), .ZN(
        n18449) );
  AOI21_X1 U20393 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n16539), .A(n18449), 
        .ZN(n18456) );
  OAI22_X1 U20394 ( .A1(n18452), .A2(n18494), .B1(n18451), .B2(n18450), .ZN(
        n18453) );
  AOI21_X1 U20395 ( .B1(n18500), .B2(n18454), .A(n18453), .ZN(n18455) );
  OAI211_X1 U20396 ( .C1(n18458), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        P2_U3033) );
  AOI21_X1 U20397 ( .B1(n18461), .B2(n18460), .A(n18459), .ZN(n18472) );
  NOR2_X1 U20398 ( .A1(n18475), .A2(n18462), .ZN(n18463) );
  AOI211_X1 U20399 ( .C1(n18466), .C2(n18465), .A(n18464), .B(n18463), .ZN(
        n18471) );
  AOI222_X1 U20400 ( .A1(n18469), .A2(n18501), .B1(n18500), .B2(n18468), .C1(
        n18467), .C2(n18481), .ZN(n18470) );
  OAI211_X1 U20401 ( .C1(n18472), .C2(n12702), .A(n18471), .B(n18470), .ZN(
        P2_U3034) );
  AOI221_X1 U20402 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12230), .C2(n18474), .A(
        n18473), .ZN(n18478) );
  OAI22_X1 U20403 ( .A1(n18490), .A2(n18476), .B1(n12688), .B2(n18475), .ZN(
        n18477) );
  NOR2_X1 U20404 ( .A1(n18478), .A2(n18477), .ZN(n18484) );
  AOI222_X1 U20405 ( .A1(n18482), .A2(n18481), .B1(n18500), .B2(n18480), .C1(
        n18501), .C2(n18479), .ZN(n18483) );
  OAI211_X1 U20406 ( .C1(n18485), .C2(n12230), .A(n18484), .B(n18483), .ZN(
        P2_U3038) );
  INV_X1 U20407 ( .A(n18486), .ZN(n18487) );
  NAND2_X1 U20408 ( .A1(n18488), .A2(n18487), .ZN(n18492) );
  OAI22_X1 U20409 ( .A1(n18491), .A2(n18490), .B1(n18489), .B2(n18492), .ZN(
        n18498) );
  INV_X1 U20410 ( .A(n18492), .ZN(n18496) );
  OAI22_X1 U20411 ( .A1(n18496), .A2(n18495), .B1(n18494), .B2(n18493), .ZN(
        n18497) );
  NOR2_X1 U20412 ( .A1(n18498), .A2(n18497), .ZN(n18505) );
  NAND2_X1 U20413 ( .A1(n18500), .A2(n18499), .ZN(n18504) );
  NAND2_X1 U20414 ( .A1(n18502), .A2(n18501), .ZN(n18503) );
  AND3_X1 U20415 ( .A1(n18505), .A2(n18504), .A3(n18503), .ZN(n18507) );
  OAI211_X1 U20416 ( .C1(n18509), .C2(n18508), .A(n18507), .B(n18506), .ZN(
        P2_U3044) );
  NAND2_X1 U20417 ( .A1(n18524), .A2(n18510), .ZN(n18526) );
  OAI21_X1 U20418 ( .B1(n18512), .B2(n18511), .A(n18532), .ZN(n18515) );
  NAND2_X1 U20419 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21665), .ZN(n18513) );
  AOI21_X1 U20420 ( .B1(n18518), .B2(n18526), .A(n18513), .ZN(n18514) );
  AOI21_X1 U20421 ( .B1(n18526), .B2(n18515), .A(n18514), .ZN(n18517) );
  NAND2_X1 U20422 ( .A1(n18517), .A2(n18516), .ZN(P2_U3177) );
  OAI22_X1 U20423 ( .A1(n18520), .A2(n18519), .B1(n18518), .B2(n18527), .ZN(
        n18522) );
  OR2_X1 U20424 ( .A1(n18522), .A2(n18521), .ZN(n18523) );
  AOI21_X1 U20425 ( .B1(n18524), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18523), 
        .ZN(n18531) );
  NOR2_X1 U20426 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18525), .ZN(n18529) );
  OAI22_X1 U20427 ( .A1(n18529), .A2(n18528), .B1(n18527), .B2(n18526), .ZN(
        n18530) );
  OAI211_X1 U20428 ( .C1(n18533), .C2(n18532), .A(n18531), .B(n18530), .ZN(
        P2_U3176) );
  NAND2_X1 U20429 ( .A1(n18535), .A2(n18534), .ZN(n18539) );
  NAND2_X1 U20430 ( .A1(n18539), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18536) );
  OAI21_X1 U20431 ( .B1(n18539), .B2(n18537), .A(n18536), .ZN(P2_U3609) );
  AOI21_X1 U20432 ( .B1(n18539), .B2(P2_FLUSH_REG_SCAN_IN), .A(n18538), .ZN(
        n18540) );
  INV_X1 U20433 ( .A(n18540), .ZN(P2_U2819) );
  INV_X1 U20434 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20014) );
  INV_X1 U20435 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18569) );
  AOI22_X1 U20436 ( .A1(n18890), .A2(n20014), .B1(n18569), .B2(U215), .ZN(U282) );
  OAI22_X1 U20437 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18890), .ZN(n18541) );
  INV_X1 U20438 ( .A(n18541), .ZN(U281) );
  OAI22_X1 U20439 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18890), .ZN(n18542) );
  INV_X1 U20440 ( .A(n18542), .ZN(U280) );
  OAI22_X1 U20441 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18890), .ZN(n18543) );
  INV_X1 U20442 ( .A(n18543), .ZN(U279) );
  OAI22_X1 U20443 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18890), .ZN(n18544) );
  INV_X1 U20444 ( .A(n18544), .ZN(U278) );
  OAI22_X1 U20445 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18890), .ZN(n18545) );
  INV_X1 U20446 ( .A(n18545), .ZN(U277) );
  OAI22_X1 U20447 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18890), .ZN(n18546) );
  INV_X1 U20448 ( .A(n18546), .ZN(U276) );
  OAI22_X1 U20449 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18890), .ZN(n18547) );
  INV_X1 U20450 ( .A(n18547), .ZN(U275) );
  OAI22_X1 U20451 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18890), .ZN(n18548) );
  INV_X1 U20452 ( .A(n18548), .ZN(U274) );
  OAI22_X1 U20453 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n18890), .ZN(n18549) );
  INV_X1 U20454 ( .A(n18549), .ZN(U273) );
  OAI22_X1 U20455 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18890), .ZN(n18550) );
  INV_X1 U20456 ( .A(n18550), .ZN(U272) );
  OAI22_X1 U20457 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18890), .ZN(n18551) );
  INV_X1 U20458 ( .A(n18551), .ZN(U271) );
  OAI22_X1 U20459 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18564), .ZN(n18552) );
  INV_X1 U20460 ( .A(n18552), .ZN(U270) );
  OAI22_X1 U20461 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18890), .ZN(n18553) );
  INV_X1 U20462 ( .A(n18553), .ZN(U269) );
  OAI22_X1 U20463 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18564), .ZN(n18554) );
  INV_X1 U20464 ( .A(n18554), .ZN(U268) );
  OAI22_X1 U20465 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18890), .ZN(n18555) );
  INV_X1 U20466 ( .A(n18555), .ZN(U267) );
  OAI22_X1 U20467 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18564), .ZN(n18556) );
  INV_X1 U20468 ( .A(n18556), .ZN(U266) );
  OAI22_X1 U20469 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18890), .ZN(n18557) );
  INV_X1 U20470 ( .A(n18557), .ZN(U265) );
  OAI22_X1 U20471 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18564), .ZN(n18558) );
  INV_X1 U20472 ( .A(n18558), .ZN(U264) );
  OAI22_X1 U20473 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18564), .ZN(n18559) );
  INV_X1 U20474 ( .A(n18559), .ZN(U263) );
  OAI22_X1 U20475 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18564), .ZN(n18560) );
  INV_X1 U20476 ( .A(n18560), .ZN(U262) );
  OAI22_X1 U20477 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18564), .ZN(n18561) );
  INV_X1 U20478 ( .A(n18561), .ZN(U261) );
  OAI22_X1 U20479 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18564), .ZN(n18562) );
  INV_X1 U20480 ( .A(n18562), .ZN(U260) );
  OAI22_X1 U20481 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18564), .ZN(n18563) );
  INV_X1 U20482 ( .A(n18563), .ZN(U259) );
  OAI22_X1 U20483 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18564), .ZN(n18565) );
  INV_X1 U20484 ( .A(n18565), .ZN(U258) );
  NOR2_X1 U20485 ( .A1(n21156), .A2(n18590), .ZN(n18634) );
  NAND2_X1 U20486 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18634), .ZN(
        n18799) );
  NOR2_X1 U20487 ( .A1(n18567), .A2(n18566), .ZN(n18685) );
  NAND2_X1 U20488 ( .A1(n18685), .A2(n20625), .ZN(n18645) );
  NAND2_X1 U20489 ( .A1(n20081), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21167) );
  AND2_X1 U20490 ( .A1(n21167), .A2(n18634), .ZN(n18896) );
  INV_X1 U20491 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20671) );
  NOR2_X2 U20492 ( .A1(n20671), .A2(n18765), .ZN(n18638) );
  NOR2_X1 U20493 ( .A1(n21153), .A2(n21156), .ZN(n18577) );
  NOR2_X1 U20494 ( .A1(n21144), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18617) );
  NAND2_X1 U20495 ( .A1(n18577), .A2(n18617), .ZN(n18902) );
  INV_X1 U20496 ( .A(n18902), .ZN(n18986) );
  AND2_X1 U20497 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18894), .ZN(n18637) );
  AOI22_X1 U20498 ( .A1(n18896), .A2(n18638), .B1(n18986), .B2(n18637), .ZN(
        n18571) );
  NAND2_X1 U20499 ( .A1(n18895), .A2(n18568), .ZN(n18576) );
  AOI21_X1 U20500 ( .B1(n21147), .B2(n18893), .A(n18576), .ZN(n18624) );
  NAND2_X1 U20501 ( .A1(n18577), .A2(n18624), .ZN(n18899) );
  NAND2_X1 U20502 ( .A1(n21147), .A2(n21144), .ZN(n21149) );
  INV_X1 U20503 ( .A(n18577), .ZN(n18575) );
  NOR2_X2 U20504 ( .A1(n21149), .A2(n18575), .ZN(n18914) );
  NOR2_X2 U20505 ( .A1(n18569), .A2(n18893), .ZN(n18642) );
  AOI22_X1 U20506 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18899), .B1(
        n18914), .B2(n18642), .ZN(n18570) );
  OAI211_X1 U20507 ( .C1(n18799), .C2(n18645), .A(n18571), .B(n18570), .ZN(
        P3_U2995) );
  NAND2_X1 U20508 ( .A1(n18634), .A2(n21144), .ZN(n18993) );
  NOR2_X1 U20509 ( .A1(n21147), .A2(n18595), .ZN(n18586) );
  NAND2_X1 U20510 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18586), .ZN(
        n18912) );
  INV_X1 U20511 ( .A(n18912), .ZN(n18919) );
  INV_X1 U20512 ( .A(n21167), .ZN(n20083) );
  AOI21_X1 U20513 ( .B1(n18902), .B2(n18993), .A(n20083), .ZN(n18903) );
  AOI22_X1 U20514 ( .A1(n18642), .A2(n18919), .B1(n18638), .B2(n18903), .ZN(
        n18574) );
  INV_X1 U20515 ( .A(n18993), .ZN(n18904) );
  INV_X1 U20516 ( .A(n18914), .ZN(n18852) );
  NAND2_X1 U20517 ( .A1(n18852), .A2(n18912), .ZN(n18582) );
  INV_X1 U20518 ( .A(n18582), .ZN(n18580) );
  OAI22_X1 U20519 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18902), .B1(n18580), 
        .B2(n18609), .ZN(n18572) );
  OAI21_X1 U20520 ( .B1(n18904), .B2(n18572), .A(n18895), .ZN(n18905) );
  AOI22_X1 U20521 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18905), .B1(
        n18914), .B2(n18637), .ZN(n18573) );
  OAI211_X1 U20522 ( .C1(n18645), .C2(n18993), .A(n18574), .B(n18573), .ZN(
        P3_U2987) );
  NAND2_X1 U20523 ( .A1(n21147), .A2(n21167), .ZN(n18631) );
  NOR2_X1 U20524 ( .A1(n18575), .A2(n18631), .ZN(n18908) );
  AOI22_X1 U20525 ( .A1(n18638), .A2(n18908), .B1(n18637), .B2(n18919), .ZN(
        n18579) );
  NOR2_X1 U20526 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18576), .ZN(
        n18633) );
  AOI22_X1 U20527 ( .A1(n18894), .A2(n18586), .B1(n18577), .B2(n18633), .ZN(
        n18909) );
  NAND2_X1 U20528 ( .A1(n21144), .A2(n18586), .ZN(n18857) );
  INV_X1 U20529 ( .A(n18857), .ZN(n18925) );
  AOI22_X1 U20530 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18909), .B1(
        n18642), .B2(n18925), .ZN(n18578) );
  OAI211_X1 U20531 ( .C1(n18645), .C2(n18902), .A(n18579), .B(n18578), .ZN(
        P3_U2979) );
  NOR2_X1 U20532 ( .A1(n20083), .A2(n18580), .ZN(n18913) );
  AOI22_X1 U20533 ( .A1(n18638), .A2(n18913), .B1(n18637), .B2(n18925), .ZN(
        n18585) );
  NAND2_X1 U20534 ( .A1(n18596), .A2(n18617), .ZN(n18923) );
  INV_X1 U20535 ( .A(n18923), .ZN(n18930) );
  NOR2_X1 U20536 ( .A1(n18925), .A2(n18930), .ZN(n18591) );
  INV_X1 U20537 ( .A(n18591), .ZN(n18583) );
  NOR2_X1 U20538 ( .A1(n18765), .A2(n18581), .ZN(n18640) );
  AOI22_X1 U20539 ( .A1(n18894), .A2(n18583), .B1(n18640), .B2(n18582), .ZN(
        n18915) );
  AOI22_X1 U20540 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18915), .B1(
        n18642), .B2(n18930), .ZN(n18584) );
  OAI211_X1 U20541 ( .C1(n18852), .C2(n18645), .A(n18585), .B(n18584), .ZN(
        P3_U2971) );
  INV_X1 U20542 ( .A(n18586), .ZN(n18587) );
  NOR2_X1 U20543 ( .A1(n20083), .A2(n18587), .ZN(n18918) );
  AOI22_X1 U20544 ( .A1(n18638), .A2(n18918), .B1(n18637), .B2(n18930), .ZN(
        n18589) );
  NAND2_X1 U20545 ( .A1(n18596), .A2(n18624), .ZN(n18920) );
  NOR2_X2 U20546 ( .A1(n21149), .A2(n18595), .ZN(n18936) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18920), .B1(
        n18642), .B2(n18936), .ZN(n18588) );
  OAI211_X1 U20548 ( .C1(n18645), .C2(n18912), .A(n18589), .B(n18588), .ZN(
        P3_U2963) );
  NOR2_X1 U20549 ( .A1(n20083), .A2(n18591), .ZN(n18924) );
  AOI22_X1 U20550 ( .A1(n18638), .A2(n18924), .B1(n18637), .B2(n18936), .ZN(
        n18594) );
  NOR2_X1 U20551 ( .A1(n18590), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18604) );
  NAND2_X1 U20552 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18604), .ZN(
        n18934) );
  INV_X1 U20553 ( .A(n18934), .ZN(n18942) );
  NOR2_X1 U20554 ( .A1(n18936), .A2(n18942), .ZN(n18599) );
  OAI21_X1 U20555 ( .B1(n18599), .B2(n18609), .A(n18591), .ZN(n18592) );
  OAI211_X1 U20556 ( .C1(n18925), .C2(n21176), .A(n18895), .B(n18592), .ZN(
        n18926) );
  AOI22_X1 U20557 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18926), .B1(
        n18642), .B2(n18942), .ZN(n18593) );
  OAI211_X1 U20558 ( .C1(n18645), .C2(n18857), .A(n18594), .B(n18593), .ZN(
        P3_U2955) );
  NAND2_X1 U20559 ( .A1(n21144), .A2(n18604), .ZN(n18940) );
  INV_X1 U20560 ( .A(n18940), .ZN(n18947) );
  NOR2_X1 U20561 ( .A1(n18595), .A2(n18631), .ZN(n18929) );
  AOI22_X1 U20562 ( .A1(n18642), .A2(n18947), .B1(n18638), .B2(n18929), .ZN(
        n18598) );
  AOI22_X1 U20563 ( .A1(n18894), .A2(n18604), .B1(n18596), .B2(n18633), .ZN(
        n18931) );
  AOI22_X1 U20564 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18931), .B1(
        n18637), .B2(n18942), .ZN(n18597) );
  OAI211_X1 U20565 ( .C1(n18645), .C2(n18923), .A(n18598), .B(n18597), .ZN(
        P3_U2947) );
  INV_X1 U20566 ( .A(n18936), .ZN(n18862) );
  NOR2_X1 U20567 ( .A1(n20083), .A2(n18599), .ZN(n18935) );
  AOI22_X1 U20568 ( .A1(n18638), .A2(n18935), .B1(n18637), .B2(n18947), .ZN(
        n18603) );
  NAND2_X1 U20569 ( .A1(n18614), .A2(n18617), .ZN(n18826) );
  INV_X1 U20570 ( .A(n18826), .ZN(n18953) );
  NOR2_X1 U20571 ( .A1(n18947), .A2(n18953), .ZN(n18608) );
  NAND2_X1 U20572 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n20081), .ZN(n18600) );
  OAI21_X1 U20573 ( .B1(n18608), .B2(n18600), .A(n18599), .ZN(n18601) );
  OAI211_X1 U20574 ( .C1(n18936), .C2(n21176), .A(n18895), .B(n18601), .ZN(
        n18937) );
  AOI22_X1 U20575 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18937), .B1(
        n18642), .B2(n18953), .ZN(n18602) );
  OAI211_X1 U20576 ( .C1(n18645), .C2(n18862), .A(n18603), .B(n18602), .ZN(
        P3_U2939) );
  INV_X1 U20577 ( .A(n18604), .ZN(n18605) );
  NOR2_X1 U20578 ( .A1(n20083), .A2(n18605), .ZN(n18941) );
  AOI22_X1 U20579 ( .A1(n18638), .A2(n18941), .B1(n18637), .B2(n18953), .ZN(
        n18607) );
  NAND2_X1 U20580 ( .A1(n18614), .A2(n18624), .ZN(n18943) );
  NOR2_X2 U20581 ( .A1(n21149), .A2(n18613), .ZN(n18959) );
  AOI22_X1 U20582 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18943), .B1(
        n18642), .B2(n18959), .ZN(n18606) );
  OAI211_X1 U20583 ( .C1(n18645), .C2(n18934), .A(n18607), .B(n18606), .ZN(
        P3_U2931) );
  NOR2_X1 U20584 ( .A1(n20083), .A2(n18608), .ZN(n18946) );
  AOI22_X1 U20585 ( .A1(n18638), .A2(n18946), .B1(n18637), .B2(n18959), .ZN(
        n18612) );
  INV_X1 U20586 ( .A(n18959), .ZN(n18951) );
  NAND2_X1 U20587 ( .A1(n21153), .A2(n21156), .ZN(n18630) );
  NOR2_X1 U20588 ( .A1(n21147), .A2(n18630), .ZN(n18622) );
  NAND2_X1 U20589 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18622), .ZN(
        n18871) );
  NAND2_X1 U20590 ( .A1(n18951), .A2(n18871), .ZN(n18619) );
  INV_X1 U20591 ( .A(n18619), .ZN(n18618) );
  OAI22_X1 U20592 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18826), .B1(n18618), 
        .B2(n18609), .ZN(n18610) );
  OAI21_X1 U20593 ( .B1(n18947), .B2(n18610), .A(n18895), .ZN(n18948) );
  INV_X1 U20594 ( .A(n18871), .ZN(n18964) );
  AOI22_X1 U20595 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18948), .B1(
        n18642), .B2(n18964), .ZN(n18611) );
  OAI211_X1 U20596 ( .C1(n18645), .C2(n18940), .A(n18612), .B(n18611), .ZN(
        P3_U2923) );
  NAND2_X1 U20597 ( .A1(n21144), .A2(n18622), .ZN(n18957) );
  INV_X1 U20598 ( .A(n18957), .ZN(n18970) );
  NOR2_X1 U20599 ( .A1(n18613), .A2(n18631), .ZN(n18952) );
  AOI22_X1 U20600 ( .A1(n18642), .A2(n18970), .B1(n18638), .B2(n18952), .ZN(
        n18616) );
  AOI22_X1 U20601 ( .A1(n18894), .A2(n18622), .B1(n18614), .B2(n18633), .ZN(
        n18954) );
  AOI22_X1 U20602 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18954), .B1(
        n18637), .B2(n18964), .ZN(n18615) );
  OAI211_X1 U20603 ( .C1(n18645), .C2(n18826), .A(n18616), .B(n18615), .ZN(
        P3_U2915) );
  INV_X1 U20604 ( .A(n18630), .ZN(n18632) );
  NAND2_X1 U20605 ( .A1(n18617), .A2(n18632), .ZN(n18968) );
  INV_X1 U20606 ( .A(n18968), .ZN(n18978) );
  NOR2_X1 U20607 ( .A1(n20083), .A2(n18618), .ZN(n18958) );
  AOI22_X1 U20608 ( .A1(n18642), .A2(n18978), .B1(n18638), .B2(n18958), .ZN(
        n18621) );
  NAND2_X1 U20609 ( .A1(n18957), .A2(n18968), .ZN(n18627) );
  AOI22_X1 U20610 ( .A1(n18894), .A2(n18627), .B1(n18640), .B2(n18619), .ZN(
        n18960) );
  AOI22_X1 U20611 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18960), .B1(
        n18637), .B2(n18970), .ZN(n18620) );
  OAI211_X1 U20612 ( .C1(n18645), .C2(n18951), .A(n18621), .B(n18620), .ZN(
        P3_U2907) );
  NOR2_X2 U20613 ( .A1(n21149), .A2(n18630), .ZN(n18988) );
  INV_X1 U20614 ( .A(n18622), .ZN(n18623) );
  NOR2_X1 U20615 ( .A1(n20083), .A2(n18623), .ZN(n18963) );
  AOI22_X1 U20616 ( .A1(n18642), .A2(n18988), .B1(n18638), .B2(n18963), .ZN(
        n18626) );
  NAND2_X1 U20617 ( .A1(n18624), .A2(n18632), .ZN(n18965) );
  AOI22_X1 U20618 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18965), .B1(
        n18637), .B2(n18978), .ZN(n18625) );
  OAI211_X1 U20619 ( .C1(n18645), .C2(n18871), .A(n18626), .B(n18625), .ZN(
        P3_U2899) );
  INV_X1 U20620 ( .A(n18799), .ZN(n18977) );
  AND2_X1 U20621 ( .A1(n21167), .A2(n18627), .ZN(n18969) );
  AOI22_X1 U20622 ( .A1(n18642), .A2(n18977), .B1(n18638), .B2(n18969), .ZN(
        n18629) );
  INV_X1 U20623 ( .A(n18988), .ZN(n18974) );
  NAND2_X1 U20624 ( .A1(n18799), .A2(n18974), .ZN(n18639) );
  AOI22_X1 U20625 ( .A1(n18894), .A2(n18639), .B1(n18640), .B2(n18627), .ZN(
        n18971) );
  AOI22_X1 U20626 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18971), .B1(
        n18637), .B2(n18988), .ZN(n18628) );
  OAI211_X1 U20627 ( .C1(n18645), .C2(n18957), .A(n18629), .B(n18628), .ZN(
        P3_U2891) );
  NOR2_X1 U20628 ( .A1(n18631), .A2(n18630), .ZN(n18975) );
  AOI22_X1 U20629 ( .A1(n18642), .A2(n18904), .B1(n18638), .B2(n18975), .ZN(
        n18636) );
  AOI22_X1 U20630 ( .A1(n18894), .A2(n18634), .B1(n18633), .B2(n18632), .ZN(
        n18979) );
  AOI22_X1 U20631 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18979), .B1(
        n18977), .B2(n18637), .ZN(n18635) );
  OAI211_X1 U20632 ( .C1(n18645), .C2(n18968), .A(n18636), .B(n18635), .ZN(
        P3_U2883) );
  AND2_X1 U20633 ( .A1(n21167), .A2(n18639), .ZN(n18984) );
  AOI22_X1 U20634 ( .A1(n18638), .A2(n18984), .B1(n18637), .B2(n18904), .ZN(
        n18644) );
  NAND2_X1 U20635 ( .A1(n18902), .A2(n18993), .ZN(n18641) );
  AOI22_X1 U20636 ( .A1(n18894), .A2(n18641), .B1(n18640), .B2(n18639), .ZN(
        n18989) );
  AOI22_X1 U20637 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18989), .B1(
        n18642), .B2(n18986), .ZN(n18643) );
  OAI211_X1 U20638 ( .C1(n18645), .C2(n18974), .A(n18644), .B(n18643), .ZN(
        P3_U2875) );
  OAI22_X1 U20639 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n18890), .ZN(n18646) );
  INV_X1 U20640 ( .A(n18646), .ZN(U257) );
  NAND2_X1 U20641 ( .A1(n18685), .A2(n20586), .ZN(n18683) );
  INV_X1 U20642 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20605) );
  NOR2_X2 U20643 ( .A1(n20605), .A2(n18765), .ZN(n18678) );
  NOR2_X2 U20644 ( .A1(n20599), .A2(n18893), .ZN(n18679) );
  AOI22_X1 U20645 ( .A1(n18896), .A2(n18678), .B1(n18986), .B2(n18679), .ZN(
        n18649) );
  NOR2_X2 U20646 ( .A1(n18647), .A2(n18893), .ZN(n18680) );
  AOI22_X1 U20647 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18899), .B1(
        n18914), .B2(n18680), .ZN(n18648) );
  OAI211_X1 U20648 ( .C1(n18799), .C2(n18683), .A(n18649), .B(n18648), .ZN(
        P3_U2994) );
  AOI22_X1 U20649 ( .A1(n18919), .A2(n18680), .B1(n18903), .B2(n18678), .ZN(
        n18651) );
  AOI22_X1 U20650 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18905), .B1(
        n18914), .B2(n18679), .ZN(n18650) );
  OAI211_X1 U20651 ( .C1(n18993), .C2(n18683), .A(n18651), .B(n18650), .ZN(
        P3_U2986) );
  AOI22_X1 U20652 ( .A1(n18919), .A2(n18679), .B1(n18908), .B2(n18678), .ZN(
        n18653) );
  AOI22_X1 U20653 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18909), .B1(
        n18925), .B2(n18680), .ZN(n18652) );
  OAI211_X1 U20654 ( .C1(n18902), .C2(n18683), .A(n18653), .B(n18652), .ZN(
        P3_U2978) );
  AOI22_X1 U20655 ( .A1(n18930), .A2(n18680), .B1(n18913), .B2(n18678), .ZN(
        n18655) );
  AOI22_X1 U20656 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18915), .B1(
        n18925), .B2(n18679), .ZN(n18654) );
  OAI211_X1 U20657 ( .C1(n18852), .C2(n18683), .A(n18655), .B(n18654), .ZN(
        P3_U2970) );
  AOI22_X1 U20658 ( .A1(n18930), .A2(n18679), .B1(n18918), .B2(n18678), .ZN(
        n18657) );
  AOI22_X1 U20659 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18920), .B1(
        n18936), .B2(n18680), .ZN(n18656) );
  OAI211_X1 U20660 ( .C1(n18912), .C2(n18683), .A(n18657), .B(n18656), .ZN(
        P3_U2962) );
  AOI22_X1 U20661 ( .A1(n18936), .A2(n18679), .B1(n18924), .B2(n18678), .ZN(
        n18659) );
  AOI22_X1 U20662 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18926), .B1(
        n18942), .B2(n18680), .ZN(n18658) );
  OAI211_X1 U20663 ( .C1(n18857), .C2(n18683), .A(n18659), .B(n18658), .ZN(
        P3_U2954) );
  AOI22_X1 U20664 ( .A1(n18929), .A2(n18678), .B1(n18947), .B2(n18680), .ZN(
        n18661) );
  AOI22_X1 U20665 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18931), .B1(
        n18942), .B2(n18679), .ZN(n18660) );
  OAI211_X1 U20666 ( .C1(n18923), .C2(n18683), .A(n18661), .B(n18660), .ZN(
        P3_U2946) );
  AOI22_X1 U20667 ( .A1(n18947), .A2(n18679), .B1(n18935), .B2(n18678), .ZN(
        n18663) );
  AOI22_X1 U20668 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18937), .B1(
        n18953), .B2(n18680), .ZN(n18662) );
  OAI211_X1 U20669 ( .C1(n18862), .C2(n18683), .A(n18663), .B(n18662), .ZN(
        P3_U2938) );
  AOI22_X1 U20670 ( .A1(n18953), .A2(n18679), .B1(n18941), .B2(n18678), .ZN(
        n18665) );
  AOI22_X1 U20671 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18943), .B1(
        n18959), .B2(n18680), .ZN(n18664) );
  OAI211_X1 U20672 ( .C1(n18934), .C2(n18683), .A(n18665), .B(n18664), .ZN(
        P3_U2930) );
  AOI22_X1 U20673 ( .A1(n18964), .A2(n18680), .B1(n18946), .B2(n18678), .ZN(
        n18667) );
  AOI22_X1 U20674 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18948), .B1(
        n18959), .B2(n18679), .ZN(n18666) );
  OAI211_X1 U20675 ( .C1(n18940), .C2(n18683), .A(n18667), .B(n18666), .ZN(
        P3_U2922) );
  AOI22_X1 U20676 ( .A1(n18970), .A2(n18680), .B1(n18952), .B2(n18678), .ZN(
        n18669) );
  AOI22_X1 U20677 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18954), .B1(
        n18964), .B2(n18679), .ZN(n18668) );
  OAI211_X1 U20678 ( .C1(n18826), .C2(n18683), .A(n18669), .B(n18668), .ZN(
        P3_U2914) );
  AOI22_X1 U20679 ( .A1(n18970), .A2(n18679), .B1(n18958), .B2(n18678), .ZN(
        n18671) );
  AOI22_X1 U20680 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18960), .B1(
        n18978), .B2(n18680), .ZN(n18670) );
  OAI211_X1 U20681 ( .C1(n18951), .C2(n18683), .A(n18671), .B(n18670), .ZN(
        P3_U2906) );
  AOI22_X1 U20682 ( .A1(n18988), .A2(n18680), .B1(n18963), .B2(n18678), .ZN(
        n18673) );
  AOI22_X1 U20683 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18965), .B1(
        n18978), .B2(n18679), .ZN(n18672) );
  OAI211_X1 U20684 ( .C1(n18871), .C2(n18683), .A(n18673), .B(n18672), .ZN(
        P3_U2898) );
  AOI22_X1 U20685 ( .A1(n18988), .A2(n18679), .B1(n18969), .B2(n18678), .ZN(
        n18675) );
  AOI22_X1 U20686 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18971), .B1(
        n18977), .B2(n18680), .ZN(n18674) );
  OAI211_X1 U20687 ( .C1(n18957), .C2(n18683), .A(n18675), .B(n18674), .ZN(
        P3_U2890) );
  AOI22_X1 U20688 ( .A1(n18904), .A2(n18680), .B1(n18975), .B2(n18678), .ZN(
        n18677) );
  AOI22_X1 U20689 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18979), .B1(
        n18977), .B2(n18679), .ZN(n18676) );
  OAI211_X1 U20690 ( .C1(n18968), .C2(n18683), .A(n18677), .B(n18676), .ZN(
        P3_U2882) );
  AOI22_X1 U20691 ( .A1(n18904), .A2(n18679), .B1(n18984), .B2(n18678), .ZN(
        n18682) );
  AOI22_X1 U20692 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18989), .B1(
        n18986), .B2(n18680), .ZN(n18681) );
  OAI211_X1 U20693 ( .C1(n18974), .C2(n18683), .A(n18682), .B(n18681), .ZN(
        P3_U2874) );
  OAI22_X1 U20694 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n18890), .ZN(n18684) );
  INV_X1 U20695 ( .A(n18684), .ZN(U256) );
  NAND2_X1 U20696 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18894), .ZN(n18707) );
  INV_X1 U20697 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20564) );
  NOR2_X2 U20698 ( .A1(n20564), .A2(n18765), .ZN(n18718) );
  NAND2_X1 U20699 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18894), .ZN(n18723) );
  INV_X1 U20700 ( .A(n18723), .ZN(n18704) );
  AOI22_X1 U20701 ( .A1(n18896), .A2(n18718), .B1(n18986), .B2(n18704), .ZN(
        n18687) );
  INV_X1 U20702 ( .A(n18685), .ZN(n18897) );
  NOR2_X2 U20703 ( .A1(n20585), .A2(n18897), .ZN(n18720) );
  AOI22_X1 U20704 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18720), .ZN(n18686) );
  OAI211_X1 U20705 ( .C1(n18852), .C2(n18707), .A(n18687), .B(n18686), .ZN(
        P3_U2993) );
  INV_X1 U20706 ( .A(n18707), .ZN(n18719) );
  AOI22_X1 U20707 ( .A1(n18919), .A2(n18719), .B1(n18903), .B2(n18718), .ZN(
        n18689) );
  AOI22_X1 U20708 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18720), .ZN(n18688) );
  OAI211_X1 U20709 ( .C1(n18852), .C2(n18723), .A(n18689), .B(n18688), .ZN(
        P3_U2985) );
  AOI22_X1 U20710 ( .A1(n18925), .A2(n18719), .B1(n18908), .B2(n18718), .ZN(
        n18691) );
  AOI22_X1 U20711 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18720), .ZN(n18690) );
  OAI211_X1 U20712 ( .C1(n18912), .C2(n18723), .A(n18691), .B(n18690), .ZN(
        P3_U2977) );
  AOI22_X1 U20713 ( .A1(n18930), .A2(n18719), .B1(n18913), .B2(n18718), .ZN(
        n18693) );
  AOI22_X1 U20714 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18720), .ZN(n18692) );
  OAI211_X1 U20715 ( .C1(n18857), .C2(n18723), .A(n18693), .B(n18692), .ZN(
        P3_U2969) );
  AOI22_X1 U20716 ( .A1(n18936), .A2(n18719), .B1(n18918), .B2(n18718), .ZN(
        n18695) );
  AOI22_X1 U20717 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18720), .ZN(n18694) );
  OAI211_X1 U20718 ( .C1(n18923), .C2(n18723), .A(n18695), .B(n18694), .ZN(
        P3_U2961) );
  AOI22_X1 U20719 ( .A1(n18936), .A2(n18704), .B1(n18924), .B2(n18718), .ZN(
        n18697) );
  AOI22_X1 U20720 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18720), .ZN(n18696) );
  OAI211_X1 U20721 ( .C1(n18934), .C2(n18707), .A(n18697), .B(n18696), .ZN(
        P3_U2953) );
  AOI22_X1 U20722 ( .A1(n18929), .A2(n18718), .B1(n18947), .B2(n18719), .ZN(
        n18699) );
  AOI22_X1 U20723 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18720), .ZN(n18698) );
  OAI211_X1 U20724 ( .C1(n18934), .C2(n18723), .A(n18699), .B(n18698), .ZN(
        P3_U2945) );
  AOI22_X1 U20725 ( .A1(n18947), .A2(n18704), .B1(n18935), .B2(n18718), .ZN(
        n18701) );
  AOI22_X1 U20726 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18720), .ZN(n18700) );
  OAI211_X1 U20727 ( .C1(n18826), .C2(n18707), .A(n18701), .B(n18700), .ZN(
        P3_U2937) );
  AOI22_X1 U20728 ( .A1(n18959), .A2(n18719), .B1(n18941), .B2(n18718), .ZN(
        n18703) );
  AOI22_X1 U20729 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18720), .ZN(n18702) );
  OAI211_X1 U20730 ( .C1(n18826), .C2(n18723), .A(n18703), .B(n18702), .ZN(
        P3_U2929) );
  AOI22_X1 U20731 ( .A1(n18959), .A2(n18704), .B1(n18946), .B2(n18718), .ZN(
        n18706) );
  AOI22_X1 U20732 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18720), .ZN(n18705) );
  OAI211_X1 U20733 ( .C1(n18871), .C2(n18707), .A(n18706), .B(n18705), .ZN(
        P3_U2921) );
  AOI22_X1 U20734 ( .A1(n18970), .A2(n18719), .B1(n18952), .B2(n18718), .ZN(
        n18709) );
  AOI22_X1 U20735 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18720), .ZN(n18708) );
  OAI211_X1 U20736 ( .C1(n18871), .C2(n18723), .A(n18709), .B(n18708), .ZN(
        P3_U2913) );
  AOI22_X1 U20737 ( .A1(n18978), .A2(n18719), .B1(n18958), .B2(n18718), .ZN(
        n18711) );
  AOI22_X1 U20738 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18720), .ZN(n18710) );
  OAI211_X1 U20739 ( .C1(n18957), .C2(n18723), .A(n18711), .B(n18710), .ZN(
        P3_U2905) );
  AOI22_X1 U20740 ( .A1(n18988), .A2(n18719), .B1(n18963), .B2(n18718), .ZN(
        n18713) );
  AOI22_X1 U20741 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18720), .ZN(n18712) );
  OAI211_X1 U20742 ( .C1(n18968), .C2(n18723), .A(n18713), .B(n18712), .ZN(
        P3_U2897) );
  AOI22_X1 U20743 ( .A1(n18977), .A2(n18719), .B1(n18969), .B2(n18718), .ZN(
        n18715) );
  AOI22_X1 U20744 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18720), .ZN(n18714) );
  OAI211_X1 U20745 ( .C1(n18974), .C2(n18723), .A(n18715), .B(n18714), .ZN(
        P3_U2889) );
  AOI22_X1 U20746 ( .A1(n18904), .A2(n18719), .B1(n18975), .B2(n18718), .ZN(
        n18717) );
  AOI22_X1 U20747 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18720), .ZN(n18716) );
  OAI211_X1 U20748 ( .C1(n18799), .C2(n18723), .A(n18717), .B(n18716), .ZN(
        P3_U2881) );
  AOI22_X1 U20749 ( .A1(n18986), .A2(n18719), .B1(n18984), .B2(n18718), .ZN(
        n18722) );
  AOI22_X1 U20750 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18720), .ZN(n18721) );
  OAI211_X1 U20751 ( .C1(n18993), .C2(n18723), .A(n18722), .B(n18721), .ZN(
        P3_U2873) );
  OAI22_X1 U20752 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n18890), .ZN(n18724) );
  INV_X1 U20753 ( .A(n18724), .ZN(U255) );
  INV_X1 U20754 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19352) );
  NOR2_X1 U20755 ( .A1(n19352), .A2(n18893), .ZN(n18754) );
  INV_X1 U20756 ( .A(n18754), .ZN(n18763) );
  NAND2_X1 U20757 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18894), .ZN(n18757) );
  INV_X1 U20758 ( .A(n18757), .ZN(n18759) );
  INV_X1 U20759 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20569) );
  NOR2_X2 U20760 ( .A1(n20569), .A2(n18765), .ZN(n18758) );
  AOI22_X1 U20761 ( .A1(n18914), .A2(n18759), .B1(n18896), .B2(n18758), .ZN(
        n18727) );
  NOR2_X2 U20762 ( .A1(n18725), .A2(n18897), .ZN(n18760) );
  AOI22_X1 U20763 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18760), .ZN(n18726) );
  OAI211_X1 U20764 ( .C1(n18902), .C2(n18763), .A(n18727), .B(n18726), .ZN(
        P3_U2992) );
  AOI22_X1 U20765 ( .A1(n18919), .A2(n18759), .B1(n18903), .B2(n18758), .ZN(
        n18729) );
  AOI22_X1 U20766 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18760), .ZN(n18728) );
  OAI211_X1 U20767 ( .C1(n18852), .C2(n18763), .A(n18729), .B(n18728), .ZN(
        P3_U2984) );
  AOI22_X1 U20768 ( .A1(n18919), .A2(n18754), .B1(n18908), .B2(n18758), .ZN(
        n18731) );
  AOI22_X1 U20769 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18760), .ZN(n18730) );
  OAI211_X1 U20770 ( .C1(n18857), .C2(n18757), .A(n18731), .B(n18730), .ZN(
        P3_U2976) );
  AOI22_X1 U20771 ( .A1(n18925), .A2(n18754), .B1(n18913), .B2(n18758), .ZN(
        n18733) );
  AOI22_X1 U20772 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18760), .ZN(n18732) );
  OAI211_X1 U20773 ( .C1(n18923), .C2(n18757), .A(n18733), .B(n18732), .ZN(
        P3_U2968) );
  AOI22_X1 U20774 ( .A1(n18936), .A2(n18759), .B1(n18918), .B2(n18758), .ZN(
        n18735) );
  AOI22_X1 U20775 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18760), .ZN(n18734) );
  OAI211_X1 U20776 ( .C1(n18923), .C2(n18763), .A(n18735), .B(n18734), .ZN(
        P3_U2960) );
  AOI22_X1 U20777 ( .A1(n18942), .A2(n18759), .B1(n18924), .B2(n18758), .ZN(
        n18737) );
  AOI22_X1 U20778 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18760), .ZN(n18736) );
  OAI211_X1 U20779 ( .C1(n18862), .C2(n18763), .A(n18737), .B(n18736), .ZN(
        P3_U2952) );
  AOI22_X1 U20780 ( .A1(n18929), .A2(n18758), .B1(n18947), .B2(n18759), .ZN(
        n18739) );
  AOI22_X1 U20781 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18760), .ZN(n18738) );
  OAI211_X1 U20782 ( .C1(n18934), .C2(n18763), .A(n18739), .B(n18738), .ZN(
        P3_U2944) );
  AOI22_X1 U20783 ( .A1(n18953), .A2(n18759), .B1(n18935), .B2(n18758), .ZN(
        n18741) );
  AOI22_X1 U20784 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18760), .ZN(n18740) );
  OAI211_X1 U20785 ( .C1(n18940), .C2(n18763), .A(n18741), .B(n18740), .ZN(
        P3_U2936) );
  AOI22_X1 U20786 ( .A1(n18959), .A2(n18759), .B1(n18941), .B2(n18758), .ZN(
        n18743) );
  AOI22_X1 U20787 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18760), .ZN(n18742) );
  OAI211_X1 U20788 ( .C1(n18826), .C2(n18763), .A(n18743), .B(n18742), .ZN(
        P3_U2928) );
  AOI22_X1 U20789 ( .A1(n18959), .A2(n18754), .B1(n18946), .B2(n18758), .ZN(
        n18745) );
  AOI22_X1 U20790 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18760), .ZN(n18744) );
  OAI211_X1 U20791 ( .C1(n18871), .C2(n18757), .A(n18745), .B(n18744), .ZN(
        P3_U2920) );
  AOI22_X1 U20792 ( .A1(n18970), .A2(n18759), .B1(n18952), .B2(n18758), .ZN(
        n18747) );
  AOI22_X1 U20793 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18760), .ZN(n18746) );
  OAI211_X1 U20794 ( .C1(n18871), .C2(n18763), .A(n18747), .B(n18746), .ZN(
        P3_U2912) );
  AOI22_X1 U20795 ( .A1(n18970), .A2(n18754), .B1(n18958), .B2(n18758), .ZN(
        n18749) );
  AOI22_X1 U20796 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18760), .ZN(n18748) );
  OAI211_X1 U20797 ( .C1(n18968), .C2(n18757), .A(n18749), .B(n18748), .ZN(
        P3_U2904) );
  AOI22_X1 U20798 ( .A1(n18988), .A2(n18759), .B1(n18963), .B2(n18758), .ZN(
        n18751) );
  AOI22_X1 U20799 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18760), .ZN(n18750) );
  OAI211_X1 U20800 ( .C1(n18968), .C2(n18763), .A(n18751), .B(n18750), .ZN(
        P3_U2896) );
  AOI22_X1 U20801 ( .A1(n18977), .A2(n18759), .B1(n18969), .B2(n18758), .ZN(
        n18753) );
  AOI22_X1 U20802 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18760), .ZN(n18752) );
  OAI211_X1 U20803 ( .C1(n18974), .C2(n18763), .A(n18753), .B(n18752), .ZN(
        P3_U2888) );
  AOI22_X1 U20804 ( .A1(n18977), .A2(n18754), .B1(n18975), .B2(n18758), .ZN(
        n18756) );
  AOI22_X1 U20805 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18760), .ZN(n18755) );
  OAI211_X1 U20806 ( .C1(n18993), .C2(n18757), .A(n18756), .B(n18755), .ZN(
        P3_U2880) );
  AOI22_X1 U20807 ( .A1(n18986), .A2(n18759), .B1(n18984), .B2(n18758), .ZN(
        n18762) );
  AOI22_X1 U20808 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18760), .ZN(n18761) );
  OAI211_X1 U20809 ( .C1(n18993), .C2(n18763), .A(n18762), .B(n18761), .ZN(
        P3_U2872) );
  OAI22_X1 U20810 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n18890), .ZN(n18764) );
  INV_X1 U20811 ( .A(n18764), .ZN(U254) );
  NAND2_X1 U20812 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18894), .ZN(n18794) );
  INV_X1 U20813 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20574) );
  NOR2_X2 U20814 ( .A1(n18765), .A2(n20574), .ZN(n18800) );
  NAND2_X1 U20815 ( .A1(n18894), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18805) );
  INV_X1 U20816 ( .A(n18805), .ZN(n18791) );
  AOI22_X1 U20817 ( .A1(n18896), .A2(n18800), .B1(n18986), .B2(n18791), .ZN(
        n18768) );
  NOR2_X2 U20818 ( .A1(n18766), .A2(n18897), .ZN(n18802) );
  AOI22_X1 U20819 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18802), .ZN(n18767) );
  OAI211_X1 U20820 ( .C1(n18852), .C2(n18794), .A(n18768), .B(n18767), .ZN(
        P3_U2991) );
  AOI22_X1 U20821 ( .A1(n18914), .A2(n18791), .B1(n18903), .B2(n18800), .ZN(
        n18770) );
  AOI22_X1 U20822 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18802), .ZN(n18769) );
  OAI211_X1 U20823 ( .C1(n18912), .C2(n18794), .A(n18770), .B(n18769), .ZN(
        P3_U2983) );
  AOI22_X1 U20824 ( .A1(n18919), .A2(n18791), .B1(n18908), .B2(n18800), .ZN(
        n18772) );
  AOI22_X1 U20825 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18802), .ZN(n18771) );
  OAI211_X1 U20826 ( .C1(n18857), .C2(n18794), .A(n18772), .B(n18771), .ZN(
        P3_U2975) );
  AOI22_X1 U20827 ( .A1(n18925), .A2(n18791), .B1(n18913), .B2(n18800), .ZN(
        n18774) );
  AOI22_X1 U20828 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18802), .ZN(n18773) );
  OAI211_X1 U20829 ( .C1(n18923), .C2(n18794), .A(n18774), .B(n18773), .ZN(
        P3_U2967) );
  AOI22_X1 U20830 ( .A1(n18930), .A2(n18791), .B1(n18918), .B2(n18800), .ZN(
        n18776) );
  AOI22_X1 U20831 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18802), .ZN(n18775) );
  OAI211_X1 U20832 ( .C1(n18862), .C2(n18794), .A(n18776), .B(n18775), .ZN(
        P3_U2959) );
  AOI22_X1 U20833 ( .A1(n18936), .A2(n18791), .B1(n18924), .B2(n18800), .ZN(
        n18778) );
  AOI22_X1 U20834 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18802), .ZN(n18777) );
  OAI211_X1 U20835 ( .C1(n18934), .C2(n18794), .A(n18778), .B(n18777), .ZN(
        P3_U2951) );
  AOI22_X1 U20836 ( .A1(n18942), .A2(n18791), .B1(n18929), .B2(n18800), .ZN(
        n18780) );
  AOI22_X1 U20837 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18802), .ZN(n18779) );
  OAI211_X1 U20838 ( .C1(n18940), .C2(n18794), .A(n18780), .B(n18779), .ZN(
        P3_U2943) );
  INV_X1 U20839 ( .A(n18794), .ZN(n18801) );
  AOI22_X1 U20840 ( .A1(n18953), .A2(n18801), .B1(n18935), .B2(n18800), .ZN(
        n18782) );
  AOI22_X1 U20841 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18802), .ZN(n18781) );
  OAI211_X1 U20842 ( .C1(n18940), .C2(n18805), .A(n18782), .B(n18781), .ZN(
        P3_U2935) );
  AOI22_X1 U20843 ( .A1(n18959), .A2(n18801), .B1(n18941), .B2(n18800), .ZN(
        n18784) );
  AOI22_X1 U20844 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18802), .ZN(n18783) );
  OAI211_X1 U20845 ( .C1(n18826), .C2(n18805), .A(n18784), .B(n18783), .ZN(
        P3_U2927) );
  AOI22_X1 U20846 ( .A1(n18964), .A2(n18801), .B1(n18946), .B2(n18800), .ZN(
        n18786) );
  AOI22_X1 U20847 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18802), .ZN(n18785) );
  OAI211_X1 U20848 ( .C1(n18951), .C2(n18805), .A(n18786), .B(n18785), .ZN(
        P3_U2919) );
  AOI22_X1 U20849 ( .A1(n18970), .A2(n18801), .B1(n18952), .B2(n18800), .ZN(
        n18788) );
  AOI22_X1 U20850 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18802), .ZN(n18787) );
  OAI211_X1 U20851 ( .C1(n18871), .C2(n18805), .A(n18788), .B(n18787), .ZN(
        P3_U2911) );
  AOI22_X1 U20852 ( .A1(n18970), .A2(n18791), .B1(n18958), .B2(n18800), .ZN(
        n18790) );
  AOI22_X1 U20853 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18802), .ZN(n18789) );
  OAI211_X1 U20854 ( .C1(n18968), .C2(n18794), .A(n18790), .B(n18789), .ZN(
        P3_U2903) );
  AOI22_X1 U20855 ( .A1(n18978), .A2(n18791), .B1(n18963), .B2(n18800), .ZN(
        n18793) );
  AOI22_X1 U20856 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18802), .ZN(n18792) );
  OAI211_X1 U20857 ( .C1(n18974), .C2(n18794), .A(n18793), .B(n18792), .ZN(
        P3_U2895) );
  AOI22_X1 U20858 ( .A1(n18977), .A2(n18801), .B1(n18969), .B2(n18800), .ZN(
        n18796) );
  AOI22_X1 U20859 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18802), .ZN(n18795) );
  OAI211_X1 U20860 ( .C1(n18974), .C2(n18805), .A(n18796), .B(n18795), .ZN(
        P3_U2887) );
  AOI22_X1 U20861 ( .A1(n18904), .A2(n18801), .B1(n18975), .B2(n18800), .ZN(
        n18798) );
  AOI22_X1 U20862 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18802), .ZN(n18797) );
  OAI211_X1 U20863 ( .C1(n18799), .C2(n18805), .A(n18798), .B(n18797), .ZN(
        P3_U2879) );
  AOI22_X1 U20864 ( .A1(n18986), .A2(n18801), .B1(n18984), .B2(n18800), .ZN(
        n18804) );
  AOI22_X1 U20865 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18802), .ZN(n18803) );
  OAI211_X1 U20866 ( .C1(n18993), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P3_U2871) );
  OAI22_X1 U20867 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n18890), .ZN(n18806) );
  INV_X1 U20868 ( .A(n18806), .ZN(U253) );
  INV_X1 U20869 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19478) );
  NOR2_X1 U20870 ( .A1(n19478), .A2(n18893), .ZN(n18842) );
  INV_X1 U20871 ( .A(n18842), .ZN(n18840) );
  AND2_X1 U20872 ( .A1(n18895), .A2(BUF2_REG_2__SCAN_IN), .ZN(n18841) );
  NAND2_X1 U20873 ( .A1(n18894), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18846) );
  INV_X1 U20874 ( .A(n18846), .ZN(n18837) );
  AOI22_X1 U20875 ( .A1(n18896), .A2(n18841), .B1(n18986), .B2(n18837), .ZN(
        n18809) );
  NOR2_X2 U20876 ( .A1(n18807), .A2(n18897), .ZN(n18843) );
  AOI22_X1 U20877 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18843), .ZN(n18808) );
  OAI211_X1 U20878 ( .C1(n18852), .C2(n18840), .A(n18809), .B(n18808), .ZN(
        P3_U2990) );
  AOI22_X1 U20879 ( .A1(n18914), .A2(n18837), .B1(n18903), .B2(n18841), .ZN(
        n18811) );
  AOI22_X1 U20880 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18843), .ZN(n18810) );
  OAI211_X1 U20881 ( .C1(n18912), .C2(n18840), .A(n18811), .B(n18810), .ZN(
        P3_U2982) );
  AOI22_X1 U20882 ( .A1(n18919), .A2(n18837), .B1(n18908), .B2(n18841), .ZN(
        n18813) );
  AOI22_X1 U20883 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18843), .ZN(n18812) );
  OAI211_X1 U20884 ( .C1(n18857), .C2(n18840), .A(n18813), .B(n18812), .ZN(
        P3_U2974) );
  AOI22_X1 U20885 ( .A1(n18925), .A2(n18837), .B1(n18913), .B2(n18841), .ZN(
        n18815) );
  AOI22_X1 U20886 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18843), .ZN(n18814) );
  OAI211_X1 U20887 ( .C1(n18923), .C2(n18840), .A(n18815), .B(n18814), .ZN(
        P3_U2966) );
  AOI22_X1 U20888 ( .A1(n18930), .A2(n18837), .B1(n18918), .B2(n18841), .ZN(
        n18817) );
  AOI22_X1 U20889 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18843), .ZN(n18816) );
  OAI211_X1 U20890 ( .C1(n18862), .C2(n18840), .A(n18817), .B(n18816), .ZN(
        P3_U2958) );
  AOI22_X1 U20891 ( .A1(n18942), .A2(n18842), .B1(n18924), .B2(n18841), .ZN(
        n18819) );
  AOI22_X1 U20892 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18843), .ZN(n18818) );
  OAI211_X1 U20893 ( .C1(n18862), .C2(n18846), .A(n18819), .B(n18818), .ZN(
        P3_U2950) );
  AOI22_X1 U20894 ( .A1(n18929), .A2(n18841), .B1(n18947), .B2(n18842), .ZN(
        n18821) );
  AOI22_X1 U20895 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18843), .ZN(n18820) );
  OAI211_X1 U20896 ( .C1(n18934), .C2(n18846), .A(n18821), .B(n18820), .ZN(
        P3_U2942) );
  AOI22_X1 U20897 ( .A1(n18953), .A2(n18842), .B1(n18935), .B2(n18841), .ZN(
        n18823) );
  AOI22_X1 U20898 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18843), .ZN(n18822) );
  OAI211_X1 U20899 ( .C1(n18940), .C2(n18846), .A(n18823), .B(n18822), .ZN(
        P3_U2934) );
  AOI22_X1 U20900 ( .A1(n18959), .A2(n18842), .B1(n18941), .B2(n18841), .ZN(
        n18825) );
  AOI22_X1 U20901 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18843), .ZN(n18824) );
  OAI211_X1 U20902 ( .C1(n18826), .C2(n18846), .A(n18825), .B(n18824), .ZN(
        P3_U2926) );
  AOI22_X1 U20903 ( .A1(n18959), .A2(n18837), .B1(n18946), .B2(n18841), .ZN(
        n18828) );
  AOI22_X1 U20904 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18843), .ZN(n18827) );
  OAI211_X1 U20905 ( .C1(n18871), .C2(n18840), .A(n18828), .B(n18827), .ZN(
        P3_U2918) );
  AOI22_X1 U20906 ( .A1(n18964), .A2(n18837), .B1(n18952), .B2(n18841), .ZN(
        n18830) );
  AOI22_X1 U20907 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18843), .ZN(n18829) );
  OAI211_X1 U20908 ( .C1(n18957), .C2(n18840), .A(n18830), .B(n18829), .ZN(
        P3_U2910) );
  AOI22_X1 U20909 ( .A1(n18978), .A2(n18842), .B1(n18958), .B2(n18841), .ZN(
        n18832) );
  AOI22_X1 U20910 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18843), .ZN(n18831) );
  OAI211_X1 U20911 ( .C1(n18957), .C2(n18846), .A(n18832), .B(n18831), .ZN(
        P3_U2902) );
  AOI22_X1 U20912 ( .A1(n18988), .A2(n18842), .B1(n18963), .B2(n18841), .ZN(
        n18834) );
  AOI22_X1 U20913 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18843), .ZN(n18833) );
  OAI211_X1 U20914 ( .C1(n18968), .C2(n18846), .A(n18834), .B(n18833), .ZN(
        P3_U2894) );
  AOI22_X1 U20915 ( .A1(n18977), .A2(n18842), .B1(n18969), .B2(n18841), .ZN(
        n18836) );
  AOI22_X1 U20916 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18843), .ZN(n18835) );
  OAI211_X1 U20917 ( .C1(n18974), .C2(n18846), .A(n18836), .B(n18835), .ZN(
        P3_U2886) );
  AOI22_X1 U20918 ( .A1(n18977), .A2(n18837), .B1(n18975), .B2(n18841), .ZN(
        n18839) );
  AOI22_X1 U20919 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18843), .ZN(n18838) );
  OAI211_X1 U20920 ( .C1(n18993), .C2(n18840), .A(n18839), .B(n18838), .ZN(
        P3_U2878) );
  AOI22_X1 U20921 ( .A1(n18986), .A2(n18842), .B1(n18984), .B2(n18841), .ZN(
        n18845) );
  AOI22_X1 U20922 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18843), .ZN(n18844) );
  OAI211_X1 U20923 ( .C1(n18993), .C2(n18846), .A(n18845), .B(n18844), .ZN(
        P3_U2870) );
  OAI22_X1 U20924 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18890), .ZN(n18847) );
  INV_X1 U20925 ( .A(n18847), .ZN(U252) );
  INV_X1 U20926 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n20630) );
  NOR2_X1 U20927 ( .A1(n20630), .A2(n18893), .ZN(n18885) );
  INV_X1 U20928 ( .A(n18885), .ZN(n18883) );
  AND2_X1 U20929 ( .A1(n18895), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18884) );
  NAND2_X1 U20930 ( .A1(n18894), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18889) );
  INV_X1 U20931 ( .A(n18889), .ZN(n18880) );
  AOI22_X1 U20932 ( .A1(n18896), .A2(n18884), .B1(n18986), .B2(n18880), .ZN(
        n18849) );
  NOR2_X2 U20933 ( .A1(n20084), .A2(n18897), .ZN(n18886) );
  AOI22_X1 U20934 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18886), .ZN(n18848) );
  OAI211_X1 U20935 ( .C1(n18852), .C2(n18883), .A(n18849), .B(n18848), .ZN(
        P3_U2989) );
  AOI22_X1 U20936 ( .A1(n18919), .A2(n18885), .B1(n18903), .B2(n18884), .ZN(
        n18851) );
  AOI22_X1 U20937 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18886), .ZN(n18850) );
  OAI211_X1 U20938 ( .C1(n18852), .C2(n18889), .A(n18851), .B(n18850), .ZN(
        P3_U2981) );
  AOI22_X1 U20939 ( .A1(n18919), .A2(n18880), .B1(n18908), .B2(n18884), .ZN(
        n18854) );
  AOI22_X1 U20940 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18886), .ZN(n18853) );
  OAI211_X1 U20941 ( .C1(n18857), .C2(n18883), .A(n18854), .B(n18853), .ZN(
        P3_U2973) );
  AOI22_X1 U20942 ( .A1(n18930), .A2(n18885), .B1(n18913), .B2(n18884), .ZN(
        n18856) );
  AOI22_X1 U20943 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18886), .ZN(n18855) );
  OAI211_X1 U20944 ( .C1(n18857), .C2(n18889), .A(n18856), .B(n18855), .ZN(
        P3_U2965) );
  AOI22_X1 U20945 ( .A1(n18930), .A2(n18880), .B1(n18918), .B2(n18884), .ZN(
        n18859) );
  AOI22_X1 U20946 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18886), .ZN(n18858) );
  OAI211_X1 U20947 ( .C1(n18862), .C2(n18883), .A(n18859), .B(n18858), .ZN(
        P3_U2957) );
  AOI22_X1 U20948 ( .A1(n18942), .A2(n18885), .B1(n18924), .B2(n18884), .ZN(
        n18861) );
  AOI22_X1 U20949 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18886), .ZN(n18860) );
  OAI211_X1 U20950 ( .C1(n18862), .C2(n18889), .A(n18861), .B(n18860), .ZN(
        P3_U2949) );
  AOI22_X1 U20951 ( .A1(n18942), .A2(n18880), .B1(n18929), .B2(n18884), .ZN(
        n18864) );
  AOI22_X1 U20952 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18886), .ZN(n18863) );
  OAI211_X1 U20953 ( .C1(n18940), .C2(n18883), .A(n18864), .B(n18863), .ZN(
        P3_U2941) );
  AOI22_X1 U20954 ( .A1(n18953), .A2(n18885), .B1(n18935), .B2(n18884), .ZN(
        n18866) );
  AOI22_X1 U20955 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18886), .ZN(n18865) );
  OAI211_X1 U20956 ( .C1(n18940), .C2(n18889), .A(n18866), .B(n18865), .ZN(
        P3_U2933) );
  AOI22_X1 U20957 ( .A1(n18953), .A2(n18880), .B1(n18941), .B2(n18884), .ZN(
        n18868) );
  AOI22_X1 U20958 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18886), .ZN(n18867) );
  OAI211_X1 U20959 ( .C1(n18951), .C2(n18883), .A(n18868), .B(n18867), .ZN(
        P3_U2925) );
  AOI22_X1 U20960 ( .A1(n18959), .A2(n18880), .B1(n18946), .B2(n18884), .ZN(
        n18870) );
  AOI22_X1 U20961 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18886), .ZN(n18869) );
  OAI211_X1 U20962 ( .C1(n18871), .C2(n18883), .A(n18870), .B(n18869), .ZN(
        P3_U2917) );
  AOI22_X1 U20963 ( .A1(n18964), .A2(n18880), .B1(n18952), .B2(n18884), .ZN(
        n18873) );
  AOI22_X1 U20964 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18886), .ZN(n18872) );
  OAI211_X1 U20965 ( .C1(n18957), .C2(n18883), .A(n18873), .B(n18872), .ZN(
        P3_U2909) );
  AOI22_X1 U20966 ( .A1(n18978), .A2(n18885), .B1(n18958), .B2(n18884), .ZN(
        n18875) );
  AOI22_X1 U20967 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18886), .ZN(n18874) );
  OAI211_X1 U20968 ( .C1(n18957), .C2(n18889), .A(n18875), .B(n18874), .ZN(
        P3_U2901) );
  AOI22_X1 U20969 ( .A1(n18988), .A2(n18885), .B1(n18963), .B2(n18884), .ZN(
        n18877) );
  AOI22_X1 U20970 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18886), .ZN(n18876) );
  OAI211_X1 U20971 ( .C1(n18968), .C2(n18889), .A(n18877), .B(n18876), .ZN(
        P3_U2893) );
  AOI22_X1 U20972 ( .A1(n18977), .A2(n18885), .B1(n18969), .B2(n18884), .ZN(
        n18879) );
  AOI22_X1 U20973 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18886), .ZN(n18878) );
  OAI211_X1 U20974 ( .C1(n18974), .C2(n18889), .A(n18879), .B(n18878), .ZN(
        P3_U2885) );
  AOI22_X1 U20975 ( .A1(n18977), .A2(n18880), .B1(n18975), .B2(n18884), .ZN(
        n18882) );
  AOI22_X1 U20976 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18886), .ZN(n18881) );
  OAI211_X1 U20977 ( .C1(n18993), .C2(n18883), .A(n18882), .B(n18881), .ZN(
        P3_U2877) );
  AOI22_X1 U20978 ( .A1(n18986), .A2(n18885), .B1(n18984), .B2(n18884), .ZN(
        n18888) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18886), .ZN(n18887) );
  OAI211_X1 U20980 ( .C1(n18993), .C2(n18889), .A(n18888), .B(n18887), .ZN(
        P3_U2869) );
  OAI22_X1 U20981 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n18890), .ZN(n18891) );
  INV_X1 U20982 ( .A(n18891), .ZN(U251) );
  NOR2_X1 U20983 ( .A1(n18893), .A2(n18892), .ZN(n18976) );
  INV_X1 U20984 ( .A(n18976), .ZN(n18992) );
  NAND2_X1 U20985 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18894), .ZN(n18982) );
  INV_X1 U20986 ( .A(n18982), .ZN(n18985) );
  AND2_X1 U20987 ( .A1(n18895), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18983) );
  AOI22_X1 U20988 ( .A1(n18914), .A2(n18985), .B1(n18896), .B2(n18983), .ZN(
        n18901) );
  NOR2_X2 U20989 ( .A1(n18898), .A2(n18897), .ZN(n18987) );
  AOI22_X1 U20990 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18899), .B1(
        n18977), .B2(n18987), .ZN(n18900) );
  OAI211_X1 U20991 ( .C1(n18902), .C2(n18992), .A(n18901), .B(n18900), .ZN(
        P3_U2988) );
  AOI22_X1 U20992 ( .A1(n18914), .A2(n18976), .B1(n18903), .B2(n18983), .ZN(
        n18907) );
  AOI22_X1 U20993 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n18987), .ZN(n18906) );
  OAI211_X1 U20994 ( .C1(n18912), .C2(n18982), .A(n18907), .B(n18906), .ZN(
        P3_U2980) );
  AOI22_X1 U20995 ( .A1(n18925), .A2(n18985), .B1(n18908), .B2(n18983), .ZN(
        n18911) );
  AOI22_X1 U20996 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18909), .B1(
        n18986), .B2(n18987), .ZN(n18910) );
  OAI211_X1 U20997 ( .C1(n18912), .C2(n18992), .A(n18911), .B(n18910), .ZN(
        P3_U2972) );
  AOI22_X1 U20998 ( .A1(n18925), .A2(n18976), .B1(n18913), .B2(n18983), .ZN(
        n18917) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18987), .ZN(n18916) );
  OAI211_X1 U21000 ( .C1(n18923), .C2(n18982), .A(n18917), .B(n18916), .ZN(
        P3_U2964) );
  AOI22_X1 U21001 ( .A1(n18936), .A2(n18985), .B1(n18918), .B2(n18983), .ZN(
        n18922) );
  AOI22_X1 U21002 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18920), .B1(
        n18919), .B2(n18987), .ZN(n18921) );
  OAI211_X1 U21003 ( .C1(n18923), .C2(n18992), .A(n18922), .B(n18921), .ZN(
        P3_U2956) );
  AOI22_X1 U21004 ( .A1(n18936), .A2(n18976), .B1(n18924), .B2(n18983), .ZN(
        n18928) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18926), .B1(
        n18925), .B2(n18987), .ZN(n18927) );
  OAI211_X1 U21006 ( .C1(n18934), .C2(n18982), .A(n18928), .B(n18927), .ZN(
        P3_U2948) );
  AOI22_X1 U21007 ( .A1(n18929), .A2(n18983), .B1(n18947), .B2(n18985), .ZN(
        n18933) );
  AOI22_X1 U21008 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18931), .B1(
        n18930), .B2(n18987), .ZN(n18932) );
  OAI211_X1 U21009 ( .C1(n18934), .C2(n18992), .A(n18933), .B(n18932), .ZN(
        P3_U2940) );
  AOI22_X1 U21010 ( .A1(n18953), .A2(n18985), .B1(n18935), .B2(n18983), .ZN(
        n18939) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18937), .B1(
        n18936), .B2(n18987), .ZN(n18938) );
  OAI211_X1 U21012 ( .C1(n18940), .C2(n18992), .A(n18939), .B(n18938), .ZN(
        P3_U2932) );
  AOI22_X1 U21013 ( .A1(n18953), .A2(n18976), .B1(n18941), .B2(n18983), .ZN(
        n18945) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18943), .B1(
        n18942), .B2(n18987), .ZN(n18944) );
  OAI211_X1 U21015 ( .C1(n18951), .C2(n18982), .A(n18945), .B(n18944), .ZN(
        P3_U2924) );
  AOI22_X1 U21016 ( .A1(n18964), .A2(n18985), .B1(n18946), .B2(n18983), .ZN(
        n18950) );
  AOI22_X1 U21017 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18987), .ZN(n18949) );
  OAI211_X1 U21018 ( .C1(n18951), .C2(n18992), .A(n18950), .B(n18949), .ZN(
        P3_U2916) );
  AOI22_X1 U21019 ( .A1(n18964), .A2(n18976), .B1(n18952), .B2(n18983), .ZN(
        n18956) );
  AOI22_X1 U21020 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18954), .B1(
        n18953), .B2(n18987), .ZN(n18955) );
  OAI211_X1 U21021 ( .C1(n18957), .C2(n18982), .A(n18956), .B(n18955), .ZN(
        P3_U2908) );
  AOI22_X1 U21022 ( .A1(n18970), .A2(n18976), .B1(n18958), .B2(n18983), .ZN(
        n18962) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18960), .B1(
        n18959), .B2(n18987), .ZN(n18961) );
  OAI211_X1 U21024 ( .C1(n18968), .C2(n18982), .A(n18962), .B(n18961), .ZN(
        P3_U2900) );
  AOI22_X1 U21025 ( .A1(n18988), .A2(n18985), .B1(n18963), .B2(n18983), .ZN(
        n18967) );
  AOI22_X1 U21026 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18965), .B1(
        n18964), .B2(n18987), .ZN(n18966) );
  OAI211_X1 U21027 ( .C1(n18968), .C2(n18992), .A(n18967), .B(n18966), .ZN(
        P3_U2892) );
  AOI22_X1 U21028 ( .A1(n18977), .A2(n18985), .B1(n18969), .B2(n18983), .ZN(
        n18973) );
  AOI22_X1 U21029 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18971), .B1(
        n18970), .B2(n18987), .ZN(n18972) );
  OAI211_X1 U21030 ( .C1(n18974), .C2(n18992), .A(n18973), .B(n18972), .ZN(
        P3_U2884) );
  AOI22_X1 U21031 ( .A1(n18977), .A2(n18976), .B1(n18975), .B2(n18983), .ZN(
        n18981) );
  AOI22_X1 U21032 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18987), .ZN(n18980) );
  OAI211_X1 U21033 ( .C1(n18993), .C2(n18982), .A(n18981), .B(n18980), .ZN(
        P3_U2876) );
  AOI22_X1 U21034 ( .A1(n18986), .A2(n18985), .B1(n18984), .B2(n18983), .ZN(
        n18991) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18989), .B1(
        n18988), .B2(n18987), .ZN(n18990) );
  OAI211_X1 U21036 ( .C1(n18993), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P3_U2868) );
  AOI22_X1 U21037 ( .A1(n18995), .A2(BUF2_REG_31__SCAN_IN), .B1(n19345), .B2(
        n18994), .ZN(n18998) );
  AOI22_X1 U21038 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19465), .B1(n18996), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18997) );
  NAND2_X1 U21039 ( .A1(n18998), .A2(n18997), .ZN(P2_U2888) );
  AOI22_X1 U21040 ( .A1(n19589), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19586), .ZN(n19000) );
  OAI21_X1 U21041 ( .B1(n19002), .B2(n19591), .A(n19000), .ZN(P2_U2966) );
  AOI22_X1 U21042 ( .A1(n19589), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19586), .ZN(n19001) );
  OAI21_X1 U21043 ( .B1(n19002), .B2(n19591), .A(n19001), .ZN(P2_U2981) );
  AOI22_X1 U21044 ( .A1(n19589), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19586), .ZN(n19003) );
  OAI21_X1 U21045 ( .B1(n19005), .B2(n19591), .A(n19003), .ZN(P2_U2965) );
  AOI22_X1 U21046 ( .A1(n19589), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n19004) );
  OAI21_X1 U21047 ( .B1(n19005), .B2(n19591), .A(n19004), .ZN(P2_U2980) );
  AOI22_X1 U21048 ( .A1(n19589), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19586), .ZN(n19006) );
  OAI21_X1 U21049 ( .B1(n19008), .B2(n19591), .A(n19006), .ZN(P2_U2964) );
  AOI22_X1 U21050 ( .A1(n19589), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n19007) );
  OAI21_X1 U21051 ( .B1(n19008), .B2(n19591), .A(n19007), .ZN(P2_U2979) );
  AOI22_X1 U21052 ( .A1(n19589), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19586), .ZN(n19009) );
  OAI21_X1 U21053 ( .B1(n19011), .B2(n19591), .A(n19009), .ZN(P2_U2963) );
  AOI22_X1 U21054 ( .A1(n19589), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19586), .ZN(n19010) );
  OAI21_X1 U21055 ( .B1(n19011), .B2(n19591), .A(n19010), .ZN(P2_U2978) );
  AOI22_X1 U21056 ( .A1(n19589), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n19586), .ZN(n19012) );
  OAI21_X1 U21057 ( .B1(n19014), .B2(n19591), .A(n19012), .ZN(P2_U2962) );
  AOI22_X1 U21058 ( .A1(n19589), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U21059 ( .B1(n19014), .B2(n19591), .A(n19013), .ZN(P2_U2977) );
  AOI22_X1 U21060 ( .A1(n19589), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n19015) );
  OAI21_X1 U21061 ( .B1(n19017), .B2(n19591), .A(n19015), .ZN(P2_U2961) );
  AOI22_X1 U21062 ( .A1(n19589), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19586), .ZN(n19016) );
  OAI21_X1 U21063 ( .B1(n19017), .B2(n19591), .A(n19016), .ZN(P2_U2976) );
  AOI22_X1 U21064 ( .A1(n19587), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19586), .ZN(n19018) );
  OAI21_X1 U21065 ( .B1(n19020), .B2(n19591), .A(n19018), .ZN(P2_U2960) );
  AOI22_X1 U21066 ( .A1(n19587), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n19019) );
  OAI21_X1 U21067 ( .B1(n19020), .B2(n19591), .A(n19019), .ZN(P2_U2975) );
  AOI22_X1 U21068 ( .A1(n19587), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n19586), .ZN(n19021) );
  OAI21_X1 U21069 ( .B1(n19029), .B2(n19591), .A(n19021), .ZN(P2_U2959) );
  AOI22_X1 U21070 ( .A1(n19589), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U21071 ( .B1(n19029), .B2(n19591), .A(n19022), .ZN(P2_U2974) );
  NAND3_X1 U21072 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19037) );
  OAI21_X1 U21073 ( .B1(n19051), .B2(n19107), .A(n19037), .ZN(n19026) );
  NAND2_X1 U21074 ( .A1(n19027), .A2(n19216), .ZN(n19024) );
  INV_X1 U21075 ( .A(n19218), .ZN(n19598) );
  OAI21_X1 U21076 ( .B1(n19200), .B2(n19598), .A(n19219), .ZN(n19023) );
  NAND2_X1 U21077 ( .A1(n19024), .A2(n19023), .ZN(n19025) );
  AND2_X1 U21078 ( .A1(n19026), .A2(n19025), .ZN(n19231) );
  OAI21_X1 U21079 ( .B1(n19027), .B2(n19598), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19028) );
  OAI21_X1 U21080 ( .B1(n19037), .B2(n13500), .A(n19028), .ZN(n19599) );
  NOR2_X2 U21081 ( .A1(n19029), .A2(n19594), .ZN(n19224) );
  NAND2_X1 U21082 ( .A1(n11858), .A2(n19596), .ZN(n19211) );
  AOI22_X1 U21083 ( .A1(n19599), .A2(n19224), .B1(n19598), .B2(n19197), .ZN(
        n19032) );
  AOI22_X1 U21084 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19592), .ZN(n19212) );
  INV_X1 U21085 ( .A(n19212), .ZN(n19189) );
  INV_X1 U21086 ( .A(n19719), .ZN(n19030) );
  AOI22_X1 U21087 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19592), .ZN(n19227) );
  INV_X1 U21088 ( .A(n19227), .ZN(n19207) );
  AOI22_X1 U21089 ( .A1(n19603), .A2(n19189), .B1(n19030), .B2(n19207), .ZN(
        n19031) );
  OAI211_X1 U21090 ( .C1(n19231), .C2(n19033), .A(n19032), .B(n19031), .ZN(
        P2_U3175) );
  INV_X1 U21091 ( .A(n19224), .ZN(n19178) );
  NAND2_X1 U21092 ( .A1(n19608), .A2(n19620), .ZN(n19036) );
  NOR2_X1 U21093 ( .A1(n19037), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19357) );
  INV_X1 U21094 ( .A(n19357), .ZN(n19607) );
  AOI21_X1 U21095 ( .B1(n19038), .B2(n19607), .A(n19164), .ZN(n19040) );
  NOR2_X1 U21096 ( .A1(n19146), .A2(n19050), .ZN(n19615) );
  OR3_X1 U21097 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19357), .A3(n19615), 
        .ZN(n19039) );
  OAI22_X1 U21098 ( .A1(n19608), .A2(n19227), .B1(n19607), .B2(n19211), .ZN(
        n19041) );
  INV_X1 U21099 ( .A(n19041), .ZN(n19047) );
  INV_X1 U21100 ( .A(n19615), .ZN(n19043) );
  AOI21_X1 U21101 ( .B1(n12190), .B2(n19216), .A(n19215), .ZN(n19042) );
  AOI21_X1 U21102 ( .B1(n19044), .B2(n19043), .A(n19042), .ZN(n19045) );
  AOI22_X1 U21103 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19189), .ZN(n19046) );
  OAI211_X1 U21104 ( .C1(n19178), .C2(n19614), .A(n19047), .B(n19046), .ZN(
        P2_U3167) );
  OAI21_X1 U21105 ( .B1(n12084), .B2(n19615), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19048) );
  OAI21_X1 U21106 ( .B1(n19050), .B2(n13500), .A(n19048), .ZN(n19616) );
  AOI22_X1 U21107 ( .A1(n19616), .A2(n19224), .B1(n19197), .B2(n19615), .ZN(
        n19057) );
  NAND2_X1 U21108 ( .A1(n19049), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19130) );
  OAI21_X1 U21109 ( .B1(n19051), .B2(n19130), .A(n19050), .ZN(n19055) );
  AOI21_X1 U21110 ( .B1(n19615), .B2(n19219), .A(n19215), .ZN(n19052) );
  OAI21_X1 U21111 ( .B1(n19053), .B2(n19202), .A(n19052), .ZN(n19054) );
  NAND2_X1 U21112 ( .A1(n19055), .A2(n19054), .ZN(n19617) );
  AOI22_X1 U21113 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19189), .ZN(n19056) );
  OAI211_X1 U21114 ( .C1(n19227), .C2(n19620), .A(n19057), .B(n19056), .ZN(
        P2_U3159) );
  AOI22_X1 U21115 ( .A1(n19622), .A2(n19224), .B1(n19621), .B2(n19197), .ZN(
        n19059) );
  AOI22_X1 U21116 ( .A1(n19630), .A2(n19189), .B1(n19623), .B2(n19207), .ZN(
        n19058) );
  OAI211_X1 U21117 ( .C1(n19626), .C2(n19060), .A(n19059), .B(n19058), .ZN(
        P2_U3151) );
  NAND3_X1 U21118 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19160), .ZN(n19069) );
  NOR2_X1 U21119 ( .A1(n19146), .A2(n19069), .ZN(n19627) );
  OAI21_X1 U21120 ( .B1(n19061), .B2(n19627), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19062) );
  OAI21_X1 U21121 ( .B1(n19069), .B2(n13500), .A(n19062), .ZN(n19628) );
  AOI22_X1 U21122 ( .A1(n19628), .A2(n19224), .B1(n19197), .B2(n19627), .ZN(
        n19068) );
  OAI21_X1 U21123 ( .B1(n19198), .B2(n19169), .A(n19069), .ZN(n19066) );
  OAI21_X1 U21124 ( .B1(n19200), .B2(n19627), .A(n19219), .ZN(n19063) );
  OAI21_X1 U21125 ( .B1(n19064), .B2(n19202), .A(n19063), .ZN(n19065) );
  NAND2_X1 U21126 ( .A1(n19066), .A2(n19065), .ZN(n19629) );
  AOI22_X1 U21127 ( .A1(n19630), .A2(n19207), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n19629), .ZN(n19067) );
  OAI211_X1 U21128 ( .C1(n19212), .C2(n19639), .A(n19068), .B(n19067), .ZN(
        P2_U3143) );
  NOR2_X1 U21129 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19069), .ZN(
        n19633) );
  INV_X1 U21130 ( .A(n19633), .ZN(n19542) );
  OAI22_X1 U21131 ( .A1(n19641), .A2(n19212), .B1(n19211), .B2(n19542), .ZN(
        n19070) );
  INV_X1 U21132 ( .A(n19070), .ZN(n19079) );
  INV_X1 U21133 ( .A(n19639), .ZN(n19366) );
  OAI21_X1 U21134 ( .B1(n19634), .B2(n19366), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19071) );
  NAND2_X1 U21135 ( .A1(n19071), .A2(n19200), .ZN(n19077) );
  NOR3_X1 U21136 ( .A1(n19159), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19093) );
  NAND2_X1 U21137 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19093), .ZN(
        n19640) );
  INV_X1 U21138 ( .A(n19640), .ZN(n19369) );
  NOR2_X1 U21139 ( .A1(n19633), .A2(n19369), .ZN(n19076) );
  INV_X1 U21140 ( .A(n19076), .ZN(n19074) );
  AOI21_X1 U21141 ( .B1(n12031), .B2(n19183), .A(n19633), .ZN(n19072) );
  NOR2_X1 U21142 ( .A1(n19072), .A2(n19594), .ZN(n19073) );
  OAI21_X1 U21143 ( .B1(n12031), .B2(n19633), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19075) );
  AOI22_X1 U21144 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19636), .B1(
        n19224), .B2(n19635), .ZN(n19078) );
  OAI211_X1 U21145 ( .C1(n19227), .C2(n19639), .A(n19079), .B(n19078), .ZN(
        P2_U3135) );
  INV_X1 U21146 ( .A(n19093), .ZN(n19087) );
  NOR2_X1 U21147 ( .A1(n13500), .A2(n19087), .ZN(n19082) );
  AOI21_X1 U21148 ( .B1(n19080), .B2(n19640), .A(n19164), .ZN(n19081) );
  NOR2_X1 U21149 ( .A1(n19082), .A2(n19081), .ZN(n19647) );
  OAI22_X1 U21150 ( .A1(n19649), .A2(n19212), .B1(n19211), .B2(n19640), .ZN(
        n19084) );
  INV_X1 U21151 ( .A(n19084), .ZN(n19092) );
  NOR2_X1 U21152 ( .A1(n19080), .A2(n19202), .ZN(n19090) );
  AOI21_X1 U21153 ( .B1(n19640), .B2(n13500), .A(n19594), .ZN(n19089) );
  NOR2_X1 U21154 ( .A1(n19085), .A2(n19130), .ZN(n19199) );
  NAND2_X1 U21155 ( .A1(n19170), .A2(n19199), .ZN(n19086) );
  NAND2_X1 U21156 ( .A1(n19087), .A2(n19086), .ZN(n19088) );
  OAI21_X1 U21157 ( .B1(n19090), .B2(n19089), .A(n19088), .ZN(n19644) );
  AOI22_X1 U21158 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19644), .B1(
        n19634), .B2(n19207), .ZN(n19091) );
  OAI211_X1 U21159 ( .C1(n19647), .C2(n19178), .A(n19092), .B(n19091), .ZN(
        P2_U3127) );
  AND2_X1 U21160 ( .A1(n19146), .A2(n19093), .ZN(n19099) );
  INV_X1 U21161 ( .A(n19099), .ZN(n19648) );
  OAI22_X1 U21162 ( .A1(n19661), .A2(n19212), .B1(n19211), .B2(n19648), .ZN(
        n19094) );
  INV_X1 U21163 ( .A(n19094), .ZN(n19103) );
  AOI21_X1 U21164 ( .B1(n19649), .B2(n19661), .A(n21639), .ZN(n19095) );
  NOR2_X1 U21165 ( .A1(n19095), .A2(n13500), .ZN(n19098) );
  NAND2_X1 U21166 ( .A1(n19159), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19128) );
  INV_X1 U21167 ( .A(n19128), .ZN(n19147) );
  AND2_X1 U21168 ( .A1(n19163), .A2(n19147), .ZN(n19655) );
  INV_X1 U21169 ( .A(n19655), .ZN(n19108) );
  OAI21_X1 U21170 ( .B1(n12087), .B2(n19164), .A(n19183), .ZN(n19096) );
  AOI21_X1 U21171 ( .B1(n19098), .B2(n19108), .A(n19096), .ZN(n19097) );
  OAI21_X1 U21172 ( .B1(n19099), .B2(n19097), .A(n19219), .ZN(n19652) );
  OAI21_X1 U21173 ( .B1(n19655), .B2(n19099), .A(n19098), .ZN(n19101) );
  OAI21_X1 U21174 ( .B1(n12087), .B2(n19099), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19100) );
  AOI22_X1 U21175 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19652), .B1(
        n19224), .B2(n19651), .ZN(n19102) );
  OAI211_X1 U21176 ( .C1(n19227), .C2(n19649), .A(n19103), .B(n19102), .ZN(
        P2_U3119) );
  NAND2_X1 U21177 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19147), .ZN(
        n19106) );
  OAI21_X1 U21178 ( .B1(n19104), .B2(n19655), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19105) );
  OAI21_X1 U21179 ( .B1(n19106), .B2(n13500), .A(n19105), .ZN(n19656) );
  AOI22_X1 U21180 ( .A1(n19656), .A2(n19224), .B1(n19655), .B2(n19197), .ZN(
        n19113) );
  OAI22_X1 U21181 ( .A1(n19131), .A2(n19107), .B1(n19128), .B2(n19179), .ZN(
        n19111) );
  OAI211_X1 U21182 ( .C1(n19109), .C2(n19202), .A(n13500), .B(n19108), .ZN(
        n19110) );
  NAND3_X1 U21183 ( .A1(n19111), .A2(n19219), .A3(n19110), .ZN(n19658) );
  AOI22_X1 U21184 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19189), .ZN(n19112) );
  OAI211_X1 U21185 ( .C1(n19227), .C2(n19661), .A(n19113), .B(n19112), .ZN(
        P2_U3111) );
  OR2_X1 U21186 ( .A1(n19114), .A2(n19128), .ZN(n19121) );
  NOR3_X2 U21187 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19179), .A3(
        n19128), .ZN(n19662) );
  OAI21_X1 U21188 ( .B1(n19116), .B2(n19662), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19115) );
  OAI21_X1 U21189 ( .B1(n13500), .B2(n19121), .A(n19115), .ZN(n19663) );
  AOI22_X1 U21190 ( .A1(n19663), .A2(n19224), .B1(n19197), .B2(n19662), .ZN(
        n19127) );
  NAND2_X1 U21191 ( .A1(n19116), .A2(n19216), .ZN(n19120) );
  INV_X1 U21192 ( .A(n19662), .ZN(n19117) );
  NAND2_X1 U21193 ( .A1(n13500), .A2(n19117), .ZN(n19118) );
  NAND2_X1 U21194 ( .A1(n19219), .A2(n19118), .ZN(n19119) );
  NAND2_X1 U21195 ( .A1(n19120), .A2(n19119), .ZN(n19123) );
  OAI221_X1 U21196 ( .B1(n21639), .B2(n19670), .C1(n21639), .C2(n19668), .A(
        n19121), .ZN(n19122) );
  NAND2_X1 U21197 ( .A1(n19123), .A2(n19122), .ZN(n19664) );
  INV_X1 U21198 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n19124) );
  OAI22_X1 U21199 ( .A1(n19670), .A2(n19212), .B1(n19557), .B2(n19124), .ZN(
        n19125) );
  INV_X1 U21200 ( .A(n19125), .ZN(n19126) );
  OAI211_X1 U21201 ( .C1(n19227), .C2(n19668), .A(n19127), .B(n19126), .ZN(
        P2_U3103) );
  NOR2_X1 U21202 ( .A1(n19195), .A2(n19128), .ZN(n19381) );
  INV_X1 U21203 ( .A(n19381), .ZN(n19669) );
  OAI22_X1 U21204 ( .A1(n19677), .A2(n19212), .B1(n19211), .B2(n19669), .ZN(
        n19129) );
  INV_X1 U21205 ( .A(n19129), .ZN(n19141) );
  OAI21_X1 U21206 ( .B1(n19131), .B2(n19130), .A(n19200), .ZN(n19139) );
  NAND2_X1 U21207 ( .A1(n19179), .A2(n19147), .ZN(n19138) );
  INV_X1 U21208 ( .A(n19138), .ZN(n19135) );
  OAI21_X1 U21209 ( .B1(n19200), .B2(n19381), .A(n19219), .ZN(n19132) );
  OAI21_X1 U21210 ( .B1(n19133), .B2(n19202), .A(n19132), .ZN(n19134) );
  OAI21_X1 U21211 ( .B1(n19139), .B2(n19135), .A(n19134), .ZN(n19673) );
  OAI21_X1 U21212 ( .B1(n19136), .B2(n19381), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19137) );
  OAI21_X1 U21213 ( .B1(n19139), .B2(n19138), .A(n19137), .ZN(n19672) );
  AOI22_X1 U21214 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19673), .B1(
        n19224), .B2(n19672), .ZN(n19140) );
  OAI211_X1 U21215 ( .C1(n19227), .C2(n19670), .A(n19141), .B(n19140), .ZN(
        P2_U3095) );
  AOI21_X1 U21216 ( .B1(n19686), .B2(n19677), .A(n21639), .ZN(n19144) );
  NOR2_X1 U21217 ( .A1(n19144), .A2(n13500), .ZN(n19151) );
  NAND2_X1 U21218 ( .A1(n19145), .A2(n19159), .ZN(n19154) );
  NAND3_X1 U21219 ( .A1(n19147), .A2(n19146), .A3(n19179), .ZN(n19676) );
  NOR2_X1 U21220 ( .A1(n19594), .A2(n19676), .ZN(n19148) );
  AOI211_X1 U21221 ( .C1(n19152), .C2(n19216), .A(n19215), .B(n19148), .ZN(
        n19149) );
  INV_X1 U21222 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n19158) );
  OAI22_X1 U21223 ( .A1(n19677), .A2(n19227), .B1(n19211), .B2(n19676), .ZN(
        n19150) );
  INV_X1 U21224 ( .A(n19150), .ZN(n19157) );
  INV_X1 U21225 ( .A(n19151), .ZN(n19155) );
  INV_X1 U21226 ( .A(n19676), .ZN(n19384) );
  OAI21_X1 U21227 ( .B1(n19152), .B2(n19384), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19153) );
  AOI22_X1 U21228 ( .A1(n19224), .A2(n19680), .B1(n19679), .B2(n19189), .ZN(
        n19156) );
  OAI211_X1 U21229 ( .C1(n19684), .C2(n19158), .A(n19157), .B(n19156), .ZN(
        P2_U3087) );
  NAND2_X1 U21230 ( .A1(n19160), .A2(n19159), .ZN(n19194) );
  OR2_X1 U21231 ( .A1(n19179), .A2(n19194), .ZN(n19171) );
  NOR2_X1 U21232 ( .A1(n13500), .A2(n19171), .ZN(n19166) );
  INV_X1 U21233 ( .A(n19194), .ZN(n19162) );
  NAND2_X1 U21234 ( .A1(n19163), .A2(n19162), .ZN(n19685) );
  AOI21_X1 U21235 ( .B1(n19161), .B2(n19685), .A(n19164), .ZN(n19165) );
  OAI22_X1 U21236 ( .A1(n19700), .A2(n19212), .B1(n19685), .B2(n19211), .ZN(
        n19168) );
  INV_X1 U21237 ( .A(n19168), .ZN(n19177) );
  NOR2_X1 U21238 ( .A1(n19170), .A2(n19169), .ZN(n19175) );
  INV_X1 U21239 ( .A(n19171), .ZN(n19174) );
  INV_X1 U21240 ( .A(n19685), .ZN(n19389) );
  OAI21_X1 U21241 ( .B1(n19200), .B2(n19389), .A(n19219), .ZN(n19172) );
  OAI21_X1 U21242 ( .B1(n19161), .B2(n19202), .A(n19172), .ZN(n19173) );
  OAI21_X1 U21243 ( .B1(n19175), .B2(n19174), .A(n19173), .ZN(n19689) );
  AOI22_X1 U21244 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19689), .B1(
        n19679), .B2(n19207), .ZN(n19176) );
  OAI211_X1 U21245 ( .C1(n19693), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        P2_U3079) );
  NOR3_X2 U21246 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19179), .A3(
        n19194), .ZN(n19694) );
  OAI21_X1 U21247 ( .B1(n19184), .B2(n19694), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19181) );
  OR2_X1 U21248 ( .A1(n19180), .A2(n19194), .ZN(n19185) );
  NAND2_X1 U21249 ( .A1(n19181), .A2(n19185), .ZN(n19695) );
  AOI22_X1 U21250 ( .A1(n19695), .A2(n19224), .B1(n19197), .B2(n19694), .ZN(
        n19191) );
  NOR2_X2 U21251 ( .A1(n19193), .A2(n19182), .ZN(n19705) );
  INV_X1 U21252 ( .A(n19705), .ZN(n19578) );
  AOI211_X1 U21253 ( .C1(n19578), .C2(n19700), .A(n13500), .B(n21639), .ZN(
        n19188) );
  AOI21_X1 U21254 ( .B1(n19184), .B2(n19183), .A(n19694), .ZN(n19186) );
  OAI21_X1 U21255 ( .B1(n19186), .B2(n19200), .A(n19185), .ZN(n19187) );
  OAI21_X1 U21256 ( .B1(n19188), .B2(n19187), .A(n19219), .ZN(n19697) );
  AOI22_X1 U21257 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19189), .ZN(n19190) );
  OAI211_X1 U21258 ( .C1(n19227), .C2(n19700), .A(n19191), .B(n19190), .ZN(
        P2_U3071) );
  NOR2_X1 U21259 ( .A1(n19194), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19205) );
  INV_X1 U21260 ( .A(n19205), .ZN(n19210) );
  NOR2_X1 U21261 ( .A1(n19195), .A2(n19194), .ZN(n19701) );
  OAI21_X1 U21262 ( .B1(n12078), .B2(n19701), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19196) );
  OAI21_X1 U21263 ( .B1(n19210), .B2(n13500), .A(n19196), .ZN(n19703) );
  AOI22_X1 U21264 ( .A1(n19703), .A2(n19224), .B1(n19197), .B2(n19701), .ZN(
        n19209) );
  AND2_X1 U21265 ( .A1(n19199), .A2(n19198), .ZN(n19206) );
  OAI21_X1 U21266 ( .B1(n19200), .B2(n19701), .A(n19219), .ZN(n19201) );
  OAI21_X1 U21267 ( .B1(n19203), .B2(n19202), .A(n19201), .ZN(n19204) );
  OAI21_X1 U21268 ( .B1(n19206), .B2(n19205), .A(n19204), .ZN(n19706) );
  AOI22_X1 U21269 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19207), .ZN(n19208) );
  OAI211_X1 U21270 ( .C1(n19212), .C2(n19711), .A(n19209), .B(n19208), .ZN(
        P2_U3063) );
  NOR2_X1 U21271 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19210), .ZN(
        n19270) );
  INV_X1 U21272 ( .A(n19270), .ZN(n19710) );
  OAI22_X1 U21273 ( .A1(n19719), .A2(n19212), .B1(n19211), .B2(n19710), .ZN(
        n19213) );
  INV_X1 U21274 ( .A(n19213), .ZN(n19226) );
  AOI21_X1 U21275 ( .B1(n19719), .B2(n19711), .A(n21639), .ZN(n19214) );
  NOR2_X1 U21276 ( .A1(n19214), .A2(n13500), .ZN(n19221) );
  AOI21_X1 U21277 ( .B1(n10961), .B2(n19216), .A(n19215), .ZN(n19217) );
  AOI21_X1 U21278 ( .B1(n19221), .B2(n19218), .A(n19217), .ZN(n19220) );
  OAI21_X1 U21279 ( .B1(n19598), .B2(n19270), .A(n19221), .ZN(n19223) );
  OAI21_X1 U21280 ( .B1(n10961), .B2(n19270), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19222) );
  AOI22_X1 U21281 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19716), .B1(
        n19224), .B2(n19715), .ZN(n19225) );
  OAI211_X1 U21282 ( .C1(n19227), .C2(n19711), .A(n19226), .B(n19225), .ZN(
        P2_U3055) );
  AOI22_X1 U21283 ( .A1(n19589), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19586), .ZN(n19228) );
  OAI21_X1 U21284 ( .B1(n19230), .B2(n19591), .A(n19228), .ZN(P2_U2958) );
  AOI22_X1 U21285 ( .A1(n19589), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U21286 ( .B1(n19230), .B2(n19591), .A(n19229), .ZN(P2_U2973) );
  INV_X1 U21287 ( .A(n19272), .ZN(n19267) );
  AOI22_X1 U21288 ( .A1(n19599), .A2(n19273), .B1(n19598), .B2(n19271), .ZN(
        n19233) );
  AOI22_X1 U21289 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19264), .ZN(n19232) );
  OAI211_X1 U21290 ( .C1(n19267), .C2(n19719), .A(n19233), .B(n19232), .ZN(
        P2_U3174) );
  INV_X1 U21291 ( .A(n19273), .ZN(n19263) );
  AOI22_X1 U21292 ( .A1(n19603), .A2(n19272), .B1(n19271), .B2(n19357), .ZN(
        n19235) );
  AOI22_X1 U21293 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19264), .ZN(n19234) );
  OAI211_X1 U21294 ( .C1(n19263), .C2(n19614), .A(n19235), .B(n19234), .ZN(
        P2_U3166) );
  AOI22_X1 U21295 ( .A1(n19616), .A2(n19273), .B1(n19271), .B2(n19615), .ZN(
        n19237) );
  AOI22_X1 U21296 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19264), .ZN(n19236) );
  OAI211_X1 U21297 ( .C1(n19267), .C2(n19620), .A(n19237), .B(n19236), .ZN(
        P2_U3158) );
  AOI22_X1 U21298 ( .A1(n19628), .A2(n19273), .B1(n19271), .B2(n19627), .ZN(
        n19239) );
  AOI22_X1 U21299 ( .A1(n19630), .A2(n19272), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n19629), .ZN(n19238) );
  OAI211_X1 U21300 ( .C1(n19276), .C2(n19639), .A(n19239), .B(n19238), .ZN(
        P2_U3142) );
  INV_X1 U21301 ( .A(n19271), .ZN(n19259) );
  OAI22_X1 U21302 ( .A1(n19641), .A2(n19276), .B1(n19259), .B2(n19542), .ZN(
        n19240) );
  INV_X1 U21303 ( .A(n19240), .ZN(n19242) );
  AOI22_X1 U21304 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19636), .B1(
        n19273), .B2(n19635), .ZN(n19241) );
  OAI211_X1 U21305 ( .C1(n19267), .C2(n19639), .A(n19242), .B(n19241), .ZN(
        P2_U3134) );
  AOI22_X1 U21306 ( .A1(n19634), .A2(n19272), .B1(n19271), .B2(n19369), .ZN(
        n19244) );
  INV_X1 U21307 ( .A(n19649), .ZN(n19643) );
  AOI22_X1 U21308 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19264), .ZN(n19243) );
  OAI211_X1 U21309 ( .C1(n19647), .C2(n19263), .A(n19244), .B(n19243), .ZN(
        P2_U3126) );
  OAI22_X1 U21310 ( .A1(n19661), .A2(n19276), .B1(n19259), .B2(n19648), .ZN(
        n19245) );
  INV_X1 U21311 ( .A(n19245), .ZN(n19247) );
  AOI22_X1 U21312 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19652), .B1(
        n19273), .B2(n19651), .ZN(n19246) );
  OAI211_X1 U21313 ( .C1(n19267), .C2(n19649), .A(n19247), .B(n19246), .ZN(
        P2_U3118) );
  AOI22_X1 U21314 ( .A1(n19656), .A2(n19273), .B1(n19271), .B2(n19655), .ZN(
        n19249) );
  AOI22_X1 U21315 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19264), .ZN(n19248) );
  OAI211_X1 U21316 ( .C1(n19267), .C2(n19661), .A(n19249), .B(n19248), .ZN(
        P2_U3110) );
  AOI22_X1 U21317 ( .A1(n19663), .A2(n19273), .B1(n19271), .B2(n19662), .ZN(
        n19253) );
  INV_X1 U21318 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n19250) );
  OAI22_X1 U21319 ( .A1(n19670), .A2(n19276), .B1(n19557), .B2(n19250), .ZN(
        n19251) );
  INV_X1 U21320 ( .A(n19251), .ZN(n19252) );
  OAI211_X1 U21321 ( .C1(n19267), .C2(n19668), .A(n19253), .B(n19252), .ZN(
        P2_U3102) );
  INV_X1 U21322 ( .A(n19670), .ZN(n19665) );
  AOI22_X1 U21323 ( .A1(n19272), .A2(n19665), .B1(n19271), .B2(n19381), .ZN(
        n19255) );
  AOI22_X1 U21324 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19673), .B1(
        n19273), .B2(n19672), .ZN(n19254) );
  OAI211_X1 U21325 ( .C1(n19276), .C2(n19677), .A(n19255), .B(n19254), .ZN(
        P2_U3094) );
  INV_X1 U21326 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n19258) );
  INV_X1 U21327 ( .A(n19677), .ZN(n19385) );
  AOI22_X1 U21328 ( .A1(n19272), .A2(n19385), .B1(n19271), .B2(n19384), .ZN(
        n19257) );
  AOI22_X1 U21329 ( .A1(n19273), .A2(n19680), .B1(n19679), .B2(n19264), .ZN(
        n19256) );
  OAI211_X1 U21330 ( .C1(n19684), .C2(n19258), .A(n19257), .B(n19256), .ZN(
        P2_U3086) );
  OAI22_X1 U21331 ( .A1(n19700), .A2(n19276), .B1(n19259), .B2(n19685), .ZN(
        n19260) );
  INV_X1 U21332 ( .A(n19260), .ZN(n19262) );
  AOI22_X1 U21333 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19689), .B1(
        n19679), .B2(n19272), .ZN(n19261) );
  OAI211_X1 U21334 ( .C1(n19693), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3078) );
  AOI22_X1 U21335 ( .A1(n19695), .A2(n19273), .B1(n19271), .B2(n19694), .ZN(
        n19266) );
  AOI22_X1 U21336 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19264), .ZN(n19265) );
  OAI211_X1 U21337 ( .C1(n19267), .C2(n19700), .A(n19266), .B(n19265), .ZN(
        P2_U3070) );
  AOI22_X1 U21338 ( .A1(n19703), .A2(n19273), .B1(n19271), .B2(n19701), .ZN(
        n19269) );
  AOI22_X1 U21339 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19272), .ZN(n19268) );
  OAI211_X1 U21340 ( .C1(n19276), .C2(n19711), .A(n19269), .B(n19268), .ZN(
        P2_U3062) );
  INV_X1 U21341 ( .A(n19711), .ZN(n19575) );
  AOI22_X1 U21342 ( .A1(n19272), .A2(n19575), .B1(n19271), .B2(n19270), .ZN(
        n19275) );
  AOI22_X1 U21343 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19273), .ZN(n19274) );
  OAI211_X1 U21344 ( .C1(n19276), .C2(n19719), .A(n19275), .B(n19274), .ZN(
        P2_U3054) );
  OAI22_X1 U21345 ( .A1(n19279), .A2(n19290), .B1(n19278), .B2(n19277), .ZN(
        n19280) );
  INV_X1 U21346 ( .A(n19280), .ZN(n19285) );
  INV_X1 U21347 ( .A(n19281), .ZN(n19282) );
  NAND3_X1 U21348 ( .A1(n19283), .A2(n19282), .A3(n19346), .ZN(n19284) );
  OAI211_X1 U21349 ( .C1(n19287), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        P2_U2914) );
  AOI22_X1 U21350 ( .A1(n19589), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n19586), .ZN(n19288) );
  OAI21_X1 U21351 ( .B1(n19290), .B2(n19591), .A(n19288), .ZN(P2_U2957) );
  AOI22_X1 U21352 ( .A1(n19589), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19289) );
  OAI21_X1 U21353 ( .B1(n19290), .B2(n19591), .A(n19289), .ZN(P2_U2972) );
  AOI22_X1 U21354 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19592), .B1(
        BUF1_REG_21__SCAN_IN), .B2(n19593), .ZN(n19342) );
  NOR2_X2 U21355 ( .A1(n19290), .A2(n19594), .ZN(n19339) );
  NAND2_X1 U21356 ( .A1(n19291), .A2(n19596), .ZN(n19336) );
  AOI22_X1 U21357 ( .A1(n19599), .A2(n19339), .B1(n19598), .B2(n19332), .ZN(
        n19293) );
  AOI22_X1 U21358 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19592), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19593), .ZN(n19337) );
  INV_X1 U21359 ( .A(n19337), .ZN(n19329) );
  AOI22_X1 U21360 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19329), .ZN(n19292) );
  OAI211_X1 U21361 ( .C1(n19342), .C2(n19719), .A(n19293), .B(n19292), .ZN(
        P2_U3173) );
  INV_X1 U21362 ( .A(n19339), .ZN(n19328) );
  OAI22_X1 U21363 ( .A1(n19620), .A2(n19337), .B1(n19336), .B2(n19607), .ZN(
        n19294) );
  INV_X1 U21364 ( .A(n19294), .ZN(n19296) );
  INV_X1 U21365 ( .A(n19342), .ZN(n19333) );
  AOI22_X1 U21366 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19611), .B1(
        n19603), .B2(n19333), .ZN(n19295) );
  OAI211_X1 U21367 ( .C1(n19328), .C2(n19614), .A(n19296), .B(n19295), .ZN(
        P2_U3165) );
  AOI22_X1 U21368 ( .A1(n19616), .A2(n19339), .B1(n19332), .B2(n19615), .ZN(
        n19298) );
  AOI22_X1 U21369 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19329), .ZN(n19297) );
  OAI211_X1 U21370 ( .C1(n19342), .C2(n19620), .A(n19298), .B(n19297), .ZN(
        P2_U3157) );
  AOI22_X1 U21371 ( .A1(n19622), .A2(n19339), .B1(n19621), .B2(n19332), .ZN(
        n19300) );
  AOI22_X1 U21372 ( .A1(n19623), .A2(n19333), .B1(n19630), .B2(n19329), .ZN(
        n19299) );
  OAI211_X1 U21373 ( .C1(n19626), .C2(n14815), .A(n19300), .B(n19299), .ZN(
        P2_U3149) );
  AOI22_X1 U21374 ( .A1(n19628), .A2(n19339), .B1(n19332), .B2(n19627), .ZN(
        n19302) );
  AOI22_X1 U21375 ( .A1(n19630), .A2(n19333), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n19629), .ZN(n19301) );
  OAI211_X1 U21376 ( .C1(n19337), .C2(n19639), .A(n19302), .B(n19301), .ZN(
        P2_U3141) );
  OAI22_X1 U21377 ( .A1(n19641), .A2(n19337), .B1(n19336), .B2(n19542), .ZN(
        n19303) );
  INV_X1 U21378 ( .A(n19303), .ZN(n19305) );
  AOI22_X1 U21379 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19636), .B1(
        n19339), .B2(n19635), .ZN(n19304) );
  OAI211_X1 U21380 ( .C1(n19342), .C2(n19639), .A(n19305), .B(n19304), .ZN(
        P2_U3133) );
  OAI22_X1 U21381 ( .A1(n19649), .A2(n19337), .B1(n19336), .B2(n19640), .ZN(
        n19306) );
  INV_X1 U21382 ( .A(n19306), .ZN(n19308) );
  AOI22_X1 U21383 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19644), .B1(
        n19634), .B2(n19333), .ZN(n19307) );
  OAI211_X1 U21384 ( .C1(n19647), .C2(n19328), .A(n19308), .B(n19307), .ZN(
        P2_U3125) );
  OAI22_X1 U21385 ( .A1(n19649), .A2(n19342), .B1(n19336), .B2(n19648), .ZN(
        n19309) );
  INV_X1 U21386 ( .A(n19309), .ZN(n19311) );
  AOI22_X1 U21387 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19652), .B1(
        n19339), .B2(n19651), .ZN(n19310) );
  OAI211_X1 U21388 ( .C1(n19337), .C2(n19661), .A(n19311), .B(n19310), .ZN(
        P2_U3117) );
  AOI22_X1 U21389 ( .A1(n19656), .A2(n19339), .B1(n19655), .B2(n19332), .ZN(
        n19313) );
  AOI22_X1 U21390 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19329), .ZN(n19312) );
  OAI211_X1 U21391 ( .C1(n19342), .C2(n19661), .A(n19313), .B(n19312), .ZN(
        P2_U3109) );
  AOI22_X1 U21392 ( .A1(n19663), .A2(n19339), .B1(n19332), .B2(n19662), .ZN(
        n19317) );
  INV_X1 U21393 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n19314) );
  OAI22_X1 U21394 ( .A1(n19670), .A2(n19337), .B1(n19557), .B2(n19314), .ZN(
        n19315) );
  INV_X1 U21395 ( .A(n19315), .ZN(n19316) );
  OAI211_X1 U21396 ( .C1(n19342), .C2(n19668), .A(n19317), .B(n19316), .ZN(
        P2_U3101) );
  OAI22_X1 U21397 ( .A1(n19677), .A2(n19337), .B1(n19336), .B2(n19669), .ZN(
        n19318) );
  INV_X1 U21398 ( .A(n19318), .ZN(n19320) );
  AOI22_X1 U21399 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19673), .B1(
        n19339), .B2(n19672), .ZN(n19319) );
  OAI211_X1 U21400 ( .C1(n19342), .C2(n19670), .A(n19320), .B(n19319), .ZN(
        P2_U3093) );
  INV_X1 U21401 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n19324) );
  OAI22_X1 U21402 ( .A1(n19677), .A2(n19342), .B1(n19336), .B2(n19676), .ZN(
        n19321) );
  INV_X1 U21403 ( .A(n19321), .ZN(n19323) );
  AOI22_X1 U21404 ( .A1(n19339), .A2(n19680), .B1(n19679), .B2(n19329), .ZN(
        n19322) );
  OAI211_X1 U21405 ( .C1(n19684), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P2_U3085) );
  OAI22_X1 U21406 ( .A1(n19700), .A2(n19337), .B1(n19336), .B2(n19685), .ZN(
        n19325) );
  INV_X1 U21407 ( .A(n19325), .ZN(n19327) );
  AOI22_X1 U21408 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19689), .B1(
        n19679), .B2(n19333), .ZN(n19326) );
  OAI211_X1 U21409 ( .C1(n19693), .C2(n19328), .A(n19327), .B(n19326), .ZN(
        P2_U3077) );
  AOI22_X1 U21410 ( .A1(n19695), .A2(n19339), .B1(n19332), .B2(n19694), .ZN(
        n19331) );
  AOI22_X1 U21411 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19329), .ZN(n19330) );
  OAI211_X1 U21412 ( .C1(n19342), .C2(n19700), .A(n19331), .B(n19330), .ZN(
        P2_U3069) );
  AOI22_X1 U21413 ( .A1(n19703), .A2(n19339), .B1(n19332), .B2(n19701), .ZN(
        n19335) );
  AOI22_X1 U21414 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19333), .ZN(n19334) );
  OAI211_X1 U21415 ( .C1(n19337), .C2(n19711), .A(n19335), .B(n19334), .ZN(
        P2_U3061) );
  OAI22_X1 U21416 ( .A1(n19719), .A2(n19337), .B1(n19336), .B2(n19710), .ZN(
        n19338) );
  INV_X1 U21417 ( .A(n19338), .ZN(n19341) );
  AOI22_X1 U21418 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19339), .ZN(n19340) );
  OAI211_X1 U21419 ( .C1(n19342), .C2(n19711), .A(n19341), .B(n19340), .ZN(
        P2_U3053) );
  INV_X1 U21420 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n22058) );
  OAI22_X1 U21421 ( .A1(n19462), .A2(n19353), .B1(n19352), .B2(n19474), .ZN(
        n19343) );
  AOI21_X1 U21422 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n19465), .A(n19343), .ZN(
        n19349) );
  AOI22_X1 U21423 ( .A1(n19347), .A2(n19346), .B1(n19345), .B2(n19344), .ZN(
        n19348) );
  OAI211_X1 U21424 ( .C1(n19463), .C2(n22058), .A(n19349), .B(n19348), .ZN(
        P2_U2899) );
  AOI22_X1 U21425 ( .A1(n19589), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19586), .ZN(n19350) );
  OAI21_X1 U21426 ( .B1(n19353), .B2(n19591), .A(n19350), .ZN(P2_U2956) );
  AOI22_X1 U21427 ( .A1(n19589), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19586), .ZN(n19351) );
  OAI21_X1 U21428 ( .B1(n19353), .B2(n19591), .A(n19351), .ZN(P2_U2971) );
  OAI22_X1 U21429 ( .A1(n22058), .A2(n19602), .B1(n19352), .B2(n19600), .ZN(
        n19397) );
  INV_X1 U21430 ( .A(n19397), .ZN(n19406) );
  NOR2_X2 U21431 ( .A1(n19353), .A2(n19594), .ZN(n19403) );
  AOI22_X1 U21432 ( .A1(n19599), .A2(n19403), .B1(n19598), .B2(n19396), .ZN(
        n19356) );
  AOI22_X1 U21433 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19592), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19593), .ZN(n19401) );
  INV_X1 U21434 ( .A(n19401), .ZN(n19393) );
  AOI22_X1 U21435 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19393), .ZN(n19355) );
  OAI211_X1 U21436 ( .C1(n19406), .C2(n19719), .A(n19356), .B(n19355), .ZN(
        P2_U3172) );
  INV_X1 U21437 ( .A(n19403), .ZN(n19392) );
  AOI22_X1 U21438 ( .A1(n19603), .A2(n19397), .B1(n19357), .B2(n19396), .ZN(
        n19359) );
  AOI22_X1 U21439 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19393), .ZN(n19358) );
  OAI211_X1 U21440 ( .C1(n19392), .C2(n19614), .A(n19359), .B(n19358), .ZN(
        P2_U3164) );
  AOI22_X1 U21441 ( .A1(n19616), .A2(n19403), .B1(n19396), .B2(n19615), .ZN(
        n19361) );
  AOI22_X1 U21442 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19393), .ZN(n19360) );
  OAI211_X1 U21443 ( .C1(n19406), .C2(n19620), .A(n19361), .B(n19360), .ZN(
        P2_U3156) );
  AOI22_X1 U21444 ( .A1(n19622), .A2(n19403), .B1(n19621), .B2(n19396), .ZN(
        n19363) );
  AOI22_X1 U21445 ( .A1(n19630), .A2(n19393), .B1(n19623), .B2(n19397), .ZN(
        n19362) );
  OAI211_X1 U21446 ( .C1(n19626), .C2(n14773), .A(n19363), .B(n19362), .ZN(
        P2_U3148) );
  AOI22_X1 U21447 ( .A1(n19628), .A2(n19403), .B1(n19396), .B2(n19627), .ZN(
        n19365) );
  AOI22_X1 U21448 ( .A1(n19630), .A2(n19397), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n19629), .ZN(n19364) );
  OAI211_X1 U21449 ( .C1(n19401), .C2(n19639), .A(n19365), .B(n19364), .ZN(
        P2_U3140) );
  AOI22_X1 U21450 ( .A1(n19366), .A2(n19397), .B1(n19396), .B2(n19633), .ZN(
        n19368) );
  AOI22_X1 U21451 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19636), .B1(
        n19403), .B2(n19635), .ZN(n19367) );
  OAI211_X1 U21452 ( .C1(n19401), .C2(n19641), .A(n19368), .B(n19367), .ZN(
        P2_U3132) );
  AOI22_X1 U21453 ( .A1(n19634), .A2(n19397), .B1(n19396), .B2(n19369), .ZN(
        n19371) );
  AOI22_X1 U21454 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19393), .ZN(n19370) );
  OAI211_X1 U21455 ( .C1(n19647), .C2(n19392), .A(n19371), .B(n19370), .ZN(
        P2_U3124) );
  INV_X1 U21456 ( .A(n19396), .ZN(n19400) );
  OAI22_X1 U21457 ( .A1(n19661), .A2(n19401), .B1(n19400), .B2(n19648), .ZN(
        n19372) );
  INV_X1 U21458 ( .A(n19372), .ZN(n19374) );
  AOI22_X1 U21459 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19652), .B1(
        n19403), .B2(n19651), .ZN(n19373) );
  OAI211_X1 U21460 ( .C1(n19406), .C2(n19649), .A(n19374), .B(n19373), .ZN(
        P2_U3116) );
  AOI22_X1 U21461 ( .A1(n19656), .A2(n19403), .B1(n19655), .B2(n19396), .ZN(
        n19376) );
  AOI22_X1 U21462 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19393), .ZN(n19375) );
  OAI211_X1 U21463 ( .C1(n19406), .C2(n19661), .A(n19376), .B(n19375), .ZN(
        P2_U3108) );
  AOI22_X1 U21464 ( .A1(n19663), .A2(n19403), .B1(n19396), .B2(n19662), .ZN(
        n19380) );
  INV_X1 U21465 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n19377) );
  OAI22_X1 U21466 ( .A1(n19670), .A2(n19401), .B1(n19557), .B2(n19377), .ZN(
        n19378) );
  INV_X1 U21467 ( .A(n19378), .ZN(n19379) );
  OAI211_X1 U21468 ( .C1(n19406), .C2(n19668), .A(n19380), .B(n19379), .ZN(
        P2_U3100) );
  AOI22_X1 U21469 ( .A1(n19397), .A2(n19665), .B1(n19396), .B2(n19381), .ZN(
        n19383) );
  AOI22_X1 U21470 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19673), .B1(
        n19403), .B2(n19672), .ZN(n19382) );
  OAI211_X1 U21471 ( .C1(n19401), .C2(n19677), .A(n19383), .B(n19382), .ZN(
        P2_U3092) );
  AOI22_X1 U21472 ( .A1(n19397), .A2(n19385), .B1(n19396), .B2(n19384), .ZN(
        n19387) );
  AOI22_X1 U21473 ( .A1(n19403), .A2(n19680), .B1(n19679), .B2(n19393), .ZN(
        n19386) );
  OAI211_X1 U21474 ( .C1(n19684), .C2(n19388), .A(n19387), .B(n19386), .ZN(
        P2_U3084) );
  AOI22_X1 U21475 ( .A1(n19397), .A2(n19679), .B1(n19396), .B2(n19389), .ZN(
        n19391) );
  INV_X1 U21476 ( .A(n19700), .ZN(n19688) );
  AOI22_X1 U21477 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19689), .B1(
        n19688), .B2(n19393), .ZN(n19390) );
  OAI211_X1 U21478 ( .C1(n19693), .C2(n19392), .A(n19391), .B(n19390), .ZN(
        P2_U3076) );
  AOI22_X1 U21479 ( .A1(n19695), .A2(n19403), .B1(n19396), .B2(n19694), .ZN(
        n19395) );
  AOI22_X1 U21480 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19393), .ZN(n19394) );
  OAI211_X1 U21481 ( .C1(n19406), .C2(n19700), .A(n19395), .B(n19394), .ZN(
        P2_U3068) );
  AOI22_X1 U21482 ( .A1(n19703), .A2(n19403), .B1(n19396), .B2(n19701), .ZN(
        n19399) );
  AOI22_X1 U21483 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19397), .ZN(n19398) );
  OAI211_X1 U21484 ( .C1(n19401), .C2(n19711), .A(n19399), .B(n19398), .ZN(
        P2_U3060) );
  OAI22_X1 U21485 ( .A1(n19719), .A2(n19401), .B1(n19710), .B2(n19400), .ZN(
        n19402) );
  INV_X1 U21486 ( .A(n19402), .ZN(n19405) );
  AOI22_X1 U21487 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19403), .ZN(n19404) );
  OAI211_X1 U21488 ( .C1(n19406), .C2(n19711), .A(n19405), .B(n19404), .ZN(
        P2_U3052) );
  AOI22_X1 U21489 ( .A1(n19589), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n19586), .ZN(n19407) );
  OAI21_X1 U21490 ( .B1(n19409), .B2(n19591), .A(n19407), .ZN(P2_U2955) );
  AOI22_X1 U21491 ( .A1(n19589), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19586), .ZN(n19408) );
  OAI21_X1 U21492 ( .B1(n19409), .B2(n19591), .A(n19408), .ZN(P2_U2970) );
  AOI22_X2 U21493 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19592), .ZN(n19456) );
  NOR2_X2 U21494 ( .A1(n19409), .A2(n19594), .ZN(n19458) );
  NAND2_X1 U21495 ( .A1(n19410), .A2(n19596), .ZN(n19455) );
  INV_X1 U21496 ( .A(n19455), .ZN(n19451) );
  AOI22_X1 U21497 ( .A1(n19599), .A2(n19458), .B1(n19598), .B2(n19451), .ZN(
        n19412) );
  AOI22_X1 U21498 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19592), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19593), .ZN(n19461) );
  INV_X1 U21499 ( .A(n19461), .ZN(n19448) );
  AOI22_X1 U21500 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19448), .ZN(n19411) );
  OAI211_X1 U21501 ( .C1(n19456), .C2(n19719), .A(n19412), .B(n19411), .ZN(
        P2_U3171) );
  INV_X1 U21502 ( .A(n19458), .ZN(n19447) );
  OAI22_X1 U21503 ( .A1(n19620), .A2(n19461), .B1(n19607), .B2(n19455), .ZN(
        n19413) );
  INV_X1 U21504 ( .A(n19413), .ZN(n19415) );
  INV_X1 U21505 ( .A(n19456), .ZN(n19452) );
  AOI22_X1 U21506 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19611), .B1(
        n19603), .B2(n19452), .ZN(n19414) );
  OAI211_X1 U21507 ( .C1(n19447), .C2(n19614), .A(n19415), .B(n19414), .ZN(
        P2_U3163) );
  AOI22_X1 U21508 ( .A1(n19616), .A2(n19458), .B1(n19451), .B2(n19615), .ZN(
        n19417) );
  AOI22_X1 U21509 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19448), .ZN(n19416) );
  OAI211_X1 U21510 ( .C1(n19456), .C2(n19620), .A(n19417), .B(n19416), .ZN(
        P2_U3155) );
  AOI22_X1 U21511 ( .A1(n19622), .A2(n19458), .B1(n19621), .B2(n19451), .ZN(
        n19419) );
  AOI22_X1 U21512 ( .A1(n19623), .A2(n19452), .B1(n19630), .B2(n19448), .ZN(
        n19418) );
  OAI211_X1 U21513 ( .C1(n19626), .C2(n14751), .A(n19419), .B(n19418), .ZN(
        P2_U3147) );
  AOI22_X1 U21514 ( .A1(n19628), .A2(n19458), .B1(n19451), .B2(n19627), .ZN(
        n19421) );
  AOI22_X1 U21515 ( .A1(n19630), .A2(n19452), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n19629), .ZN(n19420) );
  OAI211_X1 U21516 ( .C1(n19461), .C2(n19639), .A(n19421), .B(n19420), .ZN(
        P2_U3139) );
  OAI22_X1 U21517 ( .A1(n19641), .A2(n19461), .B1(n19455), .B2(n19542), .ZN(
        n19422) );
  INV_X1 U21518 ( .A(n19422), .ZN(n19424) );
  AOI22_X1 U21519 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19636), .B1(
        n19458), .B2(n19635), .ZN(n19423) );
  OAI211_X1 U21520 ( .C1(n19456), .C2(n19639), .A(n19424), .B(n19423), .ZN(
        P2_U3131) );
  OAI22_X1 U21521 ( .A1(n19641), .A2(n19456), .B1(n19455), .B2(n19640), .ZN(
        n19425) );
  INV_X1 U21522 ( .A(n19425), .ZN(n19427) );
  AOI22_X1 U21523 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19448), .ZN(n19426) );
  OAI211_X1 U21524 ( .C1(n19647), .C2(n19447), .A(n19427), .B(n19426), .ZN(
        P2_U3123) );
  OAI22_X1 U21525 ( .A1(n19649), .A2(n19456), .B1(n19455), .B2(n19648), .ZN(
        n19428) );
  INV_X1 U21526 ( .A(n19428), .ZN(n19430) );
  AOI22_X1 U21527 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19652), .B1(
        n19458), .B2(n19651), .ZN(n19429) );
  OAI211_X1 U21528 ( .C1(n19461), .C2(n19661), .A(n19430), .B(n19429), .ZN(
        P2_U3115) );
  AOI22_X1 U21529 ( .A1(n19656), .A2(n19458), .B1(n19655), .B2(n19451), .ZN(
        n19432) );
  AOI22_X1 U21530 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19448), .ZN(n19431) );
  OAI211_X1 U21531 ( .C1(n19456), .C2(n19661), .A(n19432), .B(n19431), .ZN(
        P2_U3107) );
  AOI22_X1 U21532 ( .A1(n19663), .A2(n19458), .B1(n19451), .B2(n19662), .ZN(
        n19436) );
  INV_X1 U21533 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n19433) );
  OAI22_X1 U21534 ( .A1(n19670), .A2(n19461), .B1(n19557), .B2(n19433), .ZN(
        n19434) );
  INV_X1 U21535 ( .A(n19434), .ZN(n19435) );
  OAI211_X1 U21536 ( .C1(n19456), .C2(n19668), .A(n19436), .B(n19435), .ZN(
        P2_U3099) );
  OAI22_X1 U21537 ( .A1(n19670), .A2(n19456), .B1(n19669), .B2(n19455), .ZN(
        n19437) );
  INV_X1 U21538 ( .A(n19437), .ZN(n19439) );
  AOI22_X1 U21539 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19673), .B1(
        n19458), .B2(n19672), .ZN(n19438) );
  OAI211_X1 U21540 ( .C1(n19461), .C2(n19677), .A(n19439), .B(n19438), .ZN(
        P2_U3091) );
  OAI22_X1 U21541 ( .A1(n19677), .A2(n19456), .B1(n19455), .B2(n19676), .ZN(
        n19440) );
  INV_X1 U21542 ( .A(n19440), .ZN(n19442) );
  AOI22_X1 U21543 ( .A1(n19458), .A2(n19680), .B1(n19679), .B2(n19448), .ZN(
        n19441) );
  OAI211_X1 U21544 ( .C1(n19684), .C2(n19443), .A(n19442), .B(n19441), .ZN(
        P2_U3083) );
  OAI22_X1 U21545 ( .A1(n19686), .A2(n19456), .B1(n19455), .B2(n19685), .ZN(
        n19444) );
  INV_X1 U21546 ( .A(n19444), .ZN(n19446) );
  AOI22_X1 U21547 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19689), .B1(
        n19688), .B2(n19448), .ZN(n19445) );
  OAI211_X1 U21548 ( .C1(n19693), .C2(n19447), .A(n19446), .B(n19445), .ZN(
        P2_U3075) );
  AOI22_X1 U21549 ( .A1(n19695), .A2(n19458), .B1(n19451), .B2(n19694), .ZN(
        n19450) );
  AOI22_X1 U21550 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19448), .ZN(n19449) );
  OAI211_X1 U21551 ( .C1(n19456), .C2(n19700), .A(n19450), .B(n19449), .ZN(
        P2_U3067) );
  AOI22_X1 U21552 ( .A1(n19703), .A2(n19458), .B1(n19451), .B2(n19701), .ZN(
        n19454) );
  AOI22_X1 U21553 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19452), .ZN(n19453) );
  OAI211_X1 U21554 ( .C1(n19461), .C2(n19711), .A(n19454), .B(n19453), .ZN(
        P2_U3059) );
  OAI22_X1 U21555 ( .A1(n19711), .A2(n19456), .B1(n19455), .B2(n19710), .ZN(
        n19457) );
  INV_X1 U21556 ( .A(n19457), .ZN(n19460) );
  AOI22_X1 U21557 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19458), .ZN(n19459) );
  OAI211_X1 U21558 ( .C1(n19461), .C2(n19719), .A(n19460), .B(n19459), .ZN(
        P2_U3051) );
  INV_X1 U21559 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19473) );
  INV_X1 U21560 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21963) );
  OAI22_X1 U21561 ( .A1(n19463), .A2(n21963), .B1(n19462), .B2(n19477), .ZN(
        n19464) );
  AOI21_X1 U21562 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n19465), .A(n19464), .ZN(
        n19472) );
  OAI22_X1 U21563 ( .A1(n19469), .A2(n19468), .B1(n19467), .B2(n19466), .ZN(
        n19470) );
  INV_X1 U21564 ( .A(n19470), .ZN(n19471) );
  OAI211_X1 U21565 ( .C1(n19474), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P2_U2901) );
  AOI22_X1 U21566 ( .A1(n19587), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19586), .ZN(n19475) );
  OAI21_X1 U21567 ( .B1(n19477), .B2(n19591), .A(n19475), .ZN(P2_U2954) );
  AOI22_X1 U21568 ( .A1(n19587), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19586), .ZN(n19476) );
  OAI21_X1 U21569 ( .B1(n19477), .B2(n19591), .A(n19476), .ZN(P2_U2969) );
  AOI22_X2 U21570 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n19592), .B1(
        BUF1_REG_18__SCAN_IN), .B2(n19593), .ZN(n19524) );
  NOR2_X2 U21571 ( .A1(n19477), .A2(n19594), .ZN(n19526) );
  NAND2_X1 U21572 ( .A1(n12353), .A2(n19596), .ZN(n19523) );
  AOI22_X1 U21573 ( .A1(n19599), .A2(n19526), .B1(n19598), .B2(n19519), .ZN(
        n19480) );
  INV_X1 U21574 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21961) );
  OAI22_X1 U21575 ( .A1(n21961), .A2(n19602), .B1(n19478), .B2(n19600), .ZN(
        n19520) );
  AOI22_X1 U21576 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19520), .ZN(n19479) );
  OAI211_X1 U21577 ( .C1(n19524), .C2(n19719), .A(n19480), .B(n19479), .ZN(
        P2_U3170) );
  INV_X1 U21578 ( .A(n19526), .ZN(n19516) );
  OAI22_X1 U21579 ( .A1(n19524), .A2(n19608), .B1(n19607), .B2(n19523), .ZN(
        n19481) );
  INV_X1 U21580 ( .A(n19481), .ZN(n19483) );
  AOI22_X1 U21581 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19520), .ZN(n19482) );
  OAI211_X1 U21582 ( .C1(n19516), .C2(n19614), .A(n19483), .B(n19482), .ZN(
        P2_U3162) );
  AOI22_X1 U21583 ( .A1(n19616), .A2(n19526), .B1(n19519), .B2(n19615), .ZN(
        n19485) );
  AOI22_X1 U21584 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19520), .ZN(n19484) );
  OAI211_X1 U21585 ( .C1(n19524), .C2(n19620), .A(n19485), .B(n19484), .ZN(
        P2_U3154) );
  AOI22_X1 U21586 ( .A1(n19622), .A2(n19526), .B1(n19621), .B2(n19519), .ZN(
        n19487) );
  INV_X1 U21587 ( .A(n19524), .ZN(n19513) );
  AOI22_X1 U21588 ( .A1(n19623), .A2(n19513), .B1(n19630), .B2(n19520), .ZN(
        n19486) );
  OAI211_X1 U21589 ( .C1(n19626), .C2(n14590), .A(n19487), .B(n19486), .ZN(
        P2_U3146) );
  INV_X1 U21590 ( .A(n19520), .ZN(n19529) );
  AOI22_X1 U21591 ( .A1(n19628), .A2(n19526), .B1(n19519), .B2(n19627), .ZN(
        n19489) );
  AOI22_X1 U21592 ( .A1(n19513), .A2(n19630), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n19629), .ZN(n19488) );
  OAI211_X1 U21593 ( .C1(n19529), .C2(n19639), .A(n19489), .B(n19488), .ZN(
        P2_U3138) );
  OAI22_X1 U21594 ( .A1(n19641), .A2(n19529), .B1(n19523), .B2(n19542), .ZN(
        n19490) );
  INV_X1 U21595 ( .A(n19490), .ZN(n19492) );
  AOI22_X1 U21596 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19636), .B1(
        n19526), .B2(n19635), .ZN(n19491) );
  OAI211_X1 U21597 ( .C1(n19524), .C2(n19639), .A(n19492), .B(n19491), .ZN(
        P2_U3130) );
  OAI22_X1 U21598 ( .A1(n19524), .A2(n19641), .B1(n19523), .B2(n19640), .ZN(
        n19493) );
  INV_X1 U21599 ( .A(n19493), .ZN(n19495) );
  AOI22_X1 U21600 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19520), .ZN(n19494) );
  OAI211_X1 U21601 ( .C1(n19647), .C2(n19516), .A(n19495), .B(n19494), .ZN(
        P2_U3122) );
  OAI22_X1 U21602 ( .A1(n19524), .A2(n19649), .B1(n19523), .B2(n19648), .ZN(
        n19496) );
  INV_X1 U21603 ( .A(n19496), .ZN(n19498) );
  AOI22_X1 U21604 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19652), .B1(
        n19526), .B2(n19651), .ZN(n19497) );
  OAI211_X1 U21605 ( .C1(n19529), .C2(n19661), .A(n19498), .B(n19497), .ZN(
        P2_U3114) );
  AOI22_X1 U21606 ( .A1(n19656), .A2(n19526), .B1(n19655), .B2(n19519), .ZN(
        n19500) );
  AOI22_X1 U21607 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19520), .ZN(n19499) );
  OAI211_X1 U21608 ( .C1(n19524), .C2(n19661), .A(n19500), .B(n19499), .ZN(
        P2_U3106) );
  AOI22_X1 U21609 ( .A1(n19663), .A2(n19526), .B1(n19519), .B2(n19662), .ZN(
        n19504) );
  INV_X1 U21610 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n19501) );
  OAI22_X1 U21611 ( .A1(n19670), .A2(n19529), .B1(n19557), .B2(n19501), .ZN(
        n19502) );
  INV_X1 U21612 ( .A(n19502), .ZN(n19503) );
  OAI211_X1 U21613 ( .C1(n19524), .C2(n19668), .A(n19504), .B(n19503), .ZN(
        P2_U3098) );
  OAI22_X1 U21614 ( .A1(n19677), .A2(n19529), .B1(n19523), .B2(n19669), .ZN(
        n19505) );
  INV_X1 U21615 ( .A(n19505), .ZN(n19507) );
  AOI22_X1 U21616 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19673), .B1(
        n19526), .B2(n19672), .ZN(n19506) );
  OAI211_X1 U21617 ( .C1(n19524), .C2(n19670), .A(n19507), .B(n19506), .ZN(
        P2_U3090) );
  INV_X1 U21618 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19511) );
  OAI22_X1 U21619 ( .A1(n19524), .A2(n19677), .B1(n19523), .B2(n19676), .ZN(
        n19508) );
  INV_X1 U21620 ( .A(n19508), .ZN(n19510) );
  AOI22_X1 U21621 ( .A1(n19526), .A2(n19680), .B1(n19679), .B2(n19520), .ZN(
        n19509) );
  OAI211_X1 U21622 ( .C1(n19684), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P2_U3082) );
  OAI22_X1 U21623 ( .A1(n19700), .A2(n19529), .B1(n19523), .B2(n19685), .ZN(
        n19512) );
  INV_X1 U21624 ( .A(n19512), .ZN(n19515) );
  AOI22_X1 U21625 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19689), .B1(
        n19679), .B2(n19513), .ZN(n19514) );
  OAI211_X1 U21626 ( .C1(n19693), .C2(n19516), .A(n19515), .B(n19514), .ZN(
        P2_U3074) );
  AOI22_X1 U21627 ( .A1(n19695), .A2(n19526), .B1(n19519), .B2(n19694), .ZN(
        n19518) );
  AOI22_X1 U21628 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19520), .ZN(n19517) );
  OAI211_X1 U21629 ( .C1(n19524), .C2(n19700), .A(n19518), .B(n19517), .ZN(
        P2_U3066) );
  AOI22_X1 U21630 ( .A1(n19703), .A2(n19526), .B1(n19519), .B2(n19701), .ZN(
        n19522) );
  AOI22_X1 U21631 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19706), .B1(
        n19575), .B2(n19520), .ZN(n19521) );
  OAI211_X1 U21632 ( .C1(n19524), .C2(n19578), .A(n19522), .B(n19521), .ZN(
        P2_U3058) );
  OAI22_X1 U21633 ( .A1(n19524), .A2(n19711), .B1(n19710), .B2(n19523), .ZN(
        n19525) );
  INV_X1 U21634 ( .A(n19525), .ZN(n19528) );
  AOI22_X1 U21635 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19526), .ZN(n19527) );
  OAI211_X1 U21636 ( .C1(n19529), .C2(n19719), .A(n19528), .B(n19527), .ZN(
        P2_U3050) );
  AOI22_X1 U21637 ( .A1(n19587), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n19586), .ZN(n19530) );
  OAI21_X1 U21638 ( .B1(n19532), .B2(n19591), .A(n19530), .ZN(P2_U2953) );
  AOI22_X1 U21639 ( .A1(n19587), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19586), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19531) );
  OAI21_X1 U21640 ( .B1(n19532), .B2(n19591), .A(n19531), .ZN(P2_U2968) );
  AOI22_X1 U21641 ( .A1(n19599), .A2(n19582), .B1(n19598), .B2(n19573), .ZN(
        n19534) );
  AOI22_X1 U21642 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19574), .ZN(n19533) );
  OAI211_X1 U21643 ( .C1(n19580), .C2(n19719), .A(n19534), .B(n19533), .ZN(
        P2_U3169) );
  INV_X1 U21644 ( .A(n19582), .ZN(n19570) );
  INV_X1 U21645 ( .A(n19573), .ZN(n19579) );
  OAI22_X1 U21646 ( .A1(n19608), .A2(n19580), .B1(n19579), .B2(n19607), .ZN(
        n19535) );
  INV_X1 U21647 ( .A(n19535), .ZN(n19537) );
  AOI22_X1 U21648 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19574), .ZN(n19536) );
  OAI211_X1 U21649 ( .C1(n19570), .C2(n19614), .A(n19537), .B(n19536), .ZN(
        P2_U3161) );
  AOI22_X1 U21650 ( .A1(n19616), .A2(n19582), .B1(n19573), .B2(n19615), .ZN(
        n19539) );
  AOI22_X1 U21651 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19574), .ZN(n19538) );
  OAI211_X1 U21652 ( .C1(n19580), .C2(n19620), .A(n19539), .B(n19538), .ZN(
        P2_U3153) );
  AOI22_X1 U21653 ( .A1(n19628), .A2(n19582), .B1(n19573), .B2(n19627), .ZN(
        n19541) );
  AOI22_X1 U21654 ( .A1(n19630), .A2(n19552), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n19629), .ZN(n19540) );
  OAI211_X1 U21655 ( .C1(n19585), .C2(n19639), .A(n19541), .B(n19540), .ZN(
        P2_U3137) );
  OAI22_X1 U21656 ( .A1(n19641), .A2(n19585), .B1(n19579), .B2(n19542), .ZN(
        n19543) );
  INV_X1 U21657 ( .A(n19543), .ZN(n19545) );
  AOI22_X1 U21658 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19636), .B1(
        n19582), .B2(n19635), .ZN(n19544) );
  OAI211_X1 U21659 ( .C1(n19580), .C2(n19639), .A(n19545), .B(n19544), .ZN(
        P2_U3129) );
  OAI22_X1 U21660 ( .A1(n19649), .A2(n19585), .B1(n19579), .B2(n19640), .ZN(
        n19546) );
  INV_X1 U21661 ( .A(n19546), .ZN(n19548) );
  AOI22_X1 U21662 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19644), .B1(
        n19634), .B2(n19552), .ZN(n19547) );
  OAI211_X1 U21663 ( .C1(n19647), .C2(n19570), .A(n19548), .B(n19547), .ZN(
        P2_U3121) );
  OAI22_X1 U21664 ( .A1(n19661), .A2(n19585), .B1(n19579), .B2(n19648), .ZN(
        n19549) );
  INV_X1 U21665 ( .A(n19549), .ZN(n19551) );
  AOI22_X1 U21666 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19652), .B1(
        n19582), .B2(n19651), .ZN(n19550) );
  OAI211_X1 U21667 ( .C1(n19580), .C2(n19649), .A(n19551), .B(n19550), .ZN(
        P2_U3113) );
  AOI22_X1 U21668 ( .A1(n19656), .A2(n19582), .B1(n19573), .B2(n19655), .ZN(
        n19555) );
  INV_X1 U21669 ( .A(n19661), .ZN(n19553) );
  AOI22_X1 U21670 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19658), .B1(
        n19553), .B2(n19552), .ZN(n19554) );
  OAI211_X1 U21671 ( .C1(n19585), .C2(n19668), .A(n19555), .B(n19554), .ZN(
        P2_U3105) );
  AOI22_X1 U21672 ( .A1(n19663), .A2(n19582), .B1(n19573), .B2(n19662), .ZN(
        n19560) );
  INV_X1 U21673 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n19556) );
  OAI22_X1 U21674 ( .A1(n19670), .A2(n19585), .B1(n19557), .B2(n19556), .ZN(
        n19558) );
  INV_X1 U21675 ( .A(n19558), .ZN(n19559) );
  OAI211_X1 U21676 ( .C1(n19580), .C2(n19668), .A(n19560), .B(n19559), .ZN(
        P2_U3097) );
  OAI22_X1 U21677 ( .A1(n19670), .A2(n19580), .B1(n19579), .B2(n19669), .ZN(
        n19561) );
  INV_X1 U21678 ( .A(n19561), .ZN(n19563) );
  AOI22_X1 U21679 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19673), .B1(
        n19582), .B2(n19672), .ZN(n19562) );
  OAI211_X1 U21680 ( .C1(n19585), .C2(n19677), .A(n19563), .B(n19562), .ZN(
        P2_U3089) );
  OAI22_X1 U21681 ( .A1(n19677), .A2(n19580), .B1(n19579), .B2(n19676), .ZN(
        n19564) );
  INV_X1 U21682 ( .A(n19564), .ZN(n19566) );
  AOI22_X1 U21683 ( .A1(n19582), .A2(n19680), .B1(n19679), .B2(n19574), .ZN(
        n19565) );
  OAI211_X1 U21684 ( .C1(n19684), .C2(n11142), .A(n19566), .B(n19565), .ZN(
        P2_U3081) );
  OAI22_X1 U21685 ( .A1(n19686), .A2(n19580), .B1(n19579), .B2(n19685), .ZN(
        n19567) );
  INV_X1 U21686 ( .A(n19567), .ZN(n19569) );
  AOI22_X1 U21687 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19689), .B1(
        n19688), .B2(n19574), .ZN(n19568) );
  OAI211_X1 U21688 ( .C1(n19693), .C2(n19570), .A(n19569), .B(n19568), .ZN(
        P2_U3073) );
  AOI22_X1 U21689 ( .A1(n19695), .A2(n19582), .B1(n19573), .B2(n19694), .ZN(
        n19572) );
  AOI22_X1 U21690 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19574), .ZN(n19571) );
  OAI211_X1 U21691 ( .C1(n19580), .C2(n19700), .A(n19572), .B(n19571), .ZN(
        P2_U3065) );
  AOI22_X1 U21692 ( .A1(n19703), .A2(n19582), .B1(n19573), .B2(n19701), .ZN(
        n19577) );
  AOI22_X1 U21693 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19706), .B1(
        n19575), .B2(n19574), .ZN(n19576) );
  OAI211_X1 U21694 ( .C1(n19580), .C2(n19578), .A(n19577), .B(n19576), .ZN(
        P2_U3057) );
  OAI22_X1 U21695 ( .A1(n19711), .A2(n19580), .B1(n19579), .B2(n19710), .ZN(
        n19581) );
  INV_X1 U21696 ( .A(n19581), .ZN(n19584) );
  AOI22_X1 U21697 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19582), .ZN(n19583) );
  OAI211_X1 U21698 ( .C1(n19585), .C2(n19719), .A(n19584), .B(n19583), .ZN(
        P2_U3049) );
  AOI22_X1 U21699 ( .A1(n19587), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19586), .ZN(n19588) );
  OAI21_X1 U21700 ( .B1(n19595), .B2(n19591), .A(n19588), .ZN(P2_U2952) );
  AOI22_X1 U21701 ( .A1(n19589), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19586), .ZN(n19590) );
  OAI21_X1 U21702 ( .B1(n19595), .B2(n19591), .A(n19590), .ZN(P2_U2967) );
  AOI22_X2 U21703 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19593), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19592), .ZN(n19712) );
  NOR2_X2 U21704 ( .A1(n19595), .A2(n19594), .ZN(n19714) );
  NAND2_X1 U21705 ( .A1(n19597), .A2(n19596), .ZN(n19709) );
  AOI22_X1 U21706 ( .A1(n19599), .A2(n19714), .B1(n19598), .B2(n19702), .ZN(
        n19606) );
  INV_X1 U21707 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n21714) );
  OAI22_X2 U21708 ( .A1(n21714), .A2(n19602), .B1(n19601), .B2(n19600), .ZN(
        n19696) );
  AOI22_X1 U21709 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19696), .ZN(n19605) );
  OAI211_X1 U21710 ( .C1(n19712), .C2(n19719), .A(n19606), .B(n19605), .ZN(
        P2_U3168) );
  INV_X1 U21711 ( .A(n19714), .ZN(n19692) );
  OAI22_X1 U21712 ( .A1(n19712), .A2(n19608), .B1(n19607), .B2(n19709), .ZN(
        n19609) );
  INV_X1 U21713 ( .A(n19609), .ZN(n19613) );
  AOI22_X1 U21714 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19696), .ZN(n19612) );
  OAI211_X1 U21715 ( .C1(n19692), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P2_U3160) );
  AOI22_X1 U21716 ( .A1(n19616), .A2(n19714), .B1(n19702), .B2(n19615), .ZN(
        n19619) );
  AOI22_X1 U21717 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19617), .B1(
        n19623), .B2(n19696), .ZN(n19618) );
  OAI211_X1 U21718 ( .C1(n19712), .C2(n19620), .A(n19619), .B(n19618), .ZN(
        P2_U3152) );
  AOI22_X1 U21719 ( .A1(n19622), .A2(n19714), .B1(n19621), .B2(n19702), .ZN(
        n19625) );
  INV_X1 U21720 ( .A(n19712), .ZN(n19704) );
  AOI22_X1 U21721 ( .A1(n19623), .A2(n19704), .B1(n19630), .B2(n19696), .ZN(
        n19624) );
  OAI211_X1 U21722 ( .C1(n19626), .C2(n14509), .A(n19625), .B(n19624), .ZN(
        P2_U3144) );
  INV_X1 U21723 ( .A(n19696), .ZN(n19720) );
  AOI22_X1 U21724 ( .A1(n19628), .A2(n19714), .B1(n19702), .B2(n19627), .ZN(
        n19632) );
  AOI22_X1 U21725 ( .A1(n19704), .A2(n19630), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n19629), .ZN(n19631) );
  OAI211_X1 U21726 ( .C1(n19720), .C2(n19639), .A(n19632), .B(n19631), .ZN(
        P2_U3136) );
  AOI22_X1 U21727 ( .A1(n19634), .A2(n19696), .B1(n19702), .B2(n19633), .ZN(
        n19638) );
  AOI22_X1 U21728 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19636), .B1(
        n19714), .B2(n19635), .ZN(n19637) );
  OAI211_X1 U21729 ( .C1(n19712), .C2(n19639), .A(n19638), .B(n19637), .ZN(
        P2_U3128) );
  OAI22_X1 U21730 ( .A1(n19712), .A2(n19641), .B1(n19709), .B2(n19640), .ZN(
        n19642) );
  INV_X1 U21731 ( .A(n19642), .ZN(n19646) );
  AOI22_X1 U21732 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19644), .B1(
        n19643), .B2(n19696), .ZN(n19645) );
  OAI211_X1 U21733 ( .C1(n19647), .C2(n19692), .A(n19646), .B(n19645), .ZN(
        P2_U3120) );
  OAI22_X1 U21734 ( .A1(n19712), .A2(n19649), .B1(n19709), .B2(n19648), .ZN(
        n19650) );
  INV_X1 U21735 ( .A(n19650), .ZN(n19654) );
  AOI22_X1 U21736 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19652), .B1(
        n19714), .B2(n19651), .ZN(n19653) );
  OAI211_X1 U21737 ( .C1(n19720), .C2(n19661), .A(n19654), .B(n19653), .ZN(
        P2_U3112) );
  AOI22_X1 U21738 ( .A1(n19656), .A2(n19714), .B1(n19655), .B2(n19702), .ZN(
        n19660) );
  AOI22_X1 U21739 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19658), .B1(
        n19657), .B2(n19696), .ZN(n19659) );
  OAI211_X1 U21740 ( .C1(n19712), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3104) );
  AOI22_X1 U21741 ( .A1(n19663), .A2(n19714), .B1(n19702), .B2(n19662), .ZN(
        n19667) );
  AOI22_X1 U21742 ( .A1(n19696), .A2(n19665), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n19664), .ZN(n19666) );
  OAI211_X1 U21743 ( .C1(n19712), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        P2_U3096) );
  OAI22_X1 U21744 ( .A1(n19712), .A2(n19670), .B1(n19669), .B2(n19709), .ZN(
        n19671) );
  INV_X1 U21745 ( .A(n19671), .ZN(n19675) );
  AOI22_X1 U21746 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19673), .B1(
        n19714), .B2(n19672), .ZN(n19674) );
  OAI211_X1 U21747 ( .C1(n19720), .C2(n19677), .A(n19675), .B(n19674), .ZN(
        P2_U3088) );
  INV_X1 U21748 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19683) );
  OAI22_X1 U21749 ( .A1(n19712), .A2(n19677), .B1(n19709), .B2(n19676), .ZN(
        n19678) );
  INV_X1 U21750 ( .A(n19678), .ZN(n19682) );
  AOI22_X1 U21751 ( .A1(n19714), .A2(n19680), .B1(n19679), .B2(n19696), .ZN(
        n19681) );
  OAI211_X1 U21752 ( .C1(n19684), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P2_U3080) );
  OAI22_X1 U21753 ( .A1(n19712), .A2(n19686), .B1(n19709), .B2(n19685), .ZN(
        n19687) );
  INV_X1 U21754 ( .A(n19687), .ZN(n19691) );
  AOI22_X1 U21755 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19689), .B1(
        n19688), .B2(n19696), .ZN(n19690) );
  OAI211_X1 U21756 ( .C1(n19693), .C2(n19692), .A(n19691), .B(n19690), .ZN(
        P2_U3072) );
  AOI22_X1 U21757 ( .A1(n19695), .A2(n19714), .B1(n19702), .B2(n19694), .ZN(
        n19699) );
  AOI22_X1 U21758 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19697), .B1(
        n19705), .B2(n19696), .ZN(n19698) );
  OAI211_X1 U21759 ( .C1(n19712), .C2(n19700), .A(n19699), .B(n19698), .ZN(
        P2_U3064) );
  AOI22_X1 U21760 ( .A1(n19703), .A2(n19714), .B1(n19702), .B2(n19701), .ZN(
        n19708) );
  AOI22_X1 U21761 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19706), .B1(
        n19705), .B2(n19704), .ZN(n19707) );
  OAI211_X1 U21762 ( .C1(n19720), .C2(n19711), .A(n19708), .B(n19707), .ZN(
        P2_U3056) );
  OAI22_X1 U21763 ( .A1(n19712), .A2(n19711), .B1(n19710), .B2(n19709), .ZN(
        n19713) );
  INV_X1 U21764 ( .A(n19713), .ZN(n19718) );
  AOI22_X1 U21765 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19716), .B1(
        n19715), .B2(n19714), .ZN(n19717) );
  OAI211_X1 U21766 ( .C1(n19720), .C2(n19719), .A(n19718), .B(n19717), .ZN(
        P2_U3048) );
  INV_X1 U21767 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20012) );
  INV_X1 U21768 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19721) );
  AOI222_X1 U21769 ( .A1(n20012), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20014), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19721), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19722) );
  INV_X1 U21770 ( .A(n19776), .ZN(n19774) );
  OAI22_X1 U21771 ( .A1(n19776), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n19774), .ZN(n19723) );
  INV_X1 U21772 ( .A(n19723), .ZN(U376) );
  OAI22_X1 U21773 ( .A1(n19776), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n19774), .ZN(n19724) );
  INV_X1 U21774 ( .A(n19724), .ZN(U365) );
  INV_X1 U21775 ( .A(n19776), .ZN(n19779) );
  AOI22_X1 U21776 ( .A1(n19779), .A2(n19726), .B1(n19725), .B2(n19776), .ZN(
        U354) );
  OAI22_X1 U21777 ( .A1(n19776), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n19774), .ZN(n19727) );
  INV_X1 U21778 ( .A(n19727), .ZN(U353) );
  OAI22_X1 U21779 ( .A1(n19776), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n19774), .ZN(n19728) );
  INV_X1 U21780 ( .A(n19728), .ZN(U352) );
  AOI22_X1 U21781 ( .A1(n19779), .A2(n19730), .B1(n19729), .B2(n19776), .ZN(
        U351) );
  AOI22_X1 U21782 ( .A1(n19779), .A2(n19732), .B1(n19731), .B2(n19776), .ZN(
        U350) );
  AOI22_X1 U21783 ( .A1(n19779), .A2(n19734), .B1(n19733), .B2(n19776), .ZN(
        U349) );
  AOI22_X1 U21784 ( .A1(n19779), .A2(n19736), .B1(n19735), .B2(n19776), .ZN(
        U348) );
  AOI22_X1 U21785 ( .A1(n19779), .A2(n19738), .B1(n19737), .B2(n19776), .ZN(
        U347) );
  AOI22_X1 U21786 ( .A1(n19779), .A2(n19740), .B1(n19739), .B2(n19776), .ZN(
        U375) );
  AOI22_X1 U21787 ( .A1(n19779), .A2(n19742), .B1(n19741), .B2(n19776), .ZN(
        U374) );
  AOI22_X1 U21788 ( .A1(n19779), .A2(n19744), .B1(n19743), .B2(n19776), .ZN(
        U373) );
  AOI22_X1 U21789 ( .A1(n19779), .A2(n19746), .B1(n19745), .B2(n19776), .ZN(
        U372) );
  AOI22_X1 U21790 ( .A1(n19779), .A2(n19748), .B1(n19747), .B2(n19776), .ZN(
        U371) );
  AOI22_X1 U21791 ( .A1(n19779), .A2(n19750), .B1(n19749), .B2(n19776), .ZN(
        U370) );
  AOI22_X1 U21792 ( .A1(n19779), .A2(n19752), .B1(n19751), .B2(n19776), .ZN(
        U369) );
  AOI22_X1 U21793 ( .A1(n19779), .A2(n19754), .B1(n19753), .B2(n19776), .ZN(
        U368) );
  AOI22_X1 U21794 ( .A1(n19779), .A2(n19756), .B1(n19755), .B2(n19776), .ZN(
        U367) );
  AOI22_X1 U21795 ( .A1(n19779), .A2(n19758), .B1(n19757), .B2(n19776), .ZN(
        U366) );
  AOI22_X1 U21796 ( .A1(n19779), .A2(n19760), .B1(n19759), .B2(n19776), .ZN(
        U364) );
  AOI22_X1 U21797 ( .A1(n19779), .A2(n19762), .B1(n19761), .B2(n19776), .ZN(
        U363) );
  AOI22_X1 U21798 ( .A1(n19779), .A2(n19764), .B1(n19763), .B2(n19776), .ZN(
        U362) );
  AOI22_X1 U21799 ( .A1(n19779), .A2(n19766), .B1(n19765), .B2(n19776), .ZN(
        U361) );
  AOI22_X1 U21800 ( .A1(n19779), .A2(n19768), .B1(n19767), .B2(n19776), .ZN(
        U360) );
  AOI22_X1 U21801 ( .A1(n19779), .A2(n19770), .B1(n19769), .B2(n19776), .ZN(
        U359) );
  AOI22_X1 U21802 ( .A1(n19779), .A2(n19772), .B1(n19771), .B2(n19776), .ZN(
        U358) );
  OAI22_X1 U21803 ( .A1(n19776), .A2(P3_ADDRESS_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n19774), .ZN(n19773) );
  INV_X1 U21804 ( .A(n19773), .ZN(U357) );
  OAI22_X1 U21805 ( .A1(n19776), .A2(P3_ADDRESS_REG_28__SCAN_IN), .B1(
        P2_ADDRESS_REG_28__SCAN_IN), .B2(n19774), .ZN(n19775) );
  INV_X1 U21806 ( .A(n19775), .ZN(U356) );
  AOI22_X1 U21807 ( .A1(n19779), .A2(n19778), .B1(n19777), .B2(n19776), .ZN(
        U355) );
  AOI22_X1 U21808 ( .A1(n21200), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19781) );
  OAI21_X1 U21809 ( .B1(n19782), .B2(n19815), .A(n19781), .ZN(P1_U2936) );
  AOI22_X1 U21810 ( .A1(n19797), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19783) );
  OAI21_X1 U21811 ( .B1(n19784), .B2(n19815), .A(n19783), .ZN(P1_U2935) );
  AOI22_X1 U21812 ( .A1(n19797), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19785) );
  OAI21_X1 U21813 ( .B1(n19786), .B2(n19815), .A(n19785), .ZN(P1_U2934) );
  AOI22_X1 U21814 ( .A1(n19797), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19787) );
  OAI21_X1 U21815 ( .B1(n19788), .B2(n19815), .A(n19787), .ZN(P1_U2933) );
  AOI22_X1 U21816 ( .A1(n19797), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19789) );
  OAI21_X1 U21817 ( .B1(n19790), .B2(n19815), .A(n19789), .ZN(P1_U2932) );
  AOI22_X1 U21818 ( .A1(n19797), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19791) );
  OAI21_X1 U21819 ( .B1(n19792), .B2(n19815), .A(n19791), .ZN(P1_U2931) );
  AOI22_X1 U21820 ( .A1(n19797), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19793) );
  OAI21_X1 U21821 ( .B1(n19794), .B2(n19815), .A(n19793), .ZN(P1_U2930) );
  AOI22_X1 U21822 ( .A1(n21200), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19795) );
  OAI21_X1 U21823 ( .B1(n19796), .B2(n19815), .A(n19795), .ZN(P1_U2929) );
  AOI22_X1 U21824 ( .A1(n19797), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19798) );
  OAI21_X1 U21825 ( .B1(n19799), .B2(n19815), .A(n19798), .ZN(P1_U2928) );
  AOI22_X1 U21826 ( .A1(n21200), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19800) );
  OAI21_X1 U21827 ( .B1(n19801), .B2(n19815), .A(n19800), .ZN(P1_U2927) );
  AOI22_X1 U21828 ( .A1(n21200), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19802), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19803) );
  OAI21_X1 U21829 ( .B1(n19804), .B2(n19815), .A(n19803), .ZN(P1_U2926) );
  AOI22_X1 U21830 ( .A1(n21200), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U21831 ( .B1(n19806), .B2(n19815), .A(n19805), .ZN(P1_U2925) );
  AOI22_X1 U21832 ( .A1(n21200), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U21833 ( .B1(n19808), .B2(n19815), .A(n19807), .ZN(P1_U2924) );
  AOI22_X1 U21834 ( .A1(n21200), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U21835 ( .B1(n19810), .B2(n19815), .A(n19809), .ZN(P1_U2923) );
  AOI22_X1 U21836 ( .A1(n21200), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19811) );
  OAI21_X1 U21837 ( .B1(n19812), .B2(n19815), .A(n19811), .ZN(P1_U2922) );
  AOI22_X1 U21838 ( .A1(n21200), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19813), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19814) );
  OAI21_X1 U21839 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(P1_U2921) );
  NOR2_X1 U21840 ( .A1(n11057), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19837) );
  INV_X1 U21841 ( .A(n19837), .ZN(n19841) );
  NOR2_X1 U21842 ( .A1(n12962), .A2(n11057), .ZN(n19852) );
  INV_X1 U21843 ( .A(n19852), .ZN(n19839) );
  OAI222_X1 U21844 ( .A1(n19841), .A2(n21231), .B1(n19817), .B2(n22319), .C1(
        n13784), .C2(n19839), .ZN(P1_U3197) );
  INV_X1 U21845 ( .A(n19839), .ZN(n19849) );
  AOI222_X1 U21846 ( .A1(n19837), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n19849), .ZN(n19818) );
  INV_X1 U21847 ( .A(n19818), .ZN(P1_U3198) );
  AOI222_X1 U21848 ( .A1(n19837), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n19849), .ZN(n19819) );
  INV_X1 U21849 ( .A(n19819), .ZN(P1_U3199) );
  AOI222_X1 U21850 ( .A1(n19837), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n19849), .ZN(n19820) );
  INV_X1 U21851 ( .A(n19820), .ZN(P1_U3200) );
  AOI222_X1 U21852 ( .A1(n19837), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n19849), .ZN(n19821) );
  INV_X1 U21853 ( .A(n19821), .ZN(P1_U3201) );
  AOI222_X1 U21854 ( .A1(n19837), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n19849), .ZN(n19822) );
  INV_X1 U21855 ( .A(n19822), .ZN(P1_U3202) );
  AOI222_X1 U21856 ( .A1(n19837), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n19849), .ZN(n19823) );
  INV_X1 U21857 ( .A(n19823), .ZN(P1_U3203) );
  AOI222_X1 U21858 ( .A1(n19837), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n19849), .ZN(n19824) );
  INV_X1 U21859 ( .A(n19824), .ZN(P1_U3204) );
  INV_X1 U21860 ( .A(n19841), .ZN(n19851) );
  AOI22_X1 U21861 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19851), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n11057), .ZN(n19825) );
  OAI21_X1 U21862 ( .B1(n21470), .B2(n19839), .A(n19825), .ZN(P1_U3205) );
  INV_X1 U21863 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21472) );
  AOI22_X1 U21864 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19849), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n11057), .ZN(n19826) );
  OAI21_X1 U21865 ( .B1(n21472), .B2(n19841), .A(n19826), .ZN(P1_U3206) );
  AOI222_X1 U21866 ( .A1(n19837), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n19849), .ZN(n19827) );
  INV_X1 U21867 ( .A(n19827), .ZN(P1_U3207) );
  AOI222_X1 U21868 ( .A1(n19849), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n19851), .ZN(n19828) );
  INV_X1 U21869 ( .A(n19828), .ZN(P1_U3208) );
  AOI222_X1 U21870 ( .A1(n19849), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n19851), .ZN(n19829) );
  INV_X1 U21871 ( .A(n19829), .ZN(P1_U3209) );
  AOI22_X1 U21872 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19851), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n11057), .ZN(n19830) );
  OAI21_X1 U21873 ( .B1(n21218), .B2(n19839), .A(n19830), .ZN(P1_U3210) );
  AOI22_X1 U21874 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n19852), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n11057), .ZN(n19831) );
  OAI21_X1 U21875 ( .B1(n19832), .B2(n19841), .A(n19831), .ZN(P1_U3211) );
  AOI222_X1 U21876 ( .A1(n19849), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n19851), .ZN(n19833) );
  INV_X1 U21877 ( .A(n19833), .ZN(P1_U3212) );
  AOI222_X1 U21878 ( .A1(n19851), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n19849), .ZN(n19834) );
  INV_X1 U21879 ( .A(n19834), .ZN(P1_U3213) );
  AOI222_X1 U21880 ( .A1(n19852), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n19851), .ZN(n19835) );
  INV_X1 U21881 ( .A(n19835), .ZN(P1_U3214) );
  AOI222_X1 U21882 ( .A1(n19852), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n19851), .ZN(n19836) );
  INV_X1 U21883 ( .A(n19836), .ZN(P1_U3215) );
  AOI22_X1 U21884 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19837), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n11057), .ZN(n19838) );
  OAI21_X1 U21885 ( .B1(n15655), .B2(n19839), .A(n19838), .ZN(P1_U3216) );
  AOI22_X1 U21886 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19849), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n11057), .ZN(n19840) );
  OAI21_X1 U21887 ( .B1(n21561), .B2(n19841), .A(n19840), .ZN(P1_U3217) );
  AOI222_X1 U21888 ( .A1(n19852), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n19851), .ZN(n19842) );
  INV_X1 U21889 ( .A(n19842), .ZN(P1_U3218) );
  AOI222_X1 U21890 ( .A1(n19852), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19851), .ZN(n19843) );
  INV_X1 U21891 ( .A(n19843), .ZN(P1_U3219) );
  AOI222_X1 U21892 ( .A1(n19852), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n19851), .ZN(n19844) );
  INV_X1 U21893 ( .A(n19844), .ZN(P1_U3220) );
  AOI222_X1 U21894 ( .A1(n19852), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n19851), .ZN(n19845) );
  INV_X1 U21895 ( .A(n19845), .ZN(P1_U3221) );
  AOI222_X1 U21896 ( .A1(n19849), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19851), .ZN(n19846) );
  INV_X1 U21897 ( .A(n19846), .ZN(P1_U3222) );
  AOI222_X1 U21898 ( .A1(n19851), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19849), .ZN(n19847) );
  INV_X1 U21899 ( .A(n19847), .ZN(P1_U3223) );
  AOI222_X1 U21900 ( .A1(n19852), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n19851), .ZN(n19848) );
  INV_X1 U21901 ( .A(n19848), .ZN(P1_U3224) );
  AOI222_X1 U21902 ( .A1(n19851), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n19849), .ZN(n19850) );
  INV_X1 U21903 ( .A(n19850), .ZN(P1_U3225) );
  AOI222_X1 U21904 ( .A1(n19852), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n11057), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n19851), .ZN(n19853) );
  INV_X1 U21905 ( .A(n19853), .ZN(P1_U3226) );
  OAI22_X1 U21906 ( .A1(n11057), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22319), .ZN(n19854) );
  INV_X1 U21907 ( .A(n19854), .ZN(P1_U3458) );
  NOR4_X1 U21908 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19858) );
  NOR4_X1 U21909 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19857) );
  NOR4_X1 U21910 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19856) );
  NOR4_X1 U21911 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19855) );
  NAND4_X1 U21912 ( .A1(n19858), .A2(n19857), .A3(n19856), .A4(n19855), .ZN(
        n19864) );
  NOR4_X1 U21913 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19862) );
  AOI211_X1 U21914 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19861) );
  NOR4_X1 U21915 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19860) );
  NOR4_X1 U21916 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19859) );
  NAND4_X1 U21917 ( .A1(n19862), .A2(n19861), .A3(n19860), .A4(n19859), .ZN(
        n19863) );
  NOR2_X1 U21918 ( .A1(n19864), .A2(n19863), .ZN(n19877) );
  NAND2_X1 U21919 ( .A1(n19877), .A2(n13784), .ZN(n19878) );
  INV_X1 U21920 ( .A(n19877), .ZN(n19874) );
  NOR4_X1 U21921 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .A4(
        n19874), .ZN(n19872) );
  AOI21_X1 U21922 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n19874), .A(n19872), 
        .ZN(n19865) );
  OAI21_X1 U21923 ( .B1(P1_DATAWIDTH_REG_1__SCAN_IN), .B2(n19878), .A(n19865), 
        .ZN(P1_U2808) );
  OAI22_X1 U21924 ( .A1(n11057), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22319), .ZN(n19866) );
  INV_X1 U21925 ( .A(n19866), .ZN(P1_U3459) );
  NAND3_X1 U21926 ( .A1(n19877), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U21927 ( .B1(n19877), .B2(n19868), .A(n19867), .ZN(n19870) );
  AOI211_X1 U21928 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(n19878), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19869) );
  OR2_X1 U21929 ( .A1(n19870), .A2(n19869), .ZN(P1_U3481) );
  OAI22_X1 U21930 ( .A1(n11057), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22319), .ZN(n19871) );
  INV_X1 U21931 ( .A(n19871), .ZN(P1_U3460) );
  INV_X1 U21932 ( .A(n19872), .ZN(n19873) );
  OAI221_X1 U21933 ( .B1(n19877), .B2(n19875), .C1(n19874), .C2(n13784), .A(
        n19873), .ZN(P1_U2807) );
  OAI22_X1 U21934 ( .A1(n11057), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22319), .ZN(n19876) );
  INV_X1 U21935 ( .A(n19876), .ZN(P1_U3461) );
  OAI22_X1 U21936 ( .A1(n19878), .A2(P1_REIP_REG_0__SCAN_IN), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n19877), .ZN(n19879) );
  INV_X1 U21937 ( .A(n19879), .ZN(P1_U3482) );
  INV_X1 U21938 ( .A(n19880), .ZN(n19881) );
  XNOR2_X1 U21939 ( .A(n19884), .B(n19881), .ZN(n21437) );
  AOI22_X1 U21940 ( .A1(n21441), .A2(n19889), .B1(n19888), .B2(n21437), .ZN(
        n19882) );
  OAI21_X1 U21941 ( .B1(n19892), .B2(n19883), .A(n19882), .ZN(P1_U2866) );
  INV_X1 U21942 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19891) );
  INV_X1 U21943 ( .A(n19884), .ZN(n19885) );
  AOI21_X1 U21944 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(n21419) );
  AOI22_X1 U21945 ( .A1(n21429), .A2(n19889), .B1(n19888), .B2(n21419), .ZN(
        n19890) );
  OAI21_X1 U21946 ( .B1(n19892), .B2(n19891), .A(n19890), .ZN(P1_U2867) );
  AOI22_X1 U21947 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U21948 ( .B1(n19895), .B2(n19894), .A(n19893), .ZN(n19896) );
  INV_X1 U21949 ( .A(n19896), .ZN(n21246) );
  AOI22_X1 U21950 ( .A1(n21246), .A2(n19961), .B1(n19952), .B2(n21404), .ZN(
        n19897) );
  OAI211_X1 U21951 ( .C1(n19964), .C2(n21418), .A(n19898), .B(n19897), .ZN(
        P1_U2995) );
  AOI22_X1 U21952 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U21953 ( .B1(n19899), .B2(n19901), .A(n19900), .ZN(n19902) );
  INV_X1 U21954 ( .A(n19902), .ZN(n21271) );
  AOI22_X1 U21955 ( .A1(n21271), .A2(n19961), .B1(n19952), .B2(n21429), .ZN(
        n19903) );
  OAI211_X1 U21956 ( .C1(n19964), .C2(n21422), .A(n19904), .B(n19903), .ZN(
        P1_U2994) );
  AOI22_X1 U21957 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n19910) );
  OAI21_X1 U21958 ( .B1(n19907), .B2(n19906), .A(n19905), .ZN(n19908) );
  INV_X1 U21959 ( .A(n19908), .ZN(n21259) );
  AOI22_X1 U21960 ( .A1(n21259), .A2(n19961), .B1(n19952), .B2(n21441), .ZN(
        n19909) );
  OAI211_X1 U21961 ( .C1(n19964), .C2(n21444), .A(n19910), .B(n19909), .ZN(
        P1_U2993) );
  AOI22_X1 U21962 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n19916) );
  OAI21_X1 U21963 ( .B1(n19913), .B2(n19912), .A(n19911), .ZN(n21279) );
  INV_X1 U21964 ( .A(n21279), .ZN(n19914) );
  AOI22_X1 U21965 ( .A1(n19914), .A2(n19961), .B1(n19952), .B2(n21455), .ZN(
        n19915) );
  OAI211_X1 U21966 ( .C1(n19964), .C2(n21449), .A(n19916), .B(n19915), .ZN(
        P1_U2992) );
  INV_X1 U21967 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19922) );
  NOR2_X1 U21968 ( .A1(n15692), .A2(n13221), .ZN(n19918) );
  MUX2_X1 U21969 ( .A(n19918), .B(n13221), .S(n19917), .Z(n19919) );
  XNOR2_X1 U21970 ( .A(n19919), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n21329) );
  OAI22_X1 U21971 ( .A1(n21329), .A2(n21610), .B1(n19964), .B2(n21480), .ZN(
        n19920) );
  AOI21_X1 U21972 ( .B1(n19952), .B2(n21477), .A(n19920), .ZN(n19921) );
  NAND2_X1 U21973 ( .A1(n13790), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n21324) );
  OAI211_X1 U21974 ( .C1(n19923), .C2(n19922), .A(n19921), .B(n21324), .ZN(
        P1_U2988) );
  INV_X1 U21975 ( .A(n19924), .ZN(n19929) );
  OAI21_X1 U21976 ( .B1(n13214), .B2(n13221), .A(n19925), .ZN(n19928) );
  INV_X1 U21977 ( .A(n19926), .ZN(n19927) );
  AOI21_X1 U21978 ( .B1(n19929), .B2(n19928), .A(n19927), .ZN(n21323) );
  AOI22_X1 U21979 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U21980 ( .A1(n19946), .A2(n21490), .B1(n19952), .B2(n19930), .ZN(
        n19931) );
  OAI211_X1 U21981 ( .C1(n21323), .C2(n21610), .A(n19932), .B(n19931), .ZN(
        P1_U2987) );
  INV_X1 U21982 ( .A(n19933), .ZN(n19934) );
  OAI21_X1 U21983 ( .B1(n13217), .B2(n13221), .A(n19934), .ZN(n19936) );
  AOI21_X1 U21984 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(n21341) );
  AOI22_X1 U21985 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n19939) );
  AOI22_X1 U21986 ( .A1(n21502), .A2(n19952), .B1(n19946), .B2(n21501), .ZN(
        n19938) );
  OAI211_X1 U21987 ( .C1(n21341), .C2(n21610), .A(n19939), .B(n19938), .ZN(
        P1_U2984) );
  NOR2_X1 U21988 ( .A1(n13221), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19943) );
  NOR2_X1 U21989 ( .A1(n19941), .A2(n19940), .ZN(n19942) );
  MUX2_X1 U21990 ( .A(n13221), .B(n19943), .S(n19942), .Z(n19944) );
  XNOR2_X1 U21991 ( .A(n19944), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21354) );
  AOI22_X1 U21992 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U21993 ( .A1(n19947), .A2(n19952), .B1(n19946), .B2(n19945), .ZN(
        n19948) );
  OAI211_X1 U21994 ( .C1(n21610), .C2(n21354), .A(n19949), .B(n19948), .ZN(
        P1_U2982) );
  AOI22_X1 U21995 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n19954) );
  XNOR2_X1 U21996 ( .A(n13221), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n19950) );
  XNOR2_X1 U21997 ( .A(n19951), .B(n19950), .ZN(n21375) );
  AOI22_X1 U21998 ( .A1(n21375), .A2(n19961), .B1(n19952), .B2(n21540), .ZN(
        n19953) );
  OAI211_X1 U21999 ( .C1(n19964), .C2(n21536), .A(n19954), .B(n19953), .ZN(
        P1_U2980) );
  AOI22_X1 U22000 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19955), .B1(
        n13790), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n19963) );
  NOR2_X1 U22001 ( .A1(n13221), .A2(n19958), .ZN(n19957) );
  AOI22_X1 U22002 ( .A1(n21380), .A2(n19961), .B1(n19952), .B2(n19960), .ZN(
        n19962) );
  OAI211_X1 U22003 ( .C1(n19964), .C2(n21552), .A(n19963), .B(n19962), .ZN(
        P1_U2978) );
  AND2_X1 U22004 ( .A1(n19966), .A2(n19965), .ZN(n19969) );
  OAI22_X1 U22005 ( .A1(n19969), .A2(n19968), .B1(n21614), .B2(n19967), .ZN(
        P1_U2803) );
  INV_X1 U22006 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n19971) );
  OAI21_X1 U22007 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n12962), .A(n13264), 
        .ZN(n19970) );
  AOI22_X1 U22008 ( .A1(n22319), .A2(P1_CODEFETCH_REG_SCAN_IN), .B1(n19971), 
        .B2(n19970), .ZN(P1_U2804) );
  AOI22_X1 U22009 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10962), .ZN(n19973) );
  OAI21_X1 U22010 ( .B1(n13751), .B2(n20013), .A(n19973), .ZN(U247) );
  AOI22_X1 U22011 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10962), .ZN(n19974) );
  OAI21_X1 U22012 ( .B1(n13812), .B2(n20013), .A(n19974), .ZN(U246) );
  INV_X1 U22013 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U22014 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10962), .ZN(n19975) );
  OAI21_X1 U22015 ( .B1(n19976), .B2(n20013), .A(n19975), .ZN(U245) );
  AOI22_X1 U22016 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10962), .ZN(n19977) );
  OAI21_X1 U22017 ( .B1(n14173), .B2(n20013), .A(n19977), .ZN(U244) );
  AOI22_X1 U22018 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10962), .ZN(n19978) );
  OAI21_X1 U22019 ( .B1(n14202), .B2(n20013), .A(n19978), .ZN(U243) );
  AOI22_X1 U22020 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10962), .ZN(n19979) );
  OAI21_X1 U22021 ( .B1(n16186), .B2(n20013), .A(n19979), .ZN(U242) );
  AOI22_X1 U22022 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10962), .ZN(n19980) );
  OAI21_X1 U22023 ( .B1(n13796), .B2(n20013), .A(n19980), .ZN(U241) );
  AOI22_X1 U22024 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10962), .ZN(n19981) );
  OAI21_X1 U22025 ( .B1(n13818), .B2(n20013), .A(n19981), .ZN(U240) );
  AOI22_X1 U22026 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10962), .ZN(n19982) );
  OAI21_X1 U22027 ( .B1(n19983), .B2(n20013), .A(n19982), .ZN(U239) );
  AOI22_X1 U22028 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10962), .ZN(n19984) );
  OAI21_X1 U22029 ( .B1(n19985), .B2(n20013), .A(n19984), .ZN(U238) );
  AOI22_X1 U22030 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10962), .ZN(n19986) );
  OAI21_X1 U22031 ( .B1(n19987), .B2(n20013), .A(n19986), .ZN(U237) );
  AOI22_X1 U22032 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10962), .ZN(n19988) );
  OAI21_X1 U22033 ( .B1(n19989), .B2(n20013), .A(n19988), .ZN(U236) );
  AOI22_X1 U22034 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10962), .ZN(n19990) );
  OAI21_X1 U22035 ( .B1(n14123), .B2(n20013), .A(n19990), .ZN(U235) );
  AOI22_X1 U22036 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10962), .ZN(n19991) );
  OAI21_X1 U22037 ( .B1(n19992), .B2(n20013), .A(n19991), .ZN(U234) );
  AOI22_X1 U22038 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10962), .ZN(n19993) );
  OAI21_X1 U22039 ( .B1(n19994), .B2(n20013), .A(n19993), .ZN(U233) );
  AOI22_X1 U22040 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10962), .ZN(n19995) );
  OAI21_X1 U22041 ( .B1(n13666), .B2(n20013), .A(n19995), .ZN(U232) );
  INV_X1 U22042 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21727) );
  AOI22_X1 U22043 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10962), .ZN(n19996) );
  OAI21_X1 U22044 ( .B1(n21727), .B2(n20013), .A(n19996), .ZN(U231) );
  INV_X1 U22045 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21917) );
  AOI22_X1 U22046 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10962), .ZN(n19997) );
  OAI21_X1 U22047 ( .B1(n21917), .B2(n20013), .A(n19997), .ZN(U230) );
  AOI22_X1 U22048 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10962), .ZN(n19998) );
  OAI21_X1 U22049 ( .B1(n21963), .B2(n20013), .A(n19998), .ZN(U229) );
  INV_X1 U22050 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n22011) );
  AOI22_X1 U22051 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10962), .ZN(n19999) );
  OAI21_X1 U22052 ( .B1(n22011), .B2(n20013), .A(n19999), .ZN(U228) );
  AOI22_X1 U22053 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10962), .ZN(n20000) );
  OAI21_X1 U22054 ( .B1(n22058), .B2(n20013), .A(n20000), .ZN(U227) );
  INV_X1 U22055 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n22106) );
  AOI22_X1 U22056 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10962), .ZN(n20001) );
  OAI21_X1 U22057 ( .B1(n22106), .B2(n20013), .A(n20001), .ZN(U226) );
  AOI22_X1 U22058 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10962), .ZN(n20002) );
  OAI21_X1 U22059 ( .B1(n22153), .B2(n20013), .A(n20002), .ZN(U225) );
  INV_X1 U22060 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22208) );
  AOI22_X1 U22061 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10962), .ZN(n20003) );
  OAI21_X1 U22062 ( .B1(n22208), .B2(n20013), .A(n20003), .ZN(U224) );
  AOI22_X1 U22063 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10962), .ZN(n20004) );
  OAI21_X1 U22064 ( .B1(n21714), .B2(n20013), .A(n20004), .ZN(U223) );
  INV_X1 U22065 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n21914) );
  AOI22_X1 U22066 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10962), .ZN(n20005) );
  OAI21_X1 U22067 ( .B1(n21914), .B2(n20013), .A(n20005), .ZN(U222) );
  AOI22_X1 U22068 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10962), .ZN(n20007) );
  OAI21_X1 U22069 ( .B1(n21961), .B2(n20013), .A(n20007), .ZN(U221) );
  INV_X1 U22070 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n22009) );
  AOI22_X1 U22071 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10962), .ZN(n20008) );
  OAI21_X1 U22072 ( .B1(n22009), .B2(n20013), .A(n20008), .ZN(U220) );
  INV_X1 U22073 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n22056) );
  AOI22_X1 U22074 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10962), .ZN(n20009) );
  OAI21_X1 U22075 ( .B1(n22056), .B2(n20013), .A(n20009), .ZN(U219) );
  INV_X1 U22076 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n22103) );
  AOI22_X1 U22077 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10962), .ZN(n20010) );
  OAI21_X1 U22078 ( .B1(n22103), .B2(n20013), .A(n20010), .ZN(U218) );
  AOI22_X1 U22079 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20006), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10962), .ZN(n20011) );
  OAI21_X1 U22080 ( .B1(n22151), .B2(n20013), .A(n20011), .ZN(U217) );
  OAI222_X1 U22081 ( .A1(U212), .A2(n20014), .B1(n20013), .B2(n22201), .C1(
        U214), .C2(n20012), .ZN(U216) );
  AOI22_X1 U22082 ( .A1(n22319), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20015), 
        .B2(n11057), .ZN(P1_U3483) );
  AOI21_X1 U22083 ( .B1(n21649), .B2(n21177), .A(n20016), .ZN(n20017) );
  OAI21_X1 U22084 ( .B1(n20018), .B2(n21164), .A(n20017), .ZN(n20019) );
  INV_X1 U22085 ( .A(n20019), .ZN(n20026) );
  AOI21_X1 U22086 ( .B1(n20084), .B2(n21644), .A(n20085), .ZN(n20020) );
  OAI211_X1 U22087 ( .C1(n20021), .C2(n20020), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n21649), .ZN(n20023) );
  INV_X1 U22088 ( .A(n20022), .ZN(n21179) );
  AOI21_X1 U22089 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20023), .A(n21179), 
        .ZN(n20025) );
  NAND2_X1 U22090 ( .A1(n20026), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20024) );
  OAI21_X1 U22091 ( .B1(n20026), .B2(n20025), .A(n20024), .ZN(P3_U3296) );
  NOR2_X1 U22092 ( .A1(n21165), .A2(n20027), .ZN(n20030) );
  AOI22_X1 U22093 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20075), .ZN(n20031) );
  OAI21_X1 U22094 ( .B1(n20032), .B2(n20080), .A(n20031), .ZN(P3_U2768) );
  AOI22_X1 U22095 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20075), .ZN(n20033) );
  OAI21_X1 U22096 ( .B1(n20584), .B2(n20080), .A(n20033), .ZN(P3_U2769) );
  AOI22_X1 U22097 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20075), .ZN(n20034) );
  OAI21_X1 U22098 ( .B1(n20035), .B2(n20080), .A(n20034), .ZN(P3_U2770) );
  AOI22_X1 U22099 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20075), .ZN(n20036) );
  OAI21_X1 U22100 ( .B1(n20607), .B2(n20080), .A(n20036), .ZN(P3_U2771) );
  AOI22_X1 U22101 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20075), .ZN(n20037) );
  OAI21_X1 U22102 ( .B1(n20038), .B2(n20080), .A(n20037), .ZN(P3_U2772) );
  AOI22_X1 U22103 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20075), .ZN(n20039) );
  OAI21_X1 U22104 ( .B1(n20591), .B2(n20080), .A(n20039), .ZN(P3_U2773) );
  AOI22_X1 U22105 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20075), .ZN(n20040) );
  OAI21_X1 U22106 ( .B1(n20041), .B2(n20080), .A(n20040), .ZN(P3_U2774) );
  AOI22_X1 U22107 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20075), .ZN(n20042) );
  OAI21_X1 U22108 ( .B1(n20043), .B2(n20080), .A(n20042), .ZN(P3_U2775) );
  AOI22_X1 U22109 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20044) );
  OAI21_X1 U22110 ( .B1(n20045), .B2(n20080), .A(n20044), .ZN(P3_U2776) );
  AOI22_X1 U22111 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20046) );
  OAI21_X1 U22112 ( .B1(n20626), .B2(n20080), .A(n20046), .ZN(P3_U2777) );
  AOI22_X1 U22113 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20075), .ZN(n20047) );
  OAI21_X1 U22114 ( .B1(n20048), .B2(n20080), .A(n20047), .ZN(P3_U2778) );
  AOI22_X1 U22115 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20075), .ZN(n20049) );
  OAI21_X1 U22116 ( .B1(n20655), .B2(n20080), .A(n20049), .ZN(P3_U2779) );
  AOI22_X1 U22117 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20075), .ZN(n20050) );
  OAI21_X1 U22118 ( .B1(n20051), .B2(n20080), .A(n20050), .ZN(P3_U2780) );
  AOI22_X1 U22119 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20075), .ZN(n20052) );
  OAI21_X1 U22120 ( .B1(n20643), .B2(n20080), .A(n20052), .ZN(P3_U2781) );
  AOI22_X1 U22121 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20078), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20053) );
  OAI21_X1 U22122 ( .B1(n20054), .B2(n20080), .A(n20053), .ZN(P3_U2782) );
  AOI22_X1 U22123 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20075), .ZN(n20055) );
  OAI21_X1 U22124 ( .B1(n20708), .B2(n20080), .A(n20055), .ZN(P3_U2783) );
  AOI22_X1 U22125 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20075), .ZN(n20056) );
  OAI21_X1 U22126 ( .B1(n20057), .B2(n20080), .A(n20056), .ZN(P3_U2784) );
  AOI22_X1 U22127 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20075), .ZN(n20058) );
  OAI21_X1 U22128 ( .B1(n20576), .B2(n20080), .A(n20058), .ZN(P3_U2785) );
  AOI22_X1 U22129 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20077), .ZN(n20059) );
  OAI21_X1 U22130 ( .B1(n20547), .B2(n20080), .A(n20059), .ZN(P3_U2786) );
  AOI22_X1 U22131 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20075), .ZN(n20060) );
  OAI21_X1 U22132 ( .B1(n20525), .B2(n20080), .A(n20060), .ZN(P3_U2787) );
  AOI22_X1 U22133 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20077), .ZN(n20061) );
  OAI21_X1 U22134 ( .B1(n20548), .B2(n20080), .A(n20061), .ZN(P3_U2788) );
  AOI22_X1 U22135 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20077), .ZN(n20062) );
  OAI21_X1 U22136 ( .B1(n20526), .B2(n20080), .A(n20062), .ZN(P3_U2789) );
  AOI22_X1 U22137 ( .A1(n20071), .A2(BUF2_REG_7__SCAN_IN), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20077), .ZN(n20063) );
  OAI21_X1 U22138 ( .B1(n20064), .B2(n20080), .A(n20063), .ZN(P3_U2790) );
  AOI22_X1 U22139 ( .A1(n20078), .A2(BUF2_REG_8__SCAN_IN), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20077), .ZN(n20065) );
  OAI21_X1 U22140 ( .B1(n20066), .B2(n20080), .A(n20065), .ZN(P3_U2791) );
  AOI22_X1 U22141 ( .A1(n20071), .A2(BUF2_REG_9__SCAN_IN), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20077), .ZN(n20067) );
  OAI21_X1 U22142 ( .B1(n20068), .B2(n20080), .A(n20067), .ZN(P3_U2792) );
  AOI22_X1 U22143 ( .A1(n20071), .A2(BUF2_REG_10__SCAN_IN), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20077), .ZN(n20069) );
  OAI21_X1 U22144 ( .B1(n20580), .B2(n20080), .A(n20069), .ZN(P3_U2793) );
  AOI22_X1 U22145 ( .A1(n20071), .A2(BUF2_REG_11__SCAN_IN), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20077), .ZN(n20070) );
  OAI21_X1 U22146 ( .B1(n20536), .B2(n20080), .A(n20070), .ZN(P3_U2794) );
  AOI22_X1 U22147 ( .A1(n20071), .A2(BUF2_REG_12__SCAN_IN), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20077), .ZN(n20072) );
  OAI21_X1 U22148 ( .B1(n20582), .B2(n20080), .A(n20072), .ZN(P3_U2795) );
  AOI22_X1 U22149 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20077), .ZN(n20073) );
  OAI21_X1 U22150 ( .B1(n20074), .B2(n20080), .A(n20073), .ZN(P3_U2796) );
  AOI22_X1 U22151 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20076) );
  OAI21_X1 U22152 ( .B1(n20683), .B2(n20080), .A(n20076), .ZN(P3_U2797) );
  AOI22_X1 U22153 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20078), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20077), .ZN(n20079) );
  OAI21_X1 U22154 ( .B1(n20687), .B2(n20080), .A(n20079), .ZN(P3_U2798) );
  NAND4_X1 U22155 ( .A1(n20082), .A2(n20081), .A3(n21644), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21173) );
  NOR2_X1 U22156 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21173), .ZN(
        n20193) );
  NOR2_X1 U22157 ( .A1(n20281), .A2(n20193), .ZN(n20251) );
  NOR2_X1 U22158 ( .A1(n20482), .A2(n21173), .ZN(n20495) );
  NAND2_X1 U22159 ( .A1(n21169), .A2(n20083), .ZN(n21185) );
  AOI21_X1 U22160 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20495), .A(
        n20409), .ZN(n20095) );
  INV_X1 U22161 ( .A(n21649), .ZN(n21687) );
  AOI211_X1 U22162 ( .C1(n20085), .C2(n20084), .A(n21687), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n20086) );
  INV_X1 U22163 ( .A(n20086), .ZN(n21166) );
  AOI211_X4 U22164 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20520), .A(n20086), .B(
        n20088), .ZN(n20516) );
  OAI22_X1 U22165 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20468), .B1(n20498), 
        .B2(n20098), .ZN(n20093) );
  NAND2_X1 U22166 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20520), .ZN(n20087) );
  AOI211_X4 U22167 ( .C1(n21649), .C2(n21644), .A(n20088), .B(n20087), .ZN(
        n20515) );
  NAND2_X1 U22168 ( .A1(n20089), .A2(n20720), .ZN(n20715) );
  NOR2_X1 U22169 ( .A1(n20521), .A2(n20090), .ZN(n20512) );
  INV_X1 U22170 ( .A(n20512), .ZN(n20124) );
  OAI22_X1 U22171 ( .A1(n20490), .A2(n20091), .B1(n20715), .B2(n20124), .ZN(
        n20092) );
  AOI211_X1 U22172 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n20431), .A(n20093), .B(
        n20092), .ZN(n20094) );
  OAI221_X1 U22173 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20251), .C1(
        n20096), .C2(n20095), .A(n20094), .ZN(P3_U2670) );
  AOI22_X1 U22174 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U22175 ( .B1(n20742), .B2(n21143), .A(n20729), .ZN(n20725) );
  AOI22_X1 U22176 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n20431), .B1(n20512), 
        .B2(n20725), .ZN(n20106) );
  INV_X1 U22177 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20305) );
  NAND2_X1 U22178 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20305), .ZN(
        n20212) );
  OAI21_X1 U22179 ( .B1(n20097), .B2(n20212), .A(n20495), .ZN(n20122) );
  AOI21_X1 U22180 ( .B1(n20103), .B2(n20212), .A(n20122), .ZN(n20102) );
  NAND2_X1 U22181 ( .A1(n20099), .A2(n20098), .ZN(n20100) );
  NOR3_X1 U22182 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20113) );
  AOI211_X1 U22183 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20100), .A(n20113), .B(
        n20490), .ZN(n20101) );
  AOI211_X1 U22184 ( .C1(n20281), .C2(n20103), .A(n20102), .B(n20101), .ZN(
        n20105) );
  NAND2_X1 U22185 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20111) );
  OAI211_X1 U22186 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20445), .B(n20111), .ZN(n20104) );
  NAND4_X1 U22187 ( .A1(n20107), .A2(n20106), .A3(n20105), .A4(n20104), .ZN(
        P3_U2669) );
  INV_X1 U22188 ( .A(n20121), .ZN(n20123) );
  AOI21_X1 U22189 ( .B1(n20108), .B2(n20193), .A(n20281), .ZN(n20120) );
  OAI21_X1 U22190 ( .B1(n11406), .B2(n21143), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20749) );
  NAND2_X1 U22191 ( .A1(n20109), .A2(n20749), .ZN(n20743) );
  NOR2_X1 U22192 ( .A1(n17457), .A2(n20743), .ZN(n20737) );
  NAND3_X1 U22193 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20138) );
  NAND2_X1 U22194 ( .A1(n20445), .A2(n20138), .ZN(n20110) );
  OAI22_X1 U22195 ( .A1(n20737), .A2(n20124), .B1(n20111), .B2(n20110), .ZN(
        n20118) );
  AOI21_X1 U22196 ( .B1(n20445), .B2(n20138), .A(n20431), .ZN(n20137) );
  NAND2_X1 U22197 ( .A1(n20516), .A2(P3_EBX_REG_3__SCAN_IN), .ZN(n20115) );
  NAND2_X1 U22198 ( .A1(n20113), .A2(n20112), .ZN(n20126) );
  OAI211_X1 U22199 ( .C1(n20113), .C2(n20112), .A(n20515), .B(n20126), .ZN(
        n20114) );
  OAI211_X1 U22200 ( .C1(n20137), .C2(n20116), .A(n20115), .B(n20114), .ZN(
        n20117) );
  AOI211_X1 U22201 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n20409), .A(
        n20118), .B(n20117), .ZN(n20119) );
  OAI221_X1 U22202 ( .B1(n20123), .B2(n20122), .C1(n20121), .C2(n20120), .A(
        n20119), .ZN(P3_U2668) );
  AOI21_X1 U22203 ( .B1(n11547), .B2(n21139), .A(n20124), .ZN(n20125) );
  AOI211_X1 U22204 ( .C1(n20516), .C2(P3_EBX_REG_4__SCAN_IN), .A(n10958), .B(
        n20125), .ZN(n20136) );
  NOR2_X1 U22205 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20126), .ZN(n20147) );
  AOI211_X1 U22206 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20126), .A(n20147), .B(
        n20490), .ZN(n20134) );
  AOI21_X1 U22207 ( .B1(n20127), .B2(n20193), .A(n20281), .ZN(n20132) );
  INV_X1 U22208 ( .A(n20128), .ZN(n20140) );
  OAI211_X1 U22209 ( .C1(n20212), .C2(n20140), .A(n20495), .B(n20131), .ZN(
        n20130) );
  OR3_X1 U22210 ( .A1(n20468), .A2(n20138), .A3(P3_REIP_REG_4__SCAN_IN), .ZN(
        n20129) );
  OAI211_X1 U22211 ( .C1(n20132), .C2(n20131), .A(n20130), .B(n20129), .ZN(
        n20133) );
  AOI211_X1 U22212 ( .C1(n20409), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20134), .B(n20133), .ZN(n20135) );
  OAI211_X1 U22213 ( .C1(n20137), .C2(n20825), .A(n20136), .B(n20135), .ZN(
        P3_U2667) );
  NOR2_X1 U22214 ( .A1(n20825), .A2(n20138), .ZN(n20139) );
  AOI21_X1 U22215 ( .B1(n20445), .B2(n20139), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n20144) );
  NAND2_X1 U22216 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20139), .ZN(n20164) );
  AOI21_X1 U22217 ( .B1(n20445), .B2(n20164), .A(n20431), .ZN(n20163) );
  OAI21_X1 U22218 ( .B1(n20140), .B2(n20212), .A(n20387), .ZN(n20141) );
  XOR2_X1 U22219 ( .A(n20142), .B(n20141), .Z(n20143) );
  OAI22_X1 U22220 ( .A1(n20144), .A2(n20163), .B1(n21173), .B2(n20143), .ZN(
        n20145) );
  AOI211_X1 U22221 ( .C1(n20516), .C2(P3_EBX_REG_5__SCAN_IN), .A(n10958), .B(
        n20145), .ZN(n20149) );
  NAND2_X1 U22222 ( .A1(n20147), .A2(n20146), .ZN(n20151) );
  OAI211_X1 U22223 ( .C1(n20147), .C2(n20146), .A(n20515), .B(n20151), .ZN(
        n20148) );
  OAI211_X1 U22224 ( .C1(n20500), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        P3_U2666) );
  NOR2_X1 U22225 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20151), .ZN(n20171) );
  AOI211_X1 U22226 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20151), .A(n20171), .B(
        n20490), .ZN(n20157) );
  AOI21_X1 U22227 ( .B1(n20387), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20251), .ZN(n20154) );
  OAI21_X1 U22228 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20175), .A(
        n20387), .ZN(n20160) );
  OAI21_X1 U22229 ( .B1(n21173), .B2(n20160), .A(n20153), .ZN(n20152) );
  OAI21_X1 U22230 ( .B1(n20154), .B2(n20153), .A(n20152), .ZN(n20155) );
  OAI211_X1 U22231 ( .C1(n20834), .C2(n20163), .A(n20155), .B(n21105), .ZN(
        n20156) );
  AOI211_X1 U22232 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20516), .A(n20157), .B(
        n20156), .ZN(n20158) );
  OR3_X1 U22233 ( .A1(n20468), .A2(n20164), .A3(P3_REIP_REG_6__SCAN_IN), .ZN(
        n20162) );
  OAI211_X1 U22234 ( .C1(n20500), .C2(n20159), .A(n20158), .B(n20162), .ZN(
        P3_U2665) );
  INV_X1 U22235 ( .A(n21173), .ZN(n20488) );
  XNOR2_X1 U22236 ( .A(n20161), .B(n20160), .ZN(n20169) );
  AOI21_X1 U22237 ( .B1(n20163), .B2(n20162), .A(n20165), .ZN(n20168) );
  NOR2_X1 U22238 ( .A1(n20834), .A2(n20164), .ZN(n20181) );
  NAND3_X1 U22239 ( .A1(n20445), .A2(n20181), .A3(n20165), .ZN(n20166) );
  OAI211_X1 U22240 ( .C1(n20498), .C2(n20170), .A(n21105), .B(n20166), .ZN(
        n20167) );
  AOI211_X1 U22241 ( .C1(n20488), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        n20173) );
  NAND2_X1 U22242 ( .A1(n20171), .A2(n20170), .ZN(n20179) );
  OAI211_X1 U22243 ( .C1(n20171), .C2(n20170), .A(n20515), .B(n20179), .ZN(
        n20172) );
  OAI211_X1 U22244 ( .C1(n20500), .C2(n20174), .A(n20173), .B(n20172), .ZN(
        P3_U2664) );
  NOR2_X1 U22245 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20175), .ZN(
        n20176) );
  AOI21_X1 U22246 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20176), .A(
        n20482), .ZN(n20177) );
  XNOR2_X1 U22247 ( .A(n20178), .B(n20177), .ZN(n20189) );
  NOR2_X1 U22248 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20179), .ZN(n20190) );
  AOI211_X1 U22249 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20179), .A(n20190), .B(
        n20490), .ZN(n20180) );
  AOI21_X1 U22250 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n20516), .A(n20180), .ZN(
        n20188) );
  NAND2_X1 U22251 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20181), .ZN(n20184) );
  NOR2_X1 U22252 ( .A1(n20182), .A2(n20184), .ZN(n20206) );
  OAI21_X1 U22253 ( .B1(n20206), .B2(n20468), .A(n20514), .ZN(n20202) );
  OR2_X1 U22254 ( .A1(n20468), .A2(n20206), .ZN(n20183) );
  OAI22_X1 U22255 ( .A1(n20185), .A2(n20500), .B1(n20184), .B2(n20183), .ZN(
        n20186) );
  AOI211_X1 U22256 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n20202), .A(n10958), .B(
        n20186), .ZN(n20187) );
  OAI211_X1 U22257 ( .C1(n21173), .C2(n20189), .A(n20188), .B(n20187), .ZN(
        P3_U2663) );
  NAND2_X1 U22258 ( .A1(n20190), .A2(n20192), .ZN(n20205) );
  OAI211_X1 U22259 ( .C1(n20190), .C2(n20192), .A(n20515), .B(n20205), .ZN(
        n20191) );
  OAI21_X1 U22260 ( .B1(n20192), .B2(n20498), .A(n20191), .ZN(n20198) );
  AOI21_X1 U22261 ( .B1(n20193), .B2(n20201), .A(n20281), .ZN(n20196) );
  OAI211_X1 U22262 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20214), .A(
        n20495), .B(n20195), .ZN(n20194) );
  OAI211_X1 U22263 ( .C1(n20196), .C2(n20195), .A(n21105), .B(n20194), .ZN(
        n20197) );
  AOI211_X1 U22264 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n20202), .A(n20198), .B(
        n20197), .ZN(n20200) );
  NAND3_X1 U22265 ( .A1(n20445), .A2(n20206), .A3(n20199), .ZN(n20203) );
  OAI211_X1 U22266 ( .C1(n20500), .C2(n20201), .A(n20200), .B(n20203), .ZN(
        P3_U2662) );
  INV_X1 U22267 ( .A(n20202), .ZN(n20204) );
  AOI21_X1 U22268 ( .B1(n20204), .B2(n20203), .A(n20222), .ZN(n20211) );
  NOR2_X1 U22269 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20205), .ZN(n20228) );
  AOI211_X1 U22270 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20205), .A(n20228), .B(
        n20490), .ZN(n20210) );
  INV_X1 U22271 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20208) );
  NAND2_X1 U22272 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20206), .ZN(n20221) );
  NAND2_X1 U22273 ( .A1(n20445), .A2(n20222), .ZN(n20207) );
  OAI22_X1 U22274 ( .A1(n20498), .A2(n20208), .B1(n20221), .B2(n20207), .ZN(
        n20209) );
  NOR4_X1 U22275 ( .A1(n10958), .A2(n20211), .A3(n20210), .A4(n20209), .ZN(
        n20219) );
  NOR2_X1 U22276 ( .A1(n20213), .A2(n20212), .ZN(n20237) );
  NOR2_X1 U22277 ( .A1(n20237), .A2(n20482), .ZN(n20225) );
  OR2_X1 U22278 ( .A1(n20214), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20215) );
  AOI21_X1 U22279 ( .B1(n20217), .B2(n20215), .A(n21173), .ZN(n20216) );
  OAI22_X1 U22280 ( .A1(n20217), .A2(n20225), .B1(n20281), .B2(n20216), .ZN(
        n20218) );
  OAI211_X1 U22281 ( .C1(n20500), .C2(n20220), .A(n20219), .B(n20218), .ZN(
        P3_U2661) );
  NOR2_X1 U22282 ( .A1(n20222), .A2(n20221), .ZN(n20236) );
  NAND2_X1 U22283 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20236), .ZN(n20270) );
  AOI21_X1 U22284 ( .B1(n20445), .B2(n20270), .A(n20431), .ZN(n20255) );
  NAND2_X1 U22285 ( .A1(n20445), .A2(n20236), .ZN(n20234) );
  INV_X1 U22286 ( .A(n20224), .ZN(n20226) );
  INV_X1 U22287 ( .A(n20225), .ZN(n20223) );
  OAI221_X1 U22288 ( .B1(n20226), .B2(n20225), .C1(n20224), .C2(n20223), .A(
        n20488), .ZN(n20230) );
  NAND2_X1 U22289 ( .A1(n20228), .A2(n20227), .ZN(n20242) );
  OAI211_X1 U22290 ( .C1(n20228), .C2(n20227), .A(n20515), .B(n20242), .ZN(
        n20229) );
  OAI211_X1 U22291 ( .C1(n20500), .C2(n20231), .A(n20230), .B(n20229), .ZN(
        n20232) );
  AOI211_X1 U22292 ( .C1(n20516), .C2(P3_EBX_REG_11__SCAN_IN), .A(n10958), .B(
        n20232), .ZN(n20233) );
  OAI221_X1 U22293 ( .B1(n20255), .B2(n20235), .C1(n20255), .C2(n20234), .A(
        n20233), .ZN(P3_U2660) );
  NAND3_X1 U22294 ( .A1(n20445), .A2(P3_REIP_REG_11__SCAN_IN), .A3(n20236), 
        .ZN(n20268) );
  NAND2_X1 U22295 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20237), .ZN(
        n20279) );
  NAND2_X1 U22296 ( .A1(n20387), .A2(n20279), .ZN(n20238) );
  INV_X1 U22297 ( .A(n20238), .ZN(n20240) );
  INV_X1 U22298 ( .A(n20241), .ZN(n20239) );
  AOI221_X1 U22299 ( .B1(n20241), .B2(n20240), .C1(n20239), .C2(n20238), .A(
        n21173), .ZN(n20247) );
  NOR2_X1 U22300 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20242), .ZN(n20261) );
  AOI211_X1 U22301 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20242), .A(n20261), .B(
        n20490), .ZN(n20246) );
  OAI22_X1 U22302 ( .A1(n20244), .A2(n20500), .B1(n20498), .B2(n20243), .ZN(
        n20245) );
  NOR4_X1 U22303 ( .A1(n10958), .A2(n20247), .A3(n20246), .A4(n20245), .ZN(
        n20248) );
  OAI221_X1 U22304 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n20268), .C1(n20249), 
        .C2(n20255), .A(n20248), .ZN(P3_U2659) );
  AOI22_X1 U22305 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n20264) );
  OAI21_X1 U22306 ( .B1(n20250), .B2(n20279), .A(n20387), .ZN(n20265) );
  NOR2_X1 U22307 ( .A1(n20265), .A2(n21173), .ZN(n20259) );
  AOI211_X1 U22308 ( .C1(n20387), .C2(n20252), .A(n20251), .B(n20258), .ZN(
        n20257) );
  NAND2_X1 U22309 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20269) );
  OAI21_X1 U22310 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(P3_REIP_REG_12__SCAN_IN), 
        .A(n20269), .ZN(n20253) );
  OAI22_X1 U22311 ( .A1(n20255), .A2(n20254), .B1(n20268), .B2(n20253), .ZN(
        n20256) );
  AOI211_X1 U22312 ( .C1(n20259), .C2(n20258), .A(n20257), .B(n20256), .ZN(
        n20263) );
  NAND2_X1 U22313 ( .A1(n20261), .A2(n20260), .ZN(n20267) );
  OAI211_X1 U22314 ( .C1(n20261), .C2(n20260), .A(n20515), .B(n20267), .ZN(
        n20262) );
  NAND4_X1 U22315 ( .A1(n20264), .A2(n20263), .A3(n21105), .A4(n20262), .ZN(
        P3_U2658) );
  XNOR2_X1 U22316 ( .A(n20266), .B(n20265), .ZN(n20277) );
  NOR2_X1 U22317 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20267), .ZN(n20284) );
  AOI211_X1 U22318 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20267), .A(n20284), .B(
        n20490), .ZN(n20275) );
  NOR2_X1 U22319 ( .A1(n20269), .A2(n20268), .ZN(n20278) );
  NOR3_X1 U22320 ( .A1(n20271), .A2(n20270), .A3(n20269), .ZN(n20314) );
  OAI21_X1 U22321 ( .B1(n20314), .B2(n20468), .A(n20514), .ZN(n20301) );
  OAI21_X1 U22322 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n20278), .A(n20301), 
        .ZN(n20272) );
  OAI211_X1 U22323 ( .C1(n20498), .C2(n20273), .A(n21105), .B(n20272), .ZN(
        n20274) );
  AOI211_X1 U22324 ( .C1(n20409), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20275), .B(n20274), .ZN(n20276) );
  OAI21_X1 U22325 ( .B1(n20277), .B2(n21173), .A(n20276), .ZN(P3_U2657) );
  NAND2_X1 U22326 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20278), .ZN(n20312) );
  AOI22_X1 U22327 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n20290) );
  NOR2_X1 U22328 ( .A1(n20280), .A2(n20279), .ZN(n20282) );
  AOI221_X1 U22329 ( .B1(n20282), .B2(n20488), .C1(n20286), .C2(n20488), .A(
        n20281), .ZN(n20287) );
  NAND2_X1 U22330 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20282), .ZN(
        n20324) );
  NAND2_X1 U22331 ( .A1(n20387), .A2(n20324), .ZN(n20293) );
  NAND2_X1 U22332 ( .A1(n20284), .A2(n20283), .ZN(n20291) );
  OAI211_X1 U22333 ( .C1(n20284), .C2(n20283), .A(n20515), .B(n20291), .ZN(
        n20285) );
  OAI221_X1 U22334 ( .B1(n20287), .B2(n20286), .C1(n20287), .C2(n20293), .A(
        n20285), .ZN(n20288) );
  AOI211_X1 U22335 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n20301), .A(n10958), 
        .B(n20288), .ZN(n20289) );
  OAI211_X1 U22336 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n20312), .A(n20290), 
        .B(n20289), .ZN(P3_U2656) );
  NOR2_X1 U22337 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20291), .ZN(n20309) );
  AOI211_X1 U22338 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20291), .A(n20309), .B(
        n20490), .ZN(n20292) );
  AOI211_X1 U22339 ( .C1(n20516), .C2(P3_EBX_REG_16__SCAN_IN), .A(n10958), .B(
        n20292), .ZN(n20303) );
  INV_X1 U22340 ( .A(n20293), .ZN(n20295) );
  INV_X1 U22341 ( .A(n20296), .ZN(n20294) );
  AOI221_X1 U22342 ( .B1(n20296), .B2(n20295), .C1(n20294), .C2(n20293), .A(
        n21173), .ZN(n20300) );
  AOI221_X1 U22343 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n20298), .C2(n20297), .A(n20312), .ZN(n20299) );
  AOI211_X1 U22344 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n20301), .A(n20300), 
        .B(n20299), .ZN(n20302) );
  OAI211_X1 U22345 ( .C1(n20304), .C2(n20500), .A(n20303), .B(n20302), .ZN(
        P3_U2655) );
  AOI21_X1 U22346 ( .B1(n20306), .B2(n20305), .A(n20482), .ZN(n20307) );
  XOR2_X1 U22347 ( .A(n20308), .B(n20307), .Z(n20320) );
  INV_X1 U22348 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20311) );
  NAND2_X1 U22349 ( .A1(n20309), .A2(n20311), .ZN(n20321) );
  OAI211_X1 U22350 ( .C1(n20309), .C2(n20311), .A(n20515), .B(n20321), .ZN(
        n20310) );
  OAI211_X1 U22351 ( .C1(n20498), .C2(n20311), .A(n21105), .B(n20310), .ZN(
        n20318) );
  NAND2_X1 U22352 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n20313) );
  NOR2_X1 U22353 ( .A1(n20313), .A2(n20312), .ZN(n20316) );
  NAND4_X1 U22354 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20314), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n20336) );
  AOI21_X1 U22355 ( .B1(n20445), .B2(n20336), .A(n20431), .ZN(n20335) );
  INV_X1 U22356 ( .A(n20335), .ZN(n20315) );
  MUX2_X1 U22357 ( .A(n20316), .B(n20315), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n20317) );
  AOI211_X1 U22358 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n20409), .A(
        n20318), .B(n20317), .ZN(n20319) );
  OAI21_X1 U22359 ( .B1(n21173), .B2(n20320), .A(n20319), .ZN(P3_U2654) );
  NOR2_X1 U22360 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20321), .ZN(n20343) );
  AOI211_X1 U22361 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20321), .A(n20343), .B(
        n20490), .ZN(n20323) );
  OR3_X1 U22362 ( .A1(n20468), .A2(n20336), .A3(P3_REIP_REG_18__SCAN_IN), .ZN(
        n20334) );
  OAI211_X1 U22363 ( .C1(n11093), .C2(n20500), .A(n21105), .B(n20334), .ZN(
        n20322) );
  AOI211_X1 U22364 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20516), .A(n20323), .B(
        n20322), .ZN(n20330) );
  NOR2_X1 U22365 ( .A1(n20325), .A2(n20324), .ZN(n20331) );
  OR2_X1 U22366 ( .A1(n20331), .A2(n20482), .ZN(n20327) );
  AOI21_X1 U22367 ( .B1(n20328), .B2(n20327), .A(n21173), .ZN(n20326) );
  OAI21_X1 U22368 ( .B1(n20328), .B2(n20327), .A(n20326), .ZN(n20329) );
  OAI211_X1 U22369 ( .C1(n20335), .C2(n20337), .A(n20330), .B(n20329), .ZN(
        P3_U2653) );
  NAND2_X1 U22370 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20331), .ZN(
        n20354) );
  NAND2_X1 U22371 ( .A1(n20387), .A2(n20354), .ZN(n20332) );
  XNOR2_X1 U22372 ( .A(n20333), .B(n20332), .ZN(n20342) );
  AOI21_X1 U22373 ( .B1(n20335), .B2(n20334), .A(n20338), .ZN(n20341) );
  NOR2_X1 U22374 ( .A1(n20337), .A2(n20336), .ZN(n20347) );
  NAND3_X1 U22375 ( .A1(n20445), .A2(n20347), .A3(n20338), .ZN(n20339) );
  OAI211_X1 U22376 ( .C1(n20355), .C2(n20500), .A(n21105), .B(n20339), .ZN(
        n20340) );
  AOI211_X1 U22377 ( .C1(n20488), .C2(n20342), .A(n20341), .B(n20340), .ZN(
        n20345) );
  NAND2_X1 U22378 ( .A1(n20343), .A2(n20346), .ZN(n20351) );
  OAI211_X1 U22379 ( .C1(n20343), .C2(n20346), .A(n20515), .B(n20351), .ZN(
        n20344) );
  OAI211_X1 U22380 ( .C1(n20346), .C2(n20498), .A(n20345), .B(n20344), .ZN(
        P3_U2652) );
  AOI22_X1 U22381 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n20360) );
  NAND2_X1 U22382 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20347), .ZN(n20350) );
  NOR2_X1 U22383 ( .A1(n20349), .A2(n20350), .ZN(n20377) );
  NOR2_X1 U22384 ( .A1(n20377), .A2(n20468), .ZN(n20348) );
  NOR2_X1 U22385 ( .A1(n20431), .A2(n20348), .ZN(n20376) );
  INV_X1 U22386 ( .A(n20376), .ZN(n20369) );
  OAI21_X1 U22387 ( .B1(n20468), .B2(n20350), .A(n20349), .ZN(n20353) );
  NOR2_X1 U22388 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20351), .ZN(n20364) );
  AOI211_X1 U22389 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20351), .A(n20364), .B(
        n20490), .ZN(n20352) );
  AOI21_X1 U22390 ( .B1(n20369), .B2(n20353), .A(n20352), .ZN(n20359) );
  OAI21_X1 U22391 ( .B1(n20355), .B2(n20354), .A(n20387), .ZN(n20356) );
  NAND2_X1 U22392 ( .A1(n20357), .A2(n20356), .ZN(n20361) );
  OAI211_X1 U22393 ( .C1(n20357), .C2(n20356), .A(n20488), .B(n20361), .ZN(
        n20358) );
  NAND3_X1 U22394 ( .A1(n20360), .A2(n20359), .A3(n20358), .ZN(P3_U2651) );
  NAND2_X1 U22395 ( .A1(n20387), .A2(n20361), .ZN(n20362) );
  OAI211_X1 U22396 ( .C1(n20363), .C2(n20362), .A(n20488), .B(n20380), .ZN(
        n20366) );
  NAND2_X1 U22397 ( .A1(n20364), .A2(n20372), .ZN(n20373) );
  OAI211_X1 U22398 ( .C1(n20364), .C2(n20372), .A(n20515), .B(n20373), .ZN(
        n20365) );
  OAI211_X1 U22399 ( .C1(n20500), .C2(n20367), .A(n20366), .B(n20365), .ZN(
        n20368) );
  AOI21_X1 U22400 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n20369), .A(n20368), 
        .ZN(n20371) );
  NAND3_X1 U22401 ( .A1(n20445), .A2(n20377), .A3(n20370), .ZN(n20375) );
  OAI211_X1 U22402 ( .C1(n20372), .C2(n20498), .A(n20371), .B(n20375), .ZN(
        P3_U2650) );
  NOR2_X1 U22403 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20373), .ZN(n20395) );
  AOI211_X1 U22404 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20373), .A(n20395), .B(
        n20490), .ZN(n20374) );
  AOI21_X1 U22405 ( .B1(n20409), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n20374), .ZN(n20385) );
  AOI21_X1 U22406 ( .B1(n20376), .B2(n20375), .A(n20389), .ZN(n20379) );
  NAND2_X1 U22407 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20377), .ZN(n20388) );
  NOR3_X1 U22408 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20468), .A3(n20388), 
        .ZN(n20378) );
  AOI211_X1 U22409 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20516), .A(n20379), .B(
        n20378), .ZN(n20384) );
  OAI211_X1 U22410 ( .C1(n20382), .C2(n20381), .A(n20488), .B(n20386), .ZN(
        n20383) );
  NAND3_X1 U22411 ( .A1(n20385), .A2(n20384), .A3(n20383), .ZN(P3_U2649) );
  XOR2_X1 U22412 ( .A(n20399), .B(n20400), .Z(n20393) );
  NOR2_X1 U22413 ( .A1(n20389), .A2(n20388), .ZN(n20390) );
  NAND2_X1 U22414 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20390), .ZN(n20419) );
  AOI21_X1 U22415 ( .B1(n20419), .B2(n20445), .A(n20431), .ZN(n20410) );
  AOI21_X1 U22416 ( .B1(n20445), .B2(n20390), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n20391) );
  INV_X1 U22417 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20394) );
  OAI22_X1 U22418 ( .A1(n20410), .A2(n20391), .B1(n20498), .B2(n20394), .ZN(
        n20392) );
  AOI21_X1 U22419 ( .B1(n20488), .B2(n20393), .A(n20392), .ZN(n20397) );
  NAND2_X1 U22420 ( .A1(n20395), .A2(n20394), .ZN(n20403) );
  OAI211_X1 U22421 ( .C1(n20395), .C2(n20394), .A(n20515), .B(n20403), .ZN(
        n20396) );
  OAI211_X1 U22422 ( .C1(n20500), .C2(n20398), .A(n20397), .B(n20396), .ZN(
        P3_U2648) );
  AOI22_X1 U22423 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n20408) );
  NOR2_X1 U22424 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20468), .ZN(n20416) );
  INV_X1 U22425 ( .A(n20419), .ZN(n20406) );
  NOR2_X1 U22426 ( .A1(n20402), .A2(n20401), .ZN(n20411) );
  AOI211_X1 U22427 ( .C1(n20402), .C2(n20401), .A(n20411), .B(n21173), .ZN(
        n20405) );
  NOR2_X1 U22428 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20403), .ZN(n20418) );
  AOI211_X1 U22429 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20403), .A(n20418), .B(
        n20490), .ZN(n20404) );
  AOI211_X1 U22430 ( .C1(n20416), .C2(n20406), .A(n20405), .B(n20404), .ZN(
        n20407) );
  OAI211_X1 U22431 ( .C1(n20410), .C2(n20420), .A(n20408), .B(n20407), .ZN(
        P3_U2647) );
  AOI22_X1 U22432 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20409), .B1(
        n20516), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n20425) );
  INV_X1 U22433 ( .A(n20410), .ZN(n20415) );
  AOI211_X1 U22434 ( .C1(n20413), .C2(n20412), .A(n20433), .B(n21173), .ZN(
        n20414) );
  AOI221_X1 U22435 ( .B1(n20416), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n20415), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n20414), .ZN(n20424) );
  NAND2_X1 U22436 ( .A1(n20418), .A2(n20417), .ZN(n20432) );
  OAI211_X1 U22437 ( .C1(n20418), .C2(n20417), .A(n20515), .B(n20432), .ZN(
        n20423) );
  NOR2_X1 U22438 ( .A1(n20420), .A2(n20419), .ZN(n20426) );
  NAND3_X1 U22439 ( .A1(n20445), .A2(n20426), .A3(n20421), .ZN(n20422) );
  NAND4_X1 U22440 ( .A1(n20425), .A2(n20424), .A3(n20423), .A4(n20422), .ZN(
        P3_U2646) );
  NAND2_X1 U22441 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20426), .ZN(n20427) );
  INV_X1 U22442 ( .A(n20427), .ZN(n20429) );
  NOR2_X1 U22443 ( .A1(n20428), .A2(n20427), .ZN(n20444) );
  NOR2_X1 U22444 ( .A1(n20444), .A2(n20468), .ZN(n20430) );
  AOI22_X1 U22445 ( .A1(n20516), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n20429), 
        .B2(n20430), .ZN(n20440) );
  NOR2_X1 U22446 ( .A1(n20431), .A2(n20430), .ZN(n20456) );
  INV_X1 U22447 ( .A(n20456), .ZN(n20438) );
  NOR2_X1 U22448 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20432), .ZN(n20450) );
  AOI211_X1 U22449 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20432), .A(n20450), .B(
        n20490), .ZN(n20437) );
  AOI211_X1 U22450 ( .C1(n20435), .C2(n20434), .A(n20441), .B(n21173), .ZN(
        n20436) );
  AOI211_X1 U22451 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n20438), .A(n20437), 
        .B(n20436), .ZN(n20439) );
  OAI211_X1 U22452 ( .C1(n11095), .C2(n20500), .A(n20440), .B(n20439), .ZN(
        P3_U2645) );
  NOR2_X1 U22453 ( .A1(n20441), .A2(n20482), .ZN(n20442) );
  NOR2_X1 U22454 ( .A1(n20443), .A2(n20442), .ZN(n20459) );
  AOI211_X1 U22455 ( .C1(n20443), .C2(n20442), .A(n20459), .B(n21173), .ZN(
        n20448) );
  NAND2_X1 U22456 ( .A1(n20445), .A2(n20444), .ZN(n20453) );
  OR2_X1 U22457 ( .A1(n20453), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n20455) );
  OAI21_X1 U22458 ( .B1(n20446), .B2(n20500), .A(n20455), .ZN(n20447) );
  AOI211_X1 U22459 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20516), .A(n20448), .B(
        n20447), .ZN(n20452) );
  NAND2_X1 U22460 ( .A1(n20450), .A2(n20449), .ZN(n20457) );
  OAI211_X1 U22461 ( .C1(n20450), .C2(n20449), .A(n20515), .B(n20457), .ZN(
        n20451) );
  OAI211_X1 U22462 ( .C1(n20456), .C2(n20454), .A(n20452), .B(n20451), .ZN(
        P3_U2644) );
  NOR2_X1 U22463 ( .A1(n20454), .A2(n20453), .ZN(n20484) );
  AOI22_X1 U22464 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20516), .B1(n20484), 
        .B2(n20466), .ZN(n20465) );
  NAND2_X1 U22465 ( .A1(n20456), .A2(n20455), .ZN(n20469) );
  NOR2_X1 U22466 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20457), .ZN(n20472) );
  AOI211_X1 U22467 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20457), .A(n20472), .B(
        n20490), .ZN(n20463) );
  INV_X1 U22468 ( .A(n20458), .ZN(n20461) );
  NOR2_X1 U22469 ( .A1(n20461), .A2(n20460), .ZN(n20474) );
  AOI211_X1 U22470 ( .C1(n20461), .C2(n20460), .A(n20474), .B(n21173), .ZN(
        n20462) );
  AOI211_X1 U22471 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n20469), .A(n20463), 
        .B(n20462), .ZN(n20464) );
  OAI211_X1 U22472 ( .C1(n11096), .C2(n20500), .A(n20465), .B(n20464), .ZN(
        P3_U2643) );
  NOR2_X1 U22473 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20466), .ZN(n20467) );
  AOI22_X1 U22474 ( .A1(n20516), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n20484), 
        .B2(n20467), .ZN(n20480) );
  NAND2_X1 U22475 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n20470) );
  NAND2_X1 U22476 ( .A1(n20468), .A2(n20514), .ZN(n20513) );
  AOI21_X1 U22477 ( .B1(n20470), .B2(n20513), .A(n20469), .ZN(n20486) );
  INV_X1 U22478 ( .A(n20486), .ZN(n20506) );
  INV_X1 U22479 ( .A(n20472), .ZN(n20473) );
  NAND2_X1 U22480 ( .A1(n20472), .A2(n20471), .ZN(n20489) );
  NAND2_X1 U22481 ( .A1(n20515), .A2(n20489), .ZN(n20492) );
  AOI21_X1 U22482 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n20473), .A(n20492), .ZN(
        n20478) );
  NOR2_X1 U22483 ( .A1(n20474), .A2(n20482), .ZN(n20475) );
  NOR2_X1 U22484 ( .A1(n20476), .A2(n20475), .ZN(n20483) );
  AOI211_X1 U22485 ( .C1(n20476), .C2(n20475), .A(n20483), .B(n21173), .ZN(
        n20477) );
  AOI211_X1 U22486 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n20506), .A(n20478), 
        .B(n20477), .ZN(n20479) );
  OAI211_X1 U22487 ( .C1(n20481), .C2(n20500), .A(n20480), .B(n20479), .ZN(
        P3_U2642) );
  NAND3_X1 U22488 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n20484), .ZN(n20496) );
  NOR2_X1 U22489 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20496), .ZN(n20507) );
  OAI22_X1 U22490 ( .A1(n20486), .A2(n20497), .B1(n20485), .B2(n20500), .ZN(
        n20487) );
  NOR2_X1 U22491 ( .A1(n20490), .A2(n20489), .ZN(n20505) );
  OAI21_X1 U22492 ( .B1(n20516), .B2(n20505), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20491) );
  NAND2_X1 U22493 ( .A1(n20494), .A2(n20493), .ZN(n20511) );
  INV_X1 U22494 ( .A(n20495), .ZN(n20510) );
  INV_X1 U22495 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20504) );
  NOR3_X1 U22496 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20497), .A3(n20496), 
        .ZN(n20503) );
  OAI22_X1 U22497 ( .A1(n20501), .A2(n20500), .B1(n20499), .B2(n20498), .ZN(
        n20502) );
  AOI211_X1 U22498 ( .C1(n20505), .C2(n20504), .A(n20503), .B(n20502), .ZN(
        n20509) );
  OAI21_X1 U22499 ( .B1(n20507), .B2(n20506), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n20508) );
  OAI211_X1 U22500 ( .C1(n20511), .C2(n20510), .A(n20509), .B(n20508), .ZN(
        P3_U2640) );
  AOI22_X1 U22501 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n20513), .B1(n20512), 
        .B2(n20712), .ZN(n20519) );
  NAND3_X1 U22502 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20514), .A3(
        n20730), .ZN(n20518) );
  OAI21_X1 U22503 ( .B1(n20516), .B2(n20515), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20517) );
  NAND3_X1 U22504 ( .A1(n20519), .A2(n20518), .A3(n20517), .ZN(P3_U2671) );
  NAND2_X1 U22505 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n20581) );
  NOR3_X1 U22506 ( .A1(n20522), .A2(n20521), .A3(n20520), .ZN(n20523) );
  NAND2_X1 U22507 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n20575), .ZN(n20565) );
  NAND2_X1 U22508 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20568), .ZN(n20557) );
  NAND2_X1 U22509 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n20560), .ZN(n20553) );
  NAND2_X1 U22510 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20552), .ZN(n20542) );
  NAND2_X1 U22511 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20540), .ZN(n20532) );
  NAND2_X1 U22512 ( .A1(n20532), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20531) );
  NAND2_X1 U22513 ( .A1(n20528), .A2(n20596), .ZN(n20573) );
  AOI22_X1 U22514 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20705), .B1(n20704), .B2(
        n20529), .ZN(n20530) );
  OAI221_X1 U22515 ( .B1(n20532), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20531), 
        .C2(n20686), .A(n20530), .ZN(P3_U2722) );
  INV_X1 U22516 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20535) );
  INV_X1 U22517 ( .A(n20532), .ZN(n20679) );
  AOI21_X1 U22518 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20700), .A(n20540), .ZN(
        n20534) );
  OAI222_X1 U22519 ( .A1(n20573), .A2(n20535), .B1(n20679), .B2(n20534), .C1(
        n20691), .C2(n20533), .ZN(P3_U2723) );
  INV_X1 U22520 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20541) );
  OAI21_X1 U22521 ( .B1(n20536), .B2(n20686), .A(n20542), .ZN(n20537) );
  INV_X1 U22522 ( .A(n20537), .ZN(n20539) );
  OAI222_X1 U22523 ( .A1(n20573), .A2(n20541), .B1(n20540), .B2(n20539), .C1(
        n20691), .C2(n20538), .ZN(P3_U2724) );
  NAND2_X1 U22524 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20705), .ZN(n20544) );
  OAI211_X1 U22525 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n20552), .A(n20700), .B(
        n20542), .ZN(n20543) );
  OAI211_X1 U22526 ( .C1(n20545), .C2(n20691), .A(n20544), .B(n20543), .ZN(
        P3_U2725) );
  NAND4_X1 U22527 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_7__SCAN_IN), .ZN(n20546) );
  NOR4_X4 U22528 ( .A1(n20699), .A2(n20548), .A3(n20547), .A4(n20546), .ZN(
        n20695) );
  OAI221_X1 U22529 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20695), .C1(
        P3_EAX_REG_9__SCAN_IN), .C2(P3_EAX_REG_8__SCAN_IN), .A(n20700), .ZN(
        n20551) );
  AOI22_X1 U22530 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20705), .B1(n20704), .B2(
        n20549), .ZN(n20550) );
  OAI21_X1 U22531 ( .B1(n20552), .B2(n20551), .A(n20550), .ZN(P3_U2726) );
  INV_X1 U22532 ( .A(n20553), .ZN(n20556) );
  AOI21_X1 U22533 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20700), .A(n20560), .ZN(
        n20555) );
  OAI222_X1 U22534 ( .A1(n20671), .A2(n20573), .B1(n20556), .B2(n20555), .C1(
        n20691), .C2(n20554), .ZN(P3_U2728) );
  INV_X1 U22535 ( .A(n20557), .ZN(n20563) );
  AOI21_X1 U22536 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20700), .A(n20563), .ZN(
        n20559) );
  OAI222_X1 U22537 ( .A1(n20605), .A2(n20573), .B1(n20560), .B2(n20559), .C1(
        n20691), .C2(n20558), .ZN(P3_U2729) );
  AOI21_X1 U22538 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20700), .A(n20568), .ZN(
        n20562) );
  OAI222_X1 U22539 ( .A1(n20564), .A2(n20573), .B1(n20563), .B2(n20562), .C1(
        n20691), .C2(n20561), .ZN(P3_U2730) );
  INV_X1 U22540 ( .A(n20565), .ZN(n20572) );
  AOI21_X1 U22541 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20700), .A(n20572), .ZN(
        n20567) );
  OAI222_X1 U22542 ( .A1(n20569), .A2(n20573), .B1(n20568), .B2(n20567), .C1(
        n20691), .C2(n20566), .ZN(P3_U2731) );
  AOI21_X1 U22543 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20700), .A(n20575), .ZN(
        n20571) );
  OAI222_X1 U22544 ( .A1(n20574), .A2(n20573), .B1(n20572), .B2(n20571), .C1(
        n20691), .C2(n20570), .ZN(P3_U2732) );
  AOI211_X1 U22545 ( .C1(n20699), .C2(n20576), .A(n20686), .B(n20575), .ZN(
        n20577) );
  AOI21_X1 U22546 ( .B1(n20705), .B2(BUF2_REG_2__SCAN_IN), .A(n20577), .ZN(
        n20578) );
  OAI21_X1 U22547 ( .B1(n20579), .B2(n20691), .A(n20578), .ZN(P3_U2733) );
  NOR4_X1 U22548 ( .A1(n20683), .A2(n20582), .A3(n20581), .A4(n20580), .ZN(
        n20583) );
  NOR2_X2 U22549 ( .A1(n20688), .A2(n20687), .ZN(n20685) );
  NAND2_X1 U22550 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20616), .ZN(n20612) );
  NAND2_X1 U22551 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20606), .ZN(n20592) );
  NAND2_X1 U22552 ( .A1(n20700), .A2(n20592), .ZN(n20598) );
  NAND2_X1 U22553 ( .A1(n20585), .A2(n20686), .ZN(n20672) );
  INV_X1 U22554 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20587) );
  NAND2_X1 U22555 ( .A1(n20586), .A2(n20686), .ZN(n20631) );
  OAI22_X1 U22556 ( .A1(n20588), .A2(n20691), .B1(n20587), .B2(n20631), .ZN(
        n20589) );
  AOI21_X1 U22557 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20673), .A(n20589), .ZN(
        n20590) );
  OAI221_X1 U22558 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20592), .C1(n20591), 
        .C2(n20598), .A(n20590), .ZN(P3_U2714) );
  AOI22_X1 U22559 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n20673), .ZN(n20594) );
  OAI211_X1 U22560 ( .C1(n20606), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20700), .B(
        n20592), .ZN(n20593) );
  OAI211_X1 U22561 ( .C1(n20595), .C2(n20691), .A(n20594), .B(n20593), .ZN(
        P3_U2715) );
  NAND2_X1 U22562 ( .A1(n20597), .A2(n20596), .ZN(n20707) );
  OAI21_X1 U22563 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20707), .A(n20598), .ZN(
        n20603) );
  NAND3_X1 U22564 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .ZN(n20624) );
  NOR3_X1 U22565 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20624), .A3(n20612), .ZN(
        n20602) );
  OAI22_X1 U22566 ( .A1(n20600), .A2(n20691), .B1(n20599), .B2(n20631), .ZN(
        n20601) );
  AOI211_X1 U22567 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n20603), .A(n20602), .B(
        n20601), .ZN(n20604) );
  OAI21_X1 U22568 ( .B1(n20605), .B2(n20672), .A(n20604), .ZN(P3_U2713) );
  AOI22_X1 U22569 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n20673), .ZN(n20610) );
  AOI211_X1 U22570 ( .C1(n20607), .C2(n20612), .A(n20606), .B(n20686), .ZN(
        n20608) );
  INV_X1 U22571 ( .A(n20608), .ZN(n20609) );
  OAI211_X1 U22572 ( .C1(n20611), .C2(n20691), .A(n20610), .B(n20609), .ZN(
        P3_U2716) );
  AOI22_X1 U22573 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n20673), .ZN(n20614) );
  OAI211_X1 U22574 ( .C1(n20616), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20700), .B(
        n20612), .ZN(n20613) );
  OAI211_X1 U22575 ( .C1(n20615), .C2(n20691), .A(n20614), .B(n20613), .ZN(
        P3_U2717) );
  AOI22_X1 U22576 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n20673), .ZN(n20620) );
  INV_X1 U22577 ( .A(n20675), .ZN(n20618) );
  INV_X1 U22578 ( .A(n20616), .ZN(n20617) );
  OAI211_X1 U22579 ( .C1(n20618), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20700), .B(
        n20617), .ZN(n20619) );
  OAI211_X1 U22580 ( .C1(n20621), .C2(n20691), .A(n20620), .B(n20619), .ZN(
        P3_U2718) );
  AOI22_X1 U22581 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20673), .B1(n20704), .B2(
        n20622), .ZN(n20629) );
  NAND3_X1 U22582 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n20623) );
  NOR3_X2 U22583 ( .A1(n20675), .A2(n20624), .A3(n20623), .ZN(n20668) );
  NAND2_X1 U22584 ( .A1(n20668), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20667) );
  AOI211_X1 U22585 ( .C1(n20626), .C2(n20661), .A(n20632), .B(n20686), .ZN(
        n20627) );
  INV_X1 U22586 ( .A(n20627), .ZN(n20628) );
  OAI211_X1 U22587 ( .C1(n20631), .C2(n20630), .A(n20629), .B(n20628), .ZN(
        P3_U2710) );
  AOI22_X1 U22588 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n20673), .ZN(n20634) );
  NAND2_X1 U22589 ( .A1(n20632), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20654) );
  OAI211_X1 U22590 ( .C1(n20632), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20700), .B(
        n20654), .ZN(n20633) );
  OAI211_X1 U22591 ( .C1(n20635), .C2(n20691), .A(n20634), .B(n20633), .ZN(
        P3_U2709) );
  NOR2_X2 U22592 ( .A1(n20654), .A2(n20655), .ZN(n20653) );
  NAND2_X1 U22593 ( .A1(n20653), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20649) );
  NOR2_X2 U22594 ( .A1(n20649), .A2(n20643), .ZN(n20642) );
  NAND2_X1 U22595 ( .A1(n20642), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20638) );
  NAND2_X1 U22596 ( .A1(n20638), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n20637) );
  NAND2_X1 U22597 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20674), .ZN(n20636) );
  OAI221_X1 U22598 ( .B1(n20638), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n20637), 
        .C2(n20686), .A(n20636), .ZN(P3_U2704) );
  AOI22_X1 U22599 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n20673), .ZN(n20640) );
  OAI211_X1 U22600 ( .C1(n20642), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20700), .B(
        n20638), .ZN(n20639) );
  OAI211_X1 U22601 ( .C1(n20641), .C2(n20691), .A(n20640), .B(n20639), .ZN(
        P3_U2705) );
  INV_X1 U22602 ( .A(n20642), .ZN(n20645) );
  OAI21_X1 U22603 ( .B1(n20686), .B2(n20643), .A(n20649), .ZN(n20644) );
  AOI22_X1 U22604 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20674), .B1(n20645), .B2(
        n20644), .ZN(n20648) );
  AOI22_X1 U22605 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20673), .B1(n20704), .B2(
        n20646), .ZN(n20647) );
  NAND2_X1 U22606 ( .A1(n20648), .A2(n20647), .ZN(P3_U2706) );
  AOI22_X1 U22607 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n20673), .ZN(n20651) );
  OAI211_X1 U22608 ( .C1(n20653), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20700), .B(
        n20649), .ZN(n20650) );
  OAI211_X1 U22609 ( .C1(n20652), .C2(n20691), .A(n20651), .B(n20650), .ZN(
        P3_U2707) );
  INV_X1 U22610 ( .A(n20653), .ZN(n20657) );
  OAI21_X1 U22611 ( .B1(n20686), .B2(n20655), .A(n20654), .ZN(n20656) );
  AOI22_X1 U22612 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20674), .B1(n20657), .B2(
        n20656), .ZN(n20660) );
  AOI22_X1 U22613 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20673), .B1(n20704), .B2(
        n20658), .ZN(n20659) );
  NAND2_X1 U22614 ( .A1(n20660), .A2(n20659), .ZN(P3_U2708) );
  AOI22_X1 U22615 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n20673), .ZN(n20664) );
  OAI211_X1 U22616 ( .C1(n20662), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20700), .B(
        n20661), .ZN(n20663) );
  OAI211_X1 U22617 ( .C1(n20665), .C2(n20691), .A(n20664), .B(n20663), .ZN(
        P3_U2711) );
  AOI22_X1 U22618 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n20674), .B1(n20704), .B2(
        n20666), .ZN(n20670) );
  OAI211_X1 U22619 ( .C1(n20668), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20700), .B(
        n20667), .ZN(n20669) );
  OAI211_X1 U22620 ( .C1(n20672), .C2(n20671), .A(n20670), .B(n20669), .ZN(
        P3_U2712) );
  AOI22_X1 U22621 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n20674), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n20673), .ZN(n20677) );
  OAI211_X1 U22622 ( .C1(n20685), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20700), .B(
        n20675), .ZN(n20676) );
  OAI211_X1 U22623 ( .C1(n20678), .C2(n20691), .A(n20677), .B(n20676), .ZN(
        P3_U2719) );
  NAND2_X1 U22624 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20679), .ZN(n20684) );
  NAND2_X1 U22625 ( .A1(n20700), .A2(n20688), .ZN(n20682) );
  AOI22_X1 U22626 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20705), .B1(n20704), .B2(
        n20680), .ZN(n20681) );
  OAI221_X1 U22627 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n20684), .C1(n20683), 
        .C2(n20682), .A(n20681), .ZN(P3_U2721) );
  AOI211_X1 U22628 ( .C1(n20688), .C2(n20687), .A(n20686), .B(n20685), .ZN(
        n20689) );
  AOI21_X1 U22629 ( .B1(n20705), .B2(BUF2_REG_15__SCAN_IN), .A(n20689), .ZN(
        n20690) );
  OAI21_X1 U22630 ( .B1(n20692), .B2(n20691), .A(n20690), .ZN(P3_U2720) );
  AOI22_X1 U22631 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20705), .B1(n20704), .B2(
        n20693), .ZN(n20697) );
  NAND2_X1 U22632 ( .A1(n20695), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n20694) );
  OAI211_X1 U22633 ( .C1(n20695), .C2(P3_EAX_REG_8__SCAN_IN), .A(n20700), .B(
        n20694), .ZN(n20696) );
  NAND2_X1 U22634 ( .A1(n20697), .A2(n20696), .ZN(P3_U2727) );
  AOI22_X1 U22635 ( .A1(n20705), .A2(BUF2_REG_1__SCAN_IN), .B1(n20704), .B2(
        n20698), .ZN(n20702) );
  OAI211_X1 U22636 ( .C1(n20709), .C2(P3_EAX_REG_1__SCAN_IN), .A(n20700), .B(
        n20699), .ZN(n20701) );
  NAND2_X1 U22637 ( .A1(n20702), .A2(n20701), .ZN(P3_U2734) );
  AOI22_X1 U22638 ( .A1(n20705), .A2(BUF2_REG_0__SCAN_IN), .B1(n20704), .B2(
        n20703), .ZN(n20706) );
  OAI221_X1 U22639 ( .B1(n20709), .B2(n20708), .C1(n20709), .C2(n20707), .A(
        n20706), .ZN(P3_U2735) );
  NOR2_X1 U22640 ( .A1(n20710), .A2(n20946), .ZN(n20714) );
  AOI22_X1 U22641 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20931), .B1(
        n20714), .B2(n20712), .ZN(n21148) );
  AOI222_X1 U22642 ( .A1(n20886), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21148), 
        .B2(n20757), .C1(n20712), .C2(n21178), .ZN(n20711) );
  AOI22_X1 U22643 ( .A1(n20762), .A2(n20712), .B1(n20711), .B2(n20759), .ZN(
        P3_U3290) );
  AOI211_X1 U22644 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20946), .A(
        n20713), .B(n20738), .ZN(n20722) );
  OAI22_X1 U22645 ( .A1(n20714), .A2(n20715), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20722), .ZN(n21146) );
  INV_X1 U22646 ( .A(n20715), .ZN(n20718) );
  AOI22_X1 U22647 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20716), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11497), .ZN(n20731) );
  NAND2_X1 U22648 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20732) );
  INV_X1 U22649 ( .A(n20732), .ZN(n20717) );
  AOI222_X1 U22650 ( .A1(n21146), .A2(n20757), .B1(n20718), .B2(n21178), .C1(
        n20731), .C2(n20717), .ZN(n20719) );
  AOI22_X1 U22651 ( .A1(n20762), .A2(n11406), .B1(n20719), .B2(n20759), .ZN(
        P3_U3289) );
  NAND2_X1 U22652 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20720), .ZN(
        n20735) );
  OAI33_X1 U22653 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20722), .A3(
        n11406), .B1(n21143), .B2(n20721), .B3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20728) );
  NOR2_X1 U22654 ( .A1(n20724), .A2(n20723), .ZN(n20744) );
  AOI211_X1 U22655 ( .C1(n11406), .C2(n20738), .A(n20744), .B(n20751), .ZN(
        n20726) );
  OAI22_X1 U22656 ( .A1(n20726), .A2(n20735), .B1(n21094), .B2(n20725), .ZN(
        n20727) );
  NOR2_X1 U22657 ( .A1(n20728), .A2(n20727), .ZN(n21142) );
  OAI222_X1 U22658 ( .A1(n20732), .A2(n20731), .B1(n20730), .B2(n21142), .C1(
        n20729), .C2(n20736), .ZN(n20733) );
  AOI22_X1 U22659 ( .A1(n20762), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20733), .B2(n20759), .ZN(n20734) );
  OAI21_X1 U22660 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(P3_U3288) );
  INV_X1 U22661 ( .A(n20737), .ZN(n20758) );
  NOR2_X1 U22662 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20738), .ZN(
        n20756) );
  OAI211_X1 U22663 ( .C1(n20742), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        n20745) );
  AOI22_X1 U22664 ( .A1(n21126), .A2(n20745), .B1(n20744), .B2(n20743), .ZN(
        n20754) );
  AOI222_X1 U22665 ( .A1(n20749), .A2(n20748), .B1(n20749), .B2(n20755), .C1(
        n20747), .C2(n20746), .ZN(n20750) );
  AOI21_X1 U22666 ( .B1(n20752), .B2(n20751), .A(n20750), .ZN(n20753) );
  OAI211_X1 U22667 ( .C1(n20756), .C2(n20755), .A(n20754), .B(n20753), .ZN(
        n21140) );
  AOI22_X1 U22668 ( .A1(n21178), .A2(n20758), .B1(n20757), .B2(n21140), .ZN(
        n20760) );
  AOI22_X1 U22669 ( .A1(n20762), .A2(n20761), .B1(n20760), .B2(n20759), .ZN(
        P3_U3285) );
  NAND2_X1 U22670 ( .A1(n20933), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20763) );
  AOI22_X1 U22671 ( .A1(n21126), .A2(n20764), .B1(n21103), .B2(n20763), .ZN(
        n21041) );
  AOI22_X1 U22672 ( .A1(n21126), .A2(n20769), .B1(n21103), .B2(n21053), .ZN(
        n20768) );
  AOI22_X1 U22673 ( .A1(n21063), .A2(n20766), .B1(n21125), .B2(n20765), .ZN(
        n20767) );
  NAND2_X1 U22674 ( .A1(n20946), .A2(n20886), .ZN(n21059) );
  OAI211_X1 U22675 ( .C1(n10951), .C2(n20933), .A(n21093), .B(n21059), .ZN(
        n21043) );
  AOI211_X1 U22676 ( .C1(n20946), .C2(n20769), .A(n20935), .B(n21043), .ZN(
        n20776) );
  NAND2_X1 U22677 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21105), .ZN(
        n20775) );
  AND2_X1 U22678 ( .A1(n21093), .A2(n20770), .ZN(n21054) );
  AOI22_X1 U22679 ( .A1(n21120), .A2(n20772), .B1(n20771), .B2(n21054), .ZN(
        n20774) );
  NAND2_X1 U22680 ( .A1(n10958), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n20773) );
  OAI211_X1 U22681 ( .C1(n20776), .C2(n20775), .A(n20774), .B(n20773), .ZN(
        P3_U2841) );
  NAND2_X1 U22682 ( .A1(n10951), .A2(n21094), .ZN(n21047) );
  INV_X1 U22683 ( .A(n21047), .ZN(n20777) );
  AOI221_X1 U22684 ( .B1(n20777), .B2(n20886), .C1(n20931), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n20997), .ZN(n20778) );
  AOI221_X1 U22685 ( .B1(n20965), .B2(n20780), .C1(n20847), .C2(n20779), .A(
        n20778), .ZN(n20782) );
  NAND2_X1 U22686 ( .A1(n10958), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20781) );
  OAI211_X1 U22687 ( .C1(n21022), .C2(n20886), .A(n20782), .B(n20781), .ZN(
        P3_U2862) );
  INV_X1 U22688 ( .A(n20783), .ZN(n20791) );
  AOI22_X1 U22689 ( .A1(n10958), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21006), .ZN(n20790) );
  NOR2_X1 U22690 ( .A1(n20949), .A2(n20784), .ZN(n20786) );
  AND2_X1 U22691 ( .A1(n20886), .A2(n21047), .ZN(n20785) );
  MUX2_X1 U22692 ( .A(n20786), .B(n20785), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n20788) );
  AOI22_X1 U22693 ( .A1(n21093), .A2(n20788), .B1(n20847), .B2(n20787), .ZN(
        n20789) );
  OAI211_X1 U22694 ( .C1(n20791), .C2(n20953), .A(n20790), .B(n20789), .ZN(
        P3_U2861) );
  OAI21_X1 U22695 ( .B1(n20794), .B2(n20793), .A(n20792), .ZN(n20806) );
  NAND2_X1 U22696 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20810), .ZN(
        n20802) );
  NOR2_X1 U22697 ( .A1(n11497), .A2(n20886), .ZN(n20796) );
  AOI21_X1 U22698 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21059), .A(
        n21072), .ZN(n20795) );
  AOI21_X1 U22699 ( .B1(n20796), .B2(n21126), .A(n20795), .ZN(n20800) );
  AOI22_X1 U22700 ( .A1(n21126), .A2(n20813), .B1(n20798), .B2(n20797), .ZN(
        n20799) );
  OAI221_X1 U22701 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20802), .C1(
        n20801), .C2(n20800), .A(n20799), .ZN(n20803) );
  AOI22_X1 U22702 ( .A1(n21093), .A2(n20803), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21006), .ZN(n20805) );
  OAI211_X1 U22703 ( .C1(n20953), .C2(n20806), .A(n20805), .B(n20804), .ZN(
        P3_U2860) );
  NOR2_X1 U22704 ( .A1(n11501), .A2(n21022), .ZN(n20807) );
  AOI211_X1 U22705 ( .C1(n20847), .C2(n20809), .A(n20808), .B(n20807), .ZN(
        n20816) );
  INV_X1 U22706 ( .A(n20810), .ZN(n20811) );
  NAND2_X1 U22707 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20812) );
  OAI22_X1 U22708 ( .A1(n20813), .A2(n21094), .B1(n20811), .B2(n20812), .ZN(
        n20835) );
  AOI22_X1 U22709 ( .A1(n21126), .A2(n20813), .B1(n21112), .B2(n20812), .ZN(
        n20814) );
  NAND3_X1 U22710 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20814), .A3(
        n21059), .ZN(n20818) );
  OAI211_X1 U22711 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20835), .A(
        n21093), .B(n20818), .ZN(n20815) );
  OAI211_X1 U22712 ( .C1(n20817), .C2(n20953), .A(n20816), .B(n20815), .ZN(
        P3_U2859) );
  NAND3_X1 U22713 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21085), .A3(
        n20818), .ZN(n20821) );
  NAND3_X1 U22714 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20819), .A3(
        n20835), .ZN(n20820) );
  NAND3_X1 U22715 ( .A1(n20822), .A2(n20821), .A3(n20820), .ZN(n20823) );
  AOI22_X1 U22716 ( .A1(n21093), .A2(n20823), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21006), .ZN(n20824) );
  OAI21_X1 U22717 ( .B1(n21105), .B2(n20825), .A(n20824), .ZN(P3_U2858) );
  OAI211_X1 U22718 ( .C1(n20826), .C2(n21094), .A(n21093), .B(n21059), .ZN(
        n20828) );
  OAI221_X1 U22719 ( .B1(n20828), .B2(n21112), .C1(n20828), .C2(n20827), .A(
        n21105), .ZN(n20837) );
  AND4_X1 U22720 ( .A1(n20833), .A2(n20835), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20830) );
  OAI21_X1 U22721 ( .B1(n20830), .B2(n20829), .A(n21093), .ZN(n20832) );
  NAND2_X1 U22722 ( .A1(n10958), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n20831) );
  OAI211_X1 U22723 ( .C1(n20833), .C2(n20837), .A(n20832), .B(n20831), .ZN(
        P3_U2857) );
  NOR2_X1 U22724 ( .A1(n21105), .A2(n20834), .ZN(n20841) );
  NAND2_X1 U22725 ( .A1(n20836), .A2(n20835), .ZN(n20848) );
  NOR2_X1 U22726 ( .A1(n20997), .A2(n20848), .ZN(n20839) );
  INV_X1 U22727 ( .A(n20837), .ZN(n20838) );
  MUX2_X1 U22728 ( .A(n20839), .B(n20838), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n20840) );
  AOI211_X1 U22729 ( .C1(n20847), .C2(n20842), .A(n20841), .B(n20840), .ZN(
        n20843) );
  OAI21_X1 U22730 ( .B1(n20953), .B2(n20844), .A(n20843), .ZN(P3_U2856) );
  AOI22_X1 U22731 ( .A1(n20847), .A2(n20846), .B1(n20965), .B2(n20845), .ZN(
        n20857) );
  INV_X1 U22732 ( .A(n21059), .ZN(n21114) );
  AOI211_X1 U22733 ( .C1(n21126), .C2(n20851), .A(n21114), .B(n20850), .ZN(
        n20852) );
  OAI21_X1 U22734 ( .B1(n21072), .B2(n20853), .A(n20852), .ZN(n20859) );
  NAND3_X1 U22735 ( .A1(n20877), .A2(n21093), .A3(n20859), .ZN(n20855) );
  OAI221_X1 U22736 ( .B1(n21006), .B2(n21093), .C1(n21006), .C2(n20859), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20854) );
  NAND4_X1 U22737 ( .A1(n20857), .A2(n20856), .A3(n20855), .A4(n20854), .ZN(
        P3_U2855) );
  AOI22_X1 U22738 ( .A1(n10958), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21006), .ZN(n20865) );
  NAND3_X1 U22739 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20877), .A3(
        n20858), .ZN(n20861) );
  NAND3_X1 U22740 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21085), .A3(
        n20859), .ZN(n20860) );
  OAI211_X1 U22741 ( .C1(n20862), .C2(n20993), .A(n20861), .B(n20860), .ZN(
        n20863) );
  AOI22_X1 U22742 ( .A1(n21093), .A2(n20863), .B1(n21120), .B2(n20862), .ZN(
        n20864) );
  OAI211_X1 U22743 ( .C1(n20953), .C2(n20866), .A(n20865), .B(n20864), .ZN(
        P3_U2854) );
  OAI21_X1 U22744 ( .B1(n20880), .B2(n21113), .A(n21103), .ZN(n20867) );
  OAI21_X1 U22745 ( .B1(n20868), .B2(n21094), .A(n20867), .ZN(n20889) );
  NOR2_X1 U22746 ( .A1(n21063), .A2(n21125), .ZN(n21068) );
  OAI22_X1 U22747 ( .A1(n20887), .A2(n21094), .B1(n20995), .B2(n20869), .ZN(
        n20870) );
  AOI211_X1 U22748 ( .C1(n21063), .C2(n21062), .A(n21006), .B(n20870), .ZN(
        n21117) );
  OR2_X1 U22749 ( .A1(n20886), .A2(n21113), .ZN(n20871) );
  OAI21_X1 U22750 ( .B1(n21115), .B2(n20871), .A(n20946), .ZN(n20872) );
  OAI211_X1 U22751 ( .C1(n20873), .C2(n21068), .A(n21117), .B(n20872), .ZN(
        n21107) );
  AOI211_X1 U22752 ( .C1(n20946), .C2(n20874), .A(n20889), .B(n21107), .ZN(
        n20876) );
  NOR2_X1 U22753 ( .A1(n20876), .A2(n20875), .ZN(n20882) );
  NAND2_X1 U22754 ( .A1(n20878), .A2(n20877), .ZN(n20917) );
  AOI21_X1 U22755 ( .B1(n20879), .B2(n20917), .A(n20997), .ZN(n21101) );
  INV_X1 U22756 ( .A(n21101), .ZN(n21123) );
  NOR3_X1 U22757 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n20880), .A3(
        n21123), .ZN(n20881) );
  AOI221_X1 U22758 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n10958), .C1(n20882), 
        .C2(n21105), .A(n20881), .ZN(n20883) );
  OAI21_X1 U22759 ( .B1(n20884), .B2(n21110), .A(n20883), .ZN(P3_U2851) );
  AOI22_X1 U22760 ( .A1(n10958), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n21120), 
        .B2(n20885), .ZN(n20898) );
  NOR3_X1 U22761 ( .A1(n20886), .A2(n20891), .A3(n21113), .ZN(n20888) );
  OAI22_X1 U22762 ( .A1(n10951), .A2(n20888), .B1(n20887), .B2(n21094), .ZN(
        n20902) );
  AOI211_X1 U22763 ( .C1(n21103), .C2(n20890), .A(n20889), .B(n20902), .ZN(
        n20893) );
  OAI21_X1 U22764 ( .B1(n21062), .B2(n20891), .A(n21063), .ZN(n20892) );
  OAI211_X1 U22765 ( .C1(n20894), .C2(n20995), .A(n20893), .B(n20892), .ZN(
        n21096) );
  OAI22_X1 U22766 ( .A1(n20997), .A2(n20899), .B1(n21123), .B2(n20895), .ZN(
        n20896) );
  OAI21_X1 U22767 ( .B1(n21096), .B2(n20899), .A(n20896), .ZN(n20897) );
  OAI211_X1 U22768 ( .C1(n21022), .C2(n20899), .A(n20898), .B(n20897), .ZN(
        P3_U2850) );
  NOR2_X1 U22769 ( .A1(n20919), .A2(n20917), .ZN(n20906) );
  NOR2_X1 U22770 ( .A1(n20919), .A2(n21113), .ZN(n20914) );
  OAI22_X1 U22771 ( .A1(n20931), .A2(n20914), .B1(n20900), .B2(n21094), .ZN(
        n20901) );
  AOI211_X1 U22772 ( .C1(n20903), .C2(n21047), .A(n20902), .B(n20901), .ZN(
        n20904) );
  INV_X1 U22773 ( .A(n20904), .ZN(n20905) );
  MUX2_X1 U22774 ( .A(n20906), .B(n20905), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n20907) );
  AOI21_X1 U22775 ( .B1(n21063), .B2(n20908), .A(n20907), .ZN(n20913) );
  AOI22_X1 U22776 ( .A1(n10958), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21006), .ZN(n20912) );
  AOI22_X1 U22777 ( .A1(n21120), .A2(n20910), .B1(n20965), .B2(n20909), .ZN(
        n20911) );
  OAI211_X1 U22778 ( .C1(n20913), .C2(n20997), .A(n20912), .B(n20911), .ZN(
        P3_U2848) );
  OAI221_X1 U22779 ( .B1(n21072), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n21072), .C2(n20914), .A(n21059), .ZN(n20916) );
  AOI211_X1 U22780 ( .C1(n21064), .C2(n21126), .A(n20916), .B(n20915), .ZN(
        n20926) );
  NOR4_X1 U22781 ( .A1(n20926), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20925) );
  NAND2_X1 U22782 ( .A1(n21063), .A2(n20920), .ZN(n20927) );
  OAI22_X1 U22783 ( .A1(n20995), .A2(n20922), .B1(n20921), .B2(n20927), .ZN(
        n20924) );
  AOI221_X1 U22784 ( .B1(n20925), .B2(n21093), .C1(n20924), .C2(n21093), .A(
        n20923), .ZN(n20929) );
  INV_X1 U22785 ( .A(n20926), .ZN(n21084) );
  OAI211_X1 U22786 ( .C1(n21018), .C2(n20995), .A(n21093), .B(n20927), .ZN(
        n21086) );
  OAI211_X1 U22787 ( .C1(n21084), .C2(n21086), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21105), .ZN(n20928) );
  OAI211_X1 U22788 ( .C1(n20930), .C2(n21110), .A(n20929), .B(n20928), .ZN(
        P3_U2847) );
  NAND2_X1 U22789 ( .A1(n20931), .A2(n21094), .ZN(n21102) );
  NAND2_X1 U22790 ( .A1(n20933), .A2(n20932), .ZN(n20947) );
  INV_X1 U22791 ( .A(n20947), .ZN(n20934) );
  AOI21_X1 U22792 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20934), .A(
        n10951), .ZN(n20936) );
  NAND2_X1 U22793 ( .A1(n10958), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n20940) );
  OAI211_X1 U22794 ( .C1(n21022), .C2(n20942), .A(n20941), .B(n20940), .ZN(
        P3_U2840) );
  NAND2_X1 U22795 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n20948), .ZN(
        n20943) );
  NOR4_X1 U22796 ( .A1(n20945), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n20944), .A4(n20943), .ZN(n20957) );
  AOI221_X1 U22797 ( .B1(n21103), .B2(n20947), .C1(n20946), .C2(n20947), .A(
        n21114), .ZN(n21024) );
  OAI211_X1 U22798 ( .C1(n20949), .C2(n20948), .A(n21025), .B(n21024), .ZN(
        n20961) );
  INV_X1 U22799 ( .A(n20961), .ZN(n20951) );
  OAI22_X1 U22800 ( .A1(n20951), .A2(n20963), .B1(n20993), .B2(n20950), .ZN(
        n20956) );
  OAI22_X1 U22801 ( .A1(n21110), .A2(n20954), .B1(n20953), .B2(n20952), .ZN(
        n20955) );
  AOI221_X1 U22802 ( .B1(n20957), .B2(n21093), .C1(n20956), .C2(n21093), .A(
        n20955), .ZN(n20959) );
  OAI211_X1 U22803 ( .C1(n21022), .C2(n20963), .A(n20959), .B(n20958), .ZN(
        P3_U2837) );
  INV_X1 U22804 ( .A(n20960), .ZN(n20974) );
  AOI211_X1 U22805 ( .C1(n21085), .C2(n20963), .A(n20962), .B(n20961), .ZN(
        n20967) );
  NAND2_X1 U22806 ( .A1(n21063), .A2(n20976), .ZN(n20966) );
  NAND2_X1 U22807 ( .A1(n20965), .A2(n20964), .ZN(n20982) );
  OAI221_X1 U22808 ( .B1(n20997), .B2(n20967), .C1(n20997), .C2(n20966), .A(
        n20982), .ZN(n20971) );
  INV_X1 U22809 ( .A(n21016), .ZN(n20969) );
  NOR2_X1 U22810 ( .A1(n20969), .A2(n20968), .ZN(n20970) );
  AOI222_X1 U22811 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n20971), 
        .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21006), .C1(n20971), 
        .C2(n20970), .ZN(n20973) );
  OAI211_X1 U22812 ( .C1(n20974), .C2(n21110), .A(n20973), .B(n20972), .ZN(
        P3_U2836) );
  AOI211_X1 U22813 ( .C1(n21063), .C2(n20976), .A(n20980), .B(n20975), .ZN(
        n20977) );
  OAI211_X1 U22814 ( .C1(n21072), .C2(n20978), .A(n21024), .B(n20977), .ZN(
        n20979) );
  AOI22_X1 U22815 ( .A1(n21093), .A2(n20979), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21006), .ZN(n20983) );
  AOI22_X1 U22816 ( .A1(n20983), .A2(n20982), .B1(n20981), .B2(n20980), .ZN(
        n20984) );
  AOI21_X1 U22817 ( .B1(n21120), .B2(n20985), .A(n20984), .ZN(n20987) );
  NAND2_X1 U22818 ( .A1(n20987), .A2(n20986), .ZN(P3_U2835) );
  NOR2_X1 U22819 ( .A1(n20995), .A2(n20988), .ZN(n20989) );
  AOI211_X1 U22820 ( .C1(n20991), .C2(n21063), .A(n20990), .B(n20989), .ZN(
        n21009) );
  NAND2_X1 U22821 ( .A1(n21093), .A2(n21008), .ZN(n21005) );
  AOI22_X1 U22822 ( .A1(n10958), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n21120), 
        .B2(n20992), .ZN(n21004) );
  OAI22_X1 U22823 ( .A1(n20996), .A2(n20995), .B1(n20994), .B2(n20993), .ZN(
        n21012) );
  AOI211_X1 U22824 ( .C1(n20998), .C2(n21047), .A(n20997), .B(n21012), .ZN(
        n21000) );
  NAND2_X1 U22825 ( .A1(n21000), .A2(n20999), .ZN(n21001) );
  OAI211_X1 U22826 ( .C1(n21002), .C2(n21001), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n21105), .ZN(n21003) );
  OAI211_X1 U22827 ( .C1(n21009), .C2(n21005), .A(n21004), .B(n21003), .ZN(
        P3_U2833) );
  AOI22_X1 U22828 ( .A1(n10958), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21006), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21014) );
  OAI21_X1 U22829 ( .B1(n21009), .B2(n21008), .A(n21007), .ZN(n21010) );
  OAI211_X1 U22830 ( .C1(n21012), .C2(n21011), .A(n21093), .B(n21010), .ZN(
        n21013) );
  OAI211_X1 U22831 ( .C1(n21015), .C2(n21110), .A(n21014), .B(n21013), .ZN(
        P3_U2832) );
  AOI21_X1 U22832 ( .B1(n21016), .B2(n21022), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21030) );
  NAND2_X1 U22833 ( .A1(n21019), .A2(n21017), .ZN(n21021) );
  NAND2_X1 U22834 ( .A1(n21019), .A2(n21018), .ZN(n21020) );
  AOI22_X1 U22835 ( .A1(n21063), .A2(n21021), .B1(n21125), .B2(n21020), .ZN(
        n21023) );
  NAND3_X1 U22836 ( .A1(n21024), .A2(n21023), .A3(n21022), .ZN(n21031) );
  NAND2_X1 U22837 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21025), .ZN(
        n21026) );
  OAI21_X1 U22838 ( .B1(n21031), .B2(n21026), .A(n21105), .ZN(n21037) );
  AOI21_X1 U22839 ( .B1(n21028), .B2(n21120), .A(n21027), .ZN(n21029) );
  OAI21_X1 U22840 ( .B1(n21030), .B2(n21037), .A(n21029), .ZN(P3_U2839) );
  OAI21_X1 U22841 ( .B1(n21085), .B2(n21031), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21036) );
  AOI22_X1 U22842 ( .A1(n21120), .A2(n21033), .B1(n21054), .B2(n21032), .ZN(
        n21035) );
  OAI211_X1 U22843 ( .C1(n21037), .C2(n21036), .A(n21035), .B(n21034), .ZN(
        P3_U2838) );
  AOI22_X1 U22844 ( .A1(n21063), .A2(n21039), .B1(n21125), .B2(n21038), .ZN(
        n21040) );
  NAND2_X1 U22845 ( .A1(n21041), .A2(n21040), .ZN(n21042) );
  OAI21_X1 U22846 ( .B1(n21043), .B2(n21042), .A(n21105), .ZN(n21049) );
  AOI22_X1 U22847 ( .A1(n21120), .A2(n21044), .B1(n21054), .B2(n21048), .ZN(
        n21046) );
  OAI211_X1 U22848 ( .C1(n21048), .C2(n21049), .A(n21046), .B(n21045), .ZN(
        P3_U2843) );
  NAND3_X1 U22849 ( .A1(n21048), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n21047), 
        .ZN(n21050) );
  NAND2_X1 U22850 ( .A1(n21050), .A2(n21049), .ZN(n21052) );
  OAI221_X1 U22851 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n21054), 
        .C1(n21053), .C2(n21052), .A(n21051), .ZN(n21056) );
  OAI211_X1 U22852 ( .C1(n21110), .C2(n21057), .A(n21056), .B(n21055), .ZN(
        P3_U2842) );
  NAND2_X1 U22853 ( .A1(n21058), .A2(n21101), .ZN(n21091) );
  NAND3_X1 U22854 ( .A1(n21060), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n21059), .ZN(n21070) );
  AOI211_X1 U22855 ( .C1(n21063), .C2(n21062), .A(n21065), .B(n21061), .ZN(
        n21067) );
  OAI21_X1 U22856 ( .B1(n21065), .B2(n21064), .A(n21126), .ZN(n21066) );
  OAI211_X1 U22857 ( .C1(n21068), .C2(n21067), .A(n21093), .B(n21066), .ZN(
        n21069) );
  AOI21_X1 U22858 ( .B1(n21112), .B2(n21070), .A(n21069), .ZN(n21078) );
  AOI221_X1 U22859 ( .B1(n21072), .B2(n21078), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n21078), .A(n21071), .ZN(
        n21073) );
  AOI22_X1 U22860 ( .A1(n21074), .A2(n21120), .B1(n21073), .B2(n21105), .ZN(
        n21076) );
  OAI211_X1 U22861 ( .C1(n21077), .C2(n21091), .A(n21076), .B(n21075), .ZN(
        P3_U2844) );
  NOR2_X1 U22862 ( .A1(n21090), .A2(n21091), .ZN(n21080) );
  OAI21_X1 U22863 ( .B1(n10958), .B2(n21078), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21079) );
  OAI21_X1 U22864 ( .B1(n21080), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n21079), .ZN(n21082) );
  OAI211_X1 U22865 ( .C1(n21083), .C2(n21110), .A(n21082), .B(n21081), .ZN(
        P3_U2845) );
  OAI221_X1 U22866 ( .B1(n21086), .B2(n21085), .C1(n21086), .C2(n21084), .A(
        n21105), .ZN(n21089) );
  AOI22_X1 U22867 ( .A1(n10958), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n21120), 
        .B2(n21087), .ZN(n21088) );
  OAI221_X1 U22868 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21091), 
        .C1(n21090), .C2(n21089), .A(n21088), .ZN(P3_U2846) );
  AOI22_X1 U22869 ( .A1(n10958), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21101), 
        .B2(n21092), .ZN(n21098) );
  OAI21_X1 U22870 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21094), .A(
        n21093), .ZN(n21095) );
  OAI211_X1 U22871 ( .C1(n21096), .C2(n21095), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21105), .ZN(n21097) );
  OAI211_X1 U22872 ( .C1(n21099), .C2(n21110), .A(n21098), .B(n21097), .ZN(
        P3_U2849) );
  NOR2_X1 U22873 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21115), .ZN(
        n21100) );
  AOI22_X1 U22874 ( .A1(n10958), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21101), 
        .B2(n21100), .ZN(n21109) );
  AOI22_X1 U22875 ( .A1(n21103), .A2(n21113), .B1(n21115), .B2(n21102), .ZN(
        n21104) );
  INV_X1 U22876 ( .A(n21104), .ZN(n21106) );
  OAI211_X1 U22877 ( .C1(n21107), .C2(n21106), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21105), .ZN(n21108) );
  OAI211_X1 U22878 ( .C1(n21111), .C2(n21110), .A(n21109), .B(n21108), .ZN(
        P3_U2852) );
  OAI21_X1 U22879 ( .B1(n21114), .B2(n21113), .A(n21112), .ZN(n21116) );
  AOI211_X1 U22880 ( .C1(n21117), .C2(n21116), .A(n10958), .B(n21115), .ZN(
        n21118) );
  AOI21_X1 U22881 ( .B1(n21120), .B2(n21119), .A(n21118), .ZN(n21122) );
  OAI211_X1 U22882 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21123), .A(
        n21122), .B(n21121), .ZN(P3_U2853) );
  NAND2_X1 U22883 ( .A1(n21687), .A2(n21177), .ZN(n21172) );
  INV_X1 U22884 ( .A(n21124), .ZN(n21171) );
  NOR2_X1 U22885 ( .A1(n21126), .A2(n21125), .ZN(n21128) );
  OAI222_X1 U22886 ( .A1(n21132), .A2(n21131), .B1(n21130), .B2(n21129), .C1(
        n21128), .C2(n21127), .ZN(n21190) );
  INV_X1 U22887 ( .A(n21133), .ZN(n21136) );
  AOI211_X1 U22888 ( .C1(n21136), .C2(n21649), .A(n21135), .B(n21134), .ZN(
        n21189) );
  OAI21_X1 U22889 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21189), .ZN(n21137) );
  OAI211_X1 U22890 ( .C1(n21141), .C2(n21139), .A(n21138), .B(n21137), .ZN(
        n21162) );
  AOI22_X1 U22891 ( .A1(n21151), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21140), .B2(n21141), .ZN(n21160) );
  AOI22_X1 U22892 ( .A1(n21151), .A2(n21143), .B1(n21142), .B2(n21141), .ZN(
        n21155) );
  OR3_X1 U22893 ( .A1(n21148), .A2(n21147), .A3(n21144), .ZN(n21145) );
  AOI22_X1 U22894 ( .A1(n21148), .A2(n21147), .B1(n21146), .B2(n21145), .ZN(
        n21150) );
  OAI21_X1 U22895 ( .B1(n21151), .B2(n21150), .A(n21149), .ZN(n21154) );
  AND2_X1 U22896 ( .A1(n21155), .A2(n21154), .ZN(n21152) );
  OAI221_X1 U22897 ( .B1(n21155), .B2(n21154), .C1(n21153), .C2(n21152), .A(
        n21157), .ZN(n21159) );
  AOI21_X1 U22898 ( .B1(n21157), .B2(n21156), .A(n21155), .ZN(n21158) );
  AOI222_X1 U22899 ( .A1(n21160), .A2(n21159), .B1(n21160), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21159), .C2(n21158), .ZN(
        n21161) );
  NOR4_X1 U22900 ( .A1(n21163), .A2(n21190), .A3(n21162), .A4(n21161), .ZN(
        n21187) );
  OAI211_X1 U22901 ( .C1(n21166), .C2(n21165), .A(n21164), .B(n21187), .ZN(
        n21175) );
  OAI21_X1 U22902 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21649), .A(n21175), 
        .ZN(n21181) );
  INV_X1 U22903 ( .A(n21181), .ZN(n21168) );
  NAND3_X1 U22904 ( .A1(n21169), .A2(n21168), .A3(n21167), .ZN(n21170) );
  NAND4_X1 U22905 ( .A1(n21173), .A2(n21172), .A3(n21171), .A4(n21170), .ZN(
        P3_U2997) );
  OAI221_X1 U22906 ( .B1(n21176), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21176), 
        .C2(n21175), .A(n21174), .ZN(P3_U3282) );
  AOI22_X1 U22907 ( .A1(n21179), .A2(n21178), .B1(n21687), .B2(n21177), .ZN(
        n21180) );
  INV_X1 U22908 ( .A(n21180), .ZN(n21184) );
  NOR2_X1 U22909 ( .A1(n21182), .A2(n21181), .ZN(n21183) );
  MUX2_X1 U22910 ( .A(n21184), .B(n21183), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21186) );
  OAI211_X1 U22911 ( .C1(n21187), .C2(n21188), .A(n21186), .B(n21185), .ZN(
        P3_U2996) );
  NOR2_X1 U22912 ( .A1(n21189), .A2(n21188), .ZN(n21193) );
  MUX2_X1 U22913 ( .A(P3_MORE_REG_SCAN_IN), .B(n21190), .S(n21193), .Z(
        P3_U3295) );
  OAI21_X1 U22914 ( .B1(n21193), .B2(n21192), .A(n21191), .ZN(P3_U2637) );
  AOI211_X1 U22915 ( .C1(n21195), .C2(n21881), .A(n21898), .B(n21194), .ZN(
        n21197) );
  OAI21_X1 U22916 ( .B1(n21197), .B2(n21614), .A(n21196), .ZN(n21202) );
  AOI211_X1 U22917 ( .C1(n21200), .C2(n21660), .A(n21199), .B(n21198), .ZN(
        n21201) );
  MUX2_X1 U22918 ( .A(n21202), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21201), 
        .Z(P1_U3485) );
  INV_X1 U22919 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21216) );
  NOR2_X1 U22920 ( .A1(n21216), .A2(n21203), .ZN(n21331) );
  AOI21_X1 U22921 ( .B1(n21316), .B2(n21331), .A(n21367), .ZN(n21210) );
  OAI21_X1 U22922 ( .B1(n21204), .B2(n21256), .A(n21300), .ZN(n21334) );
  AOI211_X1 U22923 ( .C1(n21206), .C2(n21205), .A(n21210), .B(n21334), .ZN(
        n21217) );
  NOR2_X1 U22924 ( .A1(n21373), .A2(n21207), .ZN(n21209) );
  AND2_X1 U22925 ( .A1(n21216), .A2(n21208), .ZN(n21221) );
  AOI211_X1 U22926 ( .C1(n21332), .C2(n21210), .A(n21209), .B(n21221), .ZN(
        n21215) );
  INV_X1 U22927 ( .A(n21211), .ZN(n21213) );
  AOI22_X1 U22928 ( .A1(n21213), .A2(n21393), .B1(n21382), .B2(n21212), .ZN(
        n21214) );
  OAI211_X1 U22929 ( .C1(n21217), .C2(n21216), .A(n21215), .B(n21214), .ZN(
        P1_U3018) );
  INV_X1 U22930 ( .A(n21217), .ZN(n21220) );
  NOR2_X1 U22931 ( .A1(n21373), .A2(n21218), .ZN(n21219) );
  AOI221_X1 U22932 ( .B1(n21221), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n21220), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n21219), .ZN(
        n21226) );
  NAND2_X1 U22933 ( .A1(n21316), .A2(n21265), .ZN(n21317) );
  NAND2_X1 U22934 ( .A1(n21222), .A2(n21317), .ZN(n21330) );
  AND2_X1 U22935 ( .A1(n21331), .A2(n21330), .ZN(n21223) );
  AOI22_X1 U22936 ( .A1(n21393), .A2(n21224), .B1(n21223), .B2(n13377), .ZN(
        n21225) );
  OAI211_X1 U22937 ( .C1(n21399), .C2(n21227), .A(n21226), .B(n21225), .ZN(
        P1_U3017) );
  NOR3_X1 U22938 ( .A1(n21228), .A2(n21230), .A3(n21256), .ZN(n21229) );
  AOI211_X1 U22939 ( .C1(n21230), .C2(n21297), .A(n21229), .B(n21312), .ZN(
        n21238) );
  NOR2_X1 U22940 ( .A1(n21373), .A2(n21231), .ZN(n21232) );
  NOR2_X1 U22941 ( .A1(n21256), .A2(n21241), .ZN(n21239) );
  AOI211_X1 U22942 ( .C1(n21382), .C2(n21233), .A(n21232), .B(n21239), .ZN(
        n21236) );
  AND2_X1 U22943 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21265), .ZN(
        n21242) );
  AOI22_X1 U22944 ( .A1(n21234), .A2(n21393), .B1(n21242), .B2(n21237), .ZN(
        n21235) );
  OAI211_X1 U22945 ( .C1(n21238), .C2(n21237), .A(n21236), .B(n21235), .ZN(
        P1_U3029) );
  NAND2_X1 U22946 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21240) );
  AOI211_X1 U22947 ( .C1(n21297), .C2(n21240), .A(n21239), .B(n21312), .ZN(
        n21252) );
  AOI22_X1 U22948 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21242), .B1(
        n21314), .B2(n21241), .ZN(n21253) );
  AOI211_X1 U22949 ( .C1(n21248), .C2(n13106), .A(n21253), .B(n21243), .ZN(
        n21245) );
  INV_X1 U22950 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21401) );
  OAI22_X1 U22951 ( .A1(n21399), .A2(n21405), .B1(n21401), .B2(n21373), .ZN(
        n21244) );
  AOI211_X1 U22952 ( .C1(n21246), .C2(n21393), .A(n21245), .B(n21244), .ZN(
        n21247) );
  OAI21_X1 U22953 ( .B1(n21252), .B2(n21248), .A(n21247), .ZN(P1_U3027) );
  AOI222_X1 U22954 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n13790), .B1(n21382), 
        .B2(n21250), .C1(n21393), .C2(n21249), .ZN(n21251) );
  OAI221_X1 U22955 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21253), .C1(
        n13106), .C2(n21252), .A(n21251), .ZN(P1_U3028) );
  INV_X1 U22956 ( .A(n21275), .ZN(n21255) );
  INV_X1 U22957 ( .A(n21254), .ZN(n21266) );
  AOI21_X1 U22958 ( .B1(n21314), .B2(n21266), .A(n21312), .ZN(n21276) );
  OAI21_X1 U22959 ( .B1(n21333), .B2(n21255), .A(n21276), .ZN(n21270) );
  AOI21_X1 U22960 ( .B1(n21265), .B2(n21264), .A(n21270), .ZN(n21263) );
  AOI22_X1 U22961 ( .A1(n13790), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n21382), 
        .B2(n21437), .ZN(n21261) );
  INV_X1 U22962 ( .A(n21265), .ZN(n21258) );
  INV_X1 U22963 ( .A(n21277), .ZN(n21257) );
  OAI22_X1 U22964 ( .A1(n21258), .A2(n21257), .B1(n21256), .B2(n21266), .ZN(
        n21293) );
  AOI22_X1 U22965 ( .A1(n21259), .A2(n21393), .B1(n21262), .B2(n21293), .ZN(
        n21260) );
  OAI211_X1 U22966 ( .C1(n21263), .C2(n21262), .A(n21261), .B(n21260), .ZN(
        P1_U3025) );
  NAND2_X1 U22967 ( .A1(n21265), .A2(n21264), .ZN(n21274) );
  NAND2_X1 U22968 ( .A1(n21314), .A2(n21266), .ZN(n21267) );
  OAI22_X1 U22969 ( .A1(n21373), .A2(n21432), .B1(n21268), .B2(n21267), .ZN(
        n21269) );
  AOI21_X1 U22970 ( .B1(n21382), .B2(n21419), .A(n21269), .ZN(n21273) );
  AOI22_X1 U22971 ( .A1(n21271), .A2(n21393), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21270), .ZN(n21272) );
  OAI211_X1 U22972 ( .C1(n21275), .C2(n21274), .A(n21273), .B(n21272), .ZN(
        P1_U3026) );
  NAND2_X1 U22973 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21293), .ZN(
        n21283) );
  OAI211_X1 U22974 ( .C1(n21333), .C2(n21277), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n21276), .ZN(n21278) );
  OAI21_X1 U22975 ( .B1(n21312), .B2(n21337), .A(n21278), .ZN(n21291) );
  OAI222_X1 U22976 ( .A1(n21458), .A2(n21399), .B1(n21373), .B2(n21453), .C1(
        n21353), .C2(n21279), .ZN(n21280) );
  INV_X1 U22977 ( .A(n21280), .ZN(n21281) );
  OAI221_X1 U22978 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21283), .C1(
        n21284), .C2(n21291), .A(n21281), .ZN(P1_U3024) );
  INV_X1 U22979 ( .A(n21282), .ZN(n21289) );
  AOI221_X1 U22980 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n21292), .C2(n21284), .A(
        n21283), .ZN(n21288) );
  OAI22_X1 U22981 ( .A1(n21286), .A2(n21399), .B1(n21285), .B2(n21373), .ZN(
        n21287) );
  AOI211_X1 U22982 ( .C1(n21289), .C2(n21393), .A(n21288), .B(n21287), .ZN(
        n21290) );
  OAI21_X1 U22983 ( .B1(n21292), .B2(n21291), .A(n21290), .ZN(P1_U3023) );
  NAND2_X1 U22984 ( .A1(n21294), .A2(n21293), .ZN(n21311) );
  AOI22_X1 U22985 ( .A1(n13790), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n21382), 
        .B2(n21464), .ZN(n21303) );
  INV_X1 U22986 ( .A(n21295), .ZN(n21301) );
  AOI22_X1 U22987 ( .A1(n21314), .A2(n21298), .B1(n21297), .B2(n21296), .ZN(
        n21299) );
  NAND2_X1 U22988 ( .A1(n21300), .A2(n21299), .ZN(n21307) );
  AOI22_X1 U22989 ( .A1(n21301), .A2(n21393), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21307), .ZN(n21302) );
  OAI211_X1 U22990 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21311), .A(
        n21303), .B(n21302), .ZN(P1_U3022) );
  OAI21_X1 U22991 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21304), .ZN(n21310) );
  AOI22_X1 U22992 ( .A1(n13790), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n21382), 
        .B2(n21305), .ZN(n21309) );
  AOI22_X1 U22993 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21307), .B1(
        n21393), .B2(n21306), .ZN(n21308) );
  OAI211_X1 U22994 ( .C1(n21311), .C2(n21310), .A(n21309), .B(n21308), .ZN(
        P1_U3021) );
  AOI21_X1 U22995 ( .B1(n21314), .B2(n21313), .A(n21312), .ZN(n21315) );
  OAI21_X1 U22996 ( .B1(n21333), .B2(n21316), .A(n21315), .ZN(n21327) );
  INV_X1 U22997 ( .A(n21327), .ZN(n21318) );
  AOI221_X1 U22998 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21318), 
        .C1(n21317), .C2(n21318), .A(n13214), .ZN(n21320) );
  INV_X1 U22999 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21487) );
  NOR2_X1 U23000 ( .A1(n21373), .A2(n21487), .ZN(n21319) );
  AOI211_X1 U23001 ( .C1(n21382), .C2(n21484), .A(n21320), .B(n21319), .ZN(
        n21322) );
  NAND3_X1 U23002 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n13214), .A3(
        n21330), .ZN(n21321) );
  OAI211_X1 U23003 ( .C1(n21323), .C2(n21353), .A(n21322), .B(n21321), .ZN(
        P1_U3019) );
  OAI21_X1 U23004 ( .B1(n21399), .B2(n21475), .A(n21324), .ZN(n21325) );
  AOI221_X1 U23005 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21327), 
        .C1(n21326), .C2(n21330), .A(n21325), .ZN(n21328) );
  OAI21_X1 U23006 ( .B1(n21329), .B2(n21353), .A(n21328), .ZN(P1_U3020) );
  NAND3_X1 U23007 ( .A1(n21331), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n21330), .ZN(n21357) );
  NOR2_X1 U23008 ( .A1(n21333), .A2(n21332), .ZN(n21335) );
  AOI211_X1 U23009 ( .C1(n21337), .C2(n21336), .A(n21335), .B(n21334), .ZN(
        n21363) );
  NAND2_X1 U23010 ( .A1(n13790), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n21338) );
  OAI221_X1 U23011 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21357), 
        .C1(n13217), .C2(n21363), .A(n21338), .ZN(n21339) );
  AOI21_X1 U23012 ( .B1(n21382), .B2(n21500), .A(n21339), .ZN(n21340) );
  OAI21_X1 U23013 ( .B1(n21341), .B2(n21353), .A(n21340), .ZN(P1_U3016) );
  NAND2_X1 U23014 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21355) );
  NOR2_X1 U23015 ( .A1(n21355), .A2(n21357), .ZN(n21350) );
  NAND2_X1 U23016 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21350), .ZN(
        n21347) );
  OAI21_X1 U23017 ( .B1(n21389), .B2(n21342), .A(n21363), .ZN(n21349) );
  NOR2_X1 U23018 ( .A1(n21373), .A2(n21535), .ZN(n21345) );
  OAI22_X1 U23019 ( .A1(n21343), .A2(n21353), .B1(n21399), .B2(n21528), .ZN(
        n21344) );
  AOI211_X1 U23020 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n21349), .A(
        n21345), .B(n21344), .ZN(n21346) );
  OAI21_X1 U23021 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21347), .A(
        n21346), .ZN(P1_U3013) );
  AOI22_X1 U23022 ( .A1(n13790), .A2(P1_REIP_REG_17__SCAN_IN), .B1(n21382), 
        .B2(n21348), .ZN(n21352) );
  OAI21_X1 U23023 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21350), .A(
        n21349), .ZN(n21351) );
  OAI211_X1 U23024 ( .C1(n21354), .C2(n21353), .A(n21352), .B(n21351), .ZN(
        P1_U3014) );
  OAI21_X1 U23025 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n21355), .ZN(n21356) );
  OAI22_X1 U23026 ( .A1(n21399), .A2(n21518), .B1(n21357), .B2(n21356), .ZN(
        n21358) );
  AOI21_X1 U23027 ( .B1(n21393), .B2(n21359), .A(n21358), .ZN(n21361) );
  NAND2_X1 U23028 ( .A1(n13790), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n21360) );
  OAI211_X1 U23029 ( .C1(n21363), .C2(n21362), .A(n21361), .B(n21360), .ZN(
        P1_U3015) );
  NOR2_X1 U23030 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21378), .ZN(
        n21365) );
  AOI22_X1 U23031 ( .A1(n13790), .A2(P1_REIP_REG_20__SCAN_IN), .B1(n21365), 
        .B2(n21364), .ZN(n21371) );
  OAI221_X1 U23032 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21367), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21366), .A(n21377), .ZN(
        n21369) );
  AOI22_X1 U23033 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21369), .B1(
        n21393), .B2(n21368), .ZN(n21370) );
  OAI211_X1 U23034 ( .C1(n21399), .C2(n21372), .A(n21371), .B(n21370), .ZN(
        P1_U3011) );
  OAI22_X1 U23035 ( .A1(n21373), .A2(n21537), .B1(n21399), .B2(n21543), .ZN(
        n21374) );
  AOI21_X1 U23036 ( .B1(n21393), .B2(n21375), .A(n21374), .ZN(n21376) );
  OAI221_X1 U23037 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21379), 
        .C1(n21378), .C2(n21377), .A(n21376), .ZN(P1_U3012) );
  AOI22_X1 U23038 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21381), .B1(
        n21393), .B2(n21380), .ZN(n21387) );
  NAND2_X1 U23039 ( .A1(n13790), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n21386) );
  NAND2_X1 U23040 ( .A1(n21382), .A2(n21550), .ZN(n21385) );
  INV_X1 U23041 ( .A(n21383), .ZN(n21384) );
  NAND4_X1 U23042 ( .A1(n21387), .A2(n21386), .A3(n21385), .A4(n21384), .ZN(
        P1_U3010) );
  NOR2_X1 U23043 ( .A1(n21389), .A2(n21388), .ZN(n21392) );
  INV_X1 U23044 ( .A(n21390), .ZN(n21391) );
  MUX2_X1 U23045 ( .A(n21392), .B(n21391), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21396) );
  AND3_X1 U23046 ( .A1(n13778), .A2(n21394), .A3(n21393), .ZN(n21395) );
  NOR2_X1 U23047 ( .A1(n21396), .A2(n21395), .ZN(n21398) );
  NAND2_X1 U23048 ( .A1(n13790), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21397) );
  OAI211_X1 U23049 ( .C1(n21400), .C2(n21399), .A(n21398), .B(n21397), .ZN(
        P1_U3030) );
  AOI21_X1 U23050 ( .B1(n21436), .B2(n21420), .A(n21435), .ZN(n21431) );
  NAND3_X1 U23051 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21402) );
  OAI21_X1 U23052 ( .B1(n21544), .B2(n21402), .A(n21401), .ZN(n21403) );
  INV_X1 U23053 ( .A(n21403), .ZN(n21415) );
  NAND2_X1 U23054 ( .A1(n21404), .A2(n21428), .ZN(n21414) );
  INV_X1 U23055 ( .A(n21405), .ZN(n21406) );
  NAND2_X1 U23056 ( .A1(n21605), .A2(n21406), .ZN(n21409) );
  NAND2_X1 U23057 ( .A1(n21597), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n21408) );
  AOI21_X1 U23058 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21519), .ZN(n21407) );
  NAND3_X1 U23059 ( .A1(n21409), .A2(n21408), .A3(n21407), .ZN(n21410) );
  AOI21_X1 U23060 ( .B1(n21412), .B2(n21411), .A(n21410), .ZN(n21413) );
  OAI211_X1 U23061 ( .C1(n21431), .C2(n21415), .A(n21414), .B(n21413), .ZN(
        n21416) );
  INV_X1 U23062 ( .A(n21416), .ZN(n21417) );
  OAI21_X1 U23063 ( .B1(n21418), .B2(n21600), .A(n21417), .ZN(P1_U2836) );
  INV_X1 U23064 ( .A(n21419), .ZN(n21426) );
  NOR3_X1 U23065 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21420), .A3(n21544), .ZN(
        n21421) );
  AOI211_X1 U23066 ( .C1(n21553), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21519), .B(n21421), .ZN(n21425) );
  INV_X1 U23067 ( .A(n21422), .ZN(n21423) );
  AOI22_X1 U23068 ( .A1(n21597), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n21423), .B2(
        n21586), .ZN(n21424) );
  OAI211_X1 U23069 ( .C1(n21592), .C2(n21426), .A(n21425), .B(n21424), .ZN(
        n21427) );
  AOI21_X1 U23070 ( .B1(n21429), .B2(n21428), .A(n21427), .ZN(n21430) );
  OAI21_X1 U23071 ( .B1(n21432), .B2(n21431), .A(n21430), .ZN(P1_U2835) );
  AND3_X1 U23072 ( .A1(n21436), .A2(n21445), .A3(n21433), .ZN(n21434) );
  AOI21_X1 U23073 ( .B1(n21597), .B2(P1_EBX_REG_6__SCAN_IN), .A(n21434), .ZN(
        n21443) );
  AOI21_X1 U23074 ( .B1(n21436), .B2(n21445), .A(n21435), .ZN(n21452) );
  INV_X1 U23075 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21439) );
  AOI22_X1 U23076 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21553), .B1(
        n21605), .B2(n21437), .ZN(n21438) );
  OAI211_X1 U23077 ( .C1(n21452), .C2(n21439), .A(n21438), .B(n21529), .ZN(
        n21440) );
  AOI21_X1 U23078 ( .B1(n21441), .B2(n21588), .A(n21440), .ZN(n21442) );
  OAI211_X1 U23079 ( .C1(n21444), .C2(n21600), .A(n21443), .B(n21442), .ZN(
        P1_U2834) );
  NAND2_X1 U23080 ( .A1(n21597), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n21448) );
  OR3_X1 U23081 ( .A1(n21544), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n21445), .ZN(
        n21447) );
  NAND2_X1 U23082 ( .A1(n21553), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n21446) );
  AND4_X1 U23083 ( .A1(n21448), .A2(n21447), .A3(n21529), .A4(n21446), .ZN(
        n21457) );
  INV_X1 U23084 ( .A(n21449), .ZN(n21450) );
  NAND2_X1 U23085 ( .A1(n21586), .A2(n21450), .ZN(n21451) );
  OAI21_X1 U23086 ( .B1(n21453), .B2(n21452), .A(n21451), .ZN(n21454) );
  AOI21_X1 U23087 ( .B1(n21455), .B2(n21588), .A(n21454), .ZN(n21456) );
  OAI211_X1 U23088 ( .C1(n21592), .C2(n21458), .A(n21457), .B(n21456), .ZN(
        P1_U2833) );
  INV_X1 U23089 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21460) );
  NAND2_X1 U23090 ( .A1(n21597), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n21459) );
  OAI211_X1 U23091 ( .C1(n21609), .C2(n21460), .A(n21459), .B(n21529), .ZN(
        n21463) );
  NOR3_X1 U23092 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21461), .A3(n21544), .ZN(
        n21462) );
  AOI211_X1 U23093 ( .C1(n21605), .C2(n21464), .A(n21463), .B(n21462), .ZN(
        n21465) );
  OAI21_X1 U23094 ( .B1(n21466), .B2(n21602), .A(n21465), .ZN(n21467) );
  AOI21_X1 U23095 ( .B1(n21468), .B2(n21586), .A(n21467), .ZN(n21469) );
  OAI21_X1 U23096 ( .B1(n21471), .B2(n21470), .A(n21469), .ZN(P1_U2831) );
  AOI22_X1 U23097 ( .A1(n21486), .A2(n21472), .B1(n21597), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n21479) );
  AOI22_X1 U23098 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n21553), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21473), .ZN(n21474) );
  OAI21_X1 U23099 ( .B1(n21592), .B2(n21475), .A(n21474), .ZN(n21476) );
  AOI211_X1 U23100 ( .C1(n21477), .C2(n21588), .A(n21519), .B(n21476), .ZN(
        n21478) );
  OAI211_X1 U23101 ( .C1(n21480), .C2(n21600), .A(n21479), .B(n21478), .ZN(
        P1_U2829) );
  INV_X1 U23102 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21482) );
  AOI21_X1 U23103 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21519), .ZN(n21481) );
  OAI21_X1 U23104 ( .B1(n21580), .B2(n21482), .A(n21481), .ZN(n21483) );
  AOI21_X1 U23105 ( .B1(n21484), .B2(n21605), .A(n21483), .ZN(n21492) );
  AOI211_X1 U23106 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n21485), .A(n21596), 
        .B(n21487), .ZN(n21489) );
  AND3_X1 U23107 ( .A1(n21487), .A2(P1_REIP_REG_11__SCAN_IN), .A3(n21486), 
        .ZN(n21488) );
  AOI211_X1 U23108 ( .C1(n21586), .C2(n21490), .A(n21489), .B(n21488), .ZN(
        n21491) );
  OAI211_X1 U23109 ( .C1(n21602), .C2(n21493), .A(n21492), .B(n21491), .ZN(
        P1_U2828) );
  NOR2_X1 U23110 ( .A1(n21495), .A2(n21494), .ZN(n21506) );
  AOI21_X1 U23111 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21507), .A(n21496), 
        .ZN(n21505) );
  INV_X1 U23112 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21498) );
  AOI21_X1 U23113 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21519), .ZN(n21497) );
  OAI21_X1 U23114 ( .B1(n21580), .B2(n21498), .A(n21497), .ZN(n21499) );
  AOI21_X1 U23115 ( .B1(n21500), .B2(n21605), .A(n21499), .ZN(n21504) );
  AOI22_X1 U23116 ( .A1(n21502), .A2(n21588), .B1(n21586), .B2(n21501), .ZN(
        n21503) );
  OAI211_X1 U23117 ( .C1(n21506), .C2(n21505), .A(n21504), .B(n21503), .ZN(
        P1_U2825) );
  AOI21_X1 U23118 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n21507), .A(n21506), 
        .ZN(n21509) );
  OAI22_X1 U23119 ( .A1(n21510), .A2(n21509), .B1(n21508), .B2(n21580), .ZN(
        n21511) );
  AOI211_X1 U23120 ( .C1(n21553), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21519), .B(n21511), .ZN(n21517) );
  INV_X1 U23121 ( .A(n21512), .ZN(n21513) );
  OAI22_X1 U23122 ( .A1(n21514), .A2(n21602), .B1(n21513), .B2(n21600), .ZN(
        n21515) );
  INV_X1 U23123 ( .A(n21515), .ZN(n21516) );
  OAI211_X1 U23124 ( .C1(n21592), .C2(n21518), .A(n21517), .B(n21516), .ZN(
        P1_U2824) );
  AOI21_X1 U23125 ( .B1(n21553), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21519), .ZN(n21520) );
  OAI21_X1 U23126 ( .B1(n21580), .B2(n21521), .A(n21520), .ZN(n21522) );
  AOI221_X1 U23127 ( .B1(n21534), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n21562), 
        .C2(n21535), .A(n21522), .ZN(n21527) );
  INV_X1 U23128 ( .A(n21523), .ZN(n21524) );
  AOI22_X1 U23129 ( .A1(n21525), .A2(n21588), .B1(n21524), .B2(n21586), .ZN(
        n21526) );
  OAI211_X1 U23130 ( .C1(n21592), .C2(n21528), .A(n21527), .B(n21526), .ZN(
        P1_U2822) );
  INV_X1 U23131 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21530) );
  OAI21_X1 U23132 ( .B1(n21609), .B2(n21530), .A(n21529), .ZN(n21533) );
  NOR2_X1 U23133 ( .A1(n21531), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n21532) );
  AOI211_X1 U23134 ( .C1(n21597), .C2(P1_EBX_REG_19__SCAN_IN), .A(n21533), .B(
        n21532), .ZN(n21542) );
  AOI21_X1 U23135 ( .B1(n21562), .B2(n21535), .A(n21534), .ZN(n21538) );
  OAI22_X1 U23136 ( .A1(n21538), .A2(n21537), .B1(n21536), .B2(n21600), .ZN(
        n21539) );
  AOI21_X1 U23137 ( .B1(n21540), .B2(n21588), .A(n21539), .ZN(n21541) );
  OAI211_X1 U23138 ( .C1(n21592), .C2(n21543), .A(n21542), .B(n21541), .ZN(
        P1_U2821) );
  NOR2_X1 U23139 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n21544), .ZN(n21560) );
  AOI22_X1 U23140 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n21559), .B1(n21545), 
        .B2(n21560), .ZN(n21547) );
  AOI22_X1 U23141 ( .A1(n21597), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21553), .ZN(n21546) );
  OAI211_X1 U23142 ( .C1(n21548), .C2(n21602), .A(n21547), .B(n21546), .ZN(
        n21549) );
  AOI21_X1 U23143 ( .B1(n21550), .B2(n21605), .A(n21549), .ZN(n21551) );
  OAI21_X1 U23144 ( .B1(n21552), .B2(n21600), .A(n21551), .ZN(P1_U2819) );
  AOI22_X1 U23145 ( .A1(n21597), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21553), .ZN(n21567) );
  INV_X1 U23146 ( .A(n21554), .ZN(n21555) );
  OAI22_X1 U23147 ( .A1(n21556), .A2(n21602), .B1(n21555), .B2(n21592), .ZN(
        n21557) );
  AOI21_X1 U23148 ( .B1(n21558), .B2(n21586), .A(n21557), .ZN(n21566) );
  OAI21_X1 U23149 ( .B1(n21560), .B2(n21559), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n21565) );
  NAND4_X1 U23150 ( .A1(n21563), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n21562), 
        .A4(n21561), .ZN(n21564) );
  NAND4_X1 U23151 ( .A1(n21567), .A2(n21566), .A3(n21565), .A4(n21564), .ZN(
        P1_U2818) );
  NOR2_X1 U23152 ( .A1(n21583), .A2(n21596), .ZN(n21584) );
  NAND2_X1 U23153 ( .A1(n21569), .A2(n21568), .ZN(n21570) );
  AOI22_X1 U23154 ( .A1(n21584), .A2(n21570), .B1(n21597), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n21577) );
  INV_X1 U23155 ( .A(n21571), .ZN(n21572) );
  OAI22_X1 U23156 ( .A1(n21573), .A2(n21602), .B1(n21572), .B2(n21600), .ZN(
        n21574) );
  AOI21_X1 U23157 ( .B1(n21575), .B2(n21605), .A(n21574), .ZN(n21576) );
  OAI211_X1 U23158 ( .C1(n15642), .C2(n21609), .A(n21577), .B(n21576), .ZN(
        P1_U2817) );
  OAI22_X1 U23159 ( .A1(n21580), .A2(n21579), .B1(n21609), .B2(n21578), .ZN(
        n21581) );
  AOI221_X1 U23160 ( .B1(n21584), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n21583), 
        .C2(n21582), .A(n21581), .ZN(n21591) );
  INV_X1 U23161 ( .A(n21585), .ZN(n21589) );
  AOI22_X1 U23162 ( .A1(n21589), .A2(n21588), .B1(n21587), .B2(n21586), .ZN(
        n21590) );
  OAI211_X1 U23163 ( .C1(n21593), .C2(n21592), .A(n21591), .B(n21590), .ZN(
        P1_U2816) );
  OAI21_X1 U23164 ( .B1(n21596), .B2(n21595), .A(n21594), .ZN(n21598) );
  AOI22_X1 U23165 ( .A1(n21599), .A2(n21598), .B1(n21597), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n21608) );
  OAI22_X1 U23166 ( .A1(n21603), .A2(n21602), .B1(n21601), .B2(n21600), .ZN(
        n21604) );
  AOI21_X1 U23167 ( .B1(n21606), .B2(n21605), .A(n21604), .ZN(n21607) );
  OAI211_X1 U23168 ( .C1(n15026), .C2(n21609), .A(n21608), .B(n21607), .ZN(
        P1_U2815) );
  OAI21_X1 U23169 ( .B1(n21612), .B2(n21611), .A(n21610), .ZN(P1_U2806) );
  NOR2_X1 U23170 ( .A1(n21614), .A2(n21613), .ZN(n21621) );
  INV_X1 U23171 ( .A(n21621), .ZN(n21616) );
  OAI22_X1 U23172 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21617), .B1(n21616), 
        .B2(n21615), .ZN(n21618) );
  NAND2_X1 U23173 ( .A1(n21619), .A2(n21618), .ZN(P1_U3163) );
  OAI21_X1 U23174 ( .B1(n21621), .B2(n21859), .A(n21620), .ZN(P1_U3466) );
  NAND2_X1 U23175 ( .A1(n21623), .A2(n21622), .ZN(n21629) );
  AOI22_X1 U23176 ( .A1(n21627), .A2(n21626), .B1(n21625), .B2(n21624), .ZN(
        n21628) );
  OAI21_X1 U23177 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21629), .A(n21628), 
        .ZN(n21630) );
  OAI21_X1 U23178 ( .B1(n21632), .B2(n21631), .A(n21630), .ZN(P1_U3161) );
  OAI21_X1 U23179 ( .B1(n21634), .B2(n21881), .A(n21633), .ZN(P1_U2805) );
  AOI21_X1 U23180 ( .B1(n21636), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21635), 
        .ZN(n21637) );
  INV_X1 U23181 ( .A(n21637), .ZN(P1_U3465) );
  INV_X1 U23182 ( .A(n21638), .ZN(n21640) );
  OAI21_X1 U23183 ( .B1(n21642), .B2(n21639), .A(n21640), .ZN(P2_U2818) );
  OAI21_X1 U23184 ( .B1(n21642), .B2(n21641), .A(n21640), .ZN(P2_U3592) );
  INV_X1 U23185 ( .A(n21643), .ZN(n21645) );
  OAI21_X1 U23186 ( .B1(n21647), .B2(n21644), .A(n21645), .ZN(P3_U2636) );
  OAI21_X1 U23187 ( .B1(n21647), .B2(n21646), .A(n21645), .ZN(P3_U3281) );
  INV_X1 U23188 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21688) );
  AOI21_X1 U23189 ( .B1(HOLD), .B2(n21648), .A(n21688), .ZN(n21650) );
  NOR2_X1 U23190 ( .A1(n21690), .A2(n21649), .ZN(n21700) );
  NOR2_X1 U23191 ( .A1(n21700), .A2(n21689), .ZN(n21704) );
  AOI21_X1 U23192 ( .B1(n21690), .B2(NA), .A(n21698), .ZN(n21702) );
  OAI22_X1 U23193 ( .A1(n18006), .A2(n21650), .B1(n21704), .B2(n21702), .ZN(
        P3_U3029) );
  NOR3_X1 U23194 ( .A1(NA), .A2(n21660), .A3(n21659), .ZN(n21653) );
  INV_X1 U23195 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21651) );
  AOI21_X1 U23196 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21651), .ZN(
        n21664) );
  AOI221_X1 U23197 ( .B1(NA), .B2(n21656), .C1(n21660), .C2(n21656), .A(n21664), .ZN(n21652) );
  AOI22_X1 U23198 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(n21653), .B1(HOLD), 
        .B2(n21652), .ZN(n21655) );
  INV_X1 U23199 ( .A(NA), .ZN(n21699) );
  OAI21_X1 U23200 ( .B1(n21659), .B2(n21660), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21661) );
  OAI211_X1 U23201 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21699), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21661), .ZN(n21654) );
  OAI21_X1 U23202 ( .B1(n21655), .B2(n13264), .A(n21654), .ZN(P1_U3196) );
  AOI22_X1 U23203 ( .A1(n21656), .A2(HOLD), .B1(P1_STATE_REG_0__SCAN_IN), .B2(
        n21664), .ZN(n21658) );
  OAI211_X1 U23204 ( .C1(n21660), .C2(n21659), .A(n21658), .B(n21657), .ZN(
        P1_U3195) );
  AOI22_X1 U23205 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(NA), .B2(
        n13264), .ZN(n21663) );
  NAND2_X1 U23206 ( .A1(n12962), .A2(n21661), .ZN(n21662) );
  OAI221_X1 U23207 ( .B1(n22319), .B2(n21664), .C1(n22319), .C2(n21663), .A(
        n21662), .ZN(P1_U3194) );
  NAND2_X1 U23208 ( .A1(n21665), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21674) );
  NAND2_X1 U23209 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21674), .ZN(n21678) );
  AOI22_X1 U23210 ( .A1(n21682), .A2(n21678), .B1(n21676), .B2(n17124), .ZN(
        n21668) );
  OAI211_X1 U23211 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(P2_STATE_REG_1__SCAN_IN), .A(HOLD), .B(n21666), .ZN(n21667) );
  OAI211_X1 U23212 ( .C1(n21699), .C2(n21679), .A(n21668), .B(n21667), .ZN(
        P2_U3209) );
  INV_X1 U23213 ( .A(HOLD), .ZN(n21697) );
  NAND2_X1 U23214 ( .A1(n21697), .A2(n21676), .ZN(n21673) );
  AOI211_X1 U23215 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21685), .B(
        n21676), .ZN(n21670) );
  AOI211_X1 U23216 ( .C1(n21671), .C2(n21673), .A(n21670), .B(n21669), .ZN(
        n21672) );
  NAND2_X1 U23217 ( .A1(n21672), .A2(n21674), .ZN(P2_U3210) );
  INV_X1 U23218 ( .A(n21673), .ZN(n21684) );
  OAI22_X1 U23219 ( .A1(NA), .A2(n21674), .B1(n21682), .B2(n21697), .ZN(n21675) );
  AOI21_X1 U23220 ( .B1(n21677), .B2(n21676), .A(n21675), .ZN(n21683) );
  INV_X1 U23221 ( .A(n21678), .ZN(n21681) );
  NOR2_X1 U23222 ( .A1(n21679), .A2(n21699), .ZN(n21680) );
  OAI33_X1 U23223 ( .A1(n21685), .A2(n21684), .A3(n21683), .B1(n21682), .B2(
        n21681), .B3(n21680), .ZN(P2_U3211) );
  AOI21_X1 U23224 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21690), .ZN(
        n21686) );
  NAND2_X1 U23225 ( .A1(n21697), .A2(n21688), .ZN(n21696) );
  AOI21_X1 U23226 ( .B1(n21686), .B2(n21696), .A(n21700), .ZN(n21694) );
  OAI21_X1 U23227 ( .B1(n21687), .B2(n21698), .A(n18006), .ZN(n21693) );
  AOI211_X1 U23228 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21689), .B(
        n21688), .ZN(n21691) );
  OAI21_X1 U23229 ( .B1(n21695), .B2(n21691), .A(n21690), .ZN(n21692) );
  OAI211_X1 U23230 ( .C1(n21695), .C2(n21694), .A(n21693), .B(n21692), .ZN(
        P3_U3030) );
  INV_X1 U23231 ( .A(n21696), .ZN(n21706) );
  OAI22_X1 U23232 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21698), .B2(n21697), .ZN(n21701)
         );
  OAI221_X1 U23233 ( .B1(n21701), .B2(n21700), .C1(n21701), .C2(n21699), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21705) );
  INV_X1 U23234 ( .A(n21702), .ZN(n21703) );
  OAI22_X1 U23235 ( .A1(n21706), .A2(n21705), .B1(n21704), .B2(n21703), .ZN(
        P3_U3031) );
  INV_X1 U23236 ( .A(n13672), .ZN(n21707) );
  INV_X1 U23237 ( .A(n22314), .ZN(n21708) );
  OR2_X1 U23238 ( .A1(n14068), .A2(n21707), .ZN(n21763) );
  OR2_X1 U23239 ( .A1(n21753), .A2(n21763), .ZN(n21725) );
  NAND3_X1 U23240 ( .A1(n21708), .A2(n21872), .A3(n21725), .ZN(n21709) );
  NAND2_X1 U23241 ( .A1(n21872), .A2(n21881), .ZN(n21847) );
  NAND2_X1 U23242 ( .A1(n21709), .A2(n21847), .ZN(n21722) );
  OR2_X1 U23243 ( .A1(n21804), .A2(n21710), .ZN(n21750) );
  NOR2_X1 U23244 ( .A1(n21750), .A2(n21884), .ZN(n21719) );
  NOR2_X1 U23245 ( .A1(n21717), .A2(n21898), .ZN(n21825) );
  INV_X1 U23246 ( .A(n21739), .ZN(n21824) );
  OR2_X1 U23247 ( .A1(n21806), .A2(n21824), .ZN(n21765) );
  INV_X1 U23248 ( .A(n21765), .ZN(n21724) );
  AOI22_X1 U23249 ( .A1(n21722), .A2(n21719), .B1(n21825), .B2(n21724), .ZN(
        n22212) );
  NAND2_X1 U23250 ( .A1(n22199), .A2(n21711), .ZN(n21862) );
  NAND2_X1 U23251 ( .A1(n19952), .A2(n15237), .ZN(n22207) );
  INV_X1 U23252 ( .A(DATAI_24_), .ZN(n21713) );
  OAI22_X1 U23253 ( .A1(n21714), .A2(n22207), .B1(n21713), .B2(n22205), .ZN(
        n21889) );
  NOR2_X2 U23254 ( .A1(n22203), .A2(n21716), .ZN(n21901) );
  NOR3_X1 U23255 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21735) );
  INV_X1 U23256 ( .A(n21735), .ZN(n21732) );
  NOR2_X1 U23257 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21732), .ZN(
        n22204) );
  AOI22_X1 U23258 ( .A1(n22314), .A2(n11069), .B1(n21901), .B2(n22204), .ZN(
        n21729) );
  INV_X1 U23259 ( .A(n21717), .ZN(n21718) );
  NOR2_X1 U23260 ( .A1(n21718), .A2(n21898), .ZN(n21852) );
  INV_X1 U23261 ( .A(n22199), .ZN(n21769) );
  NOR2_X1 U23262 ( .A1(n21852), .A2(n21769), .ZN(n21832) );
  INV_X1 U23263 ( .A(n21719), .ZN(n21721) );
  INV_X1 U23264 ( .A(n22204), .ZN(n21720) );
  AOI22_X1 U23265 ( .A1(n21722), .A2(n21721), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21720), .ZN(n21723) );
  OAI211_X1 U23266 ( .C1(n21724), .C2(n21898), .A(n21832), .B(n21723), .ZN(
        n22209) );
  OAI22_X1 U23267 ( .A1(n21727), .A2(n22207), .B1(n21726), .B2(n22205), .ZN(
        n21909) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n21909), .ZN(n21728) );
  OAI211_X1 U23269 ( .C1(n22212), .C2(n21862), .A(n21729), .B(n21728), .ZN(
        P1_U3033) );
  INV_X1 U23270 ( .A(n21909), .ZN(n21892) );
  INV_X1 U23271 ( .A(n21750), .ZN(n21731) );
  INV_X1 U23272 ( .A(n21730), .ZN(n21865) );
  NOR2_X1 U23273 ( .A1(n21864), .A2(n21732), .ZN(n22213) );
  AOI21_X1 U23274 ( .B1(n21731), .B2(n21865), .A(n22213), .ZN(n21733) );
  OAI22_X1 U23275 ( .A1(n21733), .A2(n21900), .B1(n21732), .B2(n21898), .ZN(
        n22214) );
  INV_X1 U23276 ( .A(n21862), .ZN(n21902) );
  AOI22_X1 U23277 ( .A1(n22214), .A2(n21902), .B1(n21901), .B2(n22213), .ZN(
        n21737) );
  OAI21_X1 U23278 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21859), .A(
        n22199), .ZN(n21903) );
  OAI211_X1 U23279 ( .C1(n21753), .C2(n21881), .A(n21908), .B(n21733), .ZN(
        n21734) );
  OAI211_X1 U23280 ( .C1(n21908), .C2(n21735), .A(n21869), .B(n21734), .ZN(
        n22216) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n11069), .ZN(n21736) );
  OAI211_X1 U23282 ( .C1(n21892), .C2(n22219), .A(n21737), .B(n21736), .ZN(
        P1_U3041) );
  INV_X1 U23283 ( .A(n21876), .ZN(n21822) );
  NAND3_X1 U23284 ( .A1(n22221), .A2(n22219), .A3(n21908), .ZN(n21738) );
  NAND2_X1 U23285 ( .A1(n21738), .A2(n21847), .ZN(n21741) );
  NOR2_X1 U23286 ( .A1(n21750), .A2(n21805), .ZN(n21743) );
  NOR2_X1 U23287 ( .A1(n21739), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21783) );
  AOI22_X1 U23288 ( .A1(n21741), .A2(n21743), .B1(n21825), .B2(n21783), .ZN(
        n22227) );
  INV_X1 U23289 ( .A(n21901), .ZN(n21754) );
  NOR3_X1 U23290 ( .A1(n21827), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21747) );
  NAND2_X1 U23291 ( .A1(n21864), .A2(n21747), .ZN(n22220) );
  OAI22_X1 U23292 ( .A1(n22221), .A2(n21892), .B1(n21754), .B2(n22220), .ZN(
        n21740) );
  INV_X1 U23293 ( .A(n21740), .ZN(n21746) );
  INV_X1 U23294 ( .A(n21741), .ZN(n21744) );
  NOR2_X1 U23295 ( .A1(n21783), .A2(n21898), .ZN(n21785) );
  AOI21_X1 U23296 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22220), .A(n21785), 
        .ZN(n21742) );
  OAI211_X1 U23297 ( .C1(n21744), .C2(n21743), .A(n21742), .B(n21832), .ZN(
        n22224) );
  INV_X1 U23298 ( .A(n22219), .ZN(n22223) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22224), .B1(
        n22223), .B2(n11069), .ZN(n21745) );
  OAI211_X1 U23300 ( .C1(n22227), .C2(n21862), .A(n21746), .B(n21745), .ZN(
        P1_U3049) );
  INV_X1 U23301 ( .A(n21747), .ZN(n21757) );
  AND2_X1 U23302 ( .A1(n21749), .A2(n21748), .ZN(n21894) );
  INV_X1 U23303 ( .A(n21894), .ZN(n21795) );
  OR2_X1 U23304 ( .A1(n21750), .A2(n21795), .ZN(n21751) );
  OR2_X1 U23305 ( .A1(n21864), .A2(n21757), .ZN(n22228) );
  AND2_X1 U23306 ( .A1(n21751), .A2(n22228), .ZN(n21756) );
  OAI21_X1 U23307 ( .B1(n21753), .B2(n21838), .A(n21872), .ZN(n21760) );
  OAI22_X1 U23308 ( .A1(n21898), .A2(n21757), .B1(n21756), .B2(n21760), .ZN(
        n21752) );
  INV_X1 U23309 ( .A(n21791), .ZN(n21841) );
  OAI22_X1 U23310 ( .A1(n22230), .A2(n21892), .B1(n21754), .B2(n22228), .ZN(
        n21755) );
  INV_X1 U23311 ( .A(n21755), .ZN(n21762) );
  INV_X1 U23312 ( .A(n21756), .ZN(n21759) );
  AOI21_X1 U23313 ( .B1(n21900), .B2(n21757), .A(n21903), .ZN(n21758) );
  OAI21_X1 U23314 ( .B1(n21760), .B2(n21759), .A(n21758), .ZN(n22233) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22233), .B1(
        n22232), .B2(n11069), .ZN(n21761) );
  OAI211_X1 U23316 ( .C1(n22236), .C2(n21862), .A(n21762), .B(n21761), .ZN(
        P1_U3057) );
  NOR3_X1 U23317 ( .A1(n21853), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21777) );
  INV_X1 U23318 ( .A(n21777), .ZN(n21773) );
  NOR2_X1 U23319 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21773), .ZN(
        n22238) );
  OR2_X1 U23320 ( .A1(n21850), .A2(n21764), .ZN(n21782) );
  INV_X1 U23321 ( .A(n21782), .ZN(n21767) );
  NAND2_X1 U23322 ( .A1(n21767), .A2(n21872), .ZN(n21796) );
  INV_X1 U23323 ( .A(n21852), .ZN(n21880) );
  OAI22_X1 U23324 ( .A1(n21796), .A2(n21884), .B1(n21765), .B2(n21880), .ZN(
        n22237) );
  AOI22_X1 U23325 ( .A1(n21901), .A2(n22238), .B1(n21902), .B2(n22237), .ZN(
        n21772) );
  AOI21_X1 U23326 ( .B1(n22230), .B2(n22248), .A(n21881), .ZN(n21766) );
  AOI21_X1 U23327 ( .B1(n21767), .B2(n21805), .A(n21766), .ZN(n21768) );
  NOR2_X1 U23328 ( .A1(n21768), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21770) );
  NOR2_X1 U23329 ( .A1(n21825), .A2(n21769), .ZN(n21887) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n11069), .ZN(n21771) );
  OAI211_X1 U23331 ( .C1(n21892), .C2(n22248), .A(n21772), .B(n21771), .ZN(
        P1_U3065) );
  NOR2_X1 U23332 ( .A1(n21864), .A2(n21773), .ZN(n22243) );
  INV_X1 U23333 ( .A(n22243), .ZN(n21774) );
  OAI222_X1 U23334 ( .A1(n21774), .A2(n21900), .B1(n21898), .B2(n21773), .C1(
        n21730), .C2(n21796), .ZN(n22244) );
  AOI22_X1 U23335 ( .A1(n22244), .A2(n21902), .B1(n21901), .B2(n22243), .ZN(
        n21779) );
  INV_X1 U23336 ( .A(n21792), .ZN(n21775) );
  NOR3_X1 U23337 ( .A1(n21775), .A2(n21900), .A3(n21881), .ZN(n21776) );
  OAI21_X1 U23338 ( .B1(n21777), .B2(n21776), .A(n21869), .ZN(n22245) );
  INV_X1 U23339 ( .A(n21819), .ZN(n21873) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n21909), .ZN(n21778) );
  OAI211_X1 U23341 ( .C1(n11068), .C2(n22248), .A(n21779), .B(n21778), .ZN(
        P1_U3073) );
  INV_X1 U23342 ( .A(n22250), .ZN(n21780) );
  NAND2_X1 U23343 ( .A1(n21780), .A2(n21872), .ZN(n21781) );
  OAI21_X1 U23344 ( .B1(n21781), .B2(n22257), .A(n21847), .ZN(n21787) );
  NOR2_X1 U23345 ( .A1(n21782), .A2(n21805), .ZN(n21784) );
  AOI22_X1 U23346 ( .A1(n21787), .A2(n21784), .B1(n21783), .B2(n21852), .ZN(
        n22254) );
  AOI22_X1 U23347 ( .A1(n22250), .A2(n11069), .B1(n21901), .B2(n22249), .ZN(
        n21790) );
  INV_X1 U23348 ( .A(n21784), .ZN(n21786) );
  AOI21_X1 U23349 ( .B1(n21787), .B2(n21786), .A(n21785), .ZN(n21788) );
  OAI211_X1 U23350 ( .C1(n22249), .C2(n21859), .A(n21887), .B(n21788), .ZN(
        n22251) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22251), .B1(
        n22257), .B2(n21909), .ZN(n21789) );
  OAI211_X1 U23352 ( .C1(n22254), .C2(n21862), .A(n21790), .B(n21789), .ZN(
        P1_U3081) );
  NAND2_X1 U23353 ( .A1(n21792), .A2(n21791), .ZN(n22261) );
  INV_X1 U23354 ( .A(n21793), .ZN(n22256) );
  NOR2_X1 U23355 ( .A1(n21896), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21798) );
  INV_X1 U23356 ( .A(n21798), .ZN(n21794) );
  OAI222_X1 U23357 ( .A1(n21796), .A2(n21795), .B1(n21898), .B2(n21794), .C1(
        n21793), .C2(n21900), .ZN(n22255) );
  AOI22_X1 U23358 ( .A1(n21901), .A2(n22256), .B1(n22255), .B2(n21902), .ZN(
        n21800) );
  OAI21_X1 U23359 ( .B1(n21798), .B2(n21797), .A(n21869), .ZN(n22258) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n11069), .ZN(n21799) );
  OAI211_X1 U23361 ( .C1(n21892), .C2(n22261), .A(n21800), .B(n21799), .ZN(
        P1_U3089) );
  INV_X1 U23362 ( .A(n10980), .ZN(n21801) );
  NAND2_X1 U23363 ( .A1(n21802), .A2(n21801), .ZN(n21842) );
  INV_X1 U23364 ( .A(n21842), .ZN(n21803) );
  AND2_X1 U23365 ( .A1(n21804), .A2(n21850), .ZN(n21835) );
  NOR3_X1 U23366 ( .A1(n21897), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21818) );
  INV_X1 U23367 ( .A(n21818), .ZN(n21815) );
  NOR2_X1 U23368 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21815), .ZN(
        n22262) );
  AOI21_X1 U23369 ( .B1(n21835), .B2(n21805), .A(n22262), .ZN(n21810) );
  INV_X1 U23370 ( .A(n21825), .ZN(n21808) );
  INV_X1 U23371 ( .A(n21806), .ZN(n21807) );
  NOR2_X1 U23372 ( .A1(n21807), .A2(n21824), .ZN(n21851) );
  INV_X1 U23373 ( .A(n21851), .ZN(n21855) );
  OAI22_X1 U23374 ( .A1(n21810), .A2(n21900), .B1(n21808), .B2(n21855), .ZN(
        n22263) );
  AOI22_X1 U23375 ( .A1(n22263), .A2(n21902), .B1(n21901), .B2(n22262), .ZN(
        n21814) );
  INV_X1 U23376 ( .A(n22273), .ZN(n21809) );
  OAI21_X1 U23377 ( .B1(n21809), .B2(n22264), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21811) );
  NAND2_X1 U23378 ( .A1(n21811), .A2(n21810), .ZN(n21812) );
  OAI211_X1 U23379 ( .C1(n22262), .C2(n21859), .A(n21832), .B(n21812), .ZN(
        n22265) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n11069), .ZN(n21813) );
  OAI211_X1 U23381 ( .C1(n21892), .C2(n22273), .A(n21814), .B(n21813), .ZN(
        P1_U3097) );
  NOR2_X1 U23382 ( .A1(n21864), .A2(n21815), .ZN(n22268) );
  AOI21_X1 U23383 ( .B1(n21835), .B2(n21865), .A(n22268), .ZN(n21816) );
  OAI22_X1 U23384 ( .A1(n21816), .A2(n21900), .B1(n21815), .B2(n21898), .ZN(
        n22269) );
  AOI22_X1 U23385 ( .A1(n22269), .A2(n21902), .B1(n21901), .B2(n22268), .ZN(
        n21821) );
  OAI211_X1 U23386 ( .C1(n21842), .C2(n21881), .A(n21908), .B(n21816), .ZN(
        n21817) );
  OAI211_X1 U23387 ( .C1(n21908), .C2(n21818), .A(n21869), .B(n21817), .ZN(
        n22270) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n21909), .ZN(n21820) );
  OAI211_X1 U23389 ( .C1(n11068), .C2(n22273), .A(n21821), .B(n21820), .ZN(
        P1_U3105) );
  NAND3_X1 U23390 ( .A1(n22286), .A2(n22178), .A3(n21872), .ZN(n21823) );
  NAND2_X1 U23391 ( .A1(n21823), .A2(n21847), .ZN(n21830) );
  AND2_X1 U23392 ( .A1(n21835), .A2(n21884), .ZN(n21828) );
  NAND2_X1 U23393 ( .A1(n21824), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21879) );
  INV_X1 U23394 ( .A(n21879), .ZN(n21826) );
  AOI22_X1 U23395 ( .A1(n21830), .A2(n21828), .B1(n21826), .B2(n21825), .ZN(
        n22280) );
  NOR3_X1 U23396 ( .A1(n21897), .A2(n21827), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21840) );
  NAND2_X1 U23397 ( .A1(n21864), .A2(n21840), .ZN(n22177) );
  INV_X1 U23398 ( .A(n22177), .ZN(n22274) );
  AOI22_X1 U23399 ( .A1(n22275), .A2(n11069), .B1(n21901), .B2(n22274), .ZN(
        n21834) );
  INV_X1 U23400 ( .A(n21828), .ZN(n21829) );
  AOI22_X1 U23401 ( .A1(n21830), .A2(n21829), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22177), .ZN(n21831) );
  NAND2_X1 U23402 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21879), .ZN(n21886) );
  NAND3_X1 U23403 ( .A1(n21832), .A2(n21831), .A3(n21886), .ZN(n22277) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n21909), .ZN(n21833) );
  OAI211_X1 U23405 ( .C1(n22280), .C2(n21862), .A(n21834), .B(n21833), .ZN(
        P1_U3113) );
  INV_X1 U23406 ( .A(n21840), .ZN(n21836) );
  NOR2_X1 U23407 ( .A1(n21864), .A2(n21836), .ZN(n22281) );
  AOI21_X1 U23408 ( .B1(n21835), .B2(n21894), .A(n22281), .ZN(n21837) );
  OAI22_X1 U23409 ( .A1(n21837), .A2(n21900), .B1(n21836), .B2(n21898), .ZN(
        n22282) );
  AOI22_X1 U23410 ( .A1(n22282), .A2(n21902), .B1(n21901), .B2(n22281), .ZN(
        n21844) );
  OAI211_X1 U23411 ( .C1(n21842), .C2(n21838), .A(n21908), .B(n21837), .ZN(
        n21839) );
  OAI211_X1 U23412 ( .C1(n21908), .C2(n21840), .A(n21869), .B(n21839), .ZN(
        n22283) );
  OR2_X1 U23413 ( .A1(n21842), .A2(n21841), .ZN(n21846) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n21909), .ZN(n21843) );
  OAI211_X1 U23415 ( .C1(n11068), .C2(n22286), .A(n21844), .B(n21843), .ZN(
        P1_U3121) );
  NAND3_X1 U23416 ( .A1(n21846), .A2(n21908), .A3(n22300), .ZN(n21848) );
  NAND2_X1 U23417 ( .A1(n21848), .A2(n21847), .ZN(n21857) );
  OR2_X1 U23418 ( .A1(n21850), .A2(n21849), .ZN(n21863) );
  NOR2_X1 U23419 ( .A1(n21863), .A2(n21884), .ZN(n21854) );
  AOI22_X1 U23420 ( .A1(n21857), .A2(n21854), .B1(n21852), .B2(n21851), .ZN(
        n22294) );
  INV_X1 U23421 ( .A(n22300), .ZN(n22288) );
  NOR3_X1 U23422 ( .A1(n21853), .A2(n21897), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21871) );
  INV_X1 U23423 ( .A(n21871), .ZN(n21866) );
  NOR2_X1 U23424 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21866), .ZN(
        n22287) );
  AOI22_X1 U23425 ( .A1(n22288), .A2(n21909), .B1(n21901), .B2(n22287), .ZN(
        n21861) );
  INV_X1 U23426 ( .A(n21854), .ZN(n21856) );
  AOI22_X1 U23427 ( .A1(n21857), .A2(n21856), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21855), .ZN(n21858) );
  OAI211_X1 U23428 ( .C1(n22287), .C2(n21859), .A(n21887), .B(n21858), .ZN(
        n22290) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n11069), .ZN(n21860) );
  OAI211_X1 U23430 ( .C1(n22294), .C2(n21862), .A(n21861), .B(n21860), .ZN(
        P1_U3129) );
  NOR2_X1 U23431 ( .A1(n21864), .A2(n21866), .ZN(n22295) );
  AOI21_X1 U23432 ( .B1(n21895), .B2(n21865), .A(n22295), .ZN(n21867) );
  OAI22_X1 U23433 ( .A1(n21867), .A2(n21900), .B1(n21866), .B2(n21898), .ZN(
        n22296) );
  AOI22_X1 U23434 ( .A1(n22296), .A2(n21902), .B1(n21901), .B2(n22295), .ZN(
        n21875) );
  INV_X1 U23435 ( .A(n21877), .ZN(n21868) );
  OAI21_X1 U23436 ( .B1(n21868), .B2(n21881), .A(n21867), .ZN(n21870) );
  OAI221_X1 U23437 ( .B1(n21872), .B2(n21871), .C1(n21900), .C2(n21870), .A(
        n21869), .ZN(n22297) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n21909), .ZN(n21874) );
  OAI211_X1 U23439 ( .C1(n11068), .C2(n22300), .A(n21875), .B(n21874), .ZN(
        P1_U3137) );
  NOR3_X2 U23440 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21897), .A3(
        n21896), .ZN(n22302) );
  NAND3_X1 U23441 ( .A1(n21895), .A2(n21884), .A3(n21908), .ZN(n21878) );
  OAI21_X1 U23442 ( .B1(n21880), .B2(n21879), .A(n21878), .ZN(n22301) );
  AOI22_X1 U23443 ( .A1(n21901), .A2(n22302), .B1(n21902), .B2(n22301), .ZN(
        n21891) );
  INV_X1 U23444 ( .A(n22304), .ZN(n21882) );
  AOI21_X1 U23445 ( .B1(n21882), .B2(n22318), .A(n21881), .ZN(n21883) );
  AOI21_X1 U23446 ( .B1(n21895), .B2(n21884), .A(n21883), .ZN(n21885) );
  NOR2_X1 U23447 ( .A1(n21885), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21888) );
  OAI211_X1 U23448 ( .C1(n22302), .C2(n21888), .A(n21887), .B(n21886), .ZN(
        n22305) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n11069), .ZN(n21890) );
  OAI211_X1 U23450 ( .C1(n21892), .C2(n22318), .A(n21891), .B(n21890), .ZN(
        P1_U3145) );
  NOR2_X1 U23451 ( .A1(n21893), .A2(n21897), .ZN(n22309) );
  AOI21_X1 U23452 ( .B1(n21895), .B2(n21894), .A(n22309), .ZN(n21904) );
  NOR2_X1 U23453 ( .A1(n21897), .A2(n21896), .ZN(n21907) );
  INV_X1 U23454 ( .A(n21907), .ZN(n21899) );
  OAI22_X1 U23455 ( .A1(n21904), .A2(n21900), .B1(n21899), .B2(n21898), .ZN(
        n22312) );
  AOI22_X1 U23456 ( .A1(n22312), .A2(n21902), .B1(n21901), .B2(n22309), .ZN(
        n21911) );
  AOI21_X1 U23457 ( .B1(n21905), .B2(n21904), .A(n21903), .ZN(n21906) );
  OAI21_X1 U23458 ( .B1(n21908), .B2(n21907), .A(n21906), .ZN(n22315) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n21909), .ZN(n21910) );
  OAI211_X1 U23460 ( .C1(n11068), .C2(n22318), .A(n21911), .B(n21910), .ZN(
        P1_U3153) );
  NAND2_X1 U23461 ( .A1(n22199), .A2(n21912), .ZN(n21947) );
  INV_X1 U23462 ( .A(DATAI_25_), .ZN(n21913) );
  NOR2_X2 U23463 ( .A1(n22203), .A2(n21915), .ZN(n21953) );
  AOI22_X1 U23464 ( .A1(n22314), .A2(n21950), .B1(n21953), .B2(n22204), .ZN(
        n21919) );
  OAI22_X1 U23465 ( .A1(n21917), .A2(n22207), .B1(n21916), .B2(n22205), .ZN(
        n21955) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n11061), .ZN(n21918) );
  OAI211_X1 U23467 ( .C1(n22212), .C2(n21947), .A(n21919), .B(n21918), .ZN(
        P1_U3034) );
  INV_X1 U23468 ( .A(n21947), .ZN(n21954) );
  AOI22_X1 U23469 ( .A1(n22214), .A2(n21954), .B1(n21953), .B2(n22213), .ZN(
        n21921) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n21950), .ZN(n21920) );
  OAI211_X1 U23471 ( .C1(n11060), .C2(n22219), .A(n21921), .B(n21920), .ZN(
        P1_U3042) );
  INV_X1 U23472 ( .A(n21950), .ZN(n21958) );
  INV_X1 U23473 ( .A(n21953), .ZN(n21925) );
  OAI22_X1 U23474 ( .A1(n22219), .A2(n21958), .B1(n21925), .B2(n22220), .ZN(
        n21922) );
  INV_X1 U23475 ( .A(n21922), .ZN(n21924) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22224), .B1(
        n22232), .B2(n11061), .ZN(n21923) );
  OAI211_X1 U23477 ( .C1(n22227), .C2(n21947), .A(n21924), .B(n21923), .ZN(
        P1_U3050) );
  OAI22_X1 U23478 ( .A1(n22230), .A2(n11060), .B1(n21925), .B2(n22228), .ZN(
        n21926) );
  INV_X1 U23479 ( .A(n21926), .ZN(n21928) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22233), .B1(
        n22232), .B2(n21950), .ZN(n21927) );
  OAI211_X1 U23481 ( .C1(n22236), .C2(n21947), .A(n21928), .B(n21927), .ZN(
        P1_U3058) );
  AOI22_X1 U23482 ( .A1(n21953), .A2(n22238), .B1(n21954), .B2(n22237), .ZN(
        n21930) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n21950), .ZN(n21929) );
  OAI211_X1 U23484 ( .C1(n11060), .C2(n22248), .A(n21930), .B(n21929), .ZN(
        P1_U3066) );
  AOI22_X1 U23485 ( .A1(n22244), .A2(n21954), .B1(n21953), .B2(n22243), .ZN(
        n21932) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n11061), .ZN(n21931) );
  OAI211_X1 U23487 ( .C1(n21958), .C2(n22248), .A(n21932), .B(n21931), .ZN(
        P1_U3074) );
  AOI22_X1 U23488 ( .A1(n22257), .A2(n11061), .B1(n21953), .B2(n22249), .ZN(
        n21934) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22251), .B1(
        n22250), .B2(n21950), .ZN(n21933) );
  OAI211_X1 U23490 ( .C1(n22254), .C2(n21947), .A(n21934), .B(n21933), .ZN(
        P1_U3082) );
  AOI22_X1 U23491 ( .A1(n21953), .A2(n22256), .B1(n22255), .B2(n21954), .ZN(
        n21936) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n21950), .ZN(n21935) );
  OAI211_X1 U23493 ( .C1(n11060), .C2(n22261), .A(n21936), .B(n21935), .ZN(
        P1_U3090) );
  AOI22_X1 U23494 ( .A1(n22263), .A2(n21954), .B1(n21953), .B2(n22262), .ZN(
        n21938) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n21950), .ZN(n21937) );
  OAI211_X1 U23496 ( .C1(n11060), .C2(n22273), .A(n21938), .B(n21937), .ZN(
        P1_U3098) );
  AOI22_X1 U23497 ( .A1(n22269), .A2(n21954), .B1(n21953), .B2(n22268), .ZN(
        n21940) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n11061), .ZN(n21939) );
  OAI211_X1 U23499 ( .C1(n21958), .C2(n22273), .A(n21940), .B(n21939), .ZN(
        P1_U3106) );
  AOI22_X1 U23500 ( .A1(n22275), .A2(n21950), .B1(n22274), .B2(n21953), .ZN(
        n21942) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n11061), .ZN(n21941) );
  OAI211_X1 U23502 ( .C1(n22280), .C2(n21947), .A(n21942), .B(n21941), .ZN(
        P1_U3114) );
  AOI22_X1 U23503 ( .A1(n22282), .A2(n21954), .B1(n21953), .B2(n22281), .ZN(
        n21944) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n11061), .ZN(n21943) );
  OAI211_X1 U23505 ( .C1(n21958), .C2(n22286), .A(n21944), .B(n21943), .ZN(
        P1_U3122) );
  AOI22_X1 U23506 ( .A1(n22288), .A2(n11061), .B1(n21953), .B2(n22287), .ZN(
        n21946) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n21950), .ZN(n21945) );
  OAI211_X1 U23508 ( .C1(n22294), .C2(n21947), .A(n21946), .B(n21945), .ZN(
        P1_U3130) );
  AOI22_X1 U23509 ( .A1(n22296), .A2(n21954), .B1(n21953), .B2(n22295), .ZN(
        n21949) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n11061), .ZN(n21948) );
  OAI211_X1 U23511 ( .C1(n21958), .C2(n22300), .A(n21949), .B(n21948), .ZN(
        P1_U3138) );
  AOI22_X1 U23512 ( .A1(n21953), .A2(n22302), .B1(n21954), .B2(n22301), .ZN(
        n21952) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n21950), .ZN(n21951) );
  OAI211_X1 U23514 ( .C1(n11060), .C2(n22318), .A(n21952), .B(n21951), .ZN(
        P1_U3146) );
  AOI22_X1 U23515 ( .A1(n22312), .A2(n21954), .B1(n21953), .B2(n22309), .ZN(
        n21957) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n11061), .ZN(n21956) );
  OAI211_X1 U23517 ( .C1(n21958), .C2(n22318), .A(n21957), .B(n21956), .ZN(
        P1_U3154) );
  NAND2_X1 U23518 ( .A1(n22199), .A2(n21959), .ZN(n21994) );
  NOR2_X2 U23519 ( .A1(n22203), .A2(n13056), .ZN(n22001) );
  AOI22_X1 U23520 ( .A1(n22314), .A2(n21997), .B1(n22001), .B2(n22204), .ZN(
        n21965) );
  INV_X1 U23521 ( .A(DATAI_18_), .ZN(n21962) );
  OAI22_X1 U23522 ( .A1(n21963), .A2(n22207), .B1(n21962), .B2(n22205), .ZN(
        n22003) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n22003), .ZN(n21964) );
  OAI211_X1 U23524 ( .C1(n22212), .C2(n21994), .A(n21965), .B(n21964), .ZN(
        P1_U3035) );
  INV_X1 U23525 ( .A(n22003), .ZN(n22000) );
  INV_X1 U23526 ( .A(n21994), .ZN(n22002) );
  AOI22_X1 U23527 ( .A1(n22214), .A2(n22002), .B1(n22001), .B2(n22213), .ZN(
        n21967) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n21997), .ZN(n21966) );
  OAI211_X1 U23529 ( .C1(n22000), .C2(n22219), .A(n21967), .B(n21966), .ZN(
        P1_U3043) );
  INV_X1 U23530 ( .A(n21997), .ZN(n22006) );
  INV_X1 U23531 ( .A(n22001), .ZN(n21986) );
  OAI22_X1 U23532 ( .A1(n22219), .A2(n22006), .B1(n21986), .B2(n22220), .ZN(
        n21968) );
  INV_X1 U23533 ( .A(n21968), .ZN(n21970) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22224), .B1(
        n22232), .B2(n22003), .ZN(n21969) );
  OAI211_X1 U23535 ( .C1(n22227), .C2(n21994), .A(n21970), .B(n21969), .ZN(
        P1_U3051) );
  OAI22_X1 U23536 ( .A1(n22230), .A2(n22000), .B1(n21986), .B2(n22228), .ZN(
        n21971) );
  INV_X1 U23537 ( .A(n21971), .ZN(n21973) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22233), .B1(
        n22232), .B2(n21997), .ZN(n21972) );
  OAI211_X1 U23539 ( .C1(n22236), .C2(n21994), .A(n21973), .B(n21972), .ZN(
        P1_U3059) );
  AOI22_X1 U23540 ( .A1(n22001), .A2(n22238), .B1(n22002), .B2(n22237), .ZN(
        n21975) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n21997), .ZN(n21974) );
  OAI211_X1 U23542 ( .C1(n22000), .C2(n22248), .A(n21975), .B(n21974), .ZN(
        P1_U3067) );
  AOI22_X1 U23543 ( .A1(n22244), .A2(n22002), .B1(n22001), .B2(n22243), .ZN(
        n21977) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n22003), .ZN(n21976) );
  OAI211_X1 U23545 ( .C1(n22006), .C2(n22248), .A(n21977), .B(n21976), .ZN(
        P1_U3075) );
  AOI22_X1 U23546 ( .A1(n22257), .A2(n22003), .B1(n22001), .B2(n22249), .ZN(
        n21979) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22251), .B1(
        n22250), .B2(n21997), .ZN(n21978) );
  OAI211_X1 U23548 ( .C1(n22254), .C2(n21994), .A(n21979), .B(n21978), .ZN(
        P1_U3083) );
  AOI22_X1 U23549 ( .A1(n22001), .A2(n22256), .B1(n22255), .B2(n22002), .ZN(
        n21981) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n21997), .ZN(n21980) );
  OAI211_X1 U23551 ( .C1(n22000), .C2(n22261), .A(n21981), .B(n21980), .ZN(
        P1_U3091) );
  AOI22_X1 U23552 ( .A1(n22263), .A2(n22002), .B1(n22001), .B2(n22262), .ZN(
        n21983) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n21997), .ZN(n21982) );
  OAI211_X1 U23554 ( .C1(n22000), .C2(n22273), .A(n21983), .B(n21982), .ZN(
        P1_U3099) );
  AOI22_X1 U23555 ( .A1(n22269), .A2(n22002), .B1(n22001), .B2(n22268), .ZN(
        n21985) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n22003), .ZN(n21984) );
  OAI211_X1 U23557 ( .C1(n22006), .C2(n22273), .A(n21985), .B(n21984), .ZN(
        P1_U3107) );
  OAI22_X1 U23558 ( .A1(n22286), .A2(n22000), .B1(n22177), .B2(n21986), .ZN(
        n21987) );
  INV_X1 U23559 ( .A(n21987), .ZN(n21989) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22277), .B1(
        n22275), .B2(n21997), .ZN(n21988) );
  OAI211_X1 U23561 ( .C1(n22280), .C2(n21994), .A(n21989), .B(n21988), .ZN(
        P1_U3115) );
  AOI22_X1 U23562 ( .A1(n22282), .A2(n22002), .B1(n22001), .B2(n22281), .ZN(
        n21991) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22003), .ZN(n21990) );
  OAI211_X1 U23564 ( .C1(n22006), .C2(n22286), .A(n21991), .B(n21990), .ZN(
        P1_U3123) );
  AOI22_X1 U23565 ( .A1(n22288), .A2(n22003), .B1(n22001), .B2(n22287), .ZN(
        n21993) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n21997), .ZN(n21992) );
  OAI211_X1 U23567 ( .C1(n22294), .C2(n21994), .A(n21993), .B(n21992), .ZN(
        P1_U3131) );
  AOI22_X1 U23568 ( .A1(n22296), .A2(n22002), .B1(n22001), .B2(n22295), .ZN(
        n21996) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n22003), .ZN(n21995) );
  OAI211_X1 U23570 ( .C1(n22006), .C2(n22300), .A(n21996), .B(n21995), .ZN(
        P1_U3139) );
  AOI22_X1 U23571 ( .A1(n22001), .A2(n22302), .B1(n22002), .B2(n22301), .ZN(
        n21999) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n21997), .ZN(n21998) );
  OAI211_X1 U23573 ( .C1(n22000), .C2(n22318), .A(n21999), .B(n21998), .ZN(
        P1_U3147) );
  AOI22_X1 U23574 ( .A1(n22312), .A2(n22002), .B1(n22001), .B2(n22309), .ZN(
        n22005) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22003), .ZN(n22004) );
  OAI211_X1 U23576 ( .C1(n22006), .C2(n22318), .A(n22005), .B(n22004), .ZN(
        P1_U3155) );
  NAND2_X1 U23577 ( .A1(n22199), .A2(n22007), .ZN(n22041) );
  OAI22_X1 U23578 ( .A1(n22009), .A2(n22207), .B1(n22008), .B2(n22205), .ZN(
        n22044) );
  NOR2_X2 U23579 ( .A1(n22203), .A2(n12854), .ZN(n22048) );
  AOI22_X1 U23580 ( .A1(n22314), .A2(n22044), .B1(n22048), .B2(n22204), .ZN(
        n22013) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n22050), .ZN(n22012) );
  OAI211_X1 U23582 ( .C1(n22212), .C2(n22041), .A(n22013), .B(n22012), .ZN(
        P1_U3036) );
  INV_X1 U23583 ( .A(n22050), .ZN(n22047) );
  INV_X1 U23584 ( .A(n22041), .ZN(n22049) );
  AOI22_X1 U23585 ( .A1(n22214), .A2(n22049), .B1(n22048), .B2(n22213), .ZN(
        n22015) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n22044), .ZN(n22014) );
  OAI211_X1 U23587 ( .C1(n22047), .C2(n22219), .A(n22015), .B(n22014), .ZN(
        P1_U3044) );
  INV_X1 U23588 ( .A(n22220), .ZN(n22063) );
  AOI22_X1 U23589 ( .A1(n22232), .A2(n22050), .B1(n22048), .B2(n22063), .ZN(
        n22017) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22224), .B1(
        n22223), .B2(n22044), .ZN(n22016) );
  OAI211_X1 U23591 ( .C1(n22227), .C2(n22041), .A(n22017), .B(n22016), .ZN(
        P1_U3052) );
  INV_X1 U23592 ( .A(n22044), .ZN(n22053) );
  INV_X1 U23593 ( .A(n22048), .ZN(n22033) );
  OAI22_X1 U23594 ( .A1(n22221), .A2(n22053), .B1(n22033), .B2(n22228), .ZN(
        n22018) );
  INV_X1 U23595 ( .A(n22018), .ZN(n22020) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22233), .B1(
        n22239), .B2(n22050), .ZN(n22019) );
  OAI211_X1 U23597 ( .C1(n22236), .C2(n22041), .A(n22020), .B(n22019), .ZN(
        P1_U3060) );
  AOI22_X1 U23598 ( .A1(n22048), .A2(n22238), .B1(n22049), .B2(n22237), .ZN(
        n22022) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22044), .ZN(n22021) );
  OAI211_X1 U23600 ( .C1(n22047), .C2(n22248), .A(n22022), .B(n22021), .ZN(
        P1_U3068) );
  AOI22_X1 U23601 ( .A1(n22244), .A2(n22049), .B1(n22048), .B2(n22243), .ZN(
        n22024) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n22050), .ZN(n22023) );
  OAI211_X1 U23603 ( .C1(n22053), .C2(n22248), .A(n22024), .B(n22023), .ZN(
        P1_U3076) );
  AOI22_X1 U23604 ( .A1(n22250), .A2(n22044), .B1(n22048), .B2(n22249), .ZN(
        n22026) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22251), .B1(
        n22257), .B2(n22050), .ZN(n22025) );
  OAI211_X1 U23606 ( .C1(n22254), .C2(n22041), .A(n22026), .B(n22025), .ZN(
        P1_U3084) );
  AOI22_X1 U23607 ( .A1(n22048), .A2(n22256), .B1(n22255), .B2(n22049), .ZN(
        n22028) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22044), .ZN(n22027) );
  OAI211_X1 U23609 ( .C1(n22047), .C2(n22261), .A(n22028), .B(n22027), .ZN(
        P1_U3092) );
  AOI22_X1 U23610 ( .A1(n22263), .A2(n22049), .B1(n22048), .B2(n22262), .ZN(
        n22030) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22044), .ZN(n22029) );
  OAI211_X1 U23612 ( .C1(n22047), .C2(n22273), .A(n22030), .B(n22029), .ZN(
        P1_U3100) );
  AOI22_X1 U23613 ( .A1(n22269), .A2(n22049), .B1(n22048), .B2(n22268), .ZN(
        n22032) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n22050), .ZN(n22031) );
  OAI211_X1 U23615 ( .C1(n22053), .C2(n22273), .A(n22032), .B(n22031), .ZN(
        P1_U3108) );
  OAI22_X1 U23616 ( .A1(n22178), .A2(n22053), .B1(n22177), .B2(n22033), .ZN(
        n22034) );
  INV_X1 U23617 ( .A(n22034), .ZN(n22036) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n22050), .ZN(n22035) );
  OAI211_X1 U23619 ( .C1(n22280), .C2(n22041), .A(n22036), .B(n22035), .ZN(
        P1_U3116) );
  AOI22_X1 U23620 ( .A1(n22282), .A2(n22049), .B1(n22048), .B2(n22281), .ZN(
        n22038) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22050), .ZN(n22037) );
  OAI211_X1 U23622 ( .C1(n22053), .C2(n22286), .A(n22038), .B(n22037), .ZN(
        P1_U3124) );
  AOI22_X1 U23623 ( .A1(n22288), .A2(n22050), .B1(n22048), .B2(n22287), .ZN(
        n22040) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22044), .ZN(n22039) );
  OAI211_X1 U23625 ( .C1(n22294), .C2(n22041), .A(n22040), .B(n22039), .ZN(
        P1_U3132) );
  AOI22_X1 U23626 ( .A1(n22296), .A2(n22049), .B1(n22048), .B2(n22295), .ZN(
        n22043) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n22050), .ZN(n22042) );
  OAI211_X1 U23628 ( .C1(n22053), .C2(n22300), .A(n22043), .B(n22042), .ZN(
        P1_U3140) );
  AOI22_X1 U23629 ( .A1(n22048), .A2(n22302), .B1(n22049), .B2(n22301), .ZN(
        n22046) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n22044), .ZN(n22045) );
  OAI211_X1 U23631 ( .C1(n22047), .C2(n22318), .A(n22046), .B(n22045), .ZN(
        P1_U3148) );
  AOI22_X1 U23632 ( .A1(n22312), .A2(n22049), .B1(n22048), .B2(n22309), .ZN(
        n22052) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22050), .ZN(n22051) );
  OAI211_X1 U23634 ( .C1(n22053), .C2(n22318), .A(n22052), .B(n22051), .ZN(
        P1_U3156) );
  NAND2_X1 U23635 ( .A1(n22199), .A2(n22054), .ZN(n22089) );
  OAI22_X1 U23636 ( .A1(n22056), .A2(n22207), .B1(n22055), .B2(n22205), .ZN(
        n22092) );
  NOR2_X2 U23637 ( .A1(n22203), .A2(n12970), .ZN(n22095) );
  AOI22_X1 U23638 ( .A1(n22314), .A2(n22092), .B1(n22095), .B2(n22204), .ZN(
        n22060) );
  OAI22_X1 U23639 ( .A1(n22058), .A2(n22207), .B1(n22057), .B2(n22205), .ZN(
        n22097) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n11063), .ZN(n22059) );
  OAI211_X1 U23641 ( .C1(n22212), .C2(n22089), .A(n22060), .B(n22059), .ZN(
        P1_U3037) );
  INV_X1 U23642 ( .A(n22089), .ZN(n22096) );
  AOI22_X1 U23643 ( .A1(n22214), .A2(n22096), .B1(n22095), .B2(n22213), .ZN(
        n22062) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n22092), .ZN(n22061) );
  OAI211_X1 U23645 ( .C1(n11062), .C2(n22219), .A(n22062), .B(n22061), .ZN(
        P1_U3045) );
  AOI22_X1 U23646 ( .A1(n22232), .A2(n11063), .B1(n22095), .B2(n22063), .ZN(
        n22065) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22224), .B1(
        n22223), .B2(n22092), .ZN(n22064) );
  OAI211_X1 U23648 ( .C1(n22227), .C2(n22089), .A(n22065), .B(n22064), .ZN(
        P1_U3053) );
  INV_X1 U23649 ( .A(n22092), .ZN(n22100) );
  INV_X1 U23650 ( .A(n22095), .ZN(n22081) );
  OAI22_X1 U23651 ( .A1(n22221), .A2(n22100), .B1(n22081), .B2(n22228), .ZN(
        n22066) );
  INV_X1 U23652 ( .A(n22066), .ZN(n22068) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22233), .B1(
        n22239), .B2(n11063), .ZN(n22067) );
  OAI211_X1 U23654 ( .C1(n22236), .C2(n22089), .A(n22068), .B(n22067), .ZN(
        P1_U3061) );
  AOI22_X1 U23655 ( .A1(n22095), .A2(n22238), .B1(n22096), .B2(n22237), .ZN(
        n22070) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22092), .ZN(n22069) );
  OAI211_X1 U23657 ( .C1(n11062), .C2(n22248), .A(n22070), .B(n22069), .ZN(
        P1_U3069) );
  AOI22_X1 U23658 ( .A1(n22244), .A2(n22096), .B1(n22095), .B2(n22243), .ZN(
        n22072) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n11063), .ZN(n22071) );
  OAI211_X1 U23660 ( .C1(n22100), .C2(n22248), .A(n22072), .B(n22071), .ZN(
        P1_U3077) );
  AOI22_X1 U23661 ( .A1(n22250), .A2(n22092), .B1(n22095), .B2(n22249), .ZN(
        n22074) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22251), .B1(
        n22257), .B2(n11063), .ZN(n22073) );
  OAI211_X1 U23663 ( .C1(n22254), .C2(n22089), .A(n22074), .B(n22073), .ZN(
        P1_U3085) );
  AOI22_X1 U23664 ( .A1(n22095), .A2(n22256), .B1(n22255), .B2(n22096), .ZN(
        n22076) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22092), .ZN(n22075) );
  OAI211_X1 U23666 ( .C1(n11062), .C2(n22261), .A(n22076), .B(n22075), .ZN(
        P1_U3093) );
  AOI22_X1 U23667 ( .A1(n22263), .A2(n22096), .B1(n22095), .B2(n22262), .ZN(
        n22078) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22092), .ZN(n22077) );
  OAI211_X1 U23669 ( .C1(n11062), .C2(n22273), .A(n22078), .B(n22077), .ZN(
        P1_U3101) );
  AOI22_X1 U23670 ( .A1(n22269), .A2(n22096), .B1(n22095), .B2(n22268), .ZN(
        n22080) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n11063), .ZN(n22079) );
  OAI211_X1 U23672 ( .C1(n22100), .C2(n22273), .A(n22080), .B(n22079), .ZN(
        P1_U3109) );
  OAI22_X1 U23673 ( .A1(n22178), .A2(n22100), .B1(n22177), .B2(n22081), .ZN(
        n22082) );
  INV_X1 U23674 ( .A(n22082), .ZN(n22084) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n11063), .ZN(n22083) );
  OAI211_X1 U23676 ( .C1(n22280), .C2(n22089), .A(n22084), .B(n22083), .ZN(
        P1_U3117) );
  AOI22_X1 U23677 ( .A1(n22282), .A2(n22096), .B1(n22095), .B2(n22281), .ZN(
        n22086) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n11063), .ZN(n22085) );
  OAI211_X1 U23679 ( .C1(n22100), .C2(n22286), .A(n22086), .B(n22085), .ZN(
        P1_U3125) );
  AOI22_X1 U23680 ( .A1(n22288), .A2(n11063), .B1(n22095), .B2(n22287), .ZN(
        n22088) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22092), .ZN(n22087) );
  OAI211_X1 U23682 ( .C1(n22294), .C2(n22089), .A(n22088), .B(n22087), .ZN(
        P1_U3133) );
  AOI22_X1 U23683 ( .A1(n22296), .A2(n22096), .B1(n22095), .B2(n22295), .ZN(
        n22091) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n11063), .ZN(n22090) );
  OAI211_X1 U23685 ( .C1(n22100), .C2(n22300), .A(n22091), .B(n22090), .ZN(
        P1_U3141) );
  AOI22_X1 U23686 ( .A1(n22095), .A2(n22302), .B1(n22096), .B2(n22301), .ZN(
        n22094) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n22092), .ZN(n22093) );
  OAI211_X1 U23688 ( .C1(n11062), .C2(n22318), .A(n22094), .B(n22093), .ZN(
        P1_U3149) );
  AOI22_X1 U23689 ( .A1(n22312), .A2(n22096), .B1(n22095), .B2(n22309), .ZN(
        n22099) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n11063), .ZN(n22098) );
  OAI211_X1 U23691 ( .C1(n22100), .C2(n22318), .A(n22099), .B(n22098), .ZN(
        P1_U3157) );
  NAND2_X1 U23692 ( .A1(n22199), .A2(n22101), .ZN(n22137) );
  INV_X1 U23693 ( .A(DATAI_29_), .ZN(n22102) );
  OAI22_X1 U23694 ( .A1(n22103), .A2(n22207), .B1(n22102), .B2(n22205), .ZN(
        n22140) );
  NOR2_X2 U23695 ( .A1(n22203), .A2(n22104), .ZN(n22144) );
  AOI22_X1 U23696 ( .A1(n22314), .A2(n11059), .B1(n22144), .B2(n22204), .ZN(
        n22108) );
  OAI22_X1 U23697 ( .A1(n22106), .A2(n22207), .B1(n22105), .B2(n22205), .ZN(
        n22146) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n22146), .ZN(n22107) );
  OAI211_X1 U23699 ( .C1(n22212), .C2(n22137), .A(n22108), .B(n22107), .ZN(
        P1_U3038) );
  INV_X1 U23700 ( .A(n22146), .ZN(n22143) );
  INV_X1 U23701 ( .A(n22137), .ZN(n22145) );
  AOI22_X1 U23702 ( .A1(n22214), .A2(n22145), .B1(n22144), .B2(n22213), .ZN(
        n22110) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n11059), .ZN(n22109) );
  OAI211_X1 U23704 ( .C1(n22143), .C2(n22219), .A(n22110), .B(n22109), .ZN(
        P1_U3046) );
  INV_X1 U23705 ( .A(n22144), .ZN(n22129) );
  OAI22_X1 U23706 ( .A1(n22219), .A2(n11058), .B1(n22129), .B2(n22220), .ZN(
        n22111) );
  INV_X1 U23707 ( .A(n22111), .ZN(n22113) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22224), .B1(
        n22232), .B2(n22146), .ZN(n22112) );
  OAI211_X1 U23709 ( .C1(n22227), .C2(n22137), .A(n22113), .B(n22112), .ZN(
        P1_U3054) );
  OAI22_X1 U23710 ( .A1(n22230), .A2(n22143), .B1(n22129), .B2(n22228), .ZN(
        n22114) );
  INV_X1 U23711 ( .A(n22114), .ZN(n22116) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22233), .B1(
        n22232), .B2(n11059), .ZN(n22115) );
  OAI211_X1 U23713 ( .C1(n22236), .C2(n22137), .A(n22116), .B(n22115), .ZN(
        P1_U3062) );
  AOI22_X1 U23714 ( .A1(n22144), .A2(n22238), .B1(n22145), .B2(n22237), .ZN(
        n22118) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n11059), .ZN(n22117) );
  OAI211_X1 U23716 ( .C1(n22143), .C2(n22248), .A(n22118), .B(n22117), .ZN(
        P1_U3070) );
  AOI22_X1 U23717 ( .A1(n22244), .A2(n22145), .B1(n22144), .B2(n22243), .ZN(
        n22120) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n22146), .ZN(n22119) );
  OAI211_X1 U23719 ( .C1(n11058), .C2(n22248), .A(n22120), .B(n22119), .ZN(
        P1_U3078) );
  AOI22_X1 U23720 ( .A1(n22257), .A2(n22146), .B1(n22144), .B2(n22249), .ZN(
        n22122) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22251), .B1(
        n22250), .B2(n11059), .ZN(n22121) );
  OAI211_X1 U23722 ( .C1(n22254), .C2(n22137), .A(n22122), .B(n22121), .ZN(
        P1_U3086) );
  AOI22_X1 U23723 ( .A1(n22144), .A2(n22256), .B1(n22255), .B2(n22145), .ZN(
        n22124) );
  AOI22_X1 U23724 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n11059), .ZN(n22123) );
  OAI211_X1 U23725 ( .C1(n22143), .C2(n22261), .A(n22124), .B(n22123), .ZN(
        P1_U3094) );
  AOI22_X1 U23726 ( .A1(n22263), .A2(n22145), .B1(n22144), .B2(n22262), .ZN(
        n22126) );
  AOI22_X1 U23727 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n11059), .ZN(n22125) );
  OAI211_X1 U23728 ( .C1(n22143), .C2(n22273), .A(n22126), .B(n22125), .ZN(
        P1_U3102) );
  AOI22_X1 U23729 ( .A1(n22269), .A2(n22145), .B1(n22144), .B2(n22268), .ZN(
        n22128) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n22146), .ZN(n22127) );
  OAI211_X1 U23731 ( .C1(n11058), .C2(n22273), .A(n22128), .B(n22127), .ZN(
        P1_U3110) );
  OAI22_X1 U23732 ( .A1(n22286), .A2(n22143), .B1(n22177), .B2(n22129), .ZN(
        n22130) );
  INV_X1 U23733 ( .A(n22130), .ZN(n22132) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22277), .B1(
        n22275), .B2(n11059), .ZN(n22131) );
  OAI211_X1 U23735 ( .C1(n22280), .C2(n22137), .A(n22132), .B(n22131), .ZN(
        P1_U3118) );
  AOI22_X1 U23736 ( .A1(n22282), .A2(n22145), .B1(n22144), .B2(n22281), .ZN(
        n22134) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22146), .ZN(n22133) );
  OAI211_X1 U23738 ( .C1(n11058), .C2(n22286), .A(n22134), .B(n22133), .ZN(
        P1_U3126) );
  AOI22_X1 U23739 ( .A1(n22288), .A2(n22146), .B1(n22144), .B2(n22287), .ZN(
        n22136) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n11059), .ZN(n22135) );
  OAI211_X1 U23741 ( .C1(n22294), .C2(n22137), .A(n22136), .B(n22135), .ZN(
        P1_U3134) );
  AOI22_X1 U23742 ( .A1(n22296), .A2(n22145), .B1(n22144), .B2(n22295), .ZN(
        n22139) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n22146), .ZN(n22138) );
  OAI211_X1 U23744 ( .C1(n11058), .C2(n22300), .A(n22139), .B(n22138), .ZN(
        P1_U3142) );
  AOI22_X1 U23745 ( .A1(n22144), .A2(n22302), .B1(n22145), .B2(n22301), .ZN(
        n22142) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n11059), .ZN(n22141) );
  OAI211_X1 U23747 ( .C1(n22143), .C2(n22318), .A(n22142), .B(n22141), .ZN(
        P1_U3150) );
  AOI22_X1 U23748 ( .A1(n22312), .A2(n22145), .B1(n22144), .B2(n22309), .ZN(
        n22148) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22146), .ZN(n22147) );
  OAI211_X1 U23750 ( .C1(n11058), .C2(n22318), .A(n22148), .B(n22147), .ZN(
        P1_U3158) );
  NAND2_X1 U23751 ( .A1(n22199), .A2(n22149), .ZN(n22186) );
  INV_X1 U23752 ( .A(DATAI_30_), .ZN(n22150) );
  OAI22_X1 U23753 ( .A1(n22151), .A2(n22207), .B1(n22150), .B2(n22205), .ZN(
        n22189) );
  NOR2_X2 U23754 ( .A1(n22203), .A2(n12963), .ZN(n22192) );
  AOI22_X1 U23755 ( .A1(n22314), .A2(n22189), .B1(n22192), .B2(n22204), .ZN(
        n22155) );
  OAI22_X1 U23756 ( .A1(n22153), .A2(n22207), .B1(n22152), .B2(n22205), .ZN(
        n22194) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n11065), .ZN(n22154) );
  OAI211_X1 U23758 ( .C1(n22212), .C2(n22186), .A(n22155), .B(n22154), .ZN(
        P1_U3039) );
  INV_X1 U23759 ( .A(n22186), .ZN(n22193) );
  AOI22_X1 U23760 ( .A1(n22214), .A2(n22193), .B1(n22192), .B2(n22213), .ZN(
        n22157) );
  AOI22_X1 U23761 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n22189), .ZN(n22156) );
  OAI211_X1 U23762 ( .C1(n11064), .C2(n22219), .A(n22157), .B(n22156), .ZN(
        P1_U3047) );
  INV_X1 U23763 ( .A(n22189), .ZN(n22197) );
  INV_X1 U23764 ( .A(n22192), .ZN(n22176) );
  OAI22_X1 U23765 ( .A1(n22219), .A2(n22197), .B1(n22176), .B2(n22220), .ZN(
        n22158) );
  INV_X1 U23766 ( .A(n22158), .ZN(n22160) );
  AOI22_X1 U23767 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22224), .B1(
        n22232), .B2(n11065), .ZN(n22159) );
  OAI211_X1 U23768 ( .C1(n22227), .C2(n22186), .A(n22160), .B(n22159), .ZN(
        P1_U3055) );
  OAI22_X1 U23769 ( .A1(n22221), .A2(n22197), .B1(n22176), .B2(n22228), .ZN(
        n22161) );
  INV_X1 U23770 ( .A(n22161), .ZN(n22163) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22233), .B1(
        n22239), .B2(n11065), .ZN(n22162) );
  OAI211_X1 U23772 ( .C1(n22236), .C2(n22186), .A(n22163), .B(n22162), .ZN(
        P1_U3063) );
  AOI22_X1 U23773 ( .A1(n22192), .A2(n22238), .B1(n22193), .B2(n22237), .ZN(
        n22165) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22189), .ZN(n22164) );
  OAI211_X1 U23775 ( .C1(n11064), .C2(n22248), .A(n22165), .B(n22164), .ZN(
        P1_U3071) );
  AOI22_X1 U23776 ( .A1(n22244), .A2(n22193), .B1(n22192), .B2(n22243), .ZN(
        n22167) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n11065), .ZN(n22166) );
  OAI211_X1 U23778 ( .C1(n22197), .C2(n22248), .A(n22167), .B(n22166), .ZN(
        P1_U3079) );
  AOI22_X1 U23779 ( .A1(n22257), .A2(n11065), .B1(n22192), .B2(n22249), .ZN(
        n22169) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22251), .B1(
        n22250), .B2(n22189), .ZN(n22168) );
  OAI211_X1 U23781 ( .C1(n22254), .C2(n22186), .A(n22169), .B(n22168), .ZN(
        P1_U3087) );
  AOI22_X1 U23782 ( .A1(n22192), .A2(n22256), .B1(n22255), .B2(n22193), .ZN(
        n22171) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22189), .ZN(n22170) );
  OAI211_X1 U23784 ( .C1(n11064), .C2(n22261), .A(n22171), .B(n22170), .ZN(
        P1_U3095) );
  AOI22_X1 U23785 ( .A1(n22263), .A2(n22193), .B1(n22192), .B2(n22262), .ZN(
        n22173) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22189), .ZN(n22172) );
  OAI211_X1 U23787 ( .C1(n11064), .C2(n22273), .A(n22173), .B(n22172), .ZN(
        P1_U3103) );
  AOI22_X1 U23788 ( .A1(n22269), .A2(n22193), .B1(n22192), .B2(n22268), .ZN(
        n22175) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n11065), .ZN(n22174) );
  OAI211_X1 U23790 ( .C1(n22197), .C2(n22273), .A(n22175), .B(n22174), .ZN(
        P1_U3111) );
  OAI22_X1 U23791 ( .A1(n22178), .A2(n22197), .B1(n22177), .B2(n22176), .ZN(
        n22179) );
  INV_X1 U23792 ( .A(n22179), .ZN(n22181) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n11065), .ZN(n22180) );
  OAI211_X1 U23794 ( .C1(n22280), .C2(n22186), .A(n22181), .B(n22180), .ZN(
        P1_U3119) );
  AOI22_X1 U23795 ( .A1(n22282), .A2(n22193), .B1(n22192), .B2(n22281), .ZN(
        n22183) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n11065), .ZN(n22182) );
  OAI211_X1 U23797 ( .C1(n22197), .C2(n22286), .A(n22183), .B(n22182), .ZN(
        P1_U3127) );
  AOI22_X1 U23798 ( .A1(n22288), .A2(n11065), .B1(n22192), .B2(n22287), .ZN(
        n22185) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22189), .ZN(n22184) );
  OAI211_X1 U23800 ( .C1(n22294), .C2(n22186), .A(n22185), .B(n22184), .ZN(
        P1_U3135) );
  AOI22_X1 U23801 ( .A1(n22296), .A2(n22193), .B1(n22192), .B2(n22295), .ZN(
        n22188) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n11065), .ZN(n22187) );
  OAI211_X1 U23803 ( .C1(n22197), .C2(n22300), .A(n22188), .B(n22187), .ZN(
        P1_U3143) );
  AOI22_X1 U23804 ( .A1(n22192), .A2(n22302), .B1(n22193), .B2(n22301), .ZN(
        n22191) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n22189), .ZN(n22190) );
  OAI211_X1 U23806 ( .C1(n11064), .C2(n22318), .A(n22191), .B(n22190), .ZN(
        P1_U3151) );
  AOI22_X1 U23807 ( .A1(n22312), .A2(n22193), .B1(n22192), .B2(n22309), .ZN(
        n22196) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n11065), .ZN(n22195) );
  OAI211_X1 U23809 ( .C1(n22197), .C2(n22318), .A(n22196), .B(n22195), .ZN(
        P1_U3159) );
  NAND2_X1 U23810 ( .A1(n22199), .A2(n22198), .ZN(n22293) );
  INV_X1 U23811 ( .A(DATAI_31_), .ZN(n22200) );
  OAI22_X1 U23812 ( .A1(n22201), .A2(n22207), .B1(n22200), .B2(n22205), .ZN(
        n22303) );
  NOR2_X2 U23813 ( .A1(n22203), .A2(n22202), .ZN(n22310) );
  AOI22_X1 U23814 ( .A1(n22314), .A2(n11067), .B1(n22310), .B2(n22204), .ZN(
        n22211) );
  OAI22_X1 U23815 ( .A1(n22208), .A2(n22207), .B1(n22206), .B2(n22205), .ZN(
        n22313) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22209), .B1(
        n22215), .B2(n22313), .ZN(n22210) );
  OAI211_X1 U23817 ( .C1(n22212), .C2(n22293), .A(n22211), .B(n22210), .ZN(
        P1_U3040) );
  INV_X1 U23818 ( .A(n22313), .ZN(n22308) );
  INV_X1 U23819 ( .A(n22293), .ZN(n22311) );
  AOI22_X1 U23820 ( .A1(n22214), .A2(n22311), .B1(n22310), .B2(n22213), .ZN(
        n22218) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22216), .B1(
        n22215), .B2(n11067), .ZN(n22217) );
  OAI211_X1 U23822 ( .C1(n22308), .C2(n22219), .A(n22218), .B(n22217), .ZN(
        P1_U3048) );
  INV_X1 U23823 ( .A(n22310), .ZN(n22229) );
  OAI22_X1 U23824 ( .A1(n22221), .A2(n22308), .B1(n22229), .B2(n22220), .ZN(
        n22222) );
  INV_X1 U23825 ( .A(n22222), .ZN(n22226) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22224), .B1(
        n22223), .B2(n11067), .ZN(n22225) );
  OAI211_X1 U23827 ( .C1(n22227), .C2(n22293), .A(n22226), .B(n22225), .ZN(
        P1_U3056) );
  OAI22_X1 U23828 ( .A1(n22230), .A2(n22308), .B1(n22229), .B2(n22228), .ZN(
        n22231) );
  INV_X1 U23829 ( .A(n22231), .ZN(n22235) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22233), .B1(
        n22232), .B2(n11067), .ZN(n22234) );
  OAI211_X1 U23831 ( .C1(n22236), .C2(n22293), .A(n22235), .B(n22234), .ZN(
        P1_U3064) );
  AOI22_X1 U23832 ( .A1(n22310), .A2(n22238), .B1(n22311), .B2(n22237), .ZN(
        n22242) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n11067), .ZN(n22241) );
  OAI211_X1 U23834 ( .C1(n22308), .C2(n22248), .A(n22242), .B(n22241), .ZN(
        P1_U3072) );
  AOI22_X1 U23835 ( .A1(n22244), .A2(n22311), .B1(n22310), .B2(n22243), .ZN(
        n22247) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22245), .B1(
        n22250), .B2(n22313), .ZN(n22246) );
  OAI211_X1 U23837 ( .C1(n11066), .C2(n22248), .A(n22247), .B(n22246), .ZN(
        P1_U3080) );
  AOI22_X1 U23838 ( .A1(n22257), .A2(n22313), .B1(n22310), .B2(n22249), .ZN(
        n22253) );
  AOI22_X1 U23839 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22251), .B1(
        n22250), .B2(n11067), .ZN(n22252) );
  OAI211_X1 U23840 ( .C1(n22254), .C2(n22293), .A(n22253), .B(n22252), .ZN(
        P1_U3088) );
  AOI22_X1 U23841 ( .A1(n22310), .A2(n22256), .B1(n22255), .B2(n22311), .ZN(
        n22260) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n11067), .ZN(n22259) );
  OAI211_X1 U23843 ( .C1(n22308), .C2(n22261), .A(n22260), .B(n22259), .ZN(
        P1_U3096) );
  AOI22_X1 U23844 ( .A1(n22263), .A2(n22311), .B1(n22310), .B2(n22262), .ZN(
        n22267) );
  AOI22_X1 U23845 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n11067), .ZN(n22266) );
  OAI211_X1 U23846 ( .C1(n22308), .C2(n22273), .A(n22267), .B(n22266), .ZN(
        P1_U3104) );
  AOI22_X1 U23847 ( .A1(n22269), .A2(n22311), .B1(n22310), .B2(n22268), .ZN(
        n22272) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22270), .B1(
        n22275), .B2(n22313), .ZN(n22271) );
  OAI211_X1 U23849 ( .C1(n11066), .C2(n22273), .A(n22272), .B(n22271), .ZN(
        P1_U3112) );
  AOI22_X1 U23850 ( .A1(n22275), .A2(n11067), .B1(n22274), .B2(n22310), .ZN(
        n22279) );
  AOI22_X1 U23851 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22277), .B1(
        n22276), .B2(n22313), .ZN(n22278) );
  OAI211_X1 U23852 ( .C1(n22280), .C2(n22293), .A(n22279), .B(n22278), .ZN(
        P1_U3120) );
  AOI22_X1 U23853 ( .A1(n22282), .A2(n22311), .B1(n22310), .B2(n22281), .ZN(
        n22285) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22313), .ZN(n22284) );
  OAI211_X1 U23855 ( .C1(n11066), .C2(n22286), .A(n22285), .B(n22284), .ZN(
        P1_U3128) );
  AOI22_X1 U23856 ( .A1(n22288), .A2(n22313), .B1(n22310), .B2(n22287), .ZN(
        n22292) );
  AOI22_X1 U23857 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n11067), .ZN(n22291) );
  OAI211_X1 U23858 ( .C1(n22294), .C2(n22293), .A(n22292), .B(n22291), .ZN(
        P1_U3136) );
  AOI22_X1 U23859 ( .A1(n22296), .A2(n22311), .B1(n22310), .B2(n22295), .ZN(
        n22299) );
  AOI22_X1 U23860 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22297), .B1(
        n22304), .B2(n22313), .ZN(n22298) );
  OAI211_X1 U23861 ( .C1(n11066), .C2(n22300), .A(n22299), .B(n22298), .ZN(
        P1_U3144) );
  AOI22_X1 U23862 ( .A1(n22310), .A2(n22302), .B1(n22311), .B2(n22301), .ZN(
        n22307) );
  AOI22_X1 U23863 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22305), .B1(
        n22304), .B2(n11067), .ZN(n22306) );
  OAI211_X1 U23864 ( .C1(n22308), .C2(n22318), .A(n22307), .B(n22306), .ZN(
        P1_U3152) );
  AOI22_X1 U23865 ( .A1(n22312), .A2(n22311), .B1(n22310), .B2(n22309), .ZN(
        n22317) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22315), .B1(
        n22314), .B2(n22313), .ZN(n22316) );
  OAI211_X1 U23867 ( .C1(n11066), .C2(n22318), .A(n22317), .B(n22316), .ZN(
        P1_U3160) );
  OAI22_X1 U23868 ( .A1(n11057), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22319), .ZN(n22320) );
  INV_X1 U23869 ( .A(n22320), .ZN(P1_U3486) );
  AND2_X1 U12552 ( .A1(n11886), .A2(n11084), .ZN(n12422) );
  CLKBUF_X1 U11089 ( .A(n13046), .Z(n13000) );
  CLKBUF_X1 U11143 ( .A(n14067), .Z(n10979) );
  NOR2_X2 U11181 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11260) );
  CLKBUF_X1 U11277 ( .A(n12973), .Z(n13442) );
  NOR2_X2 U11423 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14063) );
  CLKBUF_X1 U11452 ( .A(n15352), .Z(n15436) );
  CLKBUF_X1 U12042 ( .A(n17095), .Z(n17107) );
  CLKBUF_X1 U12194 ( .A(n11871), .Z(n15968) );
  CLKBUF_X2 U12277 ( .A(n11935), .Z(n11940) );
  CLKBUF_X1 U12279 ( .A(n17982), .Z(n17989) );
  CLKBUF_X1 U12843 ( .A(n20077), .Z(n20075) );
  OAI22_X1 U13377 ( .A1(n14839), .A2(n20995), .B1(n11719), .B2(n21132), .ZN(
        n21163) );
  CLKBUF_X2 U14715 ( .A(n20071), .Z(n20078) );
endmodule

